magic
tech EFS8A
magscale 1 2
timestamp 1603466439
<< viali >>
rect 20453 9469 20487 9503
rect 20177 9333 20211 9367
rect 20821 9333 20855 9367
rect 16497 8993 16531 9027
rect 23029 8993 23063 9027
rect 10057 8789 10091 8823
rect 16681 8789 16715 8823
rect 22845 8789 22879 8823
rect 16497 8585 16531 8619
rect 22661 8517 22695 8551
rect 9505 8449 9539 8483
rect 10241 8381 10275 8415
rect 10425 8381 10459 8415
rect 10793 8381 10827 8415
rect 11345 8381 11379 8415
rect 22477 8381 22511 8415
rect 9873 8313 9907 8347
rect 23029 8313 23063 8347
rect 23397 8313 23431 8347
rect 10057 8245 10091 8279
rect 10425 7973 10459 8007
rect 10793 7905 10827 7939
rect 11161 7905 11195 7939
rect 11345 7905 11379 7939
rect 11897 7905 11931 7939
rect 11897 7769 11931 7803
rect 10057 7701 10091 7735
rect 19717 7701 19751 7735
rect 9045 7497 9079 7531
rect 11345 7497 11379 7531
rect 11713 7497 11747 7531
rect 8677 7361 8711 7395
rect 9413 7293 9447 7327
rect 9781 7293 9815 7327
rect 10241 7293 10275 7327
rect 10517 7293 10551 7327
rect 10885 7293 10919 7327
rect 12081 7293 12115 7327
rect 20453 7293 20487 7327
rect 19717 7225 19751 7259
rect 19901 7225 19935 7259
rect 20085 7225 20119 7259
rect 9781 7157 9815 7191
rect 19165 7157 19199 7191
rect 19625 7157 19659 7191
rect 19993 7157 20027 7191
rect 9781 6953 9815 6987
rect 19809 6953 19843 6987
rect 21097 6953 21131 6987
rect 21281 6885 21315 6919
rect 22753 6885 22787 6919
rect 22937 6885 22971 6919
rect 9873 6817 9907 6851
rect 10333 6817 10367 6851
rect 10517 6817 10551 6851
rect 10885 6817 10919 6851
rect 21189 6817 21223 6851
rect 22845 6817 22879 6851
rect 20913 6749 20947 6783
rect 21649 6749 21683 6783
rect 22569 6749 22603 6783
rect 23305 6749 23339 6783
rect 24409 6681 24443 6715
rect 9413 6409 9447 6443
rect 9781 6409 9815 6443
rect 10517 6409 10551 6443
rect 20545 6409 20579 6443
rect 21373 6409 21407 6443
rect 22293 6409 22327 6443
rect 10793 6341 10827 6375
rect 22661 6341 22695 6375
rect 10149 6273 10183 6307
rect 24133 6273 24167 6307
rect 20913 6205 20947 6239
rect 21741 6205 21775 6239
rect 23029 6205 23063 6239
rect 24501 6205 24535 6239
rect 23397 6137 23431 6171
rect 24317 6137 24351 6171
rect 24685 6137 24719 6171
rect 25053 6137 25087 6171
rect 24593 6069 24627 6103
rect 24409 5865 24443 5899
rect 24685 5797 24719 5831
rect 3065 5117 3099 5151
rect 2973 5049 3007 5083
rect 3427 5049 3461 5083
rect 3985 4981 4019 5015
rect 25237 4777 25271 4811
rect 5870 4709 5904 4743
rect 5549 4641 5583 4675
rect 3157 4573 3191 4607
rect 6469 4437 6503 4471
rect 6009 4233 6043 4267
rect 9137 4097 9171 4131
rect 18061 4097 18095 4131
rect 20545 4097 20579 4131
rect 21005 4097 21039 4131
rect 25237 4097 25271 4131
rect 3157 4029 3191 4063
rect 5641 4029 5675 4063
rect 3065 3961 3099 3995
rect 3519 3961 3553 3995
rect 9045 3961 9079 3995
rect 9499 3961 9533 3995
rect 17785 3961 17819 3995
rect 18382 3961 18416 3995
rect 20821 3961 20855 3995
rect 21326 3961 21360 3995
rect 25558 3961 25592 3995
rect 4077 3893 4111 3927
rect 10057 3893 10091 3927
rect 18981 3893 19015 3927
rect 21925 3893 21959 3927
rect 25053 3893 25087 3927
rect 26157 3893 26191 3927
rect 2053 3689 2087 3723
rect 3249 3689 3283 3723
rect 9137 3689 9171 3723
rect 18153 3689 18187 3723
rect 24362 3621 24396 3655
rect 1409 3553 1443 3587
rect 24041 3553 24075 3587
rect 1593 3349 1627 3383
rect 24961 3349 24995 3383
rect 25237 3349 25271 3383
rect 2789 3145 2823 3179
rect 17141 3145 17175 3179
rect 22201 3145 22235 3179
rect 24409 3145 24443 3179
rect 25697 3145 25731 3179
rect 2053 3077 2087 3111
rect 21741 3077 21775 3111
rect 24133 3077 24167 3111
rect 1593 3009 1627 3043
rect 25237 3009 25271 3043
rect 1409 2941 1443 2975
rect 16497 2941 16531 2975
rect 21557 2941 21591 2975
rect 24961 2941 24995 2975
rect 25053 2941 25087 2975
rect 2421 2805 2455 2839
rect 16681 2805 16715 2839
rect 2053 2601 2087 2635
rect 2789 2601 2823 2635
rect 3525 2601 3559 2635
rect 4997 2601 5031 2635
rect 7113 2601 7147 2635
rect 7573 2601 7607 2635
rect 16773 2601 16807 2635
rect 21833 2601 21867 2635
rect 24869 2601 24903 2635
rect 26249 2601 26283 2635
rect 1593 2465 1627 2499
rect 2881 2465 2915 2499
rect 5089 2465 5123 2499
rect 5273 2465 5307 2499
rect 5733 2465 5767 2499
rect 6929 2465 6963 2499
rect 9229 2465 9263 2499
rect 9965 2465 9999 2499
rect 10425 2465 10459 2499
rect 11253 2465 11287 2499
rect 11897 2465 11931 2499
rect 15301 2465 15335 2499
rect 16313 2465 16347 2499
rect 20637 2465 20671 2499
rect 21373 2465 21407 2499
rect 24225 2465 24259 2499
rect 25237 2465 25271 2499
rect 25329 2465 25363 2499
rect 25513 2465 25547 2499
rect 26893 2465 26927 2499
rect 1409 2397 1443 2431
rect 4629 2397 4663 2431
rect 9597 2397 9631 2431
rect 9781 2397 9815 2431
rect 16129 2397 16163 2431
rect 21005 2397 21039 2431
rect 21189 2397 21223 2431
rect 25973 2397 26007 2431
rect 2329 2329 2363 2363
rect 27077 2329 27111 2363
rect 3065 2261 3099 2295
rect 11437 2261 11471 2295
rect 16037 2261 16071 2295
rect 24409 2261 24443 2295
rect 27537 2261 27571 2295
<< metal1 >>
rect 1104 13626 38824 13648
rect 1104 13574 14315 13626
rect 14367 13574 14379 13626
rect 14431 13574 14443 13626
rect 14495 13574 14507 13626
rect 14559 13574 27648 13626
rect 27700 13574 27712 13626
rect 27764 13574 27776 13626
rect 27828 13574 27840 13626
rect 27892 13574 38824 13626
rect 1104 13552 38824 13574
rect 1104 13082 38824 13104
rect 1104 13030 7648 13082
rect 7700 13030 7712 13082
rect 7764 13030 7776 13082
rect 7828 13030 7840 13082
rect 7892 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 34315 13082
rect 34367 13030 34379 13082
rect 34431 13030 34443 13082
rect 34495 13030 34507 13082
rect 34559 13030 38824 13082
rect 1104 13008 38824 13030
rect 1104 12538 38824 12560
rect 1104 12486 14315 12538
rect 14367 12486 14379 12538
rect 14431 12486 14443 12538
rect 14495 12486 14507 12538
rect 14559 12486 27648 12538
rect 27700 12486 27712 12538
rect 27764 12486 27776 12538
rect 27828 12486 27840 12538
rect 27892 12486 38824 12538
rect 1104 12464 38824 12486
rect 1104 11994 38824 12016
rect 1104 11942 7648 11994
rect 7700 11942 7712 11994
rect 7764 11942 7776 11994
rect 7828 11942 7840 11994
rect 7892 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 34315 11994
rect 34367 11942 34379 11994
rect 34431 11942 34443 11994
rect 34495 11942 34507 11994
rect 34559 11942 38824 11994
rect 1104 11920 38824 11942
rect 1104 11450 38824 11472
rect 1104 11398 14315 11450
rect 14367 11398 14379 11450
rect 14431 11398 14443 11450
rect 14495 11398 14507 11450
rect 14559 11398 27648 11450
rect 27700 11398 27712 11450
rect 27764 11398 27776 11450
rect 27828 11398 27840 11450
rect 27892 11398 38824 11450
rect 1104 11376 38824 11398
rect 26234 11228 26240 11280
rect 26292 11268 26298 11280
rect 27430 11268 27436 11280
rect 26292 11240 27436 11268
rect 26292 11228 26298 11240
rect 27430 11228 27436 11240
rect 27488 11228 27494 11280
rect 1104 10906 38824 10928
rect 1104 10854 7648 10906
rect 7700 10854 7712 10906
rect 7764 10854 7776 10906
rect 7828 10854 7840 10906
rect 7892 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 34315 10906
rect 34367 10854 34379 10906
rect 34431 10854 34443 10906
rect 34495 10854 34507 10906
rect 34559 10854 38824 10906
rect 1104 10832 38824 10854
rect 1104 10362 38824 10384
rect 1104 10310 14315 10362
rect 14367 10310 14379 10362
rect 14431 10310 14443 10362
rect 14495 10310 14507 10362
rect 14559 10310 27648 10362
rect 27700 10310 27712 10362
rect 27764 10310 27776 10362
rect 27828 10310 27840 10362
rect 27892 10310 38824 10362
rect 1104 10288 38824 10310
rect 1104 9818 38824 9840
rect 1104 9766 7648 9818
rect 7700 9766 7712 9818
rect 7764 9766 7776 9818
rect 7828 9766 7840 9818
rect 7892 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 34315 9818
rect 34367 9766 34379 9818
rect 34431 9766 34443 9818
rect 34495 9766 34507 9818
rect 34559 9766 38824 9818
rect 1104 9744 38824 9766
rect 20441 9503 20499 9509
rect 20441 9500 20453 9503
rect 20180 9472 20453 9500
rect 20180 9376 20208 9472
rect 20441 9469 20453 9472
rect 20487 9469 20499 9503
rect 20441 9463 20499 9469
rect 20162 9364 20168 9376
rect 20123 9336 20168 9364
rect 20162 9324 20168 9336
rect 20220 9324 20226 9376
rect 20806 9364 20812 9376
rect 20767 9336 20812 9364
rect 20806 9324 20812 9336
rect 20864 9324 20870 9376
rect 1104 9274 38824 9296
rect 1104 9222 14315 9274
rect 14367 9222 14379 9274
rect 14431 9222 14443 9274
rect 14495 9222 14507 9274
rect 14559 9222 27648 9274
rect 27700 9222 27712 9274
rect 27764 9222 27776 9274
rect 27828 9222 27840 9274
rect 27892 9222 38824 9274
rect 1104 9200 38824 9222
rect 16482 9024 16488 9036
rect 16443 8996 16488 9024
rect 16482 8984 16488 8996
rect 16540 8984 16546 9036
rect 23014 9024 23020 9036
rect 22975 8996 23020 9024
rect 23014 8984 23020 8996
rect 23072 8984 23078 9036
rect 10045 8823 10103 8829
rect 10045 8789 10057 8823
rect 10091 8820 10103 8823
rect 10226 8820 10232 8832
rect 10091 8792 10232 8820
rect 10091 8789 10103 8792
rect 10045 8783 10103 8789
rect 10226 8780 10232 8792
rect 10284 8780 10290 8832
rect 16666 8820 16672 8832
rect 16627 8792 16672 8820
rect 16666 8780 16672 8792
rect 16724 8780 16730 8832
rect 22830 8820 22836 8832
rect 22791 8792 22836 8820
rect 22830 8780 22836 8792
rect 22888 8780 22894 8832
rect 1104 8730 38824 8752
rect 1104 8678 7648 8730
rect 7700 8678 7712 8730
rect 7764 8678 7776 8730
rect 7828 8678 7840 8730
rect 7892 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 34315 8730
rect 34367 8678 34379 8730
rect 34431 8678 34443 8730
rect 34495 8678 34507 8730
rect 34559 8678 38824 8730
rect 1104 8656 38824 8678
rect 16482 8616 16488 8628
rect 16443 8588 16488 8616
rect 16482 8576 16488 8588
rect 16540 8576 16546 8628
rect 22554 8508 22560 8560
rect 22612 8548 22618 8560
rect 22649 8551 22707 8557
rect 22649 8548 22661 8551
rect 22612 8520 22661 8548
rect 22612 8508 22618 8520
rect 22649 8517 22661 8520
rect 22695 8517 22707 8551
rect 22649 8511 22707 8517
rect 9493 8483 9551 8489
rect 9493 8449 9505 8483
rect 9539 8480 9551 8483
rect 9539 8452 10456 8480
rect 9539 8449 9551 8452
rect 9493 8443 9551 8449
rect 10428 8424 10456 8452
rect 10226 8412 10232 8424
rect 10187 8384 10232 8412
rect 10226 8372 10232 8384
rect 10284 8372 10290 8424
rect 10410 8412 10416 8424
rect 10371 8384 10416 8412
rect 10410 8372 10416 8384
rect 10468 8372 10474 8424
rect 10502 8372 10508 8424
rect 10560 8412 10566 8424
rect 10781 8415 10839 8421
rect 10781 8412 10793 8415
rect 10560 8384 10793 8412
rect 10560 8372 10566 8384
rect 10781 8381 10793 8384
rect 10827 8381 10839 8415
rect 11330 8412 11336 8424
rect 11291 8384 11336 8412
rect 10781 8375 10839 8381
rect 11330 8372 11336 8384
rect 11388 8372 11394 8424
rect 22094 8372 22100 8424
rect 22152 8412 22158 8424
rect 22465 8415 22523 8421
rect 22465 8412 22477 8415
rect 22152 8384 22477 8412
rect 22152 8372 22158 8384
rect 22465 8381 22477 8384
rect 22511 8412 22523 8415
rect 22511 8384 23428 8412
rect 22511 8381 22523 8384
rect 22465 8375 22523 8381
rect 9861 8347 9919 8353
rect 9861 8313 9873 8347
rect 9907 8344 9919 8347
rect 10962 8344 10968 8356
rect 9907 8316 10968 8344
rect 9907 8313 9919 8316
rect 9861 8307 9919 8313
rect 10962 8304 10968 8316
rect 11020 8344 11026 8356
rect 11348 8344 11376 8372
rect 23400 8356 23428 8384
rect 23014 8344 23020 8356
rect 11020 8316 11376 8344
rect 22975 8316 23020 8344
rect 11020 8304 11026 8316
rect 23014 8304 23020 8316
rect 23072 8304 23078 8356
rect 23382 8344 23388 8356
rect 23343 8316 23388 8344
rect 23382 8304 23388 8316
rect 23440 8304 23446 8356
rect 10042 8276 10048 8288
rect 10003 8248 10048 8276
rect 10042 8236 10048 8248
rect 10100 8236 10106 8288
rect 1104 8186 38824 8208
rect 1104 8134 14315 8186
rect 14367 8134 14379 8186
rect 14431 8134 14443 8186
rect 14495 8134 14507 8186
rect 14559 8134 27648 8186
rect 27700 8134 27712 8186
rect 27764 8134 27776 8186
rect 27828 8134 27840 8186
rect 27892 8134 38824 8186
rect 1104 8112 38824 8134
rect 10410 8004 10416 8016
rect 10323 7976 10416 8004
rect 10410 7964 10416 7976
rect 10468 8004 10474 8016
rect 10468 7976 11192 8004
rect 10468 7964 10474 7976
rect 11164 7948 11192 7976
rect 10226 7896 10232 7948
rect 10284 7936 10290 7948
rect 10781 7939 10839 7945
rect 10781 7936 10793 7939
rect 10284 7908 10793 7936
rect 10284 7896 10290 7908
rect 10781 7905 10793 7908
rect 10827 7905 10839 7939
rect 11146 7936 11152 7948
rect 11107 7908 11152 7936
rect 10781 7899 10839 7905
rect 10796 7868 10824 7899
rect 11146 7896 11152 7908
rect 11204 7896 11210 7948
rect 11330 7936 11336 7948
rect 11291 7908 11336 7936
rect 11330 7896 11336 7908
rect 11388 7896 11394 7948
rect 11885 7939 11943 7945
rect 11885 7905 11897 7939
rect 11931 7936 11943 7939
rect 12066 7936 12072 7948
rect 11931 7908 12072 7936
rect 11931 7905 11943 7908
rect 11885 7899 11943 7905
rect 12066 7896 12072 7908
rect 12124 7896 12130 7948
rect 11698 7868 11704 7880
rect 10796 7840 11704 7868
rect 11698 7828 11704 7840
rect 11756 7828 11762 7880
rect 11882 7800 11888 7812
rect 11843 7772 11888 7800
rect 11882 7760 11888 7772
rect 11940 7760 11946 7812
rect 10045 7735 10103 7741
rect 10045 7701 10057 7735
rect 10091 7732 10103 7735
rect 10502 7732 10508 7744
rect 10091 7704 10508 7732
rect 10091 7701 10103 7704
rect 10045 7695 10103 7701
rect 10502 7692 10508 7704
rect 10560 7692 10566 7744
rect 19702 7732 19708 7744
rect 19663 7704 19708 7732
rect 19702 7692 19708 7704
rect 19760 7692 19766 7744
rect 1104 7642 38824 7664
rect 1104 7590 7648 7642
rect 7700 7590 7712 7642
rect 7764 7590 7776 7642
rect 7828 7590 7840 7642
rect 7892 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 34315 7642
rect 34367 7590 34379 7642
rect 34431 7590 34443 7642
rect 34495 7590 34507 7642
rect 34559 7590 38824 7642
rect 1104 7568 38824 7590
rect 9033 7531 9091 7537
rect 9033 7497 9045 7531
rect 9079 7528 9091 7531
rect 10502 7528 10508 7540
rect 9079 7500 10508 7528
rect 9079 7497 9091 7500
rect 9033 7491 9091 7497
rect 10502 7488 10508 7500
rect 10560 7528 10566 7540
rect 11330 7528 11336 7540
rect 10560 7500 11336 7528
rect 10560 7488 10566 7500
rect 11330 7488 11336 7500
rect 11388 7488 11394 7540
rect 11698 7528 11704 7540
rect 11659 7500 11704 7528
rect 11698 7488 11704 7500
rect 11756 7488 11762 7540
rect 8665 7395 8723 7401
rect 8665 7361 8677 7395
rect 8711 7392 8723 7395
rect 8711 7364 10916 7392
rect 8711 7361 8723 7364
rect 8665 7355 8723 7361
rect 9401 7327 9459 7333
rect 9401 7293 9413 7327
rect 9447 7324 9459 7327
rect 9769 7327 9827 7333
rect 9769 7324 9781 7327
rect 9447 7296 9781 7324
rect 9447 7293 9459 7296
rect 9401 7287 9459 7293
rect 9769 7293 9781 7296
rect 9815 7324 9827 7327
rect 9858 7324 9864 7336
rect 9815 7296 9864 7324
rect 9815 7293 9827 7296
rect 9769 7287 9827 7293
rect 9858 7284 9864 7296
rect 9916 7284 9922 7336
rect 10229 7327 10287 7333
rect 10229 7293 10241 7327
rect 10275 7324 10287 7327
rect 10318 7324 10324 7336
rect 10275 7296 10324 7324
rect 10275 7293 10287 7296
rect 10229 7287 10287 7293
rect 10318 7284 10324 7296
rect 10376 7284 10382 7336
rect 10502 7324 10508 7336
rect 10463 7296 10508 7324
rect 10502 7284 10508 7296
rect 10560 7284 10566 7336
rect 10888 7333 10916 7364
rect 10873 7327 10931 7333
rect 10873 7293 10885 7327
rect 10919 7324 10931 7327
rect 12066 7324 12072 7336
rect 10919 7296 12072 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 12066 7284 12072 7296
rect 12124 7284 12130 7336
rect 19242 7284 19248 7336
rect 19300 7324 19306 7336
rect 20441 7327 20499 7333
rect 20441 7324 20453 7327
rect 19300 7296 20453 7324
rect 19300 7284 19306 7296
rect 20441 7293 20453 7296
rect 20487 7293 20499 7327
rect 20441 7287 20499 7293
rect 19702 7256 19708 7268
rect 19663 7228 19708 7256
rect 19702 7216 19708 7228
rect 19760 7216 19766 7268
rect 19886 7256 19892 7268
rect 19847 7228 19892 7256
rect 19886 7216 19892 7228
rect 19944 7216 19950 7268
rect 20070 7256 20076 7268
rect 20031 7228 20076 7256
rect 20070 7216 20076 7228
rect 20128 7216 20134 7268
rect 9766 7188 9772 7200
rect 9727 7160 9772 7188
rect 9766 7148 9772 7160
rect 9824 7148 9830 7200
rect 19150 7188 19156 7200
rect 19111 7160 19156 7188
rect 19150 7148 19156 7160
rect 19208 7148 19214 7200
rect 19613 7191 19671 7197
rect 19613 7157 19625 7191
rect 19659 7188 19671 7191
rect 19981 7191 20039 7197
rect 19981 7188 19993 7191
rect 19659 7160 19993 7188
rect 19659 7157 19671 7160
rect 19613 7151 19671 7157
rect 19981 7157 19993 7160
rect 20027 7188 20039 7191
rect 20622 7188 20628 7200
rect 20027 7160 20628 7188
rect 20027 7157 20039 7160
rect 19981 7151 20039 7157
rect 20622 7148 20628 7160
rect 20680 7148 20686 7200
rect 1104 7098 38824 7120
rect 1104 7046 14315 7098
rect 14367 7046 14379 7098
rect 14431 7046 14443 7098
rect 14495 7046 14507 7098
rect 14559 7046 27648 7098
rect 27700 7046 27712 7098
rect 27764 7046 27776 7098
rect 27828 7046 27840 7098
rect 27892 7046 38824 7098
rect 1104 7024 38824 7046
rect 9766 6984 9772 6996
rect 9727 6956 9772 6984
rect 9766 6944 9772 6956
rect 9824 6944 9830 6996
rect 19797 6987 19855 6993
rect 19797 6953 19809 6987
rect 19843 6984 19855 6987
rect 19886 6984 19892 6996
rect 19843 6956 19892 6984
rect 19843 6953 19855 6956
rect 19797 6947 19855 6953
rect 19886 6944 19892 6956
rect 19944 6984 19950 6996
rect 21085 6987 21143 6993
rect 21085 6984 21097 6987
rect 19944 6956 21097 6984
rect 19944 6944 19950 6956
rect 21085 6953 21097 6956
rect 21131 6984 21143 6987
rect 21131 6956 22968 6984
rect 21131 6953 21143 6956
rect 21085 6947 21143 6953
rect 22940 6928 22968 6956
rect 9398 6876 9404 6928
rect 9456 6916 9462 6928
rect 10410 6916 10416 6928
rect 9456 6888 10416 6916
rect 9456 6876 9462 6888
rect 9858 6848 9864 6860
rect 9819 6820 9864 6848
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 10336 6857 10364 6888
rect 10410 6876 10416 6888
rect 10468 6876 10474 6928
rect 20070 6876 20076 6928
rect 20128 6916 20134 6928
rect 20806 6916 20812 6928
rect 20128 6888 20812 6916
rect 20128 6876 20134 6888
rect 20806 6876 20812 6888
rect 20864 6916 20870 6928
rect 21269 6919 21327 6925
rect 21269 6916 21281 6919
rect 20864 6888 21281 6916
rect 20864 6876 20870 6888
rect 21269 6885 21281 6888
rect 21315 6885 21327 6919
rect 22738 6916 22744 6928
rect 22699 6888 22744 6916
rect 21269 6879 21327 6885
rect 22738 6876 22744 6888
rect 22796 6876 22802 6928
rect 22922 6916 22928 6928
rect 22835 6888 22928 6916
rect 22922 6876 22928 6888
rect 22980 6876 22986 6928
rect 10321 6851 10379 6857
rect 10321 6817 10333 6851
rect 10367 6848 10379 6851
rect 10502 6848 10508 6860
rect 10367 6820 10401 6848
rect 10463 6820 10508 6848
rect 10367 6817 10379 6820
rect 10321 6811 10379 6817
rect 10502 6808 10508 6820
rect 10560 6808 10566 6860
rect 10870 6848 10876 6860
rect 10831 6820 10876 6848
rect 10870 6808 10876 6820
rect 10928 6808 10934 6860
rect 20714 6808 20720 6860
rect 20772 6848 20778 6860
rect 21177 6851 21235 6857
rect 21177 6848 21189 6851
rect 20772 6820 21189 6848
rect 20772 6808 20778 6820
rect 21177 6817 21189 6820
rect 21223 6848 21235 6851
rect 21358 6848 21364 6860
rect 21223 6820 21364 6848
rect 21223 6817 21235 6820
rect 21177 6811 21235 6817
rect 21358 6808 21364 6820
rect 21416 6848 21422 6860
rect 22002 6848 22008 6860
rect 21416 6820 22008 6848
rect 21416 6808 21422 6820
rect 22002 6808 22008 6820
rect 22060 6808 22066 6860
rect 22830 6848 22836 6860
rect 22791 6820 22836 6848
rect 22830 6808 22836 6820
rect 22888 6808 22894 6860
rect 20806 6740 20812 6792
rect 20864 6780 20870 6792
rect 20901 6783 20959 6789
rect 20901 6780 20913 6783
rect 20864 6752 20913 6780
rect 20864 6740 20870 6752
rect 20901 6749 20913 6752
rect 20947 6749 20959 6783
rect 21634 6780 21640 6792
rect 21595 6752 21640 6780
rect 20901 6743 20959 6749
rect 21634 6740 21640 6752
rect 21692 6740 21698 6792
rect 22554 6780 22560 6792
rect 22515 6752 22560 6780
rect 22554 6740 22560 6752
rect 22612 6740 22618 6792
rect 23293 6783 23351 6789
rect 23293 6749 23305 6783
rect 23339 6780 23351 6783
rect 23382 6780 23388 6792
rect 23339 6752 23388 6780
rect 23339 6749 23351 6752
rect 23293 6743 23351 6749
rect 23382 6740 23388 6752
rect 23440 6740 23446 6792
rect 24394 6712 24400 6724
rect 24355 6684 24400 6712
rect 24394 6672 24400 6684
rect 24452 6672 24458 6724
rect 1104 6554 38824 6576
rect 1104 6502 7648 6554
rect 7700 6502 7712 6554
rect 7764 6502 7776 6554
rect 7828 6502 7840 6554
rect 7892 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 34315 6554
rect 34367 6502 34379 6554
rect 34431 6502 34443 6554
rect 34495 6502 34507 6554
rect 34559 6502 38824 6554
rect 1104 6480 38824 6502
rect 9398 6440 9404 6452
rect 9359 6412 9404 6440
rect 9398 6400 9404 6412
rect 9456 6400 9462 6452
rect 9769 6443 9827 6449
rect 9769 6409 9781 6443
rect 9815 6440 9827 6443
rect 9858 6440 9864 6452
rect 9815 6412 9864 6440
rect 9815 6409 9827 6412
rect 9769 6403 9827 6409
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 10502 6440 10508 6452
rect 10463 6412 10508 6440
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 20070 6400 20076 6452
rect 20128 6440 20134 6452
rect 20533 6443 20591 6449
rect 20533 6440 20545 6443
rect 20128 6412 20545 6440
rect 20128 6400 20134 6412
rect 20533 6409 20545 6412
rect 20579 6409 20591 6443
rect 21358 6440 21364 6452
rect 21319 6412 21364 6440
rect 20533 6403 20591 6409
rect 21358 6400 21364 6412
rect 21416 6400 21422 6452
rect 22281 6443 22339 6449
rect 22281 6409 22293 6443
rect 22327 6440 22339 6443
rect 22830 6440 22836 6452
rect 22327 6412 22836 6440
rect 22327 6409 22339 6412
rect 22281 6403 22339 6409
rect 22830 6400 22836 6412
rect 22888 6400 22894 6452
rect 10410 6332 10416 6384
rect 10468 6372 10474 6384
rect 10781 6375 10839 6381
rect 10781 6372 10793 6375
rect 10468 6344 10793 6372
rect 10468 6332 10474 6344
rect 10781 6341 10793 6344
rect 10827 6341 10839 6375
rect 10781 6335 10839 6341
rect 22649 6375 22707 6381
rect 22649 6341 22661 6375
rect 22695 6372 22707 6375
rect 22738 6372 22744 6384
rect 22695 6344 22744 6372
rect 22695 6341 22707 6344
rect 22649 6335 22707 6341
rect 22738 6332 22744 6344
rect 22796 6372 22802 6384
rect 24486 6372 24492 6384
rect 22796 6344 24492 6372
rect 22796 6332 22802 6344
rect 24486 6332 24492 6344
rect 24544 6332 24550 6384
rect 10137 6307 10195 6313
rect 10137 6273 10149 6307
rect 10183 6304 10195 6307
rect 10870 6304 10876 6316
rect 10183 6276 10876 6304
rect 10183 6273 10195 6276
rect 10137 6267 10195 6273
rect 10870 6264 10876 6276
rect 10928 6264 10934 6316
rect 24118 6304 24124 6316
rect 24079 6276 24124 6304
rect 24118 6264 24124 6276
rect 24176 6264 24182 6316
rect 20898 6236 20904 6248
rect 20859 6208 20904 6236
rect 20898 6196 20904 6208
rect 20956 6196 20962 6248
rect 21729 6239 21787 6245
rect 21729 6205 21741 6239
rect 21775 6236 21787 6239
rect 22922 6236 22928 6248
rect 21775 6208 22928 6236
rect 21775 6205 21787 6208
rect 21729 6199 21787 6205
rect 22922 6196 22928 6208
rect 22980 6236 22986 6248
rect 24504 6245 24532 6332
rect 23017 6239 23075 6245
rect 23017 6236 23029 6239
rect 22980 6208 23029 6236
rect 22980 6196 22986 6208
rect 23017 6205 23029 6208
rect 23063 6236 23075 6239
rect 24489 6239 24547 6245
rect 23063 6208 24440 6236
rect 23063 6205 23075 6208
rect 23017 6199 23075 6205
rect 24412 6180 24440 6208
rect 24489 6205 24501 6239
rect 24535 6205 24547 6239
rect 24489 6199 24547 6205
rect 22554 6128 22560 6180
rect 22612 6168 22618 6180
rect 23385 6171 23443 6177
rect 23385 6168 23397 6171
rect 22612 6140 23397 6168
rect 22612 6128 22618 6140
rect 23385 6137 23397 6140
rect 23431 6168 23443 6171
rect 24302 6168 24308 6180
rect 23431 6140 24308 6168
rect 23431 6137 23443 6140
rect 23385 6131 23443 6137
rect 24302 6128 24308 6140
rect 24360 6128 24366 6180
rect 24394 6128 24400 6180
rect 24452 6168 24458 6180
rect 24673 6171 24731 6177
rect 24673 6168 24685 6171
rect 24452 6140 24685 6168
rect 24452 6128 24458 6140
rect 24673 6137 24685 6140
rect 24719 6137 24731 6171
rect 25038 6168 25044 6180
rect 24999 6140 25044 6168
rect 24673 6131 24731 6137
rect 25038 6128 25044 6140
rect 25096 6128 25102 6180
rect 24118 6060 24124 6112
rect 24176 6100 24182 6112
rect 24581 6103 24639 6109
rect 24581 6100 24593 6103
rect 24176 6072 24593 6100
rect 24176 6060 24182 6072
rect 24581 6069 24593 6072
rect 24627 6069 24639 6103
rect 24581 6063 24639 6069
rect 1104 6010 38824 6032
rect 1104 5958 14315 6010
rect 14367 5958 14379 6010
rect 14431 5958 14443 6010
rect 14495 5958 14507 6010
rect 14559 5958 27648 6010
rect 27700 5958 27712 6010
rect 27764 5958 27776 6010
rect 27828 5958 27840 6010
rect 27892 5958 38824 6010
rect 1104 5936 38824 5958
rect 24397 5899 24455 5905
rect 24397 5865 24409 5899
rect 24443 5896 24455 5899
rect 24486 5896 24492 5908
rect 24443 5868 24492 5896
rect 24443 5865 24455 5868
rect 24397 5859 24455 5865
rect 24486 5856 24492 5868
rect 24544 5856 24550 5908
rect 24302 5788 24308 5840
rect 24360 5828 24366 5840
rect 24673 5831 24731 5837
rect 24673 5828 24685 5831
rect 24360 5800 24685 5828
rect 24360 5788 24366 5800
rect 24673 5797 24685 5800
rect 24719 5797 24731 5831
rect 24673 5791 24731 5797
rect 1104 5466 38824 5488
rect 1104 5414 7648 5466
rect 7700 5414 7712 5466
rect 7764 5414 7776 5466
rect 7828 5414 7840 5466
rect 7892 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 34315 5466
rect 34367 5414 34379 5466
rect 34431 5414 34443 5466
rect 34495 5414 34507 5466
rect 34559 5414 38824 5466
rect 1104 5392 38824 5414
rect 3053 5151 3111 5157
rect 3053 5117 3065 5151
rect 3099 5148 3111 5151
rect 3142 5148 3148 5160
rect 3099 5120 3148 5148
rect 3099 5117 3111 5120
rect 3053 5111 3111 5117
rect 3142 5108 3148 5120
rect 3200 5108 3206 5160
rect 2961 5083 3019 5089
rect 2961 5049 2973 5083
rect 3007 5080 3019 5083
rect 3415 5083 3473 5089
rect 3415 5080 3427 5083
rect 3007 5052 3427 5080
rect 3007 5049 3019 5052
rect 2961 5043 3019 5049
rect 3415 5049 3427 5052
rect 3461 5080 3473 5083
rect 3510 5080 3516 5092
rect 3461 5052 3516 5080
rect 3461 5049 3473 5052
rect 3415 5043 3473 5049
rect 3510 5040 3516 5052
rect 3568 5040 3574 5092
rect 3970 5012 3976 5024
rect 3931 4984 3976 5012
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 1104 4922 38824 4944
rect 1104 4870 14315 4922
rect 14367 4870 14379 4922
rect 14431 4870 14443 4922
rect 14495 4870 14507 4922
rect 14559 4870 27648 4922
rect 27700 4870 27712 4922
rect 27764 4870 27776 4922
rect 27828 4870 27840 4922
rect 27892 4870 38824 4922
rect 1104 4848 38824 4870
rect 25038 4768 25044 4820
rect 25096 4808 25102 4820
rect 25225 4811 25283 4817
rect 25225 4808 25237 4811
rect 25096 4780 25237 4808
rect 25096 4768 25102 4780
rect 25225 4777 25237 4780
rect 25271 4777 25283 4811
rect 25225 4771 25283 4777
rect 5626 4700 5632 4752
rect 5684 4740 5690 4752
rect 5858 4743 5916 4749
rect 5858 4740 5870 4743
rect 5684 4712 5870 4740
rect 5684 4700 5690 4712
rect 5858 4709 5870 4712
rect 5904 4709 5916 4743
rect 5858 4703 5916 4709
rect 5537 4675 5595 4681
rect 5537 4641 5549 4675
rect 5583 4672 5595 4675
rect 5994 4672 6000 4684
rect 5583 4644 6000 4672
rect 5583 4641 5595 4644
rect 5537 4635 5595 4641
rect 5994 4632 6000 4644
rect 6052 4632 6058 4684
rect 3142 4604 3148 4616
rect 3103 4576 3148 4604
rect 3142 4564 3148 4576
rect 3200 4564 3206 4616
rect 5442 4428 5448 4480
rect 5500 4468 5506 4480
rect 6457 4471 6515 4477
rect 6457 4468 6469 4471
rect 5500 4440 6469 4468
rect 5500 4428 5506 4440
rect 6457 4437 6469 4440
rect 6503 4437 6515 4471
rect 6457 4431 6515 4437
rect 1104 4378 38824 4400
rect 1104 4326 7648 4378
rect 7700 4326 7712 4378
rect 7764 4326 7776 4378
rect 7828 4326 7840 4378
rect 7892 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 34315 4378
rect 34367 4326 34379 4378
rect 34431 4326 34443 4378
rect 34495 4326 34507 4378
rect 34559 4326 38824 4378
rect 1104 4304 38824 4326
rect 5994 4264 6000 4276
rect 5955 4236 6000 4264
rect 5994 4224 6000 4236
rect 6052 4224 6058 4276
rect 9122 4128 9128 4140
rect 9083 4100 9128 4128
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 18049 4131 18107 4137
rect 18049 4097 18061 4131
rect 18095 4128 18107 4131
rect 18138 4128 18144 4140
rect 18095 4100 18144 4128
rect 18095 4097 18107 4100
rect 18049 4091 18107 4097
rect 18138 4088 18144 4100
rect 18196 4128 18202 4140
rect 19242 4128 19248 4140
rect 18196 4100 19248 4128
rect 18196 4088 18202 4100
rect 19242 4088 19248 4100
rect 19300 4088 19306 4140
rect 20533 4131 20591 4137
rect 20533 4097 20545 4131
rect 20579 4128 20591 4131
rect 20993 4131 21051 4137
rect 20993 4128 21005 4131
rect 20579 4100 21005 4128
rect 20579 4097 20591 4100
rect 20533 4091 20591 4097
rect 20993 4097 21005 4100
rect 21039 4128 21051 4131
rect 21634 4128 21640 4140
rect 21039 4100 21640 4128
rect 21039 4097 21051 4100
rect 20993 4091 21051 4097
rect 21634 4088 21640 4100
rect 21692 4088 21698 4140
rect 25038 4088 25044 4140
rect 25096 4128 25102 4140
rect 25225 4131 25283 4137
rect 25225 4128 25237 4131
rect 25096 4100 25237 4128
rect 25096 4088 25102 4100
rect 25225 4097 25237 4100
rect 25271 4097 25283 4131
rect 25225 4091 25283 4097
rect 3145 4063 3203 4069
rect 3145 4029 3157 4063
rect 3191 4060 3203 4063
rect 3234 4060 3240 4072
rect 3191 4032 3240 4060
rect 3191 4029 3203 4032
rect 3145 4023 3203 4029
rect 3234 4020 3240 4032
rect 3292 4020 3298 4072
rect 5626 4060 5632 4072
rect 5587 4032 5632 4060
rect 5626 4020 5632 4032
rect 5684 4020 5690 4072
rect 3510 4001 3516 4004
rect 3053 3995 3111 4001
rect 3053 3961 3065 3995
rect 3099 3992 3111 3995
rect 3507 3992 3516 4001
rect 3099 3964 3516 3992
rect 3099 3961 3111 3964
rect 3053 3955 3111 3961
rect 3507 3955 3516 3964
rect 3510 3952 3516 3955
rect 3568 3952 3574 4004
rect 9490 4001 9496 4004
rect 9033 3995 9091 4001
rect 9033 3961 9045 3995
rect 9079 3992 9091 3995
rect 9487 3992 9496 4001
rect 9079 3964 9496 3992
rect 9079 3961 9091 3964
rect 9033 3955 9091 3961
rect 9487 3955 9496 3964
rect 9490 3952 9496 3955
rect 9548 3952 9554 4004
rect 17770 3992 17776 4004
rect 17731 3964 17776 3992
rect 17770 3952 17776 3964
rect 17828 3992 17834 4004
rect 21358 4001 21364 4004
rect 18370 3995 18428 4001
rect 18370 3992 18382 3995
rect 17828 3964 18382 3992
rect 17828 3952 17834 3964
rect 18370 3961 18382 3964
rect 18416 3992 18428 3995
rect 20809 3995 20867 4001
rect 20809 3992 20821 3995
rect 18416 3964 20821 3992
rect 18416 3961 18428 3964
rect 18370 3955 18428 3961
rect 20809 3961 20821 3964
rect 20855 3992 20867 3995
rect 21314 3995 21364 4001
rect 21314 3992 21326 3995
rect 20855 3964 21326 3992
rect 20855 3961 20867 3964
rect 20809 3955 20867 3961
rect 21314 3961 21326 3964
rect 21360 3961 21364 3995
rect 21314 3955 21364 3961
rect 21358 3952 21364 3955
rect 21416 3992 21422 4004
rect 25590 4001 25596 4004
rect 25546 3995 25596 4001
rect 25546 3992 25558 3995
rect 21416 3964 21462 3992
rect 25056 3964 25558 3992
rect 21416 3952 21422 3964
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 4065 3927 4123 3933
rect 4065 3924 4077 3927
rect 2832 3896 4077 3924
rect 2832 3884 2838 3896
rect 4065 3893 4077 3896
rect 4111 3893 4123 3927
rect 10042 3924 10048 3936
rect 10003 3896 10048 3924
rect 4065 3887 4123 3893
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 18966 3924 18972 3936
rect 18927 3896 18972 3924
rect 18966 3884 18972 3896
rect 19024 3884 19030 3936
rect 21910 3924 21916 3936
rect 21871 3896 21916 3924
rect 21910 3884 21916 3896
rect 21968 3884 21974 3936
rect 24302 3884 24308 3936
rect 24360 3924 24366 3936
rect 25056 3933 25084 3964
rect 25546 3961 25558 3964
rect 25592 3961 25596 3995
rect 25546 3955 25596 3961
rect 25590 3952 25596 3955
rect 25648 3992 25654 4004
rect 25648 3964 25694 3992
rect 25648 3952 25654 3964
rect 25041 3927 25099 3933
rect 25041 3924 25053 3927
rect 24360 3896 25053 3924
rect 24360 3884 24366 3896
rect 25041 3893 25053 3896
rect 25087 3893 25099 3927
rect 26142 3924 26148 3936
rect 26103 3896 26148 3924
rect 25041 3887 25099 3893
rect 26142 3884 26148 3896
rect 26200 3884 26206 3936
rect 1104 3834 38824 3856
rect 1104 3782 14315 3834
rect 14367 3782 14379 3834
rect 14431 3782 14443 3834
rect 14495 3782 14507 3834
rect 14559 3782 27648 3834
rect 27700 3782 27712 3834
rect 27764 3782 27776 3834
rect 27828 3782 27840 3834
rect 27892 3782 38824 3834
rect 1104 3760 38824 3782
rect 2038 3720 2044 3732
rect 1999 3692 2044 3720
rect 2038 3680 2044 3692
rect 2096 3680 2102 3732
rect 3234 3720 3240 3732
rect 3195 3692 3240 3720
rect 3234 3680 3240 3692
rect 3292 3680 3298 3732
rect 9122 3720 9128 3732
rect 9083 3692 9128 3720
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 18138 3720 18144 3732
rect 18099 3692 18144 3720
rect 18138 3680 18144 3692
rect 18196 3680 18202 3732
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3584 1455 3587
rect 2056 3584 2084 3680
rect 24302 3612 24308 3664
rect 24360 3661 24366 3664
rect 24360 3655 24408 3661
rect 24360 3621 24362 3655
rect 24396 3621 24408 3655
rect 24360 3615 24408 3621
rect 24360 3612 24366 3615
rect 1443 3556 2084 3584
rect 1443 3553 1455 3556
rect 1397 3547 1455 3553
rect 23474 3544 23480 3596
rect 23532 3584 23538 3596
rect 24029 3587 24087 3593
rect 24029 3584 24041 3587
rect 23532 3556 24041 3584
rect 23532 3544 23538 3556
rect 24029 3553 24041 3556
rect 24075 3584 24087 3587
rect 24210 3584 24216 3596
rect 24075 3556 24216 3584
rect 24075 3553 24087 3556
rect 24029 3547 24087 3553
rect 24210 3544 24216 3556
rect 24268 3544 24274 3596
rect 1581 3383 1639 3389
rect 1581 3349 1593 3383
rect 1627 3380 1639 3383
rect 3694 3380 3700 3392
rect 1627 3352 3700 3380
rect 1627 3349 1639 3352
rect 1581 3343 1639 3349
rect 3694 3340 3700 3352
rect 3752 3340 3758 3392
rect 24949 3383 25007 3389
rect 24949 3349 24961 3383
rect 24995 3380 25007 3383
rect 25222 3380 25228 3392
rect 24995 3352 25228 3380
rect 24995 3349 25007 3352
rect 24949 3343 25007 3349
rect 25222 3340 25228 3352
rect 25280 3340 25286 3392
rect 1104 3290 38824 3312
rect 1104 3238 7648 3290
rect 7700 3238 7712 3290
rect 7764 3238 7776 3290
rect 7828 3238 7840 3290
rect 7892 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 34315 3290
rect 34367 3238 34379 3290
rect 34431 3238 34443 3290
rect 34495 3238 34507 3290
rect 34559 3238 38824 3290
rect 1104 3216 38824 3238
rect 2777 3179 2835 3185
rect 2777 3145 2789 3179
rect 2823 3176 2835 3179
rect 3970 3176 3976 3188
rect 2823 3148 3976 3176
rect 2823 3145 2835 3148
rect 2777 3139 2835 3145
rect 2038 3108 2044 3120
rect 1999 3080 2044 3108
rect 2038 3068 2044 3080
rect 2096 3068 2102 3120
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3040 1639 3043
rect 2792 3040 2820 3139
rect 3970 3136 3976 3148
rect 4028 3136 4034 3188
rect 16758 3136 16764 3188
rect 16816 3176 16822 3188
rect 17126 3176 17132 3188
rect 16816 3148 17132 3176
rect 16816 3136 16822 3148
rect 17126 3136 17132 3148
rect 17184 3136 17190 3188
rect 22186 3176 22192 3188
rect 22147 3148 22192 3176
rect 22186 3136 22192 3148
rect 22244 3136 22250 3188
rect 24210 3136 24216 3188
rect 24268 3176 24274 3188
rect 24397 3179 24455 3185
rect 24397 3176 24409 3179
rect 24268 3148 24409 3176
rect 24268 3136 24274 3148
rect 24397 3145 24409 3148
rect 24443 3145 24455 3179
rect 25682 3176 25688 3188
rect 25643 3148 25688 3176
rect 24397 3139 24455 3145
rect 25682 3136 25688 3148
rect 25740 3136 25746 3188
rect 21726 3108 21732 3120
rect 21687 3080 21732 3108
rect 21726 3068 21732 3080
rect 21784 3068 21790 3120
rect 24121 3111 24179 3117
rect 24121 3077 24133 3111
rect 24167 3108 24179 3111
rect 24302 3108 24308 3120
rect 24167 3080 24308 3108
rect 24167 3077 24179 3080
rect 24121 3071 24179 3077
rect 24302 3068 24308 3080
rect 24360 3068 24366 3120
rect 25222 3040 25228 3052
rect 1627 3012 2820 3040
rect 25183 3012 25228 3040
rect 1627 3009 1639 3012
rect 1581 3003 1639 3009
rect 25222 3000 25228 3012
rect 25280 3000 25286 3052
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2972 1455 2975
rect 16485 2975 16543 2981
rect 1443 2944 2452 2972
rect 1443 2941 1455 2944
rect 1397 2935 1455 2941
rect 2424 2848 2452 2944
rect 16485 2941 16497 2975
rect 16531 2972 16543 2975
rect 16758 2972 16764 2984
rect 16531 2944 16764 2972
rect 16531 2941 16543 2944
rect 16485 2935 16543 2941
rect 16758 2932 16764 2944
rect 16816 2932 16822 2984
rect 21545 2975 21603 2981
rect 21545 2941 21557 2975
rect 21591 2972 21603 2975
rect 21818 2972 21824 2984
rect 21591 2944 21824 2972
rect 21591 2941 21603 2944
rect 21545 2935 21603 2941
rect 21818 2932 21824 2944
rect 21876 2972 21882 2984
rect 22186 2972 22192 2984
rect 21876 2944 22192 2972
rect 21876 2932 21882 2944
rect 22186 2932 22192 2944
rect 22244 2932 22250 2984
rect 24949 2975 25007 2981
rect 24949 2941 24961 2975
rect 24995 2972 25007 2975
rect 25038 2972 25044 2984
rect 24995 2944 25044 2972
rect 24995 2941 25007 2944
rect 24949 2935 25007 2941
rect 25038 2932 25044 2944
rect 25096 2932 25102 2984
rect 2406 2836 2412 2848
rect 2367 2808 2412 2836
rect 2406 2796 2412 2808
rect 2464 2796 2470 2848
rect 16666 2836 16672 2848
rect 16627 2808 16672 2836
rect 16666 2796 16672 2808
rect 16724 2796 16730 2848
rect 1104 2746 38824 2768
rect 1104 2694 14315 2746
rect 14367 2694 14379 2746
rect 14431 2694 14443 2746
rect 14495 2694 14507 2746
rect 14559 2694 27648 2746
rect 27700 2694 27712 2746
rect 27764 2694 27776 2746
rect 27828 2694 27840 2746
rect 27892 2694 38824 2746
rect 1104 2672 38824 2694
rect 2041 2635 2099 2641
rect 2041 2601 2053 2635
rect 2087 2632 2099 2635
rect 2130 2632 2136 2644
rect 2087 2604 2136 2632
rect 2087 2601 2099 2604
rect 2041 2595 2099 2601
rect 2130 2592 2136 2604
rect 2188 2592 2194 2644
rect 2774 2632 2780 2644
rect 2735 2604 2780 2632
rect 2774 2592 2780 2604
rect 2832 2592 2838 2644
rect 3510 2632 3516 2644
rect 3471 2604 3516 2632
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 4982 2632 4988 2644
rect 4943 2604 4988 2632
rect 4982 2592 4988 2604
rect 5040 2632 5046 2644
rect 7098 2632 7104 2644
rect 5040 2604 5120 2632
rect 7059 2604 7104 2632
rect 5040 2592 5046 2604
rect 1581 2499 1639 2505
rect 1581 2465 1593 2499
rect 1627 2496 1639 2499
rect 2792 2496 2820 2592
rect 1627 2468 2820 2496
rect 2869 2499 2927 2505
rect 1627 2465 1639 2468
rect 1581 2459 1639 2465
rect 2869 2465 2881 2499
rect 2915 2496 2927 2499
rect 3528 2496 3556 2592
rect 5092 2505 5120 2604
rect 7098 2592 7104 2604
rect 7156 2592 7162 2644
rect 7558 2632 7564 2644
rect 7519 2604 7564 2632
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 16758 2632 16764 2644
rect 16719 2604 16764 2632
rect 16758 2592 16764 2604
rect 16816 2592 16822 2644
rect 21818 2632 21824 2644
rect 21779 2604 21824 2632
rect 21818 2592 21824 2604
rect 21876 2592 21882 2644
rect 24857 2635 24915 2641
rect 24857 2601 24869 2635
rect 24903 2632 24915 2635
rect 25682 2632 25688 2644
rect 24903 2604 25688 2632
rect 24903 2601 24915 2604
rect 24857 2595 24915 2601
rect 2915 2468 3556 2496
rect 5077 2499 5135 2505
rect 2915 2465 2927 2468
rect 2869 2459 2927 2465
rect 5077 2465 5089 2499
rect 5123 2465 5135 2499
rect 5077 2459 5135 2465
rect 5261 2499 5319 2505
rect 5261 2465 5273 2499
rect 5307 2496 5319 2499
rect 5442 2496 5448 2508
rect 5307 2468 5448 2496
rect 5307 2465 5319 2468
rect 5261 2459 5319 2465
rect 1394 2428 1400 2440
rect 1355 2400 1400 2428
rect 1394 2388 1400 2400
rect 1452 2388 1458 2440
rect 4617 2431 4675 2437
rect 4617 2397 4629 2431
rect 4663 2428 4675 2431
rect 5276 2428 5304 2459
rect 5442 2456 5448 2468
rect 5500 2456 5506 2508
rect 5721 2499 5779 2505
rect 5721 2465 5733 2499
rect 5767 2496 5779 2499
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 5767 2468 6929 2496
rect 5767 2465 5779 2468
rect 5721 2459 5779 2465
rect 6917 2465 6929 2468
rect 6963 2496 6975 2499
rect 7576 2496 7604 2592
rect 6963 2468 7604 2496
rect 9217 2499 9275 2505
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 9217 2465 9229 2499
rect 9263 2496 9275 2499
rect 9953 2499 10011 2505
rect 9953 2496 9965 2499
rect 9263 2468 9965 2496
rect 9263 2465 9275 2468
rect 9217 2459 9275 2465
rect 9953 2465 9965 2468
rect 9999 2496 10011 2499
rect 10042 2496 10048 2508
rect 9999 2468 10048 2496
rect 9999 2465 10011 2468
rect 9953 2459 10011 2465
rect 10042 2456 10048 2468
rect 10100 2456 10106 2508
rect 10413 2499 10471 2505
rect 10413 2465 10425 2499
rect 10459 2496 10471 2499
rect 11241 2499 11299 2505
rect 11241 2496 11253 2499
rect 10459 2468 11253 2496
rect 10459 2465 10471 2468
rect 10413 2459 10471 2465
rect 11241 2465 11253 2468
rect 11287 2496 11299 2499
rect 11882 2496 11888 2508
rect 11287 2468 11888 2496
rect 11287 2465 11299 2468
rect 11241 2459 11299 2465
rect 11882 2456 11888 2468
rect 11940 2456 11946 2508
rect 15289 2499 15347 2505
rect 15289 2465 15301 2499
rect 15335 2496 15347 2499
rect 16298 2496 16304 2508
rect 15335 2468 16304 2496
rect 15335 2465 15347 2468
rect 15289 2459 15347 2465
rect 16298 2456 16304 2468
rect 16356 2456 16362 2508
rect 20625 2499 20683 2505
rect 20625 2465 20637 2499
rect 20671 2496 20683 2499
rect 21361 2499 21419 2505
rect 21361 2496 21373 2499
rect 20671 2468 21373 2496
rect 20671 2465 20683 2468
rect 20625 2459 20683 2465
rect 21361 2465 21373 2468
rect 21407 2496 21419 2499
rect 21910 2496 21916 2508
rect 21407 2468 21916 2496
rect 21407 2465 21419 2468
rect 21361 2459 21419 2465
rect 21910 2456 21916 2468
rect 21968 2456 21974 2508
rect 24213 2499 24271 2505
rect 24213 2465 24225 2499
rect 24259 2496 24271 2499
rect 24872 2496 24900 2595
rect 25682 2592 25688 2604
rect 25740 2592 25746 2644
rect 26142 2592 26148 2644
rect 26200 2632 26206 2644
rect 26237 2635 26295 2641
rect 26237 2632 26249 2635
rect 26200 2604 26249 2632
rect 26200 2592 26206 2604
rect 26237 2601 26249 2604
rect 26283 2601 26295 2635
rect 26237 2595 26295 2601
rect 24259 2468 24900 2496
rect 25225 2499 25283 2505
rect 24259 2465 24271 2468
rect 24213 2459 24271 2465
rect 25225 2465 25237 2499
rect 25271 2496 25283 2499
rect 25314 2496 25320 2508
rect 25271 2468 25320 2496
rect 25271 2465 25283 2468
rect 25225 2459 25283 2465
rect 25314 2456 25320 2468
rect 25372 2456 25378 2508
rect 25501 2499 25559 2505
rect 25501 2465 25513 2499
rect 25547 2496 25559 2499
rect 26160 2496 26188 2592
rect 25547 2468 26188 2496
rect 26881 2499 26939 2505
rect 25547 2465 25559 2468
rect 25501 2459 25559 2465
rect 26881 2465 26893 2499
rect 26927 2496 26939 2499
rect 27522 2496 27528 2508
rect 26927 2468 27528 2496
rect 26927 2465 26939 2468
rect 26881 2459 26939 2465
rect 4663 2400 5304 2428
rect 9585 2431 9643 2437
rect 4663 2397 4675 2400
rect 4617 2391 4675 2397
rect 9585 2397 9597 2431
rect 9631 2428 9643 2431
rect 9766 2428 9772 2440
rect 9631 2400 9772 2428
rect 9631 2397 9643 2400
rect 9585 2391 9643 2397
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 16117 2431 16175 2437
rect 16117 2397 16129 2431
rect 16163 2397 16175 2431
rect 16117 2391 16175 2397
rect 20993 2431 21051 2437
rect 20993 2397 21005 2431
rect 21039 2428 21051 2431
rect 21174 2428 21180 2440
rect 21039 2400 21180 2428
rect 21039 2397 21051 2400
rect 20993 2391 21051 2397
rect 1412 2360 1440 2388
rect 2317 2363 2375 2369
rect 2317 2360 2329 2363
rect 1412 2332 2329 2360
rect 2317 2329 2329 2332
rect 2363 2329 2375 2363
rect 2317 2323 2375 2329
rect 3050 2292 3056 2304
rect 3011 2264 3056 2292
rect 3050 2252 3056 2264
rect 3108 2252 3114 2304
rect 11422 2292 11428 2304
rect 11383 2264 11428 2292
rect 11422 2252 11428 2264
rect 11480 2252 11486 2304
rect 16022 2292 16028 2304
rect 15983 2264 16028 2292
rect 16022 2252 16028 2264
rect 16080 2292 16086 2304
rect 16132 2292 16160 2391
rect 21174 2388 21180 2400
rect 21232 2388 21238 2440
rect 25961 2431 26019 2437
rect 25961 2397 25973 2431
rect 26007 2428 26019 2431
rect 26896 2428 26924 2459
rect 27522 2456 27528 2468
rect 27580 2456 27586 2508
rect 26007 2400 26924 2428
rect 26007 2397 26019 2400
rect 25961 2391 26019 2397
rect 27062 2360 27068 2372
rect 27023 2332 27068 2360
rect 27062 2320 27068 2332
rect 27120 2320 27126 2372
rect 24394 2292 24400 2304
rect 16080 2264 16160 2292
rect 24355 2264 24400 2292
rect 16080 2252 16086 2264
rect 24394 2252 24400 2264
rect 24452 2252 24458 2304
rect 27522 2292 27528 2304
rect 27483 2264 27528 2292
rect 27522 2252 27528 2264
rect 27580 2252 27586 2304
rect 1104 2202 38824 2224
rect 1104 2150 7648 2202
rect 7700 2150 7712 2202
rect 7764 2150 7776 2202
rect 7828 2150 7840 2202
rect 7892 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 34315 2202
rect 34367 2150 34379 2202
rect 34431 2150 34443 2202
rect 34495 2150 34507 2202
rect 34559 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 14315 13574 14367 13626
rect 14379 13574 14431 13626
rect 14443 13574 14495 13626
rect 14507 13574 14559 13626
rect 27648 13574 27700 13626
rect 27712 13574 27764 13626
rect 27776 13574 27828 13626
rect 27840 13574 27892 13626
rect 7648 13030 7700 13082
rect 7712 13030 7764 13082
rect 7776 13030 7828 13082
rect 7840 13030 7892 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 34315 13030 34367 13082
rect 34379 13030 34431 13082
rect 34443 13030 34495 13082
rect 34507 13030 34559 13082
rect 14315 12486 14367 12538
rect 14379 12486 14431 12538
rect 14443 12486 14495 12538
rect 14507 12486 14559 12538
rect 27648 12486 27700 12538
rect 27712 12486 27764 12538
rect 27776 12486 27828 12538
rect 27840 12486 27892 12538
rect 7648 11942 7700 11994
rect 7712 11942 7764 11994
rect 7776 11942 7828 11994
rect 7840 11942 7892 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 34315 11942 34367 11994
rect 34379 11942 34431 11994
rect 34443 11942 34495 11994
rect 34507 11942 34559 11994
rect 14315 11398 14367 11450
rect 14379 11398 14431 11450
rect 14443 11398 14495 11450
rect 14507 11398 14559 11450
rect 27648 11398 27700 11450
rect 27712 11398 27764 11450
rect 27776 11398 27828 11450
rect 27840 11398 27892 11450
rect 26240 11228 26292 11280
rect 27436 11228 27488 11280
rect 7648 10854 7700 10906
rect 7712 10854 7764 10906
rect 7776 10854 7828 10906
rect 7840 10854 7892 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 34315 10854 34367 10906
rect 34379 10854 34431 10906
rect 34443 10854 34495 10906
rect 34507 10854 34559 10906
rect 14315 10310 14367 10362
rect 14379 10310 14431 10362
rect 14443 10310 14495 10362
rect 14507 10310 14559 10362
rect 27648 10310 27700 10362
rect 27712 10310 27764 10362
rect 27776 10310 27828 10362
rect 27840 10310 27892 10362
rect 7648 9766 7700 9818
rect 7712 9766 7764 9818
rect 7776 9766 7828 9818
rect 7840 9766 7892 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 34315 9766 34367 9818
rect 34379 9766 34431 9818
rect 34443 9766 34495 9818
rect 34507 9766 34559 9818
rect 20168 9367 20220 9376
rect 20168 9333 20177 9367
rect 20177 9333 20211 9367
rect 20211 9333 20220 9367
rect 20168 9324 20220 9333
rect 20812 9367 20864 9376
rect 20812 9333 20821 9367
rect 20821 9333 20855 9367
rect 20855 9333 20864 9367
rect 20812 9324 20864 9333
rect 14315 9222 14367 9274
rect 14379 9222 14431 9274
rect 14443 9222 14495 9274
rect 14507 9222 14559 9274
rect 27648 9222 27700 9274
rect 27712 9222 27764 9274
rect 27776 9222 27828 9274
rect 27840 9222 27892 9274
rect 16488 9027 16540 9036
rect 16488 8993 16497 9027
rect 16497 8993 16531 9027
rect 16531 8993 16540 9027
rect 16488 8984 16540 8993
rect 23020 9027 23072 9036
rect 23020 8993 23029 9027
rect 23029 8993 23063 9027
rect 23063 8993 23072 9027
rect 23020 8984 23072 8993
rect 10232 8780 10284 8832
rect 16672 8823 16724 8832
rect 16672 8789 16681 8823
rect 16681 8789 16715 8823
rect 16715 8789 16724 8823
rect 16672 8780 16724 8789
rect 22836 8823 22888 8832
rect 22836 8789 22845 8823
rect 22845 8789 22879 8823
rect 22879 8789 22888 8823
rect 22836 8780 22888 8789
rect 7648 8678 7700 8730
rect 7712 8678 7764 8730
rect 7776 8678 7828 8730
rect 7840 8678 7892 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 34315 8678 34367 8730
rect 34379 8678 34431 8730
rect 34443 8678 34495 8730
rect 34507 8678 34559 8730
rect 16488 8619 16540 8628
rect 16488 8585 16497 8619
rect 16497 8585 16531 8619
rect 16531 8585 16540 8619
rect 16488 8576 16540 8585
rect 22560 8508 22612 8560
rect 10232 8415 10284 8424
rect 10232 8381 10241 8415
rect 10241 8381 10275 8415
rect 10275 8381 10284 8415
rect 10232 8372 10284 8381
rect 10416 8415 10468 8424
rect 10416 8381 10425 8415
rect 10425 8381 10459 8415
rect 10459 8381 10468 8415
rect 10416 8372 10468 8381
rect 10508 8372 10560 8424
rect 11336 8415 11388 8424
rect 11336 8381 11345 8415
rect 11345 8381 11379 8415
rect 11379 8381 11388 8415
rect 11336 8372 11388 8381
rect 22100 8372 22152 8424
rect 10968 8304 11020 8356
rect 23020 8347 23072 8356
rect 23020 8313 23029 8347
rect 23029 8313 23063 8347
rect 23063 8313 23072 8347
rect 23020 8304 23072 8313
rect 23388 8347 23440 8356
rect 23388 8313 23397 8347
rect 23397 8313 23431 8347
rect 23431 8313 23440 8347
rect 23388 8304 23440 8313
rect 10048 8279 10100 8288
rect 10048 8245 10057 8279
rect 10057 8245 10091 8279
rect 10091 8245 10100 8279
rect 10048 8236 10100 8245
rect 14315 8134 14367 8186
rect 14379 8134 14431 8186
rect 14443 8134 14495 8186
rect 14507 8134 14559 8186
rect 27648 8134 27700 8186
rect 27712 8134 27764 8186
rect 27776 8134 27828 8186
rect 27840 8134 27892 8186
rect 10416 8007 10468 8016
rect 10416 7973 10425 8007
rect 10425 7973 10459 8007
rect 10459 7973 10468 8007
rect 10416 7964 10468 7973
rect 10232 7896 10284 7948
rect 11152 7939 11204 7948
rect 11152 7905 11161 7939
rect 11161 7905 11195 7939
rect 11195 7905 11204 7939
rect 11152 7896 11204 7905
rect 11336 7939 11388 7948
rect 11336 7905 11345 7939
rect 11345 7905 11379 7939
rect 11379 7905 11388 7939
rect 11336 7896 11388 7905
rect 12072 7896 12124 7948
rect 11704 7828 11756 7880
rect 11888 7803 11940 7812
rect 11888 7769 11897 7803
rect 11897 7769 11931 7803
rect 11931 7769 11940 7803
rect 11888 7760 11940 7769
rect 10508 7692 10560 7744
rect 19708 7735 19760 7744
rect 19708 7701 19717 7735
rect 19717 7701 19751 7735
rect 19751 7701 19760 7735
rect 19708 7692 19760 7701
rect 7648 7590 7700 7642
rect 7712 7590 7764 7642
rect 7776 7590 7828 7642
rect 7840 7590 7892 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 34315 7590 34367 7642
rect 34379 7590 34431 7642
rect 34443 7590 34495 7642
rect 34507 7590 34559 7642
rect 10508 7488 10560 7540
rect 11336 7531 11388 7540
rect 11336 7497 11345 7531
rect 11345 7497 11379 7531
rect 11379 7497 11388 7531
rect 11336 7488 11388 7497
rect 11704 7531 11756 7540
rect 11704 7497 11713 7531
rect 11713 7497 11747 7531
rect 11747 7497 11756 7531
rect 11704 7488 11756 7497
rect 9864 7284 9916 7336
rect 10324 7284 10376 7336
rect 10508 7327 10560 7336
rect 10508 7293 10517 7327
rect 10517 7293 10551 7327
rect 10551 7293 10560 7327
rect 10508 7284 10560 7293
rect 12072 7327 12124 7336
rect 12072 7293 12081 7327
rect 12081 7293 12115 7327
rect 12115 7293 12124 7327
rect 12072 7284 12124 7293
rect 19248 7284 19300 7336
rect 19708 7259 19760 7268
rect 19708 7225 19717 7259
rect 19717 7225 19751 7259
rect 19751 7225 19760 7259
rect 19708 7216 19760 7225
rect 19892 7259 19944 7268
rect 19892 7225 19901 7259
rect 19901 7225 19935 7259
rect 19935 7225 19944 7259
rect 19892 7216 19944 7225
rect 20076 7259 20128 7268
rect 20076 7225 20085 7259
rect 20085 7225 20119 7259
rect 20119 7225 20128 7259
rect 20076 7216 20128 7225
rect 9772 7191 9824 7200
rect 9772 7157 9781 7191
rect 9781 7157 9815 7191
rect 9815 7157 9824 7191
rect 9772 7148 9824 7157
rect 19156 7191 19208 7200
rect 19156 7157 19165 7191
rect 19165 7157 19199 7191
rect 19199 7157 19208 7191
rect 19156 7148 19208 7157
rect 20628 7148 20680 7200
rect 14315 7046 14367 7098
rect 14379 7046 14431 7098
rect 14443 7046 14495 7098
rect 14507 7046 14559 7098
rect 27648 7046 27700 7098
rect 27712 7046 27764 7098
rect 27776 7046 27828 7098
rect 27840 7046 27892 7098
rect 9772 6987 9824 6996
rect 9772 6953 9781 6987
rect 9781 6953 9815 6987
rect 9815 6953 9824 6987
rect 9772 6944 9824 6953
rect 19892 6944 19944 6996
rect 9404 6876 9456 6928
rect 9864 6851 9916 6860
rect 9864 6817 9873 6851
rect 9873 6817 9907 6851
rect 9907 6817 9916 6851
rect 9864 6808 9916 6817
rect 10416 6876 10468 6928
rect 20076 6876 20128 6928
rect 20812 6876 20864 6928
rect 22744 6919 22796 6928
rect 22744 6885 22753 6919
rect 22753 6885 22787 6919
rect 22787 6885 22796 6919
rect 22744 6876 22796 6885
rect 22928 6919 22980 6928
rect 22928 6885 22937 6919
rect 22937 6885 22971 6919
rect 22971 6885 22980 6919
rect 22928 6876 22980 6885
rect 10508 6851 10560 6860
rect 10508 6817 10517 6851
rect 10517 6817 10551 6851
rect 10551 6817 10560 6851
rect 10508 6808 10560 6817
rect 10876 6851 10928 6860
rect 10876 6817 10885 6851
rect 10885 6817 10919 6851
rect 10919 6817 10928 6851
rect 10876 6808 10928 6817
rect 20720 6808 20772 6860
rect 21364 6808 21416 6860
rect 22008 6808 22060 6860
rect 22836 6851 22888 6860
rect 22836 6817 22845 6851
rect 22845 6817 22879 6851
rect 22879 6817 22888 6851
rect 22836 6808 22888 6817
rect 20812 6740 20864 6792
rect 21640 6783 21692 6792
rect 21640 6749 21649 6783
rect 21649 6749 21683 6783
rect 21683 6749 21692 6783
rect 21640 6740 21692 6749
rect 22560 6783 22612 6792
rect 22560 6749 22569 6783
rect 22569 6749 22603 6783
rect 22603 6749 22612 6783
rect 22560 6740 22612 6749
rect 23388 6740 23440 6792
rect 24400 6715 24452 6724
rect 24400 6681 24409 6715
rect 24409 6681 24443 6715
rect 24443 6681 24452 6715
rect 24400 6672 24452 6681
rect 7648 6502 7700 6554
rect 7712 6502 7764 6554
rect 7776 6502 7828 6554
rect 7840 6502 7892 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 34315 6502 34367 6554
rect 34379 6502 34431 6554
rect 34443 6502 34495 6554
rect 34507 6502 34559 6554
rect 9404 6443 9456 6452
rect 9404 6409 9413 6443
rect 9413 6409 9447 6443
rect 9447 6409 9456 6443
rect 9404 6400 9456 6409
rect 9864 6400 9916 6452
rect 10508 6443 10560 6452
rect 10508 6409 10517 6443
rect 10517 6409 10551 6443
rect 10551 6409 10560 6443
rect 10508 6400 10560 6409
rect 20076 6400 20128 6452
rect 21364 6443 21416 6452
rect 21364 6409 21373 6443
rect 21373 6409 21407 6443
rect 21407 6409 21416 6443
rect 21364 6400 21416 6409
rect 22836 6400 22888 6452
rect 10416 6332 10468 6384
rect 22744 6332 22796 6384
rect 24492 6332 24544 6384
rect 10876 6264 10928 6316
rect 24124 6307 24176 6316
rect 24124 6273 24133 6307
rect 24133 6273 24167 6307
rect 24167 6273 24176 6307
rect 24124 6264 24176 6273
rect 20904 6239 20956 6248
rect 20904 6205 20913 6239
rect 20913 6205 20947 6239
rect 20947 6205 20956 6239
rect 20904 6196 20956 6205
rect 22928 6196 22980 6248
rect 22560 6128 22612 6180
rect 24308 6171 24360 6180
rect 24308 6137 24317 6171
rect 24317 6137 24351 6171
rect 24351 6137 24360 6171
rect 24308 6128 24360 6137
rect 24400 6128 24452 6180
rect 25044 6171 25096 6180
rect 25044 6137 25053 6171
rect 25053 6137 25087 6171
rect 25087 6137 25096 6171
rect 25044 6128 25096 6137
rect 24124 6060 24176 6112
rect 14315 5958 14367 6010
rect 14379 5958 14431 6010
rect 14443 5958 14495 6010
rect 14507 5958 14559 6010
rect 27648 5958 27700 6010
rect 27712 5958 27764 6010
rect 27776 5958 27828 6010
rect 27840 5958 27892 6010
rect 24492 5856 24544 5908
rect 24308 5788 24360 5840
rect 7648 5414 7700 5466
rect 7712 5414 7764 5466
rect 7776 5414 7828 5466
rect 7840 5414 7892 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 34315 5414 34367 5466
rect 34379 5414 34431 5466
rect 34443 5414 34495 5466
rect 34507 5414 34559 5466
rect 3148 5108 3200 5160
rect 3516 5040 3568 5092
rect 3976 5015 4028 5024
rect 3976 4981 3985 5015
rect 3985 4981 4019 5015
rect 4019 4981 4028 5015
rect 3976 4972 4028 4981
rect 14315 4870 14367 4922
rect 14379 4870 14431 4922
rect 14443 4870 14495 4922
rect 14507 4870 14559 4922
rect 27648 4870 27700 4922
rect 27712 4870 27764 4922
rect 27776 4870 27828 4922
rect 27840 4870 27892 4922
rect 25044 4768 25096 4820
rect 5632 4700 5684 4752
rect 6000 4632 6052 4684
rect 3148 4607 3200 4616
rect 3148 4573 3157 4607
rect 3157 4573 3191 4607
rect 3191 4573 3200 4607
rect 3148 4564 3200 4573
rect 5448 4428 5500 4480
rect 7648 4326 7700 4378
rect 7712 4326 7764 4378
rect 7776 4326 7828 4378
rect 7840 4326 7892 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 34315 4326 34367 4378
rect 34379 4326 34431 4378
rect 34443 4326 34495 4378
rect 34507 4326 34559 4378
rect 6000 4267 6052 4276
rect 6000 4233 6009 4267
rect 6009 4233 6043 4267
rect 6043 4233 6052 4267
rect 6000 4224 6052 4233
rect 9128 4131 9180 4140
rect 9128 4097 9137 4131
rect 9137 4097 9171 4131
rect 9171 4097 9180 4131
rect 9128 4088 9180 4097
rect 18144 4088 18196 4140
rect 19248 4088 19300 4140
rect 21640 4088 21692 4140
rect 25044 4088 25096 4140
rect 3240 4020 3292 4072
rect 5632 4063 5684 4072
rect 5632 4029 5641 4063
rect 5641 4029 5675 4063
rect 5675 4029 5684 4063
rect 5632 4020 5684 4029
rect 3516 3995 3568 4004
rect 3516 3961 3519 3995
rect 3519 3961 3553 3995
rect 3553 3961 3568 3995
rect 3516 3952 3568 3961
rect 9496 3995 9548 4004
rect 9496 3961 9499 3995
rect 9499 3961 9533 3995
rect 9533 3961 9548 3995
rect 9496 3952 9548 3961
rect 17776 3995 17828 4004
rect 17776 3961 17785 3995
rect 17785 3961 17819 3995
rect 17819 3961 17828 3995
rect 17776 3952 17828 3961
rect 21364 3952 21416 4004
rect 2780 3884 2832 3936
rect 10048 3927 10100 3936
rect 10048 3893 10057 3927
rect 10057 3893 10091 3927
rect 10091 3893 10100 3927
rect 10048 3884 10100 3893
rect 18972 3927 19024 3936
rect 18972 3893 18981 3927
rect 18981 3893 19015 3927
rect 19015 3893 19024 3927
rect 18972 3884 19024 3893
rect 21916 3927 21968 3936
rect 21916 3893 21925 3927
rect 21925 3893 21959 3927
rect 21959 3893 21968 3927
rect 21916 3884 21968 3893
rect 24308 3884 24360 3936
rect 25596 3952 25648 4004
rect 26148 3927 26200 3936
rect 26148 3893 26157 3927
rect 26157 3893 26191 3927
rect 26191 3893 26200 3927
rect 26148 3884 26200 3893
rect 14315 3782 14367 3834
rect 14379 3782 14431 3834
rect 14443 3782 14495 3834
rect 14507 3782 14559 3834
rect 27648 3782 27700 3834
rect 27712 3782 27764 3834
rect 27776 3782 27828 3834
rect 27840 3782 27892 3834
rect 2044 3723 2096 3732
rect 2044 3689 2053 3723
rect 2053 3689 2087 3723
rect 2087 3689 2096 3723
rect 2044 3680 2096 3689
rect 3240 3723 3292 3732
rect 3240 3689 3249 3723
rect 3249 3689 3283 3723
rect 3283 3689 3292 3723
rect 3240 3680 3292 3689
rect 9128 3723 9180 3732
rect 9128 3689 9137 3723
rect 9137 3689 9171 3723
rect 9171 3689 9180 3723
rect 9128 3680 9180 3689
rect 18144 3723 18196 3732
rect 18144 3689 18153 3723
rect 18153 3689 18187 3723
rect 18187 3689 18196 3723
rect 18144 3680 18196 3689
rect 24308 3612 24360 3664
rect 23480 3544 23532 3596
rect 24216 3544 24268 3596
rect 3700 3340 3752 3392
rect 25228 3383 25280 3392
rect 25228 3349 25237 3383
rect 25237 3349 25271 3383
rect 25271 3349 25280 3383
rect 25228 3340 25280 3349
rect 7648 3238 7700 3290
rect 7712 3238 7764 3290
rect 7776 3238 7828 3290
rect 7840 3238 7892 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 34315 3238 34367 3290
rect 34379 3238 34431 3290
rect 34443 3238 34495 3290
rect 34507 3238 34559 3290
rect 2044 3111 2096 3120
rect 2044 3077 2053 3111
rect 2053 3077 2087 3111
rect 2087 3077 2096 3111
rect 2044 3068 2096 3077
rect 3976 3136 4028 3188
rect 16764 3136 16816 3188
rect 17132 3179 17184 3188
rect 17132 3145 17141 3179
rect 17141 3145 17175 3179
rect 17175 3145 17184 3179
rect 17132 3136 17184 3145
rect 22192 3179 22244 3188
rect 22192 3145 22201 3179
rect 22201 3145 22235 3179
rect 22235 3145 22244 3179
rect 22192 3136 22244 3145
rect 24216 3136 24268 3188
rect 25688 3179 25740 3188
rect 25688 3145 25697 3179
rect 25697 3145 25731 3179
rect 25731 3145 25740 3179
rect 25688 3136 25740 3145
rect 21732 3111 21784 3120
rect 21732 3077 21741 3111
rect 21741 3077 21775 3111
rect 21775 3077 21784 3111
rect 21732 3068 21784 3077
rect 24308 3068 24360 3120
rect 25228 3043 25280 3052
rect 25228 3009 25237 3043
rect 25237 3009 25271 3043
rect 25271 3009 25280 3043
rect 25228 3000 25280 3009
rect 16764 2932 16816 2984
rect 21824 2932 21876 2984
rect 22192 2932 22244 2984
rect 25044 2975 25096 2984
rect 25044 2941 25053 2975
rect 25053 2941 25087 2975
rect 25087 2941 25096 2975
rect 25044 2932 25096 2941
rect 2412 2839 2464 2848
rect 2412 2805 2421 2839
rect 2421 2805 2455 2839
rect 2455 2805 2464 2839
rect 2412 2796 2464 2805
rect 16672 2839 16724 2848
rect 16672 2805 16681 2839
rect 16681 2805 16715 2839
rect 16715 2805 16724 2839
rect 16672 2796 16724 2805
rect 14315 2694 14367 2746
rect 14379 2694 14431 2746
rect 14443 2694 14495 2746
rect 14507 2694 14559 2746
rect 27648 2694 27700 2746
rect 27712 2694 27764 2746
rect 27776 2694 27828 2746
rect 27840 2694 27892 2746
rect 2136 2592 2188 2644
rect 2780 2635 2832 2644
rect 2780 2601 2789 2635
rect 2789 2601 2823 2635
rect 2823 2601 2832 2635
rect 2780 2592 2832 2601
rect 3516 2635 3568 2644
rect 3516 2601 3525 2635
rect 3525 2601 3559 2635
rect 3559 2601 3568 2635
rect 3516 2592 3568 2601
rect 4988 2635 5040 2644
rect 4988 2601 4997 2635
rect 4997 2601 5031 2635
rect 5031 2601 5040 2635
rect 7104 2635 7156 2644
rect 4988 2592 5040 2601
rect 7104 2601 7113 2635
rect 7113 2601 7147 2635
rect 7147 2601 7156 2635
rect 7104 2592 7156 2601
rect 7564 2635 7616 2644
rect 7564 2601 7573 2635
rect 7573 2601 7607 2635
rect 7607 2601 7616 2635
rect 7564 2592 7616 2601
rect 16764 2635 16816 2644
rect 16764 2601 16773 2635
rect 16773 2601 16807 2635
rect 16807 2601 16816 2635
rect 16764 2592 16816 2601
rect 21824 2635 21876 2644
rect 21824 2601 21833 2635
rect 21833 2601 21867 2635
rect 21867 2601 21876 2635
rect 21824 2592 21876 2601
rect 1400 2431 1452 2440
rect 1400 2397 1409 2431
rect 1409 2397 1443 2431
rect 1443 2397 1452 2431
rect 1400 2388 1452 2397
rect 5448 2456 5500 2508
rect 10048 2456 10100 2508
rect 11888 2499 11940 2508
rect 11888 2465 11897 2499
rect 11897 2465 11931 2499
rect 11931 2465 11940 2499
rect 11888 2456 11940 2465
rect 16304 2499 16356 2508
rect 16304 2465 16313 2499
rect 16313 2465 16347 2499
rect 16347 2465 16356 2499
rect 16304 2456 16356 2465
rect 21916 2456 21968 2508
rect 25688 2592 25740 2644
rect 26148 2592 26200 2644
rect 25320 2499 25372 2508
rect 25320 2465 25329 2499
rect 25329 2465 25363 2499
rect 25363 2465 25372 2499
rect 25320 2456 25372 2465
rect 9772 2431 9824 2440
rect 9772 2397 9781 2431
rect 9781 2397 9815 2431
rect 9815 2397 9824 2431
rect 9772 2388 9824 2397
rect 21180 2431 21232 2440
rect 3056 2295 3108 2304
rect 3056 2261 3065 2295
rect 3065 2261 3099 2295
rect 3099 2261 3108 2295
rect 3056 2252 3108 2261
rect 11428 2295 11480 2304
rect 11428 2261 11437 2295
rect 11437 2261 11471 2295
rect 11471 2261 11480 2295
rect 11428 2252 11480 2261
rect 16028 2295 16080 2304
rect 16028 2261 16037 2295
rect 16037 2261 16071 2295
rect 16071 2261 16080 2295
rect 21180 2397 21189 2431
rect 21189 2397 21223 2431
rect 21223 2397 21232 2431
rect 21180 2388 21232 2397
rect 27528 2456 27580 2508
rect 27068 2363 27120 2372
rect 27068 2329 27077 2363
rect 27077 2329 27111 2363
rect 27111 2329 27120 2363
rect 27068 2320 27120 2329
rect 24400 2295 24452 2304
rect 16028 2252 16080 2261
rect 24400 2261 24409 2295
rect 24409 2261 24443 2295
rect 24443 2261 24452 2295
rect 24400 2252 24452 2261
rect 27528 2295 27580 2304
rect 27528 2261 27537 2295
rect 27537 2261 27571 2295
rect 27571 2261 27580 2295
rect 27528 2252 27580 2261
rect 7648 2150 7700 2202
rect 7712 2150 7764 2202
rect 7776 2150 7828 2202
rect 7840 2150 7892 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
rect 34315 2150 34367 2202
rect 34379 2150 34431 2202
rect 34443 2150 34495 2202
rect 34507 2150 34559 2202
<< metal2 >>
rect 2502 15520 2558 16000
rect 7470 15520 7526 16000
rect 12438 15520 12494 16000
rect 17498 15520 17554 16000
rect 22466 15520 22522 16000
rect 27434 15520 27490 16000
rect 32494 15520 32550 16000
rect 37462 15520 37518 16000
rect 2516 15450 2544 15520
rect 2056 15422 2544 15450
rect 2056 3738 2084 15422
rect 7484 11234 7512 15520
rect 7622 13084 7918 13104
rect 7678 13082 7702 13084
rect 7758 13082 7782 13084
rect 7838 13082 7862 13084
rect 7700 13030 7702 13082
rect 7764 13030 7776 13082
rect 7838 13030 7840 13082
rect 7678 13028 7702 13030
rect 7758 13028 7782 13030
rect 7838 13028 7862 13030
rect 7622 13008 7918 13028
rect 7622 11996 7918 12016
rect 7678 11994 7702 11996
rect 7758 11994 7782 11996
rect 7838 11994 7862 11996
rect 7700 11942 7702 11994
rect 7764 11942 7776 11994
rect 7838 11942 7840 11994
rect 7678 11940 7702 11942
rect 7758 11940 7782 11942
rect 7838 11940 7862 11942
rect 7622 11920 7918 11940
rect 7024 11206 7512 11234
rect 5998 7304 6054 7313
rect 5998 7239 6054 7248
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 3160 4622 3188 5102
rect 3516 5092 3568 5098
rect 3516 5034 3568 5040
rect 3148 4616 3200 4622
rect 3146 4584 3148 4593
rect 3200 4584 3202 4593
rect 3146 4519 3202 4528
rect 3240 4072 3292 4078
rect 3528 4049 3556 5034
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3240 4014 3292 4020
rect 3514 4040 3570 4049
rect 2780 3936 2832 3942
rect 3252 3913 3280 4014
rect 3514 3975 3516 3984
rect 3568 3975 3570 3984
rect 3516 3946 3568 3952
rect 2780 3878 2832 3884
rect 3238 3904 3294 3913
rect 2044 3732 2096 3738
rect 2044 3674 2096 3680
rect 2056 3210 2084 3674
rect 2056 3182 2176 3210
rect 2044 3120 2096 3126
rect 2042 3088 2044 3097
rect 2096 3088 2098 3097
rect 2042 3023 2098 3032
rect 2148 2650 2176 3182
rect 2412 2848 2464 2854
rect 2410 2816 2412 2825
rect 2464 2816 2466 2825
rect 2410 2751 2466 2760
rect 2792 2650 2820 3878
rect 3238 3839 3294 3848
rect 3252 3738 3280 3839
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3700 3392 3752 3398
rect 3700 3334 3752 3340
rect 3514 3088 3570 3097
rect 3514 3023 3570 3032
rect 3528 2650 3556 3023
rect 2136 2644 2188 2650
rect 2136 2586 2188 2592
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 1400 2440 1452 2446
rect 1400 2382 1452 2388
rect 1412 1578 1440 2382
rect 3056 2304 3108 2310
rect 3056 2246 3108 2252
rect 1228 1550 1440 1578
rect 1228 480 1256 1550
rect 3068 1465 3096 2246
rect 3054 1456 3110 1465
rect 3054 1391 3110 1400
rect 3712 480 3740 3334
rect 3988 3194 4016 4966
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 4986 2952 5042 2961
rect 4986 2887 5042 2896
rect 5000 2650 5028 2887
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 5460 2514 5488 4422
rect 5644 4078 5672 4694
rect 6012 4690 6040 7239
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 6012 4282 6040 4626
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 5632 4072 5684 4078
rect 5630 4040 5632 4049
rect 5684 4040 5686 4049
rect 5630 3975 5686 3984
rect 7024 3097 7052 11206
rect 7622 10908 7918 10928
rect 7678 10906 7702 10908
rect 7758 10906 7782 10908
rect 7838 10906 7862 10908
rect 7700 10854 7702 10906
rect 7764 10854 7776 10906
rect 7838 10854 7840 10906
rect 7678 10852 7702 10854
rect 7758 10852 7782 10854
rect 7838 10852 7862 10854
rect 7622 10832 7918 10852
rect 7622 9820 7918 9840
rect 7678 9818 7702 9820
rect 7758 9818 7782 9820
rect 7838 9818 7862 9820
rect 7700 9766 7702 9818
rect 7764 9766 7776 9818
rect 7838 9766 7840 9818
rect 7678 9764 7702 9766
rect 7758 9764 7782 9766
rect 7838 9764 7862 9766
rect 7622 9744 7918 9764
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 7622 8732 7918 8752
rect 7678 8730 7702 8732
rect 7758 8730 7782 8732
rect 7838 8730 7862 8732
rect 7700 8678 7702 8730
rect 7764 8678 7776 8730
rect 7838 8678 7840 8730
rect 7678 8676 7702 8678
rect 7758 8676 7782 8678
rect 7838 8676 7862 8678
rect 7622 8656 7918 8676
rect 10244 8430 10272 8774
rect 11150 8664 11206 8673
rect 11150 8599 11206 8608
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 7622 7644 7918 7664
rect 7678 7642 7702 7644
rect 7758 7642 7782 7644
rect 7838 7642 7862 7644
rect 7700 7590 7702 7642
rect 7764 7590 7776 7642
rect 7838 7590 7840 7642
rect 7678 7588 7702 7590
rect 7758 7588 7782 7590
rect 7838 7588 7862 7590
rect 7622 7568 7918 7588
rect 9864 7336 9916 7342
rect 9770 7304 9826 7313
rect 9864 7278 9916 7284
rect 9770 7239 9826 7248
rect 9784 7206 9812 7239
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 9404 6928 9456 6934
rect 9404 6870 9456 6876
rect 7622 6556 7918 6576
rect 7678 6554 7702 6556
rect 7758 6554 7782 6556
rect 7838 6554 7862 6556
rect 7700 6502 7702 6554
rect 7764 6502 7776 6554
rect 7838 6502 7840 6554
rect 7678 6500 7702 6502
rect 7758 6500 7782 6502
rect 7838 6500 7862 6502
rect 7622 6480 7918 6500
rect 9416 6458 9444 6870
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9126 5672 9182 5681
rect 9126 5607 9182 5616
rect 7622 5468 7918 5488
rect 7678 5466 7702 5468
rect 7758 5466 7782 5468
rect 7838 5466 7862 5468
rect 7700 5414 7702 5466
rect 7764 5414 7776 5466
rect 7838 5414 7840 5466
rect 7678 5412 7702 5414
rect 7758 5412 7782 5414
rect 7838 5412 7862 5414
rect 7622 5392 7918 5412
rect 7622 4380 7918 4400
rect 7678 4378 7702 4380
rect 7758 4378 7782 4380
rect 7838 4378 7862 4380
rect 7700 4326 7702 4378
rect 7764 4326 7776 4378
rect 7838 4326 7840 4378
rect 7678 4324 7702 4326
rect 7758 4324 7782 4326
rect 7838 4324 7862 4326
rect 7622 4304 7918 4324
rect 9140 4146 9168 5607
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9140 3738 9168 4082
rect 9494 4040 9550 4049
rect 9494 3975 9496 3984
rect 9548 3975 9550 3984
rect 9496 3946 9548 3952
rect 9784 3913 9812 6938
rect 9876 6866 9904 7278
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9876 6458 9904 6802
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9876 6225 9904 6394
rect 9862 6216 9918 6225
rect 9862 6151 9918 6160
rect 10060 4593 10088 8230
rect 10244 7954 10272 8366
rect 10428 8022 10456 8366
rect 10416 8016 10468 8022
rect 10416 7958 10468 7964
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 10428 7426 10456 7958
rect 10520 7750 10548 8366
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10520 7546 10548 7686
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10336 7398 10456 7426
rect 10336 7342 10364 7398
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 10428 6934 10456 7398
rect 10520 7342 10548 7482
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10416 6928 10468 6934
rect 10416 6870 10468 6876
rect 10428 6390 10456 6870
rect 10520 6866 10548 7278
rect 10980 6882 11008 8298
rect 11164 7954 11192 8599
rect 11334 8528 11390 8537
rect 11334 8463 11390 8472
rect 11348 8430 11376 8463
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 11348 7721 11376 7890
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11334 7712 11390 7721
rect 11334 7647 11390 7656
rect 11348 7546 11376 7647
rect 11716 7585 11744 7822
rect 11888 7812 11940 7818
rect 11888 7754 11940 7760
rect 11702 7576 11758 7585
rect 11336 7540 11388 7546
rect 11702 7511 11704 7520
rect 11336 7482 11388 7488
rect 11756 7511 11758 7520
rect 11704 7482 11756 7488
rect 10888 6866 11008 6882
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10876 6860 11008 6866
rect 10928 6854 11008 6860
rect 10876 6802 10928 6808
rect 10520 6458 10548 6802
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10416 6384 10468 6390
rect 10416 6326 10468 6332
rect 10888 6322 10916 6802
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 11900 5681 11928 7754
rect 12084 7342 12112 7890
rect 12072 7336 12124 7342
rect 12070 7304 12072 7313
rect 12124 7304 12126 7313
rect 12070 7239 12126 7248
rect 11886 5672 11942 5681
rect 11886 5607 11942 5616
rect 10046 4584 10102 4593
rect 10046 4519 10102 4528
rect 10048 3936 10100 3942
rect 9770 3904 9826 3913
rect 10048 3878 10100 3884
rect 9770 3839 9826 3848
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 7622 3292 7918 3312
rect 7678 3290 7702 3292
rect 7758 3290 7782 3292
rect 7838 3290 7862 3292
rect 7700 3238 7702 3290
rect 7764 3238 7776 3290
rect 7838 3238 7840 3290
rect 7678 3236 7702 3238
rect 7758 3236 7782 3238
rect 7838 3236 7862 3238
rect 7622 3216 7918 3236
rect 7010 3088 7066 3097
rect 7010 3023 7066 3032
rect 6182 2816 6238 2825
rect 6182 2751 6238 2760
rect 7102 2816 7158 2825
rect 7102 2751 7158 2760
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 6196 480 6224 2751
rect 7116 2650 7144 2751
rect 7562 2680 7618 2689
rect 7104 2644 7156 2650
rect 7562 2615 7564 2624
rect 7104 2586 7156 2592
rect 7616 2615 7618 2624
rect 7564 2586 7616 2592
rect 10060 2514 10088 3878
rect 11150 2952 11206 2961
rect 11150 2887 11206 2896
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 9772 2440 9824 2446
rect 9770 2408 9772 2417
rect 9824 2408 9826 2417
rect 9770 2343 9826 2352
rect 7622 2204 7918 2224
rect 7678 2202 7702 2204
rect 7758 2202 7782 2204
rect 7838 2202 7862 2204
rect 7700 2150 7702 2202
rect 7764 2150 7776 2202
rect 7838 2150 7840 2202
rect 7678 2148 7702 2150
rect 7758 2148 7782 2150
rect 7838 2148 7862 2150
rect 7622 2128 7918 2148
rect 8666 1456 8722 1465
rect 8666 1391 8722 1400
rect 8680 480 8708 1391
rect 11164 480 11192 2887
rect 12452 2689 12480 15520
rect 17512 15450 17540 15520
rect 22480 15450 22508 15520
rect 16868 15422 17540 15450
rect 22204 15422 22508 15450
rect 14289 13628 14585 13648
rect 14345 13626 14369 13628
rect 14425 13626 14449 13628
rect 14505 13626 14529 13628
rect 14367 13574 14369 13626
rect 14431 13574 14443 13626
rect 14505 13574 14507 13626
rect 14345 13572 14369 13574
rect 14425 13572 14449 13574
rect 14505 13572 14529 13574
rect 14289 13552 14585 13572
rect 14289 12540 14585 12560
rect 14345 12538 14369 12540
rect 14425 12538 14449 12540
rect 14505 12538 14529 12540
rect 14367 12486 14369 12538
rect 14431 12486 14443 12538
rect 14505 12486 14507 12538
rect 14345 12484 14369 12486
rect 14425 12484 14449 12486
rect 14505 12484 14529 12486
rect 14289 12464 14585 12484
rect 14289 11452 14585 11472
rect 14345 11450 14369 11452
rect 14425 11450 14449 11452
rect 14505 11450 14529 11452
rect 14367 11398 14369 11450
rect 14431 11398 14443 11450
rect 14505 11398 14507 11450
rect 14345 11396 14369 11398
rect 14425 11396 14449 11398
rect 14505 11396 14529 11398
rect 14289 11376 14585 11396
rect 14289 10364 14585 10384
rect 14345 10362 14369 10364
rect 14425 10362 14449 10364
rect 14505 10362 14529 10364
rect 14367 10310 14369 10362
rect 14431 10310 14443 10362
rect 14505 10310 14507 10362
rect 14345 10308 14369 10310
rect 14425 10308 14449 10310
rect 14505 10308 14529 10310
rect 14289 10288 14585 10308
rect 14289 9276 14585 9296
rect 14345 9274 14369 9276
rect 14425 9274 14449 9276
rect 14505 9274 14529 9276
rect 14367 9222 14369 9274
rect 14431 9222 14443 9274
rect 14505 9222 14507 9274
rect 14345 9220 14369 9222
rect 14425 9220 14449 9222
rect 14505 9220 14529 9222
rect 14289 9200 14585 9220
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 16500 8634 16528 8978
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16684 8673 16712 8774
rect 16670 8664 16726 8673
rect 16488 8628 16540 8634
rect 16670 8599 16726 8608
rect 16488 8570 16540 8576
rect 16500 8401 16528 8570
rect 16486 8392 16542 8401
rect 16486 8327 16542 8336
rect 14289 8188 14585 8208
rect 14345 8186 14369 8188
rect 14425 8186 14449 8188
rect 14505 8186 14529 8188
rect 14367 8134 14369 8186
rect 14431 8134 14443 8186
rect 14505 8134 14507 8186
rect 14345 8132 14369 8134
rect 14425 8132 14449 8134
rect 14505 8132 14529 8134
rect 14289 8112 14585 8132
rect 14289 7100 14585 7120
rect 14345 7098 14369 7100
rect 14425 7098 14449 7100
rect 14505 7098 14529 7100
rect 14367 7046 14369 7098
rect 14431 7046 14443 7098
rect 14505 7046 14507 7098
rect 14345 7044 14369 7046
rect 14425 7044 14449 7046
rect 14505 7044 14529 7046
rect 14289 7024 14585 7044
rect 14289 6012 14585 6032
rect 14345 6010 14369 6012
rect 14425 6010 14449 6012
rect 14505 6010 14529 6012
rect 14367 5958 14369 6010
rect 14431 5958 14443 6010
rect 14505 5958 14507 6010
rect 14345 5956 14369 5958
rect 14425 5956 14449 5958
rect 14505 5956 14529 5958
rect 14289 5936 14585 5956
rect 14289 4924 14585 4944
rect 14345 4922 14369 4924
rect 14425 4922 14449 4924
rect 14505 4922 14529 4924
rect 14367 4870 14369 4922
rect 14431 4870 14443 4922
rect 14505 4870 14507 4922
rect 14345 4868 14369 4870
rect 14425 4868 14449 4870
rect 14505 4868 14529 4870
rect 14289 4848 14585 4868
rect 14289 3836 14585 3856
rect 14345 3834 14369 3836
rect 14425 3834 14449 3836
rect 14505 3834 14529 3836
rect 14367 3782 14369 3834
rect 14431 3782 14443 3834
rect 14505 3782 14507 3834
rect 14345 3780 14369 3782
rect 14425 3780 14449 3782
rect 14505 3780 14529 3782
rect 14289 3760 14585 3780
rect 16302 3360 16358 3369
rect 16302 3295 16358 3304
rect 13634 2816 13690 2825
rect 13634 2751 13690 2760
rect 12438 2680 12494 2689
rect 12438 2615 12494 2624
rect 11886 2544 11942 2553
rect 11886 2479 11888 2488
rect 11940 2479 11942 2488
rect 11888 2450 11940 2456
rect 11428 2304 11480 2310
rect 11428 2246 11480 2252
rect 11440 1465 11468 2246
rect 11426 1456 11482 1465
rect 11426 1391 11482 1400
rect 13648 480 13676 2751
rect 14289 2748 14585 2768
rect 14345 2746 14369 2748
rect 14425 2746 14449 2748
rect 14505 2746 14529 2748
rect 14367 2694 14369 2746
rect 14431 2694 14443 2746
rect 14505 2694 14507 2746
rect 14345 2692 14369 2694
rect 14425 2692 14449 2694
rect 14505 2692 14529 2694
rect 14289 2672 14585 2692
rect 16316 2514 16344 3295
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 16776 2990 16804 3130
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 16672 2848 16724 2854
rect 16670 2816 16672 2825
rect 16724 2816 16726 2825
rect 16670 2751 16726 2760
rect 16776 2650 16804 2926
rect 16764 2644 16816 2650
rect 16764 2586 16816 2592
rect 16868 2553 16896 15422
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 20812 9376 20864 9382
rect 20812 9318 20864 9324
rect 20180 8537 20208 9318
rect 20166 8528 20222 8537
rect 20166 8463 20222 8472
rect 19890 8392 19946 8401
rect 19890 8327 19946 8336
rect 19708 7744 19760 7750
rect 19708 7686 19760 7692
rect 19720 7449 19748 7686
rect 19706 7440 19762 7449
rect 19706 7375 19762 7384
rect 19248 7336 19300 7342
rect 19248 7278 19300 7284
rect 19156 7200 19208 7206
rect 19156 7142 19208 7148
rect 19168 7041 19196 7142
rect 19154 7032 19210 7041
rect 19154 6967 19210 6976
rect 19260 4146 19288 7278
rect 19720 7274 19748 7375
rect 19904 7274 19932 8327
rect 19708 7268 19760 7274
rect 19708 7210 19760 7216
rect 19892 7268 19944 7274
rect 19892 7210 19944 7216
rect 20076 7268 20128 7274
rect 20076 7210 20128 7216
rect 19720 7177 19748 7210
rect 19706 7168 19762 7177
rect 19706 7103 19762 7112
rect 19904 7002 19932 7210
rect 20088 7041 20116 7210
rect 20628 7200 20680 7206
rect 20680 7148 20760 7154
rect 20628 7142 20760 7148
rect 20640 7126 20760 7142
rect 20074 7032 20130 7041
rect 19892 6996 19944 7002
rect 20074 6967 20130 6976
rect 19892 6938 19944 6944
rect 20088 6934 20116 6967
rect 20076 6928 20128 6934
rect 20076 6870 20128 6876
rect 20088 6458 20116 6870
rect 20732 6866 20760 7126
rect 20824 6934 20852 9318
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 22100 8424 22152 8430
rect 22100 8366 22152 8372
rect 22112 7834 22140 8366
rect 22020 7806 22140 7834
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 20812 6928 20864 6934
rect 20812 6870 20864 6876
rect 22020 6866 22048 7806
rect 22204 7698 22232 15422
rect 27448 11286 27476 15520
rect 27622 13628 27918 13648
rect 27678 13626 27702 13628
rect 27758 13626 27782 13628
rect 27838 13626 27862 13628
rect 27700 13574 27702 13626
rect 27764 13574 27776 13626
rect 27838 13574 27840 13626
rect 27678 13572 27702 13574
rect 27758 13572 27782 13574
rect 27838 13572 27862 13574
rect 27622 13552 27918 13572
rect 27622 12540 27918 12560
rect 27678 12538 27702 12540
rect 27758 12538 27782 12540
rect 27838 12538 27862 12540
rect 27700 12486 27702 12538
rect 27764 12486 27776 12538
rect 27838 12486 27840 12538
rect 27678 12484 27702 12486
rect 27758 12484 27782 12486
rect 27838 12484 27862 12486
rect 27622 12464 27918 12484
rect 27622 11452 27918 11472
rect 27678 11450 27702 11452
rect 27758 11450 27782 11452
rect 27838 11450 27862 11452
rect 27700 11398 27702 11450
rect 27764 11398 27776 11450
rect 27838 11398 27840 11450
rect 27678 11396 27702 11398
rect 27758 11396 27782 11398
rect 27838 11396 27862 11398
rect 27622 11376 27918 11396
rect 26240 11280 26292 11286
rect 26240 11222 26292 11228
rect 27436 11280 27488 11286
rect 27436 11222 27488 11228
rect 25686 10568 25742 10577
rect 25686 10503 25742 10512
rect 23020 9036 23072 9042
rect 23020 8978 23072 8984
rect 22836 8832 22888 8838
rect 22836 8774 22888 8780
rect 22560 8560 22612 8566
rect 22560 8502 22612 8508
rect 22742 8528 22798 8537
rect 22112 7670 22232 7698
rect 20720 6860 20772 6866
rect 20720 6802 20772 6808
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 22008 6860 22060 6866
rect 22008 6802 22060 6808
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 20824 6338 20852 6734
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 21376 6458 21404 6802
rect 21640 6792 21692 6798
rect 21640 6734 21692 6740
rect 21364 6452 21416 6458
rect 21364 6394 21416 6400
rect 20824 6310 20944 6338
rect 20916 6254 20944 6310
rect 20904 6248 20956 6254
rect 20902 6216 20904 6225
rect 20956 6216 20958 6225
rect 20902 6151 20958 6160
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 21652 4146 21680 6734
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 21640 4140 21692 4146
rect 21640 4082 21692 4088
rect 17774 4040 17830 4049
rect 17774 3975 17776 3984
rect 17828 3975 17830 3984
rect 17776 3946 17828 3952
rect 18156 3738 18184 4082
rect 21364 4004 21416 4010
rect 21364 3946 21416 3952
rect 18972 3936 19024 3942
rect 18972 3878 19024 3884
rect 18144 3732 18196 3738
rect 18144 3674 18196 3680
rect 17130 3496 17186 3505
rect 17130 3431 17186 3440
rect 17144 3194 17172 3431
rect 18984 3369 19012 3878
rect 21376 3777 21404 3946
rect 21916 3936 21968 3942
rect 21916 3878 21968 3884
rect 21362 3768 21418 3777
rect 21362 3703 21418 3712
rect 18970 3360 19026 3369
rect 18970 3295 19026 3304
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 21732 3120 21784 3126
rect 21730 3088 21732 3097
rect 21784 3088 21786 3097
rect 21730 3023 21786 3032
rect 21824 2984 21876 2990
rect 21824 2926 21876 2932
rect 21836 2650 21864 2926
rect 21824 2644 21876 2650
rect 21824 2586 21876 2592
rect 16854 2544 16910 2553
rect 16304 2508 16356 2514
rect 21928 2514 21956 3878
rect 22112 3505 22140 7670
rect 22572 7313 22600 8502
rect 22742 8463 22798 8472
rect 22558 7304 22614 7313
rect 22558 7239 22614 7248
rect 22572 6798 22600 7239
rect 22756 6934 22784 8463
rect 22848 7449 22876 8774
rect 23032 8362 23060 8978
rect 24490 8392 24546 8401
rect 23020 8356 23072 8362
rect 23020 8298 23072 8304
rect 23388 8356 23440 8362
rect 24490 8327 24546 8336
rect 23388 8298 23440 8304
rect 22834 7440 22890 7449
rect 22834 7375 22890 7384
rect 22744 6928 22796 6934
rect 22744 6870 22796 6876
rect 22560 6792 22612 6798
rect 22560 6734 22612 6740
rect 22572 6186 22600 6734
rect 22756 6390 22784 6870
rect 22848 6866 22876 7375
rect 22928 6928 22980 6934
rect 22928 6870 22980 6876
rect 22836 6860 22888 6866
rect 22836 6802 22888 6808
rect 22848 6458 22876 6802
rect 22836 6452 22888 6458
rect 22836 6394 22888 6400
rect 22744 6384 22796 6390
rect 22744 6326 22796 6332
rect 22940 6254 22968 6870
rect 22928 6248 22980 6254
rect 23032 6225 23060 8298
rect 23400 7857 23428 8298
rect 23386 7848 23442 7857
rect 23386 7783 23442 7792
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 24398 6760 24454 6769
rect 22928 6190 22980 6196
rect 23018 6216 23074 6225
rect 22560 6180 22612 6186
rect 23018 6151 23074 6160
rect 22560 6122 22612 6128
rect 23400 3618 23428 6734
rect 24398 6695 24400 6704
rect 24452 6695 24454 6704
rect 24400 6666 24452 6672
rect 24124 6316 24176 6322
rect 24124 6258 24176 6264
rect 24136 6225 24164 6258
rect 24122 6216 24178 6225
rect 24412 6186 24440 6666
rect 24504 6390 24532 8327
rect 24492 6384 24544 6390
rect 24492 6326 24544 6332
rect 24122 6151 24178 6160
rect 24308 6180 24360 6186
rect 24136 6118 24164 6151
rect 24308 6122 24360 6128
rect 24400 6180 24452 6186
rect 24400 6122 24452 6128
rect 24124 6112 24176 6118
rect 24124 6054 24176 6060
rect 24320 5846 24348 6122
rect 24504 5914 24532 6326
rect 25044 6180 25096 6186
rect 25044 6122 25096 6128
rect 24492 5908 24544 5914
rect 24492 5850 24544 5856
rect 24308 5840 24360 5846
rect 24308 5782 24360 5788
rect 25056 4826 25084 6122
rect 25044 4820 25096 4826
rect 25044 4762 25096 4768
rect 25056 4146 25084 4762
rect 25044 4140 25096 4146
rect 25044 4082 25096 4088
rect 25594 4040 25650 4049
rect 25594 3975 25596 3984
rect 25648 3975 25650 3984
rect 25596 3946 25648 3952
rect 24308 3936 24360 3942
rect 24308 3878 24360 3884
rect 24320 3777 24348 3878
rect 24306 3768 24362 3777
rect 24306 3703 24362 3712
rect 24320 3670 24348 3703
rect 24308 3664 24360 3670
rect 23400 3602 23520 3618
rect 24308 3606 24360 3612
rect 23400 3596 23532 3602
rect 23400 3590 23480 3596
rect 23480 3538 23532 3544
rect 24216 3596 24268 3602
rect 24216 3538 24268 3544
rect 22098 3496 22154 3505
rect 22098 3431 22154 3440
rect 22190 3224 22246 3233
rect 24228 3194 24256 3538
rect 22190 3159 22192 3168
rect 22244 3159 22246 3168
rect 24216 3188 24268 3194
rect 22192 3130 22244 3136
rect 24216 3130 24268 3136
rect 22204 2990 22232 3130
rect 24320 3126 24348 3606
rect 25228 3392 25280 3398
rect 25228 3334 25280 3340
rect 24308 3120 24360 3126
rect 24308 3062 24360 3068
rect 25240 3058 25268 3334
rect 25700 3194 25728 10503
rect 26148 3936 26200 3942
rect 26148 3878 26200 3884
rect 25688 3188 25740 3194
rect 25688 3130 25740 3136
rect 25228 3052 25280 3058
rect 25228 2994 25280 3000
rect 22192 2984 22244 2990
rect 25044 2984 25096 2990
rect 22192 2926 22244 2932
rect 25042 2952 25044 2961
rect 25096 2952 25098 2961
rect 25042 2887 25098 2896
rect 23662 2816 23718 2825
rect 23662 2751 23718 2760
rect 16854 2479 16910 2488
rect 21916 2508 21968 2514
rect 16304 2450 16356 2456
rect 21916 2450 21968 2456
rect 21180 2440 21232 2446
rect 16210 2408 16266 2417
rect 16210 2343 16266 2352
rect 21178 2408 21180 2417
rect 21232 2408 21234 2417
rect 21178 2343 21234 2352
rect 16028 2304 16080 2310
rect 16026 2272 16028 2281
rect 16080 2272 16082 2281
rect 16026 2207 16082 2216
rect 16224 480 16252 2343
rect 20810 2272 20866 2281
rect 20810 2207 20866 2216
rect 20824 1986 20852 2207
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 20824 1958 21220 1986
rect 18694 1456 18750 1465
rect 18694 1391 18750 1400
rect 18708 480 18736 1391
rect 21192 480 21220 1958
rect 23676 480 23704 2751
rect 25700 2650 25728 3130
rect 26160 2650 26188 3878
rect 26252 3233 26280 11222
rect 32508 10577 32536 15520
rect 35162 14648 35218 14657
rect 35162 14583 35218 14592
rect 34289 13084 34585 13104
rect 34345 13082 34369 13084
rect 34425 13082 34449 13084
rect 34505 13082 34529 13084
rect 34367 13030 34369 13082
rect 34431 13030 34443 13082
rect 34505 13030 34507 13082
rect 34345 13028 34369 13030
rect 34425 13028 34449 13030
rect 34505 13028 34529 13030
rect 34289 13008 34585 13028
rect 34289 11996 34585 12016
rect 34345 11994 34369 11996
rect 34425 11994 34449 11996
rect 34505 11994 34529 11996
rect 34367 11942 34369 11994
rect 34431 11942 34443 11994
rect 34505 11942 34507 11994
rect 34345 11940 34369 11942
rect 34425 11940 34449 11942
rect 34505 11940 34529 11942
rect 34289 11920 34585 11940
rect 34289 10908 34585 10928
rect 34345 10906 34369 10908
rect 34425 10906 34449 10908
rect 34505 10906 34529 10908
rect 34367 10854 34369 10906
rect 34431 10854 34443 10906
rect 34505 10854 34507 10906
rect 34345 10852 34369 10854
rect 34425 10852 34449 10854
rect 34505 10852 34529 10854
rect 34289 10832 34585 10852
rect 32494 10568 32550 10577
rect 32494 10503 32550 10512
rect 27622 10364 27918 10384
rect 27678 10362 27702 10364
rect 27758 10362 27782 10364
rect 27838 10362 27862 10364
rect 27700 10310 27702 10362
rect 27764 10310 27776 10362
rect 27838 10310 27840 10362
rect 27678 10308 27702 10310
rect 27758 10308 27782 10310
rect 27838 10308 27862 10310
rect 27622 10288 27918 10308
rect 34289 9820 34585 9840
rect 34345 9818 34369 9820
rect 34425 9818 34449 9820
rect 34505 9818 34529 9820
rect 34367 9766 34369 9818
rect 34431 9766 34443 9818
rect 34505 9766 34507 9818
rect 34345 9764 34369 9766
rect 34425 9764 34449 9766
rect 34505 9764 34529 9766
rect 34289 9744 34585 9764
rect 30930 9344 30986 9353
rect 27622 9276 27918 9296
rect 30930 9279 30986 9288
rect 27678 9274 27702 9276
rect 27758 9274 27782 9276
rect 27838 9274 27862 9276
rect 27700 9222 27702 9274
rect 27764 9222 27776 9274
rect 27838 9222 27840 9274
rect 27678 9220 27702 9222
rect 27758 9220 27782 9222
rect 27838 9220 27862 9222
rect 27622 9200 27918 9220
rect 30944 8537 30972 9279
rect 34289 8732 34585 8752
rect 34345 8730 34369 8732
rect 34425 8730 34449 8732
rect 34505 8730 34529 8732
rect 34367 8678 34369 8730
rect 34431 8678 34443 8730
rect 34505 8678 34507 8730
rect 34345 8676 34369 8678
rect 34425 8676 34449 8678
rect 34505 8676 34529 8678
rect 34289 8656 34585 8676
rect 30930 8528 30986 8537
rect 30930 8463 30986 8472
rect 27622 8188 27918 8208
rect 27678 8186 27702 8188
rect 27758 8186 27782 8188
rect 27838 8186 27862 8188
rect 27700 8134 27702 8186
rect 27764 8134 27776 8186
rect 27838 8134 27840 8186
rect 27678 8132 27702 8134
rect 27758 8132 27782 8134
rect 27838 8132 27862 8134
rect 27622 8112 27918 8132
rect 34289 7644 34585 7664
rect 34345 7642 34369 7644
rect 34425 7642 34449 7644
rect 34505 7642 34529 7644
rect 34367 7590 34369 7642
rect 34431 7590 34443 7642
rect 34505 7590 34507 7642
rect 34345 7588 34369 7590
rect 34425 7588 34449 7590
rect 34505 7588 34529 7590
rect 34289 7568 34585 7588
rect 27622 7100 27918 7120
rect 27678 7098 27702 7100
rect 27758 7098 27782 7100
rect 27838 7098 27862 7100
rect 27700 7046 27702 7098
rect 27764 7046 27776 7098
rect 27838 7046 27840 7098
rect 27678 7044 27702 7046
rect 27758 7044 27782 7046
rect 27838 7044 27862 7046
rect 27622 7024 27918 7044
rect 34610 6760 34666 6769
rect 34610 6695 34666 6704
rect 34289 6556 34585 6576
rect 34345 6554 34369 6556
rect 34425 6554 34449 6556
rect 34505 6554 34529 6556
rect 34367 6502 34369 6554
rect 34431 6502 34443 6554
rect 34505 6502 34507 6554
rect 34345 6500 34369 6502
rect 34425 6500 34449 6502
rect 34505 6500 34529 6502
rect 34289 6480 34585 6500
rect 27622 6012 27918 6032
rect 27678 6010 27702 6012
rect 27758 6010 27782 6012
rect 27838 6010 27862 6012
rect 27700 5958 27702 6010
rect 27764 5958 27776 6010
rect 27838 5958 27840 6010
rect 27678 5956 27702 5958
rect 27758 5956 27782 5958
rect 27838 5956 27862 5958
rect 27622 5936 27918 5956
rect 34289 5468 34585 5488
rect 34345 5466 34369 5468
rect 34425 5466 34449 5468
rect 34505 5466 34529 5468
rect 34367 5414 34369 5466
rect 34431 5414 34443 5466
rect 34505 5414 34507 5466
rect 34345 5412 34369 5414
rect 34425 5412 34449 5414
rect 34505 5412 34529 5414
rect 34289 5392 34585 5412
rect 27622 4924 27918 4944
rect 27678 4922 27702 4924
rect 27758 4922 27782 4924
rect 27838 4922 27862 4924
rect 27700 4870 27702 4922
rect 27764 4870 27776 4922
rect 27838 4870 27840 4922
rect 27678 4868 27702 4870
rect 27758 4868 27782 4870
rect 27838 4868 27862 4870
rect 27622 4848 27918 4868
rect 34289 4380 34585 4400
rect 34345 4378 34369 4380
rect 34425 4378 34449 4380
rect 34505 4378 34529 4380
rect 34367 4326 34369 4378
rect 34431 4326 34443 4378
rect 34505 4326 34507 4378
rect 34345 4324 34369 4326
rect 34425 4324 34449 4326
rect 34505 4324 34529 4326
rect 34289 4304 34585 4324
rect 27622 3836 27918 3856
rect 27678 3834 27702 3836
rect 27758 3834 27782 3836
rect 27838 3834 27862 3836
rect 27700 3782 27702 3834
rect 27764 3782 27776 3834
rect 27838 3782 27840 3834
rect 27678 3780 27702 3782
rect 27758 3780 27782 3782
rect 27838 3780 27862 3782
rect 27622 3760 27918 3780
rect 34289 3292 34585 3312
rect 34345 3290 34369 3292
rect 34425 3290 34449 3292
rect 34505 3290 34529 3292
rect 34367 3238 34369 3290
rect 34431 3238 34443 3290
rect 34505 3238 34507 3290
rect 34345 3236 34369 3238
rect 34425 3236 34449 3238
rect 34505 3236 34529 3238
rect 26238 3224 26294 3233
rect 34289 3216 34585 3236
rect 26238 3159 26294 3168
rect 28722 3088 28778 3097
rect 28722 3023 28778 3032
rect 27622 2748 27918 2768
rect 27678 2746 27702 2748
rect 27758 2746 27782 2748
rect 27838 2746 27862 2748
rect 27700 2694 27702 2746
rect 27764 2694 27776 2746
rect 27838 2694 27840 2746
rect 27678 2692 27702 2694
rect 27758 2692 27782 2694
rect 27838 2692 27862 2694
rect 27622 2672 27918 2692
rect 25688 2644 25740 2650
rect 25688 2586 25740 2592
rect 26148 2644 26200 2650
rect 26148 2586 26200 2592
rect 25318 2544 25374 2553
rect 25318 2479 25320 2488
rect 25372 2479 25374 2488
rect 27528 2508 27580 2514
rect 25320 2450 25372 2456
rect 27528 2450 27580 2456
rect 26146 2408 26202 2417
rect 26146 2343 26202 2352
rect 27066 2408 27122 2417
rect 27066 2343 27068 2352
rect 24400 2304 24452 2310
rect 24398 2272 24400 2281
rect 24452 2272 24454 2281
rect 24398 2207 24454 2216
rect 26160 480 26188 2343
rect 27120 2343 27122 2352
rect 27068 2314 27120 2320
rect 27540 2310 27568 2450
rect 27528 2304 27580 2310
rect 27528 2246 27580 2252
rect 27540 2009 27568 2246
rect 27526 2000 27582 2009
rect 27526 1935 27582 1944
rect 28736 480 28764 3023
rect 31206 2952 31262 2961
rect 31206 2887 31262 2896
rect 31220 480 31248 2887
rect 33690 2272 33746 2281
rect 33690 2207 33746 2216
rect 33704 480 33732 2207
rect 34289 2204 34585 2224
rect 34345 2202 34369 2204
rect 34425 2202 34449 2204
rect 34505 2202 34529 2204
rect 34367 2150 34369 2202
rect 34431 2150 34443 2202
rect 34505 2150 34507 2202
rect 34345 2148 34369 2150
rect 34425 2148 34449 2150
rect 34505 2148 34529 2150
rect 34289 2128 34585 2148
rect 34624 1329 34652 6695
rect 35176 4049 35204 14583
rect 35622 11928 35678 11937
rect 35622 11863 35678 11872
rect 35636 7857 35664 11863
rect 35622 7848 35678 7857
rect 35622 7783 35678 7792
rect 35162 4040 35218 4049
rect 35162 3975 35218 3984
rect 36174 2544 36230 2553
rect 36174 2479 36230 2488
rect 34610 1320 34666 1329
rect 34610 1255 34666 1264
rect 36188 480 36216 2479
rect 37476 2009 37504 15520
rect 38658 2408 38714 2417
rect 38658 2343 38714 2352
rect 37462 2000 37518 2009
rect 37462 1935 37518 1944
rect 38672 480 38700 2343
rect 1214 0 1270 480
rect 3698 0 3754 480
rect 6182 0 6238 480
rect 8666 0 8722 480
rect 11150 0 11206 480
rect 13634 0 13690 480
rect 16210 0 16266 480
rect 18694 0 18750 480
rect 21178 0 21234 480
rect 23662 0 23718 480
rect 26146 0 26202 480
rect 28722 0 28778 480
rect 31206 0 31262 480
rect 33690 0 33746 480
rect 36174 0 36230 480
rect 38658 0 38714 480
<< via2 >>
rect 7622 13082 7678 13084
rect 7702 13082 7758 13084
rect 7782 13082 7838 13084
rect 7862 13082 7918 13084
rect 7622 13030 7648 13082
rect 7648 13030 7678 13082
rect 7702 13030 7712 13082
rect 7712 13030 7758 13082
rect 7782 13030 7828 13082
rect 7828 13030 7838 13082
rect 7862 13030 7892 13082
rect 7892 13030 7918 13082
rect 7622 13028 7678 13030
rect 7702 13028 7758 13030
rect 7782 13028 7838 13030
rect 7862 13028 7918 13030
rect 7622 11994 7678 11996
rect 7702 11994 7758 11996
rect 7782 11994 7838 11996
rect 7862 11994 7918 11996
rect 7622 11942 7648 11994
rect 7648 11942 7678 11994
rect 7702 11942 7712 11994
rect 7712 11942 7758 11994
rect 7782 11942 7828 11994
rect 7828 11942 7838 11994
rect 7862 11942 7892 11994
rect 7892 11942 7918 11994
rect 7622 11940 7678 11942
rect 7702 11940 7758 11942
rect 7782 11940 7838 11942
rect 7862 11940 7918 11942
rect 5998 7248 6054 7304
rect 3146 4564 3148 4584
rect 3148 4564 3200 4584
rect 3200 4564 3202 4584
rect 3146 4528 3202 4564
rect 3514 4004 3570 4040
rect 3514 3984 3516 4004
rect 3516 3984 3568 4004
rect 3568 3984 3570 4004
rect 2042 3068 2044 3088
rect 2044 3068 2096 3088
rect 2096 3068 2098 3088
rect 2042 3032 2098 3068
rect 2410 2796 2412 2816
rect 2412 2796 2464 2816
rect 2464 2796 2466 2816
rect 2410 2760 2466 2796
rect 3238 3848 3294 3904
rect 3514 3032 3570 3088
rect 3054 1400 3110 1456
rect 4986 2896 5042 2952
rect 5630 4020 5632 4040
rect 5632 4020 5684 4040
rect 5684 4020 5686 4040
rect 5630 3984 5686 4020
rect 7622 10906 7678 10908
rect 7702 10906 7758 10908
rect 7782 10906 7838 10908
rect 7862 10906 7918 10908
rect 7622 10854 7648 10906
rect 7648 10854 7678 10906
rect 7702 10854 7712 10906
rect 7712 10854 7758 10906
rect 7782 10854 7828 10906
rect 7828 10854 7838 10906
rect 7862 10854 7892 10906
rect 7892 10854 7918 10906
rect 7622 10852 7678 10854
rect 7702 10852 7758 10854
rect 7782 10852 7838 10854
rect 7862 10852 7918 10854
rect 7622 9818 7678 9820
rect 7702 9818 7758 9820
rect 7782 9818 7838 9820
rect 7862 9818 7918 9820
rect 7622 9766 7648 9818
rect 7648 9766 7678 9818
rect 7702 9766 7712 9818
rect 7712 9766 7758 9818
rect 7782 9766 7828 9818
rect 7828 9766 7838 9818
rect 7862 9766 7892 9818
rect 7892 9766 7918 9818
rect 7622 9764 7678 9766
rect 7702 9764 7758 9766
rect 7782 9764 7838 9766
rect 7862 9764 7918 9766
rect 7622 8730 7678 8732
rect 7702 8730 7758 8732
rect 7782 8730 7838 8732
rect 7862 8730 7918 8732
rect 7622 8678 7648 8730
rect 7648 8678 7678 8730
rect 7702 8678 7712 8730
rect 7712 8678 7758 8730
rect 7782 8678 7828 8730
rect 7828 8678 7838 8730
rect 7862 8678 7892 8730
rect 7892 8678 7918 8730
rect 7622 8676 7678 8678
rect 7702 8676 7758 8678
rect 7782 8676 7838 8678
rect 7862 8676 7918 8678
rect 11150 8608 11206 8664
rect 7622 7642 7678 7644
rect 7702 7642 7758 7644
rect 7782 7642 7838 7644
rect 7862 7642 7918 7644
rect 7622 7590 7648 7642
rect 7648 7590 7678 7642
rect 7702 7590 7712 7642
rect 7712 7590 7758 7642
rect 7782 7590 7828 7642
rect 7828 7590 7838 7642
rect 7862 7590 7892 7642
rect 7892 7590 7918 7642
rect 7622 7588 7678 7590
rect 7702 7588 7758 7590
rect 7782 7588 7838 7590
rect 7862 7588 7918 7590
rect 9770 7248 9826 7304
rect 7622 6554 7678 6556
rect 7702 6554 7758 6556
rect 7782 6554 7838 6556
rect 7862 6554 7918 6556
rect 7622 6502 7648 6554
rect 7648 6502 7678 6554
rect 7702 6502 7712 6554
rect 7712 6502 7758 6554
rect 7782 6502 7828 6554
rect 7828 6502 7838 6554
rect 7862 6502 7892 6554
rect 7892 6502 7918 6554
rect 7622 6500 7678 6502
rect 7702 6500 7758 6502
rect 7782 6500 7838 6502
rect 7862 6500 7918 6502
rect 9126 5616 9182 5672
rect 7622 5466 7678 5468
rect 7702 5466 7758 5468
rect 7782 5466 7838 5468
rect 7862 5466 7918 5468
rect 7622 5414 7648 5466
rect 7648 5414 7678 5466
rect 7702 5414 7712 5466
rect 7712 5414 7758 5466
rect 7782 5414 7828 5466
rect 7828 5414 7838 5466
rect 7862 5414 7892 5466
rect 7892 5414 7918 5466
rect 7622 5412 7678 5414
rect 7702 5412 7758 5414
rect 7782 5412 7838 5414
rect 7862 5412 7918 5414
rect 7622 4378 7678 4380
rect 7702 4378 7758 4380
rect 7782 4378 7838 4380
rect 7862 4378 7918 4380
rect 7622 4326 7648 4378
rect 7648 4326 7678 4378
rect 7702 4326 7712 4378
rect 7712 4326 7758 4378
rect 7782 4326 7828 4378
rect 7828 4326 7838 4378
rect 7862 4326 7892 4378
rect 7892 4326 7918 4378
rect 7622 4324 7678 4326
rect 7702 4324 7758 4326
rect 7782 4324 7838 4326
rect 7862 4324 7918 4326
rect 9494 4004 9550 4040
rect 9494 3984 9496 4004
rect 9496 3984 9548 4004
rect 9548 3984 9550 4004
rect 9862 6160 9918 6216
rect 11334 8472 11390 8528
rect 11334 7656 11390 7712
rect 11702 7540 11758 7576
rect 11702 7520 11704 7540
rect 11704 7520 11756 7540
rect 11756 7520 11758 7540
rect 12070 7284 12072 7304
rect 12072 7284 12124 7304
rect 12124 7284 12126 7304
rect 12070 7248 12126 7284
rect 11886 5616 11942 5672
rect 10046 4528 10102 4584
rect 9770 3848 9826 3904
rect 7622 3290 7678 3292
rect 7702 3290 7758 3292
rect 7782 3290 7838 3292
rect 7862 3290 7918 3292
rect 7622 3238 7648 3290
rect 7648 3238 7678 3290
rect 7702 3238 7712 3290
rect 7712 3238 7758 3290
rect 7782 3238 7828 3290
rect 7828 3238 7838 3290
rect 7862 3238 7892 3290
rect 7892 3238 7918 3290
rect 7622 3236 7678 3238
rect 7702 3236 7758 3238
rect 7782 3236 7838 3238
rect 7862 3236 7918 3238
rect 7010 3032 7066 3088
rect 6182 2760 6238 2816
rect 7102 2760 7158 2816
rect 7562 2644 7618 2680
rect 7562 2624 7564 2644
rect 7564 2624 7616 2644
rect 7616 2624 7618 2644
rect 11150 2896 11206 2952
rect 9770 2388 9772 2408
rect 9772 2388 9824 2408
rect 9824 2388 9826 2408
rect 9770 2352 9826 2388
rect 7622 2202 7678 2204
rect 7702 2202 7758 2204
rect 7782 2202 7838 2204
rect 7862 2202 7918 2204
rect 7622 2150 7648 2202
rect 7648 2150 7678 2202
rect 7702 2150 7712 2202
rect 7712 2150 7758 2202
rect 7782 2150 7828 2202
rect 7828 2150 7838 2202
rect 7862 2150 7892 2202
rect 7892 2150 7918 2202
rect 7622 2148 7678 2150
rect 7702 2148 7758 2150
rect 7782 2148 7838 2150
rect 7862 2148 7918 2150
rect 8666 1400 8722 1456
rect 14289 13626 14345 13628
rect 14369 13626 14425 13628
rect 14449 13626 14505 13628
rect 14529 13626 14585 13628
rect 14289 13574 14315 13626
rect 14315 13574 14345 13626
rect 14369 13574 14379 13626
rect 14379 13574 14425 13626
rect 14449 13574 14495 13626
rect 14495 13574 14505 13626
rect 14529 13574 14559 13626
rect 14559 13574 14585 13626
rect 14289 13572 14345 13574
rect 14369 13572 14425 13574
rect 14449 13572 14505 13574
rect 14529 13572 14585 13574
rect 14289 12538 14345 12540
rect 14369 12538 14425 12540
rect 14449 12538 14505 12540
rect 14529 12538 14585 12540
rect 14289 12486 14315 12538
rect 14315 12486 14345 12538
rect 14369 12486 14379 12538
rect 14379 12486 14425 12538
rect 14449 12486 14495 12538
rect 14495 12486 14505 12538
rect 14529 12486 14559 12538
rect 14559 12486 14585 12538
rect 14289 12484 14345 12486
rect 14369 12484 14425 12486
rect 14449 12484 14505 12486
rect 14529 12484 14585 12486
rect 14289 11450 14345 11452
rect 14369 11450 14425 11452
rect 14449 11450 14505 11452
rect 14529 11450 14585 11452
rect 14289 11398 14315 11450
rect 14315 11398 14345 11450
rect 14369 11398 14379 11450
rect 14379 11398 14425 11450
rect 14449 11398 14495 11450
rect 14495 11398 14505 11450
rect 14529 11398 14559 11450
rect 14559 11398 14585 11450
rect 14289 11396 14345 11398
rect 14369 11396 14425 11398
rect 14449 11396 14505 11398
rect 14529 11396 14585 11398
rect 14289 10362 14345 10364
rect 14369 10362 14425 10364
rect 14449 10362 14505 10364
rect 14529 10362 14585 10364
rect 14289 10310 14315 10362
rect 14315 10310 14345 10362
rect 14369 10310 14379 10362
rect 14379 10310 14425 10362
rect 14449 10310 14495 10362
rect 14495 10310 14505 10362
rect 14529 10310 14559 10362
rect 14559 10310 14585 10362
rect 14289 10308 14345 10310
rect 14369 10308 14425 10310
rect 14449 10308 14505 10310
rect 14529 10308 14585 10310
rect 14289 9274 14345 9276
rect 14369 9274 14425 9276
rect 14449 9274 14505 9276
rect 14529 9274 14585 9276
rect 14289 9222 14315 9274
rect 14315 9222 14345 9274
rect 14369 9222 14379 9274
rect 14379 9222 14425 9274
rect 14449 9222 14495 9274
rect 14495 9222 14505 9274
rect 14529 9222 14559 9274
rect 14559 9222 14585 9274
rect 14289 9220 14345 9222
rect 14369 9220 14425 9222
rect 14449 9220 14505 9222
rect 14529 9220 14585 9222
rect 16670 8608 16726 8664
rect 16486 8336 16542 8392
rect 14289 8186 14345 8188
rect 14369 8186 14425 8188
rect 14449 8186 14505 8188
rect 14529 8186 14585 8188
rect 14289 8134 14315 8186
rect 14315 8134 14345 8186
rect 14369 8134 14379 8186
rect 14379 8134 14425 8186
rect 14449 8134 14495 8186
rect 14495 8134 14505 8186
rect 14529 8134 14559 8186
rect 14559 8134 14585 8186
rect 14289 8132 14345 8134
rect 14369 8132 14425 8134
rect 14449 8132 14505 8134
rect 14529 8132 14585 8134
rect 14289 7098 14345 7100
rect 14369 7098 14425 7100
rect 14449 7098 14505 7100
rect 14529 7098 14585 7100
rect 14289 7046 14315 7098
rect 14315 7046 14345 7098
rect 14369 7046 14379 7098
rect 14379 7046 14425 7098
rect 14449 7046 14495 7098
rect 14495 7046 14505 7098
rect 14529 7046 14559 7098
rect 14559 7046 14585 7098
rect 14289 7044 14345 7046
rect 14369 7044 14425 7046
rect 14449 7044 14505 7046
rect 14529 7044 14585 7046
rect 14289 6010 14345 6012
rect 14369 6010 14425 6012
rect 14449 6010 14505 6012
rect 14529 6010 14585 6012
rect 14289 5958 14315 6010
rect 14315 5958 14345 6010
rect 14369 5958 14379 6010
rect 14379 5958 14425 6010
rect 14449 5958 14495 6010
rect 14495 5958 14505 6010
rect 14529 5958 14559 6010
rect 14559 5958 14585 6010
rect 14289 5956 14345 5958
rect 14369 5956 14425 5958
rect 14449 5956 14505 5958
rect 14529 5956 14585 5958
rect 14289 4922 14345 4924
rect 14369 4922 14425 4924
rect 14449 4922 14505 4924
rect 14529 4922 14585 4924
rect 14289 4870 14315 4922
rect 14315 4870 14345 4922
rect 14369 4870 14379 4922
rect 14379 4870 14425 4922
rect 14449 4870 14495 4922
rect 14495 4870 14505 4922
rect 14529 4870 14559 4922
rect 14559 4870 14585 4922
rect 14289 4868 14345 4870
rect 14369 4868 14425 4870
rect 14449 4868 14505 4870
rect 14529 4868 14585 4870
rect 14289 3834 14345 3836
rect 14369 3834 14425 3836
rect 14449 3834 14505 3836
rect 14529 3834 14585 3836
rect 14289 3782 14315 3834
rect 14315 3782 14345 3834
rect 14369 3782 14379 3834
rect 14379 3782 14425 3834
rect 14449 3782 14495 3834
rect 14495 3782 14505 3834
rect 14529 3782 14559 3834
rect 14559 3782 14585 3834
rect 14289 3780 14345 3782
rect 14369 3780 14425 3782
rect 14449 3780 14505 3782
rect 14529 3780 14585 3782
rect 16302 3304 16358 3360
rect 13634 2760 13690 2816
rect 12438 2624 12494 2680
rect 11886 2508 11942 2544
rect 11886 2488 11888 2508
rect 11888 2488 11940 2508
rect 11940 2488 11942 2508
rect 11426 1400 11482 1456
rect 14289 2746 14345 2748
rect 14369 2746 14425 2748
rect 14449 2746 14505 2748
rect 14529 2746 14585 2748
rect 14289 2694 14315 2746
rect 14315 2694 14345 2746
rect 14369 2694 14379 2746
rect 14379 2694 14425 2746
rect 14449 2694 14495 2746
rect 14495 2694 14505 2746
rect 14529 2694 14559 2746
rect 14559 2694 14585 2746
rect 14289 2692 14345 2694
rect 14369 2692 14425 2694
rect 14449 2692 14505 2694
rect 14529 2692 14585 2694
rect 16670 2796 16672 2816
rect 16672 2796 16724 2816
rect 16724 2796 16726 2816
rect 16670 2760 16726 2796
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 20166 8472 20222 8528
rect 19890 8336 19946 8392
rect 19706 7384 19762 7440
rect 19154 6976 19210 7032
rect 19706 7112 19762 7168
rect 20074 6976 20130 7032
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 27622 13626 27678 13628
rect 27702 13626 27758 13628
rect 27782 13626 27838 13628
rect 27862 13626 27918 13628
rect 27622 13574 27648 13626
rect 27648 13574 27678 13626
rect 27702 13574 27712 13626
rect 27712 13574 27758 13626
rect 27782 13574 27828 13626
rect 27828 13574 27838 13626
rect 27862 13574 27892 13626
rect 27892 13574 27918 13626
rect 27622 13572 27678 13574
rect 27702 13572 27758 13574
rect 27782 13572 27838 13574
rect 27862 13572 27918 13574
rect 27622 12538 27678 12540
rect 27702 12538 27758 12540
rect 27782 12538 27838 12540
rect 27862 12538 27918 12540
rect 27622 12486 27648 12538
rect 27648 12486 27678 12538
rect 27702 12486 27712 12538
rect 27712 12486 27758 12538
rect 27782 12486 27828 12538
rect 27828 12486 27838 12538
rect 27862 12486 27892 12538
rect 27892 12486 27918 12538
rect 27622 12484 27678 12486
rect 27702 12484 27758 12486
rect 27782 12484 27838 12486
rect 27862 12484 27918 12486
rect 27622 11450 27678 11452
rect 27702 11450 27758 11452
rect 27782 11450 27838 11452
rect 27862 11450 27918 11452
rect 27622 11398 27648 11450
rect 27648 11398 27678 11450
rect 27702 11398 27712 11450
rect 27712 11398 27758 11450
rect 27782 11398 27828 11450
rect 27828 11398 27838 11450
rect 27862 11398 27892 11450
rect 27892 11398 27918 11450
rect 27622 11396 27678 11398
rect 27702 11396 27758 11398
rect 27782 11396 27838 11398
rect 27862 11396 27918 11398
rect 25686 10512 25742 10568
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 20902 6196 20904 6216
rect 20904 6196 20956 6216
rect 20956 6196 20958 6216
rect 20902 6160 20958 6196
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 17774 4004 17830 4040
rect 17774 3984 17776 4004
rect 17776 3984 17828 4004
rect 17828 3984 17830 4004
rect 17130 3440 17186 3496
rect 21362 3712 21418 3768
rect 18970 3304 19026 3360
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 21730 3068 21732 3088
rect 21732 3068 21784 3088
rect 21784 3068 21786 3088
rect 21730 3032 21786 3068
rect 16854 2488 16910 2544
rect 22742 8472 22798 8528
rect 22558 7248 22614 7304
rect 24490 8336 24546 8392
rect 22834 7384 22890 7440
rect 23386 7792 23442 7848
rect 23018 6160 23074 6216
rect 24398 6724 24454 6760
rect 24398 6704 24400 6724
rect 24400 6704 24452 6724
rect 24452 6704 24454 6724
rect 24122 6160 24178 6216
rect 25594 4004 25650 4040
rect 25594 3984 25596 4004
rect 25596 3984 25648 4004
rect 25648 3984 25650 4004
rect 24306 3712 24362 3768
rect 22098 3440 22154 3496
rect 22190 3188 22246 3224
rect 22190 3168 22192 3188
rect 22192 3168 22244 3188
rect 22244 3168 22246 3188
rect 25042 2932 25044 2952
rect 25044 2932 25096 2952
rect 25096 2932 25098 2952
rect 25042 2896 25098 2932
rect 23662 2760 23718 2816
rect 16210 2352 16266 2408
rect 21178 2388 21180 2408
rect 21180 2388 21232 2408
rect 21232 2388 21234 2408
rect 21178 2352 21234 2388
rect 16026 2252 16028 2272
rect 16028 2252 16080 2272
rect 16080 2252 16082 2272
rect 16026 2216 16082 2252
rect 20810 2216 20866 2272
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 18694 1400 18750 1456
rect 35162 14592 35218 14648
rect 34289 13082 34345 13084
rect 34369 13082 34425 13084
rect 34449 13082 34505 13084
rect 34529 13082 34585 13084
rect 34289 13030 34315 13082
rect 34315 13030 34345 13082
rect 34369 13030 34379 13082
rect 34379 13030 34425 13082
rect 34449 13030 34495 13082
rect 34495 13030 34505 13082
rect 34529 13030 34559 13082
rect 34559 13030 34585 13082
rect 34289 13028 34345 13030
rect 34369 13028 34425 13030
rect 34449 13028 34505 13030
rect 34529 13028 34585 13030
rect 34289 11994 34345 11996
rect 34369 11994 34425 11996
rect 34449 11994 34505 11996
rect 34529 11994 34585 11996
rect 34289 11942 34315 11994
rect 34315 11942 34345 11994
rect 34369 11942 34379 11994
rect 34379 11942 34425 11994
rect 34449 11942 34495 11994
rect 34495 11942 34505 11994
rect 34529 11942 34559 11994
rect 34559 11942 34585 11994
rect 34289 11940 34345 11942
rect 34369 11940 34425 11942
rect 34449 11940 34505 11942
rect 34529 11940 34585 11942
rect 34289 10906 34345 10908
rect 34369 10906 34425 10908
rect 34449 10906 34505 10908
rect 34529 10906 34585 10908
rect 34289 10854 34315 10906
rect 34315 10854 34345 10906
rect 34369 10854 34379 10906
rect 34379 10854 34425 10906
rect 34449 10854 34495 10906
rect 34495 10854 34505 10906
rect 34529 10854 34559 10906
rect 34559 10854 34585 10906
rect 34289 10852 34345 10854
rect 34369 10852 34425 10854
rect 34449 10852 34505 10854
rect 34529 10852 34585 10854
rect 32494 10512 32550 10568
rect 27622 10362 27678 10364
rect 27702 10362 27758 10364
rect 27782 10362 27838 10364
rect 27862 10362 27918 10364
rect 27622 10310 27648 10362
rect 27648 10310 27678 10362
rect 27702 10310 27712 10362
rect 27712 10310 27758 10362
rect 27782 10310 27828 10362
rect 27828 10310 27838 10362
rect 27862 10310 27892 10362
rect 27892 10310 27918 10362
rect 27622 10308 27678 10310
rect 27702 10308 27758 10310
rect 27782 10308 27838 10310
rect 27862 10308 27918 10310
rect 34289 9818 34345 9820
rect 34369 9818 34425 9820
rect 34449 9818 34505 9820
rect 34529 9818 34585 9820
rect 34289 9766 34315 9818
rect 34315 9766 34345 9818
rect 34369 9766 34379 9818
rect 34379 9766 34425 9818
rect 34449 9766 34495 9818
rect 34495 9766 34505 9818
rect 34529 9766 34559 9818
rect 34559 9766 34585 9818
rect 34289 9764 34345 9766
rect 34369 9764 34425 9766
rect 34449 9764 34505 9766
rect 34529 9764 34585 9766
rect 30930 9288 30986 9344
rect 27622 9274 27678 9276
rect 27702 9274 27758 9276
rect 27782 9274 27838 9276
rect 27862 9274 27918 9276
rect 27622 9222 27648 9274
rect 27648 9222 27678 9274
rect 27702 9222 27712 9274
rect 27712 9222 27758 9274
rect 27782 9222 27828 9274
rect 27828 9222 27838 9274
rect 27862 9222 27892 9274
rect 27892 9222 27918 9274
rect 27622 9220 27678 9222
rect 27702 9220 27758 9222
rect 27782 9220 27838 9222
rect 27862 9220 27918 9222
rect 34289 8730 34345 8732
rect 34369 8730 34425 8732
rect 34449 8730 34505 8732
rect 34529 8730 34585 8732
rect 34289 8678 34315 8730
rect 34315 8678 34345 8730
rect 34369 8678 34379 8730
rect 34379 8678 34425 8730
rect 34449 8678 34495 8730
rect 34495 8678 34505 8730
rect 34529 8678 34559 8730
rect 34559 8678 34585 8730
rect 34289 8676 34345 8678
rect 34369 8676 34425 8678
rect 34449 8676 34505 8678
rect 34529 8676 34585 8678
rect 30930 8472 30986 8528
rect 27622 8186 27678 8188
rect 27702 8186 27758 8188
rect 27782 8186 27838 8188
rect 27862 8186 27918 8188
rect 27622 8134 27648 8186
rect 27648 8134 27678 8186
rect 27702 8134 27712 8186
rect 27712 8134 27758 8186
rect 27782 8134 27828 8186
rect 27828 8134 27838 8186
rect 27862 8134 27892 8186
rect 27892 8134 27918 8186
rect 27622 8132 27678 8134
rect 27702 8132 27758 8134
rect 27782 8132 27838 8134
rect 27862 8132 27918 8134
rect 34289 7642 34345 7644
rect 34369 7642 34425 7644
rect 34449 7642 34505 7644
rect 34529 7642 34585 7644
rect 34289 7590 34315 7642
rect 34315 7590 34345 7642
rect 34369 7590 34379 7642
rect 34379 7590 34425 7642
rect 34449 7590 34495 7642
rect 34495 7590 34505 7642
rect 34529 7590 34559 7642
rect 34559 7590 34585 7642
rect 34289 7588 34345 7590
rect 34369 7588 34425 7590
rect 34449 7588 34505 7590
rect 34529 7588 34585 7590
rect 27622 7098 27678 7100
rect 27702 7098 27758 7100
rect 27782 7098 27838 7100
rect 27862 7098 27918 7100
rect 27622 7046 27648 7098
rect 27648 7046 27678 7098
rect 27702 7046 27712 7098
rect 27712 7046 27758 7098
rect 27782 7046 27828 7098
rect 27828 7046 27838 7098
rect 27862 7046 27892 7098
rect 27892 7046 27918 7098
rect 27622 7044 27678 7046
rect 27702 7044 27758 7046
rect 27782 7044 27838 7046
rect 27862 7044 27918 7046
rect 34610 6704 34666 6760
rect 34289 6554 34345 6556
rect 34369 6554 34425 6556
rect 34449 6554 34505 6556
rect 34529 6554 34585 6556
rect 34289 6502 34315 6554
rect 34315 6502 34345 6554
rect 34369 6502 34379 6554
rect 34379 6502 34425 6554
rect 34449 6502 34495 6554
rect 34495 6502 34505 6554
rect 34529 6502 34559 6554
rect 34559 6502 34585 6554
rect 34289 6500 34345 6502
rect 34369 6500 34425 6502
rect 34449 6500 34505 6502
rect 34529 6500 34585 6502
rect 27622 6010 27678 6012
rect 27702 6010 27758 6012
rect 27782 6010 27838 6012
rect 27862 6010 27918 6012
rect 27622 5958 27648 6010
rect 27648 5958 27678 6010
rect 27702 5958 27712 6010
rect 27712 5958 27758 6010
rect 27782 5958 27828 6010
rect 27828 5958 27838 6010
rect 27862 5958 27892 6010
rect 27892 5958 27918 6010
rect 27622 5956 27678 5958
rect 27702 5956 27758 5958
rect 27782 5956 27838 5958
rect 27862 5956 27918 5958
rect 34289 5466 34345 5468
rect 34369 5466 34425 5468
rect 34449 5466 34505 5468
rect 34529 5466 34585 5468
rect 34289 5414 34315 5466
rect 34315 5414 34345 5466
rect 34369 5414 34379 5466
rect 34379 5414 34425 5466
rect 34449 5414 34495 5466
rect 34495 5414 34505 5466
rect 34529 5414 34559 5466
rect 34559 5414 34585 5466
rect 34289 5412 34345 5414
rect 34369 5412 34425 5414
rect 34449 5412 34505 5414
rect 34529 5412 34585 5414
rect 27622 4922 27678 4924
rect 27702 4922 27758 4924
rect 27782 4922 27838 4924
rect 27862 4922 27918 4924
rect 27622 4870 27648 4922
rect 27648 4870 27678 4922
rect 27702 4870 27712 4922
rect 27712 4870 27758 4922
rect 27782 4870 27828 4922
rect 27828 4870 27838 4922
rect 27862 4870 27892 4922
rect 27892 4870 27918 4922
rect 27622 4868 27678 4870
rect 27702 4868 27758 4870
rect 27782 4868 27838 4870
rect 27862 4868 27918 4870
rect 34289 4378 34345 4380
rect 34369 4378 34425 4380
rect 34449 4378 34505 4380
rect 34529 4378 34585 4380
rect 34289 4326 34315 4378
rect 34315 4326 34345 4378
rect 34369 4326 34379 4378
rect 34379 4326 34425 4378
rect 34449 4326 34495 4378
rect 34495 4326 34505 4378
rect 34529 4326 34559 4378
rect 34559 4326 34585 4378
rect 34289 4324 34345 4326
rect 34369 4324 34425 4326
rect 34449 4324 34505 4326
rect 34529 4324 34585 4326
rect 27622 3834 27678 3836
rect 27702 3834 27758 3836
rect 27782 3834 27838 3836
rect 27862 3834 27918 3836
rect 27622 3782 27648 3834
rect 27648 3782 27678 3834
rect 27702 3782 27712 3834
rect 27712 3782 27758 3834
rect 27782 3782 27828 3834
rect 27828 3782 27838 3834
rect 27862 3782 27892 3834
rect 27892 3782 27918 3834
rect 27622 3780 27678 3782
rect 27702 3780 27758 3782
rect 27782 3780 27838 3782
rect 27862 3780 27918 3782
rect 34289 3290 34345 3292
rect 34369 3290 34425 3292
rect 34449 3290 34505 3292
rect 34529 3290 34585 3292
rect 34289 3238 34315 3290
rect 34315 3238 34345 3290
rect 34369 3238 34379 3290
rect 34379 3238 34425 3290
rect 34449 3238 34495 3290
rect 34495 3238 34505 3290
rect 34529 3238 34559 3290
rect 34559 3238 34585 3290
rect 34289 3236 34345 3238
rect 34369 3236 34425 3238
rect 34449 3236 34505 3238
rect 34529 3236 34585 3238
rect 26238 3168 26294 3224
rect 28722 3032 28778 3088
rect 27622 2746 27678 2748
rect 27702 2746 27758 2748
rect 27782 2746 27838 2748
rect 27862 2746 27918 2748
rect 27622 2694 27648 2746
rect 27648 2694 27678 2746
rect 27702 2694 27712 2746
rect 27712 2694 27758 2746
rect 27782 2694 27828 2746
rect 27828 2694 27838 2746
rect 27862 2694 27892 2746
rect 27892 2694 27918 2746
rect 27622 2692 27678 2694
rect 27702 2692 27758 2694
rect 27782 2692 27838 2694
rect 27862 2692 27918 2694
rect 25318 2508 25374 2544
rect 25318 2488 25320 2508
rect 25320 2488 25372 2508
rect 25372 2488 25374 2508
rect 26146 2352 26202 2408
rect 27066 2372 27122 2408
rect 27066 2352 27068 2372
rect 27068 2352 27120 2372
rect 27120 2352 27122 2372
rect 24398 2252 24400 2272
rect 24400 2252 24452 2272
rect 24452 2252 24454 2272
rect 24398 2216 24454 2252
rect 27526 1944 27582 2000
rect 31206 2896 31262 2952
rect 33690 2216 33746 2272
rect 34289 2202 34345 2204
rect 34369 2202 34425 2204
rect 34449 2202 34505 2204
rect 34529 2202 34585 2204
rect 34289 2150 34315 2202
rect 34315 2150 34345 2202
rect 34369 2150 34379 2202
rect 34379 2150 34425 2202
rect 34449 2150 34495 2202
rect 34495 2150 34505 2202
rect 34529 2150 34559 2202
rect 34559 2150 34585 2202
rect 34289 2148 34345 2150
rect 34369 2148 34425 2150
rect 34449 2148 34505 2150
rect 34529 2148 34585 2150
rect 35622 11872 35678 11928
rect 35622 7792 35678 7848
rect 35162 3984 35218 4040
rect 36174 2488 36230 2544
rect 34610 1264 34666 1320
rect 38658 2352 38714 2408
rect 37462 1944 37518 2000
<< metal3 >>
rect 35157 14650 35223 14653
rect 39520 14650 40000 14680
rect 35157 14648 40000 14650
rect 35157 14592 35162 14648
rect 35218 14592 40000 14648
rect 35157 14590 40000 14592
rect 35157 14587 35223 14590
rect 39520 14560 40000 14590
rect 14277 13632 14597 13633
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 13567 14597 13568
rect 27610 13632 27930 13633
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 13567 27930 13568
rect 7610 13088 7930 13089
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7930 13088
rect 7610 13023 7930 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 34277 13088 34597 13089
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 13023 34597 13024
rect 14277 12544 14597 12545
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 12479 14597 12480
rect 27610 12544 27930 12545
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 12479 27930 12480
rect 7610 12000 7930 12001
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7930 12000
rect 7610 11935 7930 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 34277 12000 34597 12001
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 34277 11935 34597 11936
rect 35617 11930 35683 11933
rect 39520 11930 40000 11960
rect 35617 11928 40000 11930
rect 35617 11872 35622 11928
rect 35678 11872 40000 11928
rect 35617 11870 40000 11872
rect 35617 11867 35683 11870
rect 39520 11840 40000 11870
rect 14277 11456 14597 11457
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 11391 14597 11392
rect 27610 11456 27930 11457
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 11391 27930 11392
rect 7610 10912 7930 10913
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7930 10912
rect 7610 10847 7930 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 34277 10912 34597 10913
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 10847 34597 10848
rect 25681 10570 25747 10573
rect 32489 10570 32555 10573
rect 25681 10568 32555 10570
rect 25681 10512 25686 10568
rect 25742 10512 32494 10568
rect 32550 10512 32555 10568
rect 25681 10510 32555 10512
rect 25681 10507 25747 10510
rect 32489 10507 32555 10510
rect 14277 10368 14597 10369
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 10303 14597 10304
rect 27610 10368 27930 10369
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 10303 27930 10304
rect 7610 9824 7930 9825
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7930 9824
rect 7610 9759 7930 9760
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 34277 9824 34597 9825
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 9759 34597 9760
rect 30925 9346 30991 9349
rect 39520 9346 40000 9376
rect 30925 9344 40000 9346
rect 30925 9288 30930 9344
rect 30986 9288 40000 9344
rect 30925 9286 40000 9288
rect 30925 9283 30991 9286
rect 14277 9280 14597 9281
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 9215 14597 9216
rect 27610 9280 27930 9281
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 39520 9256 40000 9286
rect 27610 9215 27930 9216
rect 7610 8736 7930 8737
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7930 8736
rect 7610 8671 7930 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 34277 8736 34597 8737
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 8671 34597 8672
rect 11145 8666 11211 8669
rect 16665 8666 16731 8669
rect 11145 8664 16731 8666
rect 11145 8608 11150 8664
rect 11206 8608 16670 8664
rect 16726 8608 16731 8664
rect 11145 8606 16731 8608
rect 11145 8603 11211 8606
rect 16665 8603 16731 8606
rect 11329 8530 11395 8533
rect 20161 8530 20227 8533
rect 22737 8530 22803 8533
rect 30925 8530 30991 8533
rect 11329 8528 22803 8530
rect 11329 8472 11334 8528
rect 11390 8472 20166 8528
rect 20222 8472 22742 8528
rect 22798 8472 22803 8528
rect 11329 8470 22803 8472
rect 11329 8467 11395 8470
rect 20161 8467 20227 8470
rect 22737 8467 22803 8470
rect 26190 8528 30991 8530
rect 26190 8472 30930 8528
rect 30986 8472 30991 8528
rect 26190 8470 30991 8472
rect 16481 8394 16547 8397
rect 19885 8394 19951 8397
rect 16481 8392 19951 8394
rect 16481 8336 16486 8392
rect 16542 8336 19890 8392
rect 19946 8336 19951 8392
rect 16481 8334 19951 8336
rect 16481 8331 16547 8334
rect 19885 8331 19951 8334
rect 24485 8394 24551 8397
rect 26190 8394 26250 8470
rect 30925 8467 30991 8470
rect 24485 8392 26250 8394
rect 24485 8336 24490 8392
rect 24546 8336 26250 8392
rect 24485 8334 26250 8336
rect 24485 8331 24551 8334
rect 14277 8192 14597 8193
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 8127 14597 8128
rect 27610 8192 27930 8193
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 8127 27930 8128
rect 23381 7850 23447 7853
rect 35617 7850 35683 7853
rect 23381 7848 35683 7850
rect 23381 7792 23386 7848
rect 23442 7792 35622 7848
rect 35678 7792 35683 7848
rect 23381 7790 35683 7792
rect 23381 7787 23447 7790
rect 35617 7787 35683 7790
rect 11329 7714 11395 7717
rect 11329 7712 17234 7714
rect 11329 7656 11334 7712
rect 11390 7656 17234 7712
rect 11329 7654 17234 7656
rect 11329 7651 11395 7654
rect 7610 7648 7930 7649
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7930 7648
rect 7610 7583 7930 7584
rect 11697 7578 11763 7581
rect 11697 7576 17050 7578
rect 11697 7520 11702 7576
rect 11758 7520 17050 7576
rect 11697 7518 17050 7520
rect 11697 7515 11763 7518
rect 5993 7306 6059 7309
rect 9765 7306 9831 7309
rect 5993 7304 9831 7306
rect 5993 7248 5998 7304
rect 6054 7248 9770 7304
rect 9826 7248 9831 7304
rect 5993 7246 9831 7248
rect 5993 7243 6059 7246
rect 9765 7243 9831 7246
rect 12065 7306 12131 7309
rect 12065 7304 16912 7306
rect 12065 7248 12070 7304
rect 12126 7248 16912 7304
rect 12065 7246 16912 7248
rect 12065 7243 12131 7246
rect 14277 7104 14597 7105
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 7039 14597 7040
rect 16852 7034 16912 7246
rect 16990 7170 17050 7518
rect 17174 7306 17234 7654
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 34277 7648 34597 7649
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 7583 34597 7584
rect 19701 7442 19767 7445
rect 22829 7442 22895 7445
rect 19701 7440 22895 7442
rect 19701 7384 19706 7440
rect 19762 7384 22834 7440
rect 22890 7384 22895 7440
rect 19701 7382 22895 7384
rect 19701 7379 19767 7382
rect 22829 7379 22895 7382
rect 22553 7306 22619 7309
rect 17174 7304 22619 7306
rect 17174 7248 22558 7304
rect 22614 7248 22619 7304
rect 17174 7246 22619 7248
rect 22553 7243 22619 7246
rect 19701 7170 19767 7173
rect 16990 7168 19767 7170
rect 16990 7112 19706 7168
rect 19762 7112 19767 7168
rect 16990 7110 19767 7112
rect 19701 7107 19767 7110
rect 27610 7104 27930 7105
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 7039 27930 7040
rect 19149 7034 19215 7037
rect 20069 7034 20135 7037
rect 16852 7032 20135 7034
rect 16852 6976 19154 7032
rect 19210 6976 20074 7032
rect 20130 6976 20135 7032
rect 16852 6974 20135 6976
rect 19149 6971 19215 6974
rect 20069 6971 20135 6974
rect 24393 6762 24459 6765
rect 34605 6762 34671 6765
rect 24393 6760 34671 6762
rect 24393 6704 24398 6760
rect 24454 6704 34610 6760
rect 34666 6704 34671 6760
rect 24393 6702 34671 6704
rect 24393 6699 24459 6702
rect 34605 6699 34671 6702
rect 39520 6626 40000 6656
rect 35574 6566 40000 6626
rect 7610 6560 7930 6561
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7930 6560
rect 7610 6495 7930 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 34277 6560 34597 6561
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 6495 34597 6496
rect 9857 6218 9923 6221
rect 20897 6218 20963 6221
rect 23013 6218 23079 6221
rect 24117 6218 24183 6221
rect 35574 6218 35634 6566
rect 39520 6536 40000 6566
rect 9857 6216 35634 6218
rect 9857 6160 9862 6216
rect 9918 6160 20902 6216
rect 20958 6160 23018 6216
rect 23074 6160 24122 6216
rect 24178 6160 35634 6216
rect 9857 6158 35634 6160
rect 9857 6155 9923 6158
rect 20897 6155 20963 6158
rect 23013 6155 23079 6158
rect 24117 6155 24183 6158
rect 14277 6016 14597 6017
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 5951 14597 5952
rect 27610 6016 27930 6017
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 5951 27930 5952
rect 9121 5674 9187 5677
rect 11881 5674 11947 5677
rect 9121 5672 11947 5674
rect 9121 5616 9126 5672
rect 9182 5616 11886 5672
rect 11942 5616 11947 5672
rect 9121 5614 11947 5616
rect 9121 5611 9187 5614
rect 11881 5611 11947 5614
rect 7610 5472 7930 5473
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7930 5472
rect 7610 5407 7930 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 34277 5472 34597 5473
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 5407 34597 5408
rect 14277 4928 14597 4929
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 4863 14597 4864
rect 27610 4928 27930 4929
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 4863 27930 4864
rect 3141 4586 3207 4589
rect 10041 4586 10107 4589
rect 3141 4584 10107 4586
rect 3141 4528 3146 4584
rect 3202 4528 10046 4584
rect 10102 4528 10107 4584
rect 3141 4526 10107 4528
rect 3141 4523 3207 4526
rect 10041 4523 10107 4526
rect 7610 4384 7930 4385
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7930 4384
rect 7610 4319 7930 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 34277 4384 34597 4385
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 4319 34597 4320
rect 3509 4042 3575 4045
rect 5625 4042 5691 4045
rect 9489 4042 9555 4045
rect 17769 4042 17835 4045
rect 3509 4040 17835 4042
rect 3509 3984 3514 4040
rect 3570 3984 5630 4040
rect 5686 3984 9494 4040
rect 9550 3984 17774 4040
rect 17830 3984 17835 4040
rect 3509 3982 17835 3984
rect 3509 3979 3575 3982
rect 5625 3979 5691 3982
rect 9489 3979 9555 3982
rect 17769 3979 17835 3982
rect 25589 4042 25655 4045
rect 35157 4042 35223 4045
rect 25589 4040 35223 4042
rect 25589 3984 25594 4040
rect 25650 3984 35162 4040
rect 35218 3984 35223 4040
rect 25589 3982 35223 3984
rect 25589 3979 25655 3982
rect 35157 3979 35223 3982
rect 3233 3906 3299 3909
rect 9765 3906 9831 3909
rect 3233 3904 9831 3906
rect 3233 3848 3238 3904
rect 3294 3848 9770 3904
rect 9826 3848 9831 3904
rect 3233 3846 9831 3848
rect 3233 3843 3299 3846
rect 9765 3843 9831 3846
rect 14277 3840 14597 3841
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 3775 14597 3776
rect 27610 3840 27930 3841
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 39520 3816 40000 3936
rect 27610 3775 27930 3776
rect 21357 3770 21423 3773
rect 24301 3770 24367 3773
rect 21357 3768 24367 3770
rect 21357 3712 21362 3768
rect 21418 3712 24306 3768
rect 24362 3712 24367 3768
rect 21357 3710 24367 3712
rect 21357 3707 21423 3710
rect 24301 3707 24367 3710
rect 17125 3498 17191 3501
rect 22093 3498 22159 3501
rect 17125 3496 22159 3498
rect 17125 3440 17130 3496
rect 17186 3440 22098 3496
rect 22154 3440 22159 3496
rect 17125 3438 22159 3440
rect 17125 3435 17191 3438
rect 22093 3435 22159 3438
rect 16297 3362 16363 3365
rect 18965 3362 19031 3365
rect 16297 3360 19031 3362
rect 16297 3304 16302 3360
rect 16358 3304 18970 3360
rect 19026 3304 19031 3360
rect 16297 3302 19031 3304
rect 16297 3299 16363 3302
rect 18965 3299 19031 3302
rect 7610 3296 7930 3297
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7930 3296
rect 7610 3231 7930 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 34277 3296 34597 3297
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 3231 34597 3232
rect 22185 3226 22251 3229
rect 26233 3226 26299 3229
rect 22185 3224 26299 3226
rect 22185 3168 22190 3224
rect 22246 3168 26238 3224
rect 26294 3168 26299 3224
rect 22185 3166 26299 3168
rect 22185 3163 22251 3166
rect 26233 3163 26299 3166
rect 2037 3090 2103 3093
rect 3509 3090 3575 3093
rect 7005 3090 7071 3093
rect 2037 3088 7071 3090
rect 2037 3032 2042 3088
rect 2098 3032 3514 3088
rect 3570 3032 7010 3088
rect 7066 3032 7071 3088
rect 2037 3030 7071 3032
rect 2037 3027 2103 3030
rect 3509 3027 3575 3030
rect 7005 3027 7071 3030
rect 21725 3090 21791 3093
rect 28717 3090 28783 3093
rect 21725 3088 28783 3090
rect 21725 3032 21730 3088
rect 21786 3032 28722 3088
rect 28778 3032 28783 3088
rect 21725 3030 28783 3032
rect 21725 3027 21791 3030
rect 28717 3027 28783 3030
rect 4981 2954 5047 2957
rect 11145 2954 11211 2957
rect 4981 2952 11211 2954
rect 4981 2896 4986 2952
rect 5042 2896 11150 2952
rect 11206 2896 11211 2952
rect 4981 2894 11211 2896
rect 4981 2891 5047 2894
rect 11145 2891 11211 2894
rect 25037 2954 25103 2957
rect 31201 2954 31267 2957
rect 25037 2952 31267 2954
rect 25037 2896 25042 2952
rect 25098 2896 31206 2952
rect 31262 2896 31267 2952
rect 25037 2894 31267 2896
rect 25037 2891 25103 2894
rect 31201 2891 31267 2894
rect 2405 2818 2471 2821
rect 6177 2818 6243 2821
rect 2405 2816 6243 2818
rect 2405 2760 2410 2816
rect 2466 2760 6182 2816
rect 6238 2760 6243 2816
rect 2405 2758 6243 2760
rect 2405 2755 2471 2758
rect 6177 2755 6243 2758
rect 7097 2818 7163 2821
rect 13629 2818 13695 2821
rect 7097 2816 13695 2818
rect 7097 2760 7102 2816
rect 7158 2760 13634 2816
rect 13690 2760 13695 2816
rect 7097 2758 13695 2760
rect 7097 2755 7163 2758
rect 13629 2755 13695 2758
rect 16665 2818 16731 2821
rect 23657 2818 23723 2821
rect 16665 2816 23723 2818
rect 16665 2760 16670 2816
rect 16726 2760 23662 2816
rect 23718 2760 23723 2816
rect 16665 2758 23723 2760
rect 16665 2755 16731 2758
rect 23657 2755 23723 2758
rect 14277 2752 14597 2753
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2687 14597 2688
rect 27610 2752 27930 2753
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2687 27930 2688
rect 7557 2682 7623 2685
rect 12433 2682 12499 2685
rect 7557 2680 12499 2682
rect 7557 2624 7562 2680
rect 7618 2624 12438 2680
rect 12494 2624 12499 2680
rect 7557 2622 12499 2624
rect 7557 2619 7623 2622
rect 12433 2619 12499 2622
rect 11881 2546 11947 2549
rect 16849 2546 16915 2549
rect 11881 2544 16915 2546
rect 11881 2488 11886 2544
rect 11942 2488 16854 2544
rect 16910 2488 16915 2544
rect 11881 2486 16915 2488
rect 11881 2483 11947 2486
rect 16849 2483 16915 2486
rect 25313 2546 25379 2549
rect 36169 2546 36235 2549
rect 25313 2544 36235 2546
rect 25313 2488 25318 2544
rect 25374 2488 36174 2544
rect 36230 2488 36235 2544
rect 25313 2486 36235 2488
rect 25313 2483 25379 2486
rect 36169 2483 36235 2486
rect 9765 2410 9831 2413
rect 16205 2410 16271 2413
rect 9765 2408 16271 2410
rect 9765 2352 9770 2408
rect 9826 2352 16210 2408
rect 16266 2352 16271 2408
rect 9765 2350 16271 2352
rect 9765 2347 9831 2350
rect 16205 2347 16271 2350
rect 21173 2410 21239 2413
rect 26141 2410 26207 2413
rect 21173 2408 26207 2410
rect 21173 2352 21178 2408
rect 21234 2352 26146 2408
rect 26202 2352 26207 2408
rect 21173 2350 26207 2352
rect 21173 2347 21239 2350
rect 26141 2347 26207 2350
rect 27061 2410 27127 2413
rect 38653 2410 38719 2413
rect 27061 2408 38719 2410
rect 27061 2352 27066 2408
rect 27122 2352 38658 2408
rect 38714 2352 38719 2408
rect 27061 2350 38719 2352
rect 27061 2347 27127 2350
rect 38653 2347 38719 2350
rect 16021 2274 16087 2277
rect 20805 2274 20871 2277
rect 16021 2272 20871 2274
rect 16021 2216 16026 2272
rect 16082 2216 20810 2272
rect 20866 2216 20871 2272
rect 16021 2214 20871 2216
rect 16021 2211 16087 2214
rect 20805 2211 20871 2214
rect 24393 2274 24459 2277
rect 33685 2274 33751 2277
rect 24393 2272 33751 2274
rect 24393 2216 24398 2272
rect 24454 2216 33690 2272
rect 33746 2216 33751 2272
rect 24393 2214 33751 2216
rect 24393 2211 24459 2214
rect 33685 2211 33751 2214
rect 7610 2208 7930 2209
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7930 2208
rect 7610 2143 7930 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 34277 2208 34597 2209
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2143 34597 2144
rect 27521 2002 27587 2005
rect 37457 2002 37523 2005
rect 27521 2000 37523 2002
rect 27521 1944 27526 2000
rect 27582 1944 37462 2000
rect 37518 1944 37523 2000
rect 27521 1942 37523 1944
rect 27521 1939 27587 1942
rect 37457 1939 37523 1942
rect 3049 1458 3115 1461
rect 8661 1458 8727 1461
rect 3049 1456 8727 1458
rect 3049 1400 3054 1456
rect 3110 1400 8666 1456
rect 8722 1400 8727 1456
rect 3049 1398 8727 1400
rect 3049 1395 3115 1398
rect 8661 1395 8727 1398
rect 11421 1458 11487 1461
rect 18689 1458 18755 1461
rect 11421 1456 18755 1458
rect 11421 1400 11426 1456
rect 11482 1400 18694 1456
rect 18750 1400 18755 1456
rect 11421 1398 18755 1400
rect 11421 1395 11487 1398
rect 18689 1395 18755 1398
rect 34605 1322 34671 1325
rect 39520 1322 40000 1352
rect 34605 1320 40000 1322
rect 34605 1264 34610 1320
rect 34666 1264 40000 1320
rect 34605 1262 40000 1264
rect 34605 1259 34671 1262
rect 39520 1232 40000 1262
<< via3 >>
rect 14285 13628 14349 13632
rect 14285 13572 14289 13628
rect 14289 13572 14345 13628
rect 14345 13572 14349 13628
rect 14285 13568 14349 13572
rect 14365 13628 14429 13632
rect 14365 13572 14369 13628
rect 14369 13572 14425 13628
rect 14425 13572 14429 13628
rect 14365 13568 14429 13572
rect 14445 13628 14509 13632
rect 14445 13572 14449 13628
rect 14449 13572 14505 13628
rect 14505 13572 14509 13628
rect 14445 13568 14509 13572
rect 14525 13628 14589 13632
rect 14525 13572 14529 13628
rect 14529 13572 14585 13628
rect 14585 13572 14589 13628
rect 14525 13568 14589 13572
rect 27618 13628 27682 13632
rect 27618 13572 27622 13628
rect 27622 13572 27678 13628
rect 27678 13572 27682 13628
rect 27618 13568 27682 13572
rect 27698 13628 27762 13632
rect 27698 13572 27702 13628
rect 27702 13572 27758 13628
rect 27758 13572 27762 13628
rect 27698 13568 27762 13572
rect 27778 13628 27842 13632
rect 27778 13572 27782 13628
rect 27782 13572 27838 13628
rect 27838 13572 27842 13628
rect 27778 13568 27842 13572
rect 27858 13628 27922 13632
rect 27858 13572 27862 13628
rect 27862 13572 27918 13628
rect 27918 13572 27922 13628
rect 27858 13568 27922 13572
rect 7618 13084 7682 13088
rect 7618 13028 7622 13084
rect 7622 13028 7678 13084
rect 7678 13028 7682 13084
rect 7618 13024 7682 13028
rect 7698 13084 7762 13088
rect 7698 13028 7702 13084
rect 7702 13028 7758 13084
rect 7758 13028 7762 13084
rect 7698 13024 7762 13028
rect 7778 13084 7842 13088
rect 7778 13028 7782 13084
rect 7782 13028 7838 13084
rect 7838 13028 7842 13084
rect 7778 13024 7842 13028
rect 7858 13084 7922 13088
rect 7858 13028 7862 13084
rect 7862 13028 7918 13084
rect 7918 13028 7922 13084
rect 7858 13024 7922 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 34285 13084 34349 13088
rect 34285 13028 34289 13084
rect 34289 13028 34345 13084
rect 34345 13028 34349 13084
rect 34285 13024 34349 13028
rect 34365 13084 34429 13088
rect 34365 13028 34369 13084
rect 34369 13028 34425 13084
rect 34425 13028 34429 13084
rect 34365 13024 34429 13028
rect 34445 13084 34509 13088
rect 34445 13028 34449 13084
rect 34449 13028 34505 13084
rect 34505 13028 34509 13084
rect 34445 13024 34509 13028
rect 34525 13084 34589 13088
rect 34525 13028 34529 13084
rect 34529 13028 34585 13084
rect 34585 13028 34589 13084
rect 34525 13024 34589 13028
rect 14285 12540 14349 12544
rect 14285 12484 14289 12540
rect 14289 12484 14345 12540
rect 14345 12484 14349 12540
rect 14285 12480 14349 12484
rect 14365 12540 14429 12544
rect 14365 12484 14369 12540
rect 14369 12484 14425 12540
rect 14425 12484 14429 12540
rect 14365 12480 14429 12484
rect 14445 12540 14509 12544
rect 14445 12484 14449 12540
rect 14449 12484 14505 12540
rect 14505 12484 14509 12540
rect 14445 12480 14509 12484
rect 14525 12540 14589 12544
rect 14525 12484 14529 12540
rect 14529 12484 14585 12540
rect 14585 12484 14589 12540
rect 14525 12480 14589 12484
rect 27618 12540 27682 12544
rect 27618 12484 27622 12540
rect 27622 12484 27678 12540
rect 27678 12484 27682 12540
rect 27618 12480 27682 12484
rect 27698 12540 27762 12544
rect 27698 12484 27702 12540
rect 27702 12484 27758 12540
rect 27758 12484 27762 12540
rect 27698 12480 27762 12484
rect 27778 12540 27842 12544
rect 27778 12484 27782 12540
rect 27782 12484 27838 12540
rect 27838 12484 27842 12540
rect 27778 12480 27842 12484
rect 27858 12540 27922 12544
rect 27858 12484 27862 12540
rect 27862 12484 27918 12540
rect 27918 12484 27922 12540
rect 27858 12480 27922 12484
rect 7618 11996 7682 12000
rect 7618 11940 7622 11996
rect 7622 11940 7678 11996
rect 7678 11940 7682 11996
rect 7618 11936 7682 11940
rect 7698 11996 7762 12000
rect 7698 11940 7702 11996
rect 7702 11940 7758 11996
rect 7758 11940 7762 11996
rect 7698 11936 7762 11940
rect 7778 11996 7842 12000
rect 7778 11940 7782 11996
rect 7782 11940 7838 11996
rect 7838 11940 7842 11996
rect 7778 11936 7842 11940
rect 7858 11996 7922 12000
rect 7858 11940 7862 11996
rect 7862 11940 7918 11996
rect 7918 11940 7922 11996
rect 7858 11936 7922 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 34285 11996 34349 12000
rect 34285 11940 34289 11996
rect 34289 11940 34345 11996
rect 34345 11940 34349 11996
rect 34285 11936 34349 11940
rect 34365 11996 34429 12000
rect 34365 11940 34369 11996
rect 34369 11940 34425 11996
rect 34425 11940 34429 11996
rect 34365 11936 34429 11940
rect 34445 11996 34509 12000
rect 34445 11940 34449 11996
rect 34449 11940 34505 11996
rect 34505 11940 34509 11996
rect 34445 11936 34509 11940
rect 34525 11996 34589 12000
rect 34525 11940 34529 11996
rect 34529 11940 34585 11996
rect 34585 11940 34589 11996
rect 34525 11936 34589 11940
rect 14285 11452 14349 11456
rect 14285 11396 14289 11452
rect 14289 11396 14345 11452
rect 14345 11396 14349 11452
rect 14285 11392 14349 11396
rect 14365 11452 14429 11456
rect 14365 11396 14369 11452
rect 14369 11396 14425 11452
rect 14425 11396 14429 11452
rect 14365 11392 14429 11396
rect 14445 11452 14509 11456
rect 14445 11396 14449 11452
rect 14449 11396 14505 11452
rect 14505 11396 14509 11452
rect 14445 11392 14509 11396
rect 14525 11452 14589 11456
rect 14525 11396 14529 11452
rect 14529 11396 14585 11452
rect 14585 11396 14589 11452
rect 14525 11392 14589 11396
rect 27618 11452 27682 11456
rect 27618 11396 27622 11452
rect 27622 11396 27678 11452
rect 27678 11396 27682 11452
rect 27618 11392 27682 11396
rect 27698 11452 27762 11456
rect 27698 11396 27702 11452
rect 27702 11396 27758 11452
rect 27758 11396 27762 11452
rect 27698 11392 27762 11396
rect 27778 11452 27842 11456
rect 27778 11396 27782 11452
rect 27782 11396 27838 11452
rect 27838 11396 27842 11452
rect 27778 11392 27842 11396
rect 27858 11452 27922 11456
rect 27858 11396 27862 11452
rect 27862 11396 27918 11452
rect 27918 11396 27922 11452
rect 27858 11392 27922 11396
rect 7618 10908 7682 10912
rect 7618 10852 7622 10908
rect 7622 10852 7678 10908
rect 7678 10852 7682 10908
rect 7618 10848 7682 10852
rect 7698 10908 7762 10912
rect 7698 10852 7702 10908
rect 7702 10852 7758 10908
rect 7758 10852 7762 10908
rect 7698 10848 7762 10852
rect 7778 10908 7842 10912
rect 7778 10852 7782 10908
rect 7782 10852 7838 10908
rect 7838 10852 7842 10908
rect 7778 10848 7842 10852
rect 7858 10908 7922 10912
rect 7858 10852 7862 10908
rect 7862 10852 7918 10908
rect 7918 10852 7922 10908
rect 7858 10848 7922 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 34285 10908 34349 10912
rect 34285 10852 34289 10908
rect 34289 10852 34345 10908
rect 34345 10852 34349 10908
rect 34285 10848 34349 10852
rect 34365 10908 34429 10912
rect 34365 10852 34369 10908
rect 34369 10852 34425 10908
rect 34425 10852 34429 10908
rect 34365 10848 34429 10852
rect 34445 10908 34509 10912
rect 34445 10852 34449 10908
rect 34449 10852 34505 10908
rect 34505 10852 34509 10908
rect 34445 10848 34509 10852
rect 34525 10908 34589 10912
rect 34525 10852 34529 10908
rect 34529 10852 34585 10908
rect 34585 10852 34589 10908
rect 34525 10848 34589 10852
rect 14285 10364 14349 10368
rect 14285 10308 14289 10364
rect 14289 10308 14345 10364
rect 14345 10308 14349 10364
rect 14285 10304 14349 10308
rect 14365 10364 14429 10368
rect 14365 10308 14369 10364
rect 14369 10308 14425 10364
rect 14425 10308 14429 10364
rect 14365 10304 14429 10308
rect 14445 10364 14509 10368
rect 14445 10308 14449 10364
rect 14449 10308 14505 10364
rect 14505 10308 14509 10364
rect 14445 10304 14509 10308
rect 14525 10364 14589 10368
rect 14525 10308 14529 10364
rect 14529 10308 14585 10364
rect 14585 10308 14589 10364
rect 14525 10304 14589 10308
rect 27618 10364 27682 10368
rect 27618 10308 27622 10364
rect 27622 10308 27678 10364
rect 27678 10308 27682 10364
rect 27618 10304 27682 10308
rect 27698 10364 27762 10368
rect 27698 10308 27702 10364
rect 27702 10308 27758 10364
rect 27758 10308 27762 10364
rect 27698 10304 27762 10308
rect 27778 10364 27842 10368
rect 27778 10308 27782 10364
rect 27782 10308 27838 10364
rect 27838 10308 27842 10364
rect 27778 10304 27842 10308
rect 27858 10364 27922 10368
rect 27858 10308 27862 10364
rect 27862 10308 27918 10364
rect 27918 10308 27922 10364
rect 27858 10304 27922 10308
rect 7618 9820 7682 9824
rect 7618 9764 7622 9820
rect 7622 9764 7678 9820
rect 7678 9764 7682 9820
rect 7618 9760 7682 9764
rect 7698 9820 7762 9824
rect 7698 9764 7702 9820
rect 7702 9764 7758 9820
rect 7758 9764 7762 9820
rect 7698 9760 7762 9764
rect 7778 9820 7842 9824
rect 7778 9764 7782 9820
rect 7782 9764 7838 9820
rect 7838 9764 7842 9820
rect 7778 9760 7842 9764
rect 7858 9820 7922 9824
rect 7858 9764 7862 9820
rect 7862 9764 7918 9820
rect 7918 9764 7922 9820
rect 7858 9760 7922 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 34285 9820 34349 9824
rect 34285 9764 34289 9820
rect 34289 9764 34345 9820
rect 34345 9764 34349 9820
rect 34285 9760 34349 9764
rect 34365 9820 34429 9824
rect 34365 9764 34369 9820
rect 34369 9764 34425 9820
rect 34425 9764 34429 9820
rect 34365 9760 34429 9764
rect 34445 9820 34509 9824
rect 34445 9764 34449 9820
rect 34449 9764 34505 9820
rect 34505 9764 34509 9820
rect 34445 9760 34509 9764
rect 34525 9820 34589 9824
rect 34525 9764 34529 9820
rect 34529 9764 34585 9820
rect 34585 9764 34589 9820
rect 34525 9760 34589 9764
rect 14285 9276 14349 9280
rect 14285 9220 14289 9276
rect 14289 9220 14345 9276
rect 14345 9220 14349 9276
rect 14285 9216 14349 9220
rect 14365 9276 14429 9280
rect 14365 9220 14369 9276
rect 14369 9220 14425 9276
rect 14425 9220 14429 9276
rect 14365 9216 14429 9220
rect 14445 9276 14509 9280
rect 14445 9220 14449 9276
rect 14449 9220 14505 9276
rect 14505 9220 14509 9276
rect 14445 9216 14509 9220
rect 14525 9276 14589 9280
rect 14525 9220 14529 9276
rect 14529 9220 14585 9276
rect 14585 9220 14589 9276
rect 14525 9216 14589 9220
rect 27618 9276 27682 9280
rect 27618 9220 27622 9276
rect 27622 9220 27678 9276
rect 27678 9220 27682 9276
rect 27618 9216 27682 9220
rect 27698 9276 27762 9280
rect 27698 9220 27702 9276
rect 27702 9220 27758 9276
rect 27758 9220 27762 9276
rect 27698 9216 27762 9220
rect 27778 9276 27842 9280
rect 27778 9220 27782 9276
rect 27782 9220 27838 9276
rect 27838 9220 27842 9276
rect 27778 9216 27842 9220
rect 27858 9276 27922 9280
rect 27858 9220 27862 9276
rect 27862 9220 27918 9276
rect 27918 9220 27922 9276
rect 27858 9216 27922 9220
rect 7618 8732 7682 8736
rect 7618 8676 7622 8732
rect 7622 8676 7678 8732
rect 7678 8676 7682 8732
rect 7618 8672 7682 8676
rect 7698 8732 7762 8736
rect 7698 8676 7702 8732
rect 7702 8676 7758 8732
rect 7758 8676 7762 8732
rect 7698 8672 7762 8676
rect 7778 8732 7842 8736
rect 7778 8676 7782 8732
rect 7782 8676 7838 8732
rect 7838 8676 7842 8732
rect 7778 8672 7842 8676
rect 7858 8732 7922 8736
rect 7858 8676 7862 8732
rect 7862 8676 7918 8732
rect 7918 8676 7922 8732
rect 7858 8672 7922 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 34285 8732 34349 8736
rect 34285 8676 34289 8732
rect 34289 8676 34345 8732
rect 34345 8676 34349 8732
rect 34285 8672 34349 8676
rect 34365 8732 34429 8736
rect 34365 8676 34369 8732
rect 34369 8676 34425 8732
rect 34425 8676 34429 8732
rect 34365 8672 34429 8676
rect 34445 8732 34509 8736
rect 34445 8676 34449 8732
rect 34449 8676 34505 8732
rect 34505 8676 34509 8732
rect 34445 8672 34509 8676
rect 34525 8732 34589 8736
rect 34525 8676 34529 8732
rect 34529 8676 34585 8732
rect 34585 8676 34589 8732
rect 34525 8672 34589 8676
rect 14285 8188 14349 8192
rect 14285 8132 14289 8188
rect 14289 8132 14345 8188
rect 14345 8132 14349 8188
rect 14285 8128 14349 8132
rect 14365 8188 14429 8192
rect 14365 8132 14369 8188
rect 14369 8132 14425 8188
rect 14425 8132 14429 8188
rect 14365 8128 14429 8132
rect 14445 8188 14509 8192
rect 14445 8132 14449 8188
rect 14449 8132 14505 8188
rect 14505 8132 14509 8188
rect 14445 8128 14509 8132
rect 14525 8188 14589 8192
rect 14525 8132 14529 8188
rect 14529 8132 14585 8188
rect 14585 8132 14589 8188
rect 14525 8128 14589 8132
rect 27618 8188 27682 8192
rect 27618 8132 27622 8188
rect 27622 8132 27678 8188
rect 27678 8132 27682 8188
rect 27618 8128 27682 8132
rect 27698 8188 27762 8192
rect 27698 8132 27702 8188
rect 27702 8132 27758 8188
rect 27758 8132 27762 8188
rect 27698 8128 27762 8132
rect 27778 8188 27842 8192
rect 27778 8132 27782 8188
rect 27782 8132 27838 8188
rect 27838 8132 27842 8188
rect 27778 8128 27842 8132
rect 27858 8188 27922 8192
rect 27858 8132 27862 8188
rect 27862 8132 27918 8188
rect 27918 8132 27922 8188
rect 27858 8128 27922 8132
rect 7618 7644 7682 7648
rect 7618 7588 7622 7644
rect 7622 7588 7678 7644
rect 7678 7588 7682 7644
rect 7618 7584 7682 7588
rect 7698 7644 7762 7648
rect 7698 7588 7702 7644
rect 7702 7588 7758 7644
rect 7758 7588 7762 7644
rect 7698 7584 7762 7588
rect 7778 7644 7842 7648
rect 7778 7588 7782 7644
rect 7782 7588 7838 7644
rect 7838 7588 7842 7644
rect 7778 7584 7842 7588
rect 7858 7644 7922 7648
rect 7858 7588 7862 7644
rect 7862 7588 7918 7644
rect 7918 7588 7922 7644
rect 7858 7584 7922 7588
rect 14285 7100 14349 7104
rect 14285 7044 14289 7100
rect 14289 7044 14345 7100
rect 14345 7044 14349 7100
rect 14285 7040 14349 7044
rect 14365 7100 14429 7104
rect 14365 7044 14369 7100
rect 14369 7044 14425 7100
rect 14425 7044 14429 7100
rect 14365 7040 14429 7044
rect 14445 7100 14509 7104
rect 14445 7044 14449 7100
rect 14449 7044 14505 7100
rect 14505 7044 14509 7100
rect 14445 7040 14509 7044
rect 14525 7100 14589 7104
rect 14525 7044 14529 7100
rect 14529 7044 14585 7100
rect 14585 7044 14589 7100
rect 14525 7040 14589 7044
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 34285 7644 34349 7648
rect 34285 7588 34289 7644
rect 34289 7588 34345 7644
rect 34345 7588 34349 7644
rect 34285 7584 34349 7588
rect 34365 7644 34429 7648
rect 34365 7588 34369 7644
rect 34369 7588 34425 7644
rect 34425 7588 34429 7644
rect 34365 7584 34429 7588
rect 34445 7644 34509 7648
rect 34445 7588 34449 7644
rect 34449 7588 34505 7644
rect 34505 7588 34509 7644
rect 34445 7584 34509 7588
rect 34525 7644 34589 7648
rect 34525 7588 34529 7644
rect 34529 7588 34585 7644
rect 34585 7588 34589 7644
rect 34525 7584 34589 7588
rect 27618 7100 27682 7104
rect 27618 7044 27622 7100
rect 27622 7044 27678 7100
rect 27678 7044 27682 7100
rect 27618 7040 27682 7044
rect 27698 7100 27762 7104
rect 27698 7044 27702 7100
rect 27702 7044 27758 7100
rect 27758 7044 27762 7100
rect 27698 7040 27762 7044
rect 27778 7100 27842 7104
rect 27778 7044 27782 7100
rect 27782 7044 27838 7100
rect 27838 7044 27842 7100
rect 27778 7040 27842 7044
rect 27858 7100 27922 7104
rect 27858 7044 27862 7100
rect 27862 7044 27918 7100
rect 27918 7044 27922 7100
rect 27858 7040 27922 7044
rect 7618 6556 7682 6560
rect 7618 6500 7622 6556
rect 7622 6500 7678 6556
rect 7678 6500 7682 6556
rect 7618 6496 7682 6500
rect 7698 6556 7762 6560
rect 7698 6500 7702 6556
rect 7702 6500 7758 6556
rect 7758 6500 7762 6556
rect 7698 6496 7762 6500
rect 7778 6556 7842 6560
rect 7778 6500 7782 6556
rect 7782 6500 7838 6556
rect 7838 6500 7842 6556
rect 7778 6496 7842 6500
rect 7858 6556 7922 6560
rect 7858 6500 7862 6556
rect 7862 6500 7918 6556
rect 7918 6500 7922 6556
rect 7858 6496 7922 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 34285 6556 34349 6560
rect 34285 6500 34289 6556
rect 34289 6500 34345 6556
rect 34345 6500 34349 6556
rect 34285 6496 34349 6500
rect 34365 6556 34429 6560
rect 34365 6500 34369 6556
rect 34369 6500 34425 6556
rect 34425 6500 34429 6556
rect 34365 6496 34429 6500
rect 34445 6556 34509 6560
rect 34445 6500 34449 6556
rect 34449 6500 34505 6556
rect 34505 6500 34509 6556
rect 34445 6496 34509 6500
rect 34525 6556 34589 6560
rect 34525 6500 34529 6556
rect 34529 6500 34585 6556
rect 34585 6500 34589 6556
rect 34525 6496 34589 6500
rect 14285 6012 14349 6016
rect 14285 5956 14289 6012
rect 14289 5956 14345 6012
rect 14345 5956 14349 6012
rect 14285 5952 14349 5956
rect 14365 6012 14429 6016
rect 14365 5956 14369 6012
rect 14369 5956 14425 6012
rect 14425 5956 14429 6012
rect 14365 5952 14429 5956
rect 14445 6012 14509 6016
rect 14445 5956 14449 6012
rect 14449 5956 14505 6012
rect 14505 5956 14509 6012
rect 14445 5952 14509 5956
rect 14525 6012 14589 6016
rect 14525 5956 14529 6012
rect 14529 5956 14585 6012
rect 14585 5956 14589 6012
rect 14525 5952 14589 5956
rect 27618 6012 27682 6016
rect 27618 5956 27622 6012
rect 27622 5956 27678 6012
rect 27678 5956 27682 6012
rect 27618 5952 27682 5956
rect 27698 6012 27762 6016
rect 27698 5956 27702 6012
rect 27702 5956 27758 6012
rect 27758 5956 27762 6012
rect 27698 5952 27762 5956
rect 27778 6012 27842 6016
rect 27778 5956 27782 6012
rect 27782 5956 27838 6012
rect 27838 5956 27842 6012
rect 27778 5952 27842 5956
rect 27858 6012 27922 6016
rect 27858 5956 27862 6012
rect 27862 5956 27918 6012
rect 27918 5956 27922 6012
rect 27858 5952 27922 5956
rect 7618 5468 7682 5472
rect 7618 5412 7622 5468
rect 7622 5412 7678 5468
rect 7678 5412 7682 5468
rect 7618 5408 7682 5412
rect 7698 5468 7762 5472
rect 7698 5412 7702 5468
rect 7702 5412 7758 5468
rect 7758 5412 7762 5468
rect 7698 5408 7762 5412
rect 7778 5468 7842 5472
rect 7778 5412 7782 5468
rect 7782 5412 7838 5468
rect 7838 5412 7842 5468
rect 7778 5408 7842 5412
rect 7858 5468 7922 5472
rect 7858 5412 7862 5468
rect 7862 5412 7918 5468
rect 7918 5412 7922 5468
rect 7858 5408 7922 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 34285 5468 34349 5472
rect 34285 5412 34289 5468
rect 34289 5412 34345 5468
rect 34345 5412 34349 5468
rect 34285 5408 34349 5412
rect 34365 5468 34429 5472
rect 34365 5412 34369 5468
rect 34369 5412 34425 5468
rect 34425 5412 34429 5468
rect 34365 5408 34429 5412
rect 34445 5468 34509 5472
rect 34445 5412 34449 5468
rect 34449 5412 34505 5468
rect 34505 5412 34509 5468
rect 34445 5408 34509 5412
rect 34525 5468 34589 5472
rect 34525 5412 34529 5468
rect 34529 5412 34585 5468
rect 34585 5412 34589 5468
rect 34525 5408 34589 5412
rect 14285 4924 14349 4928
rect 14285 4868 14289 4924
rect 14289 4868 14345 4924
rect 14345 4868 14349 4924
rect 14285 4864 14349 4868
rect 14365 4924 14429 4928
rect 14365 4868 14369 4924
rect 14369 4868 14425 4924
rect 14425 4868 14429 4924
rect 14365 4864 14429 4868
rect 14445 4924 14509 4928
rect 14445 4868 14449 4924
rect 14449 4868 14505 4924
rect 14505 4868 14509 4924
rect 14445 4864 14509 4868
rect 14525 4924 14589 4928
rect 14525 4868 14529 4924
rect 14529 4868 14585 4924
rect 14585 4868 14589 4924
rect 14525 4864 14589 4868
rect 27618 4924 27682 4928
rect 27618 4868 27622 4924
rect 27622 4868 27678 4924
rect 27678 4868 27682 4924
rect 27618 4864 27682 4868
rect 27698 4924 27762 4928
rect 27698 4868 27702 4924
rect 27702 4868 27758 4924
rect 27758 4868 27762 4924
rect 27698 4864 27762 4868
rect 27778 4924 27842 4928
rect 27778 4868 27782 4924
rect 27782 4868 27838 4924
rect 27838 4868 27842 4924
rect 27778 4864 27842 4868
rect 27858 4924 27922 4928
rect 27858 4868 27862 4924
rect 27862 4868 27918 4924
rect 27918 4868 27922 4924
rect 27858 4864 27922 4868
rect 7618 4380 7682 4384
rect 7618 4324 7622 4380
rect 7622 4324 7678 4380
rect 7678 4324 7682 4380
rect 7618 4320 7682 4324
rect 7698 4380 7762 4384
rect 7698 4324 7702 4380
rect 7702 4324 7758 4380
rect 7758 4324 7762 4380
rect 7698 4320 7762 4324
rect 7778 4380 7842 4384
rect 7778 4324 7782 4380
rect 7782 4324 7838 4380
rect 7838 4324 7842 4380
rect 7778 4320 7842 4324
rect 7858 4380 7922 4384
rect 7858 4324 7862 4380
rect 7862 4324 7918 4380
rect 7918 4324 7922 4380
rect 7858 4320 7922 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 34285 4380 34349 4384
rect 34285 4324 34289 4380
rect 34289 4324 34345 4380
rect 34345 4324 34349 4380
rect 34285 4320 34349 4324
rect 34365 4380 34429 4384
rect 34365 4324 34369 4380
rect 34369 4324 34425 4380
rect 34425 4324 34429 4380
rect 34365 4320 34429 4324
rect 34445 4380 34509 4384
rect 34445 4324 34449 4380
rect 34449 4324 34505 4380
rect 34505 4324 34509 4380
rect 34445 4320 34509 4324
rect 34525 4380 34589 4384
rect 34525 4324 34529 4380
rect 34529 4324 34585 4380
rect 34585 4324 34589 4380
rect 34525 4320 34589 4324
rect 14285 3836 14349 3840
rect 14285 3780 14289 3836
rect 14289 3780 14345 3836
rect 14345 3780 14349 3836
rect 14285 3776 14349 3780
rect 14365 3836 14429 3840
rect 14365 3780 14369 3836
rect 14369 3780 14425 3836
rect 14425 3780 14429 3836
rect 14365 3776 14429 3780
rect 14445 3836 14509 3840
rect 14445 3780 14449 3836
rect 14449 3780 14505 3836
rect 14505 3780 14509 3836
rect 14445 3776 14509 3780
rect 14525 3836 14589 3840
rect 14525 3780 14529 3836
rect 14529 3780 14585 3836
rect 14585 3780 14589 3836
rect 14525 3776 14589 3780
rect 27618 3836 27682 3840
rect 27618 3780 27622 3836
rect 27622 3780 27678 3836
rect 27678 3780 27682 3836
rect 27618 3776 27682 3780
rect 27698 3836 27762 3840
rect 27698 3780 27702 3836
rect 27702 3780 27758 3836
rect 27758 3780 27762 3836
rect 27698 3776 27762 3780
rect 27778 3836 27842 3840
rect 27778 3780 27782 3836
rect 27782 3780 27838 3836
rect 27838 3780 27842 3836
rect 27778 3776 27842 3780
rect 27858 3836 27922 3840
rect 27858 3780 27862 3836
rect 27862 3780 27918 3836
rect 27918 3780 27922 3836
rect 27858 3776 27922 3780
rect 7618 3292 7682 3296
rect 7618 3236 7622 3292
rect 7622 3236 7678 3292
rect 7678 3236 7682 3292
rect 7618 3232 7682 3236
rect 7698 3292 7762 3296
rect 7698 3236 7702 3292
rect 7702 3236 7758 3292
rect 7758 3236 7762 3292
rect 7698 3232 7762 3236
rect 7778 3292 7842 3296
rect 7778 3236 7782 3292
rect 7782 3236 7838 3292
rect 7838 3236 7842 3292
rect 7778 3232 7842 3236
rect 7858 3292 7922 3296
rect 7858 3236 7862 3292
rect 7862 3236 7918 3292
rect 7918 3236 7922 3292
rect 7858 3232 7922 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 34285 3292 34349 3296
rect 34285 3236 34289 3292
rect 34289 3236 34345 3292
rect 34345 3236 34349 3292
rect 34285 3232 34349 3236
rect 34365 3292 34429 3296
rect 34365 3236 34369 3292
rect 34369 3236 34425 3292
rect 34425 3236 34429 3292
rect 34365 3232 34429 3236
rect 34445 3292 34509 3296
rect 34445 3236 34449 3292
rect 34449 3236 34505 3292
rect 34505 3236 34509 3292
rect 34445 3232 34509 3236
rect 34525 3292 34589 3296
rect 34525 3236 34529 3292
rect 34529 3236 34585 3292
rect 34585 3236 34589 3292
rect 34525 3232 34589 3236
rect 14285 2748 14349 2752
rect 14285 2692 14289 2748
rect 14289 2692 14345 2748
rect 14345 2692 14349 2748
rect 14285 2688 14349 2692
rect 14365 2748 14429 2752
rect 14365 2692 14369 2748
rect 14369 2692 14425 2748
rect 14425 2692 14429 2748
rect 14365 2688 14429 2692
rect 14445 2748 14509 2752
rect 14445 2692 14449 2748
rect 14449 2692 14505 2748
rect 14505 2692 14509 2748
rect 14445 2688 14509 2692
rect 14525 2748 14589 2752
rect 14525 2692 14529 2748
rect 14529 2692 14585 2748
rect 14585 2692 14589 2748
rect 14525 2688 14589 2692
rect 27618 2748 27682 2752
rect 27618 2692 27622 2748
rect 27622 2692 27678 2748
rect 27678 2692 27682 2748
rect 27618 2688 27682 2692
rect 27698 2748 27762 2752
rect 27698 2692 27702 2748
rect 27702 2692 27758 2748
rect 27758 2692 27762 2748
rect 27698 2688 27762 2692
rect 27778 2748 27842 2752
rect 27778 2692 27782 2748
rect 27782 2692 27838 2748
rect 27838 2692 27842 2748
rect 27778 2688 27842 2692
rect 27858 2748 27922 2752
rect 27858 2692 27862 2748
rect 27862 2692 27918 2748
rect 27918 2692 27922 2748
rect 27858 2688 27922 2692
rect 7618 2204 7682 2208
rect 7618 2148 7622 2204
rect 7622 2148 7678 2204
rect 7678 2148 7682 2204
rect 7618 2144 7682 2148
rect 7698 2204 7762 2208
rect 7698 2148 7702 2204
rect 7702 2148 7758 2204
rect 7758 2148 7762 2204
rect 7698 2144 7762 2148
rect 7778 2204 7842 2208
rect 7778 2148 7782 2204
rect 7782 2148 7838 2204
rect 7838 2148 7842 2204
rect 7778 2144 7842 2148
rect 7858 2204 7922 2208
rect 7858 2148 7862 2204
rect 7862 2148 7918 2204
rect 7918 2148 7922 2204
rect 7858 2144 7922 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
rect 34285 2204 34349 2208
rect 34285 2148 34289 2204
rect 34289 2148 34345 2204
rect 34345 2148 34349 2204
rect 34285 2144 34349 2148
rect 34365 2204 34429 2208
rect 34365 2148 34369 2204
rect 34369 2148 34425 2204
rect 34425 2148 34429 2204
rect 34365 2144 34429 2148
rect 34445 2204 34509 2208
rect 34445 2148 34449 2204
rect 34449 2148 34505 2204
rect 34505 2148 34509 2204
rect 34445 2144 34509 2148
rect 34525 2204 34589 2208
rect 34525 2148 34529 2204
rect 34529 2148 34585 2204
rect 34585 2148 34589 2204
rect 34525 2144 34589 2148
<< metal4 >>
rect 7610 13088 7931 13648
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7931 13088
rect 7610 12000 7931 13024
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7931 12000
rect 7610 10912 7931 11936
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7931 10912
rect 7610 9824 7931 10848
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7931 9824
rect 7610 8736 7931 9760
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7931 8736
rect 7610 7648 7931 8672
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7931 7648
rect 7610 6560 7931 7584
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7931 6560
rect 7610 5472 7931 6496
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7931 5472
rect 7610 4384 7931 5408
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7931 4384
rect 7610 3296 7931 4320
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7931 3296
rect 7610 2208 7931 3232
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7931 2208
rect 7610 2128 7931 2144
rect 14277 13632 14597 13648
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 12544 14597 13568
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 11456 14597 12480
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 10368 14597 11392
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 9280 14597 10304
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 8192 14597 9216
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 7104 14597 8128
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 6016 14597 7040
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 4928 14597 5952
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 3840 14597 4864
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 2752 14597 3776
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2128 14597 2688
rect 20944 13088 21264 13648
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 2208 21264 3232
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
rect 27610 13632 27930 13648
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 12544 27930 13568
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 11456 27930 12480
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 10368 27930 11392
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 9280 27930 10304
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 27610 8192 27930 9216
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 7104 27930 8128
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 6016 27930 7040
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 4928 27930 5952
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 3840 27930 4864
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 2752 27930 3776
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2128 27930 2688
rect 34277 13088 34597 13648
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 12000 34597 13024
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 34277 10912 34597 11936
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 9824 34597 10848
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 8736 34597 9760
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 7648 34597 8672
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 6560 34597 7584
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 5472 34597 6496
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 4384 34597 5408
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 3296 34597 4320
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 2208 34597 3232
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2128 34597 2144
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 774 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_15 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_11
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_11
timestamp 1586364061
transform 1 0 2116 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2668 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 2300 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _20_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_42 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__20__A
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_19 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_31
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_36 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4416 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_39
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_43
timestamp 1586364061
transform 1 0 5060 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _21_
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_43
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_55
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__21__A
timestamp 1586364061
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_59
timestamp 1586364061
transform 1 0 6532 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_67
timestamp 1586364061
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_71
timestamp 1586364061
transform 1 0 7636 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_1_55 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_83
timestamp 1586364061
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_44
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_102
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _22_
timestamp 1586364061
transform 1 0 11224 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_45
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_56
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__22__A
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_114
timestamp 1586364061
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_46
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_160
timestamp 1586364061
transform 1 0 15824 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 774 592
use scs8hd_buf_2  _23_
timestamp 1586364061
transform 1 0 16468 0 1 2720
box -38 -48 406 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 16100 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__23__A
timestamp 1586364061
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_171
timestamp 1586364061
transform 1 0 16836 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_47
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_57
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_183
timestamp 1586364061
transform 1 0 17940 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _16_
timestamp 1586364061
transform 1 0 21528 0 1 2720
box -38 -48 406 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_48
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__16__A
timestamp 1586364061
transform 1 0 22080 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_226
timestamp 1586364061
transform 1 0 21896 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_226
timestamp 1586364061
transform 1 0 21896 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_230
timestamp 1586364061
transform 1 0 22264 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_49
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_58
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 24012 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_238
timestamp 1586364061
transform 1 0 23000 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_246
timestamp 1586364061
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_242
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_255
timestamp 1586364061
transform 1 0 24564 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_251
timestamp 1586364061
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_255
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__17__A
timestamp 1586364061
transform 1 0 24748 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _17_
timestamp 1586364061
transform 1 0 24196 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_259
timestamp 1586364061
transform 1 0 24932 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 25300 0 -1 2720
box -38 -48 774 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 25024 0 1 2720
box -38 -48 774 592
use scs8hd_buf_2  _18_
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_50
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_271
timestamp 1586364061
transform 1 0 26036 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_275
timestamp 1586364061
transform 1 0 26404 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_284
timestamp 1586364061
transform 1 0 27232 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_268
timestamp 1586364061
transform 1 0 25760 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_280
timestamp 1586364061
transform 1 0 26864 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__18__A
timestamp 1586364061
transform 1 0 27416 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_288
timestamp 1586364061
transform 1 0 27600 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_0_300
timestamp 1586364061
transform 1 0 28704 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_292
timestamp 1586364061
transform 1 0 27968 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_51
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_59
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_308
timestamp 1586364061
transform 1 0 29440 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_311
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_304
timestamp 1586364061
transform 1 0 29072 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_306
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_318
timestamp 1586364061
transform 1 0 30360 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_323
timestamp 1586364061
transform 1 0 30820 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_335
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_330
timestamp 1586364061
transform 1 0 31464 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_52
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_342
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_354
timestamp 1586364061
transform 1 0 33672 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_342
timestamp 1586364061
transform 1 0 32568 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_354
timestamp 1586364061
transform 1 0 33672 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_53
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_60
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_366
timestamp 1586364061
transform 1 0 34776 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_373
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_367
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_385
timestamp 1586364061
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_379
timestamp 1586364061
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_391
timestamp 1586364061
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_54
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_397
timestamp 1586364061
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_3  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_403
timestamp 1586364061
transform 1 0 38180 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _19_
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__19__A
timestamp 1586364061
transform 1 0 1932 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_7
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_11
timestamp 1586364061
transform 1 0 2116 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_61
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3128 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_19
timestamp 1586364061
transform 1 0 2852 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_6  FILLER_2_24
timestamp 1586364061
transform 1 0 3312 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_30
timestamp 1586364061
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_86
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_89
timestamp 1586364061
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_62
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_63
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_186
timestamp 1586364061
transform 1 0 18216 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_64
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_198
timestamp 1586364061
transform 1 0 19320 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_210
timestamp 1586364061
transform 1 0 20424 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24012 0 -1 3808
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_2_247
timestamp 1586364061
transform 1 0 23828 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 25208 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_260
timestamp 1586364061
transform 1 0 25024 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_264
timestamp 1586364061
transform 1 0 25392 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_272
timestamp 1586364061
transform 1 0 26128 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_288
timestamp 1586364061
transform 1 0 27600 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_300
timestamp 1586364061
transform 1 0 28704 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_312
timestamp 1586364061
transform 1 0 29808 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_324
timestamp 1586364061
transform 1 0 30912 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_337
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_349
timestamp 1586364061
transform 1 0 33212 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_361
timestamp 1586364061
transform 1 0 34316 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_373
timestamp 1586364061
transform 1 0 35420 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_385
timestamp 1586364061
transform 1 0 36524 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_406
timestamp 1586364061
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3128 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2944 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_33
timestamp 1586364061
transform 1 0 4140 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5520 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_45
timestamp 1586364061
transform 1 0 5244 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_50
timestamp 1586364061
transform 1 0 5704 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_3_54
timestamp 1586364061
transform 1 0 6072 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_60
timestamp 1586364061
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9108 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8924 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_3_82
timestamp 1586364061
transform 1 0 8648 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_195
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20792 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20424 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_207
timestamp 1586364061
transform 1 0 20148 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_212
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20976 0 1 3808
box -38 -48 1050 592
use scs8hd_decap_12  FILLER_3_227
timestamp 1586364061
transform 1 0 21988 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_239
timestamp 1586364061
transform 1 0 23092 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_243
timestamp 1586364061
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_273
timestamp 1586364061
transform 1 0 26220 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_285
timestamp 1586364061
transform 1 0 27324 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_297
timestamp 1586364061
transform 1 0 28428 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_306
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_318
timestamp 1586364061
transform 1 0 30360 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_330
timestamp 1586364061
transform 1 0 31464 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_342
timestamp 1586364061
transform 1 0 32568 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_354
timestamp 1586364061
transform 1 0 33672 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_367
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_379
timestamp 1586364061
transform 1 0 35972 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_391
timestamp 1586364061
transform 1 0 37076 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_403
timestamp 1586364061
transform 1 0 38180 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3036 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5520 0 -1 4896
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_59
timestamp 1586364061
transform 1 0 6532 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_71
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_83
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_91
timestamp 1586364061
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25208 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_259
timestamp 1586364061
transform 1 0 24932 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_264
timestamp 1586364061
transform 1 0 25392 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_272
timestamp 1586364061
transform 1 0 26128 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_288
timestamp 1586364061
transform 1 0 27600 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_300
timestamp 1586364061
transform 1 0 28704 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_312
timestamp 1586364061
transform 1 0 29808 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_324
timestamp 1586364061
transform 1 0 30912 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_337
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_349
timestamp 1586364061
transform 1 0 33212 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_361
timestamp 1586364061
transform 1 0 34316 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_373
timestamp 1586364061
transform 1 0 35420 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_385
timestamp 1586364061
transform 1 0 36524 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_406
timestamp 1586364061
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3036 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_32
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_44
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_56
timestamp 1586364061
transform 1 0 6256 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_60
timestamp 1586364061
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_281
timestamp 1586364061
transform 1 0 26956 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_293
timestamp 1586364061
transform 1 0 28060 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_306
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_318
timestamp 1586364061
transform 1 0 30360 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_330
timestamp 1586364061
transform 1 0 31464 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_342
timestamp 1586364061
transform 1 0 32568 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_354
timestamp 1586364061
transform 1 0 33672 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_367
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_379
timestamp 1586364061
transform 1 0 35972 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_391
timestamp 1586364061
transform 1 0 37076 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_5_403
timestamp 1586364061
transform 1 0 38180 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__15__B
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_91
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__15__D
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__15__A
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_103
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_99
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__12__B
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__15__C
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_107
timestamp 1586364061
transform 1 0 10948 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_119
timestamp 1586364061
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__09__D
timestamp 1586364061
transform 1 0 20516 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_213
timestamp 1586364061
transform 1 0 20700 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_221
timestamp 1586364061
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_217
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__C
timestamp 1586364061
transform 1 0 21252 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__A
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_231
timestamp 1586364061
transform 1 0 22356 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_225
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__07__C
timestamp 1586364061
transform 1 0 22172 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__B
timestamp 1586364061
transform 1 0 21620 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_239
timestamp 1586364061
transform 1 0 23092 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_235
timestamp 1586364061
transform 1 0 22724 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__07__D
timestamp 1586364061
transform 1 0 22908 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__07__B
timestamp 1586364061
transform 1 0 22540 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_249
timestamp 1586364061
transform 1 0 24012 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_243
timestamp 1586364061
transform 1 0 23460 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__07__A
timestamp 1586364061
transform 1 0 23276 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_and4_4  _05_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24288 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__05__C
timestamp 1586364061
transform 1 0 24104 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__05__B
timestamp 1586364061
transform 1 0 24288 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__05__A
timestamp 1586364061
transform 1 0 24656 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_254
timestamp 1586364061
transform 1 0 24472 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_258
timestamp 1586364061
transform 1 0 24840 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_261
timestamp 1586364061
transform 1 0 25116 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_270
timestamp 1586364061
transform 1 0 25944 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_274
timestamp 1586364061
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_273
timestamp 1586364061
transform 1 0 26220 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_285
timestamp 1586364061
transform 1 0 27324 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_288
timestamp 1586364061
transform 1 0 27600 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_300
timestamp 1586364061
transform 1 0 28704 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_297
timestamp 1586364061
transform 1 0 28428 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_312
timestamp 1586364061
transform 1 0 29808 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_306
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_318
timestamp 1586364061
transform 1 0 30360 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_324
timestamp 1586364061
transform 1 0 30912 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_337
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_330
timestamp 1586364061
transform 1 0 31464 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_349
timestamp 1586364061
transform 1 0 33212 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_342
timestamp 1586364061
transform 1 0 32568 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_354
timestamp 1586364061
transform 1 0 33672 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_361
timestamp 1586364061
transform 1 0 34316 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_373
timestamp 1586364061
transform 1 0 35420 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_367
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_385
timestamp 1586364061
transform 1 0 36524 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_379
timestamp 1586364061
transform 1 0 35972 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_391
timestamp 1586364061
transform 1 0 37076 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_398
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_406
timestamp 1586364061
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_403
timestamp 1586364061
transform 1 0 38180 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use scs8hd_nor4_4  _15_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_110
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_122
timestamp 1586364061
transform 1 0 12328 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_134
timestamp 1586364061
transform 1 0 13432 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_8_146
timestamp 1586364061
transform 1 0 14536 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_152
timestamp 1586364061
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__10__B
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_204
timestamp 1586364061
transform 1 0 19872 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_212
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_and4_4  _09_
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_224
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 774 592
use scs8hd_and4_4  _07_
timestamp 1586364061
transform 1 0 22540 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_1  FILLER_8_232
timestamp 1586364061
transform 1 0 22448 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_242
timestamp 1586364061
transform 1 0 23368 0 -1 7072
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__05__D
timestamp 1586364061
transform 1 0 24288 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_250
timestamp 1586364061
transform 1 0 24104 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_254
timestamp 1586364061
transform 1 0 24472 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_266
timestamp 1586364061
transform 1 0 25576 0 -1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_274
timestamp 1586364061
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_288
timestamp 1586364061
transform 1 0 27600 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_300
timestamp 1586364061
transform 1 0 28704 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_312
timestamp 1586364061
transform 1 0 29808 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_324
timestamp 1586364061
transform 1 0 30912 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_337
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_349
timestamp 1586364061
transform 1 0 33212 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_361
timestamp 1586364061
transform 1 0 34316 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_373
timestamp 1586364061
transform 1 0 35420 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_385
timestamp 1586364061
transform 1 0 36524 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_406
timestamp 1586364061
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__13__A
timestamp 1586364061
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__13__C
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__13__D
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_80
timestamp 1586364061
transform 1 0 8464 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_83
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_87
timestamp 1586364061
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _13_
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__12__C
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__12__A
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__12__D
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_108
timestamp 1586364061
transform 1 0 11040 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_112
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_116
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_120
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__10__D
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_and4_4  _10_
timestamp 1586364061
transform 1 0 19688 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__10__C
timestamp 1586364061
transform 1 0 19504 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_198
timestamp 1586364061
transform 1 0 19320 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_211
timestamp 1586364061
transform 1 0 20516 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_223
timestamp 1586364061
transform 1 0 21620 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_9_235
timestamp 1586364061
transform 1 0 22724 0 1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_9_243
timestamp 1586364061
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_281
timestamp 1586364061
transform 1 0 26956 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_293
timestamp 1586364061
transform 1 0 28060 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_306
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_318
timestamp 1586364061
transform 1 0 30360 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_330
timestamp 1586364061
transform 1 0 31464 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_342
timestamp 1586364061
transform 1 0 32568 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_354
timestamp 1586364061
transform 1 0 33672 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_367
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_379
timestamp 1586364061
transform 1 0 35972 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_391
timestamp 1586364061
transform 1 0 37076 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_9_403
timestamp 1586364061
transform 1 0 38180 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use scs8hd_nor4_4  _12_
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__14__C
timestamp 1586364061
transform 1 0 9936 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__13__B
timestamp 1586364061
transform 1 0 10304 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_98
timestamp 1586364061
transform 1 0 10120 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_119
timestamp 1586364061
transform 1 0 12052 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_131
timestamp 1586364061
transform 1 0 13156 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_143
timestamp 1586364061
transform 1 0 14260 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_151
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__10__A
timestamp 1586364061
transform 1 0 19688 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_204
timestamp 1586364061
transform 1 0 19872 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_212
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_288
timestamp 1586364061
transform 1 0 27600 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_300
timestamp 1586364061
transform 1 0 28704 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_312
timestamp 1586364061
transform 1 0 29808 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_324
timestamp 1586364061
transform 1 0 30912 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_337
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_349
timestamp 1586364061
transform 1 0 33212 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_361
timestamp 1586364061
transform 1 0 34316 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_373
timestamp 1586364061
transform 1 0 35420 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_385
timestamp 1586364061
transform 1 0 36524 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_398
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_406
timestamp 1586364061
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 406 592
use scs8hd_nor4_4  _14_
timestamp 1586364061
transform 1 0 9936 0 1 8160
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__14__D
timestamp 1586364061
transform 1 0 9752 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__14__B
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_92
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_11_113
timestamp 1586364061
transform 1 0 11500 0 1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_11_121
timestamp 1586364061
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__11__A
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_165
timestamp 1586364061
transform 1 0 16284 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_168
timestamp 1586364061
transform 1 0 16560 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_11_180
timestamp 1586364061
transform 1 0 17664 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use scs8hd_buf_1  _04_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__06__A
timestamp 1586364061
transform 1 0 22908 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__04__A
timestamp 1586364061
transform 1 0 23276 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_235
timestamp 1586364061
transform 1 0 22724 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_239
timestamp 1586364061
transform 1 0 23092 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_243
timestamp 1586364061
transform 1 0 23460 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_281
timestamp 1586364061
transform 1 0 26956 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_293
timestamp 1586364061
transform 1 0 28060 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_306
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_318
timestamp 1586364061
transform 1 0 30360 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_330
timestamp 1586364061
transform 1 0 31464 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_342
timestamp 1586364061
transform 1 0 32568 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_354
timestamp 1586364061
transform 1 0 33672 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_367
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_379
timestamp 1586364061
transform 1 0 35972 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_391
timestamp 1586364061
transform 1 0 37076 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_11_403
timestamp 1586364061
transform 1 0 38180 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__14__A
timestamp 1586364061
transform 1 0 9936 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_98
timestamp 1586364061
transform 1 0 10120 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_110
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_122
timestamp 1586364061
transform 1 0 12328 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_134
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_12_146
timestamp 1586364061
transform 1 0 14536 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_152
timestamp 1586364061
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_inv_8  _11_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_12  FILLER_12_175
timestamp 1586364061
transform 1 0 17204 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_187
timestamp 1586364061
transform 1 0 18308 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_199
timestamp 1586364061
transform 1 0 19412 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_12_211
timestamp 1586364061
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_8  _06_
timestamp 1586364061
transform 1 0 22356 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_240
timestamp 1586364061
transform 1 0 23184 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_252
timestamp 1586364061
transform 1 0 24288 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_264
timestamp 1586364061
transform 1 0 25392 0 -1 9248
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_272
timestamp 1586364061
transform 1 0 26128 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_288
timestamp 1586364061
transform 1 0 27600 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_300
timestamp 1586364061
transform 1 0 28704 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_312
timestamp 1586364061
transform 1 0 29808 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_324
timestamp 1586364061
transform 1 0 30912 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_337
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_349
timestamp 1586364061
transform 1 0 33212 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_361
timestamp 1586364061
transform 1 0 34316 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_373
timestamp 1586364061
transform 1 0 35420 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_385
timestamp 1586364061
transform 1 0 36524 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_398
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_406
timestamp 1586364061
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_8  _08_
timestamp 1586364061
transform 1 0 20332 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__08__A
timestamp 1586364061
transform 1 0 20148 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_204
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_218
timestamp 1586364061
transform 1 0 21160 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_230
timestamp 1586364061
transform 1 0 22264 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_242
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_281
timestamp 1586364061
transform 1 0 26956 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_293
timestamp 1586364061
transform 1 0 28060 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_288
timestamp 1586364061
transform 1 0 27600 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_300
timestamp 1586364061
transform 1 0 28704 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_306
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_318
timestamp 1586364061
transform 1 0 30360 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_312
timestamp 1586364061
transform 1 0 29808 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_330
timestamp 1586364061
transform 1 0 31464 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_324
timestamp 1586364061
transform 1 0 30912 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_337
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_342
timestamp 1586364061
transform 1 0 32568 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_354
timestamp 1586364061
transform 1 0 33672 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_349
timestamp 1586364061
transform 1 0 33212 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_367
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_361
timestamp 1586364061
transform 1 0 34316 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_373
timestamp 1586364061
transform 1 0 35420 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_379
timestamp 1586364061
transform 1 0 35972 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_391
timestamp 1586364061
transform 1 0 37076 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_385
timestamp 1586364061
transform 1 0 36524 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_403
timestamp 1586364061
transform 1 0 38180 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_398
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_406
timestamp 1586364061
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_281
timestamp 1586364061
transform 1 0 26956 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_293
timestamp 1586364061
transform 1 0 28060 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_306
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_318
timestamp 1586364061
transform 1 0 30360 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_330
timestamp 1586364061
transform 1 0 31464 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_342
timestamp 1586364061
transform 1 0 32568 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_354
timestamp 1586364061
transform 1 0 33672 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_367
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_379
timestamp 1586364061
transform 1 0 35972 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_391
timestamp 1586364061
transform 1 0 37076 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_403
timestamp 1586364061
transform 1 0 38180 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_178
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_288
timestamp 1586364061
transform 1 0 27600 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_300
timestamp 1586364061
transform 1 0 28704 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_312
timestamp 1586364061
transform 1 0 29808 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_324
timestamp 1586364061
transform 1 0 30912 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_337
timestamp 1586364061
transform 1 0 32108 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_349
timestamp 1586364061
transform 1 0 33212 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_361
timestamp 1586364061
transform 1 0 34316 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_373
timestamp 1586364061
transform 1 0 35420 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_385
timestamp 1586364061
transform 1 0 36524 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_398
timestamp 1586364061
transform 1 0 37720 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_406
timestamp 1586364061
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_281
timestamp 1586364061
transform 1 0 26956 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_293
timestamp 1586364061
transform 1 0 28060 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_306
timestamp 1586364061
transform 1 0 29256 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_318
timestamp 1586364061
transform 1 0 30360 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_330
timestamp 1586364061
transform 1 0 31464 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_342
timestamp 1586364061
transform 1 0 32568 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_354
timestamp 1586364061
transform 1 0 33672 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_367
timestamp 1586364061
transform 1 0 34868 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_379
timestamp 1586364061
transform 1 0 35972 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_391
timestamp 1586364061
transform 1 0 37076 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_403
timestamp 1586364061
transform 1 0 38180 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_288
timestamp 1586364061
transform 1 0 27600 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_300
timestamp 1586364061
transform 1 0 28704 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_312
timestamp 1586364061
transform 1 0 29808 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_324
timestamp 1586364061
transform 1 0 30912 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_337
timestamp 1586364061
transform 1 0 32108 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_349
timestamp 1586364061
transform 1 0 33212 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_361
timestamp 1586364061
transform 1 0 34316 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_373
timestamp 1586364061
transform 1 0 35420 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_385
timestamp 1586364061
transform 1 0 36524 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_398
timestamp 1586364061
transform 1 0 37720 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_406
timestamp 1586364061
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_63
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_75
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_94
timestamp 1586364061
transform 1 0 9752 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_118
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15364 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_156
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_230
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_242
timestamp 1586364061
transform 1 0 23368 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_249
timestamp 1586364061
transform 1 0 24012 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_261
timestamp 1586364061
transform 1 0 25116 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 26772 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_281
timestamp 1586364061
transform 1 0 26956 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_273
timestamp 1586364061
transform 1 0 26220 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_280
timestamp 1586364061
transform 1 0 26864 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_293
timestamp 1586364061
transform 1 0 28060 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_292
timestamp 1586364061
transform 1 0 27968 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 29624 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_306
timestamp 1586364061
transform 1 0 29256 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_318
timestamp 1586364061
transform 1 0 30360 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_304
timestamp 1586364061
transform 1 0 29072 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_311
timestamp 1586364061
transform 1 0 29716 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_330
timestamp 1586364061
transform 1 0 31464 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_323
timestamp 1586364061
transform 1 0 30820 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_335
timestamp 1586364061
transform 1 0 31924 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 32476 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_342
timestamp 1586364061
transform 1 0 32568 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_354
timestamp 1586364061
transform 1 0 33672 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_342
timestamp 1586364061
transform 1 0 32568 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_354
timestamp 1586364061
transform 1 0 33672 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 35328 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_367
timestamp 1586364061
transform 1 0 34868 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_366
timestamp 1586364061
transform 1 0 34776 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_373
timestamp 1586364061
transform 1 0 35420 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_379
timestamp 1586364061
transform 1 0 35972 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_391
timestamp 1586364061
transform 1 0 37076 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_385
timestamp 1586364061
transform 1 0 36524 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 38180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_403
timestamp 1586364061
transform 1 0 38180 0 1 12512
box -38 -48 406 592
use scs8hd_decap_6  FILLER_20_397
timestamp 1586364061
transform 1 0 37628 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  FILLER_20_404
timestamp 1586364061
transform 1 0 38272 0 -1 13600
box -38 -48 314 592
<< labels >>
rlabel metal3 s 39520 3816 40000 3936 6 address[0]
port 0 nsew default input
rlabel metal3 s 39520 6536 40000 6656 6 address[1]
port 1 nsew default input
rlabel metal3 s 39520 9256 40000 9376 6 address[2]
port 2 nsew default input
rlabel metal3 s 39520 11840 40000 11960 6 address[3]
port 3 nsew default input
rlabel metal2 s 1214 0 1270 480 6 bottom_width_0_height_0__pin_0_
port 4 nsew default input
rlabel metal2 s 26146 0 26202 480 6 bottom_width_0_height_0__pin_10_
port 5 nsew default input
rlabel metal2 s 28722 0 28778 480 6 bottom_width_0_height_0__pin_11_
port 6 nsew default tristate
rlabel metal2 s 31206 0 31262 480 6 bottom_width_0_height_0__pin_12_
port 7 nsew default input
rlabel metal2 s 33690 0 33746 480 6 bottom_width_0_height_0__pin_13_
port 8 nsew default tristate
rlabel metal2 s 36174 0 36230 480 6 bottom_width_0_height_0__pin_14_
port 9 nsew default input
rlabel metal2 s 38658 0 38714 480 6 bottom_width_0_height_0__pin_15_
port 10 nsew default tristate
rlabel metal2 s 3698 0 3754 480 6 bottom_width_0_height_0__pin_1_
port 11 nsew default tristate
rlabel metal2 s 6182 0 6238 480 6 bottom_width_0_height_0__pin_2_
port 12 nsew default input
rlabel metal2 s 8666 0 8722 480 6 bottom_width_0_height_0__pin_3_
port 13 nsew default tristate
rlabel metal2 s 11150 0 11206 480 6 bottom_width_0_height_0__pin_4_
port 14 nsew default input
rlabel metal2 s 13634 0 13690 480 6 bottom_width_0_height_0__pin_5_
port 15 nsew default tristate
rlabel metal2 s 16210 0 16266 480 6 bottom_width_0_height_0__pin_6_
port 16 nsew default input
rlabel metal2 s 18694 0 18750 480 6 bottom_width_0_height_0__pin_7_
port 17 nsew default tristate
rlabel metal2 s 21178 0 21234 480 6 bottom_width_0_height_0__pin_8_
port 18 nsew default input
rlabel metal2 s 23662 0 23718 480 6 bottom_width_0_height_0__pin_9_
port 19 nsew default tristate
rlabel metal3 s 39520 14560 40000 14680 6 data_in
port 20 nsew default input
rlabel metal3 s 39520 1232 40000 1352 6 enable
port 21 nsew default input
rlabel metal2 s 2502 15520 2558 16000 6 gfpga_pad_GPIO_PAD[0]
port 22 nsew default bidirectional
rlabel metal2 s 7470 15520 7526 16000 6 gfpga_pad_GPIO_PAD[1]
port 23 nsew default bidirectional
rlabel metal2 s 12438 15520 12494 16000 6 gfpga_pad_GPIO_PAD[2]
port 24 nsew default bidirectional
rlabel metal2 s 17498 15520 17554 16000 6 gfpga_pad_GPIO_PAD[3]
port 25 nsew default bidirectional
rlabel metal2 s 22466 15520 22522 16000 6 gfpga_pad_GPIO_PAD[4]
port 26 nsew default bidirectional
rlabel metal2 s 27434 15520 27490 16000 6 gfpga_pad_GPIO_PAD[5]
port 27 nsew default bidirectional
rlabel metal2 s 32494 15520 32550 16000 6 gfpga_pad_GPIO_PAD[6]
port 28 nsew default bidirectional
rlabel metal2 s 37462 15520 37518 16000 6 gfpga_pad_GPIO_PAD[7]
port 29 nsew default bidirectional
rlabel metal4 s 7611 2128 7931 13648 6 vpwr
port 30 nsew default input
rlabel metal4 s 14277 2128 14597 13648 6 vgnd
port 31 nsew default input
<< end >>
