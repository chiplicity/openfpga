magic
tech EFS8A
magscale 1 2
timestamp 1604399598
<< locali >>
rect 12449 19295 12483 19329
rect 12391 19261 12483 19295
rect 14565 13855 14599 13957
rect 13645 12087 13679 12393
rect 12449 11543 12483 11713
rect 3985 8279 4019 8381
rect 2605 7191 2639 7497
rect 8401 7259 8435 7429
<< viali >>
rect 1409 25313 1443 25347
rect 2513 25313 2547 25347
rect 1593 25177 1627 25211
rect 2053 25109 2087 25143
rect 2329 25109 2363 25143
rect 2697 25109 2731 25143
rect 3065 25109 3099 25143
rect 2421 24905 2455 24939
rect 2053 24769 2087 24803
rect 3249 24769 3283 24803
rect 1409 24701 1443 24735
rect 3065 24701 3099 24735
rect 3617 24701 3651 24735
rect 15945 24701 15979 24735
rect 16497 24701 16531 24735
rect 2973 24633 3007 24667
rect 1593 24565 1627 24599
rect 2605 24565 2639 24599
rect 7481 24565 7515 24599
rect 16129 24565 16163 24599
rect 1961 24361 1995 24395
rect 2881 24361 2915 24395
rect 6377 24361 6411 24395
rect 7849 24361 7883 24395
rect 14289 24361 14323 24395
rect 15485 24361 15519 24395
rect 16681 24361 16715 24395
rect 18889 24361 18923 24395
rect 21097 24361 21131 24395
rect 6285 24293 6319 24327
rect 1409 24225 1443 24259
rect 2789 24225 2823 24259
rect 4445 24225 4479 24259
rect 12081 24225 12115 24259
rect 14105 24225 14139 24259
rect 15301 24225 15335 24259
rect 16497 24225 16531 24259
rect 17601 24225 17635 24259
rect 18705 24225 18739 24259
rect 20913 24225 20947 24259
rect 3065 24157 3099 24191
rect 4537 24157 4571 24191
rect 4721 24157 4755 24191
rect 6561 24157 6595 24191
rect 7941 24157 7975 24191
rect 8125 24157 8159 24191
rect 2421 24089 2455 24123
rect 3801 24089 3835 24123
rect 5917 24089 5951 24123
rect 12265 24089 12299 24123
rect 17785 24089 17819 24123
rect 2237 24021 2271 24055
rect 3433 24021 3467 24055
rect 4077 24021 4111 24055
rect 5273 24021 5307 24055
rect 6929 24021 6963 24055
rect 7389 24021 7423 24055
rect 7481 24021 7515 24055
rect 2053 23817 2087 23851
rect 2145 23817 2179 23851
rect 3157 23817 3191 23851
rect 3617 23817 3651 23851
rect 5457 23817 5491 23851
rect 6009 23817 6043 23851
rect 6377 23817 6411 23851
rect 9137 23817 9171 23851
rect 10333 23817 10367 23851
rect 12633 23817 12667 23851
rect 13093 23817 13127 23851
rect 14473 23817 14507 23851
rect 17049 23817 17083 23851
rect 18245 23817 18279 23851
rect 19625 23817 19659 23851
rect 21373 23817 21407 23851
rect 23857 23817 23891 23851
rect 14013 23749 14047 23783
rect 15117 23749 15151 23783
rect 2697 23681 2731 23715
rect 2513 23613 2547 23647
rect 2605 23613 2639 23647
rect 4077 23613 4111 23647
rect 6837 23613 6871 23647
rect 10149 23613 10183 23647
rect 10701 23613 10735 23647
rect 11253 23613 11287 23647
rect 11805 23613 11839 23647
rect 12449 23613 12483 23647
rect 13829 23613 13863 23647
rect 14933 23613 14967 23647
rect 16865 23613 16899 23647
rect 17785 23613 17819 23647
rect 18061 23613 18095 23647
rect 19441 23613 19475 23647
rect 19993 23613 20027 23647
rect 21189 23613 21223 23647
rect 21741 23613 21775 23647
rect 23673 23613 23707 23647
rect 24225 23613 24259 23647
rect 3985 23545 4019 23579
rect 4344 23545 4378 23579
rect 7104 23545 7138 23579
rect 1685 23477 1719 23511
rect 8217 23477 8251 23511
rect 8769 23477 8803 23511
rect 11437 23477 11471 23511
rect 12173 23477 12207 23511
rect 13645 23477 13679 23511
rect 14749 23477 14783 23511
rect 15485 23477 15519 23511
rect 16589 23477 16623 23511
rect 17509 23477 17543 23511
rect 18613 23477 18647 23511
rect 18981 23477 19015 23511
rect 20913 23477 20947 23511
rect 2145 23273 2179 23307
rect 3157 23273 3191 23307
rect 5273 23273 5307 23307
rect 9873 23273 9907 23307
rect 12725 23273 12759 23307
rect 14105 23273 14139 23307
rect 17233 23273 17267 23307
rect 18337 23273 18371 23307
rect 21097 23273 21131 23307
rect 22385 23273 22419 23307
rect 4353 23205 4387 23239
rect 6644 23205 6678 23239
rect 5181 23137 5215 23171
rect 6009 23137 6043 23171
rect 9689 23137 9723 23171
rect 12541 23137 12575 23171
rect 15301 23137 15335 23171
rect 17049 23137 17083 23171
rect 18153 23137 18187 23171
rect 20913 23137 20947 23171
rect 22201 23137 22235 23171
rect 2237 23069 2271 23103
rect 2421 23069 2455 23103
rect 5457 23069 5491 23103
rect 6377 23069 6411 23103
rect 13553 23069 13587 23103
rect 1685 23001 1719 23035
rect 4721 23001 4755 23035
rect 1777 22933 1811 22967
rect 2881 22933 2915 22967
rect 3801 22933 3835 22967
rect 4813 22933 4847 22967
rect 7757 22933 7791 22967
rect 8493 22933 8527 22967
rect 14473 22933 14507 22967
rect 15485 22933 15519 22967
rect 2053 22729 2087 22763
rect 2605 22729 2639 22763
rect 4905 22729 4939 22763
rect 6193 22729 6227 22763
rect 15761 22729 15795 22763
rect 16865 22729 16899 22763
rect 17141 22729 17175 22763
rect 20913 22729 20947 22763
rect 6837 22661 6871 22695
rect 8401 22661 8435 22695
rect 12909 22661 12943 22695
rect 2697 22593 2731 22627
rect 5641 22593 5675 22627
rect 5825 22593 5859 22627
rect 7481 22593 7515 22627
rect 8953 22593 8987 22627
rect 14565 22593 14599 22627
rect 1409 22525 1443 22559
rect 2964 22525 2998 22559
rect 5549 22525 5583 22559
rect 12173 22525 12207 22559
rect 12725 22525 12759 22559
rect 13277 22525 13311 22559
rect 15577 22525 15611 22559
rect 16129 22525 16163 22559
rect 16681 22525 16715 22559
rect 22201 22525 22235 22559
rect 6561 22457 6595 22491
rect 7297 22457 7331 22491
rect 8861 22457 8895 22491
rect 13921 22457 13955 22491
rect 14381 22457 14415 22491
rect 17601 22457 17635 22491
rect 1593 22389 1627 22423
rect 4077 22389 4111 22423
rect 5181 22389 5215 22423
rect 7205 22389 7239 22423
rect 7849 22389 7883 22423
rect 8217 22389 8251 22423
rect 8769 22389 8803 22423
rect 9781 22389 9815 22423
rect 9965 22389 9999 22423
rect 14013 22389 14047 22423
rect 14473 22389 14507 22423
rect 15393 22389 15427 22423
rect 18245 22389 18279 22423
rect 4077 22185 4111 22219
rect 5641 22185 5675 22219
rect 6285 22185 6319 22219
rect 7941 22185 7975 22219
rect 8493 22185 8527 22219
rect 13829 22185 13863 22219
rect 4445 22117 4479 22151
rect 1409 22049 1443 22083
rect 1676 22049 1710 22083
rect 3893 22049 3927 22083
rect 4537 22049 4571 22083
rect 5273 22049 5307 22083
rect 6745 22049 6779 22083
rect 6837 22049 6871 22083
rect 10885 22049 10919 22083
rect 13737 22049 13771 22083
rect 15557 22049 15591 22083
rect 4629 21981 4663 22015
rect 7021 21981 7055 22015
rect 10977 21981 11011 22015
rect 11161 21981 11195 22015
rect 13921 21981 13955 22015
rect 15301 21981 15335 22015
rect 2789 21913 2823 21947
rect 6377 21913 6411 21947
rect 10517 21913 10551 21947
rect 12541 21913 12575 21947
rect 16681 21913 16715 21947
rect 3525 21845 3559 21879
rect 7389 21845 7423 21879
rect 7757 21845 7791 21879
rect 9045 21845 9079 21879
rect 10333 21845 10367 21879
rect 11529 21845 11563 21879
rect 13277 21845 13311 21879
rect 13369 21845 13403 21879
rect 14473 21845 14507 21879
rect 4721 21641 4755 21675
rect 6469 21641 6503 21675
rect 10609 21641 10643 21675
rect 13553 21641 13587 21675
rect 15577 21641 15611 21675
rect 10241 21573 10275 21607
rect 1685 21505 1719 21539
rect 2145 21505 2179 21539
rect 2237 21505 2271 21539
rect 5457 21505 5491 21539
rect 7665 21505 7699 21539
rect 8033 21505 8067 21539
rect 9505 21505 9539 21539
rect 11437 21505 11471 21539
rect 13001 21505 13035 21539
rect 4445 21437 4479 21471
rect 5273 21437 5307 21471
rect 11253 21437 11287 21471
rect 11805 21437 11839 21471
rect 14197 21437 14231 21471
rect 16129 21437 16163 21471
rect 2482 21369 2516 21403
rect 6101 21369 6135 21403
rect 7389 21369 7423 21403
rect 8401 21369 8435 21403
rect 8861 21369 8895 21403
rect 9413 21369 9447 21403
rect 12265 21369 12299 21403
rect 12817 21369 12851 21403
rect 14464 21369 14498 21403
rect 3617 21301 3651 21335
rect 4905 21301 4939 21335
rect 5365 21301 5399 21335
rect 7021 21301 7055 21335
rect 7481 21301 7515 21335
rect 8953 21301 8987 21335
rect 9321 21301 9355 21335
rect 10793 21301 10827 21335
rect 11161 21301 11195 21335
rect 12449 21301 12483 21335
rect 12909 21301 12943 21335
rect 14105 21301 14139 21335
rect 2329 21097 2363 21131
rect 2421 21097 2455 21131
rect 3525 21097 3559 21131
rect 5733 21097 5767 21131
rect 5917 21097 5951 21131
rect 6285 21097 6319 21131
rect 7481 21097 7515 21131
rect 7849 21097 7883 21131
rect 9045 21097 9079 21131
rect 11621 21097 11655 21131
rect 12725 21097 12759 21131
rect 13553 21097 13587 21131
rect 15577 21097 15611 21131
rect 2881 21029 2915 21063
rect 3801 21029 3835 21063
rect 4813 21029 4847 21063
rect 7389 21029 7423 21063
rect 9934 21029 9968 21063
rect 13461 21029 13495 21063
rect 1409 20961 1443 20995
rect 2789 20961 2823 20995
rect 4721 20961 4755 20995
rect 12165 20961 12199 20995
rect 13093 20961 13127 20995
rect 13921 20961 13955 20995
rect 2973 20893 3007 20927
rect 4905 20893 4939 20927
rect 6377 20893 6411 20927
rect 6469 20893 6503 20927
rect 7941 20893 7975 20927
rect 8125 20893 8159 20927
rect 9689 20893 9723 20927
rect 14013 20893 14047 20927
rect 14197 20893 14231 20927
rect 1961 20825 1995 20859
rect 1593 20757 1627 20791
rect 4353 20757 4387 20791
rect 5365 20757 5399 20791
rect 7021 20757 7055 20791
rect 8493 20757 8527 20791
rect 11069 20757 11103 20791
rect 12357 20757 12391 20791
rect 2145 20553 2179 20587
rect 5549 20553 5583 20587
rect 6285 20553 6319 20587
rect 7205 20553 7239 20587
rect 8769 20553 8803 20587
rect 9321 20553 9355 20587
rect 11253 20553 11287 20587
rect 14381 20553 14415 20587
rect 14749 20553 14783 20587
rect 15209 20553 15243 20587
rect 1409 20349 1443 20383
rect 2513 20349 2547 20383
rect 3341 20349 3375 20383
rect 3433 20349 3467 20383
rect 7389 20349 7423 20383
rect 9873 20349 9907 20383
rect 10129 20349 10163 20383
rect 12449 20349 12483 20383
rect 12716 20349 12750 20383
rect 2881 20281 2915 20315
rect 3678 20281 3712 20315
rect 7656 20281 7690 20315
rect 12265 20281 12299 20315
rect 1593 20213 1627 20247
rect 4813 20213 4847 20247
rect 6009 20213 6043 20247
rect 9781 20213 9815 20247
rect 11897 20213 11931 20247
rect 13829 20213 13863 20247
rect 1961 20009 1995 20043
rect 2421 20009 2455 20043
rect 3525 20009 3559 20043
rect 6009 20009 6043 20043
rect 6929 20009 6963 20043
rect 8585 20009 8619 20043
rect 9321 20009 9355 20043
rect 10333 20009 10367 20043
rect 13553 20009 13587 20043
rect 4344 19941 4378 19975
rect 10784 19941 10818 19975
rect 12541 19941 12575 19975
rect 1409 19873 1443 19907
rect 2513 19873 2547 19907
rect 4084 19873 4118 19907
rect 13461 19873 13495 19907
rect 13921 19873 13955 19907
rect 7021 19805 7055 19839
rect 7113 19805 7147 19839
rect 8125 19805 8159 19839
rect 9965 19805 9999 19839
rect 10517 19805 10551 19839
rect 14013 19805 14047 19839
rect 14105 19805 14139 19839
rect 2697 19737 2731 19771
rect 3065 19737 3099 19771
rect 11897 19737 11931 19771
rect 13093 19737 13127 19771
rect 14565 19737 14599 19771
rect 1593 19669 1627 19703
rect 3801 19669 3835 19703
rect 5457 19669 5491 19703
rect 6561 19669 6595 19703
rect 7757 19669 7791 19703
rect 8401 19669 8435 19703
rect 2329 19465 2363 19499
rect 6193 19465 6227 19499
rect 7021 19465 7055 19499
rect 7665 19465 7699 19499
rect 10609 19465 10643 19499
rect 12633 19465 12667 19499
rect 15577 19465 15611 19499
rect 4445 19329 4479 19363
rect 8309 19329 8343 19363
rect 9873 19329 9907 19363
rect 11437 19329 11471 19363
rect 12449 19329 12483 19363
rect 13185 19329 13219 19363
rect 1409 19261 1443 19295
rect 2513 19261 2547 19295
rect 3709 19261 3743 19295
rect 4169 19261 4203 19295
rect 5365 19261 5399 19295
rect 5825 19261 5859 19295
rect 6653 19261 6687 19295
rect 9597 19261 9631 19295
rect 9689 19261 9723 19295
rect 11161 19261 11195 19295
rect 11253 19261 11287 19295
rect 11897 19261 11931 19295
rect 12265 19261 12299 19295
rect 12357 19261 12391 19295
rect 13001 19261 13035 19295
rect 14105 19261 14139 19295
rect 14197 19261 14231 19295
rect 14464 19261 14498 19295
rect 4905 19193 4939 19227
rect 8125 19193 8159 19227
rect 9137 19193 9171 19227
rect 1593 19125 1627 19159
rect 2053 19125 2087 19159
rect 2697 19125 2731 19159
rect 3157 19125 3191 19159
rect 3801 19125 3835 19159
rect 4261 19125 4295 19159
rect 5181 19125 5215 19159
rect 7573 19125 7607 19159
rect 8033 19125 8067 19159
rect 8677 19125 8711 19159
rect 9229 19125 9263 19159
rect 10793 19125 10827 19159
rect 13093 19125 13127 19159
rect 13737 19125 13771 19159
rect 3893 18921 3927 18955
rect 4537 18921 4571 18955
rect 4997 18921 5031 18955
rect 6101 18921 6135 18955
rect 7205 18921 7239 18955
rect 8125 18921 8159 18955
rect 9045 18921 9079 18955
rect 10793 18921 10827 18955
rect 11253 18921 11287 18955
rect 14105 18921 14139 18955
rect 15301 18921 15335 18955
rect 3525 18853 3559 18887
rect 4353 18853 4387 18887
rect 4905 18853 4939 18887
rect 11713 18853 11747 18887
rect 12173 18853 12207 18887
rect 1409 18785 1443 18819
rect 2513 18785 2547 18819
rect 6469 18785 6503 18819
rect 6561 18785 6595 18819
rect 8033 18785 8067 18819
rect 10057 18785 10091 18819
rect 11161 18785 11195 18819
rect 12992 18785 13026 18819
rect 5089 18717 5123 18751
rect 6653 18717 6687 18751
rect 8217 18717 8251 18751
rect 10149 18717 10183 18751
rect 10333 18717 10367 18751
rect 12725 18717 12759 18751
rect 2421 18649 2455 18683
rect 7481 18649 7515 18683
rect 1593 18581 1627 18615
rect 2053 18581 2087 18615
rect 2697 18581 2731 18615
rect 3157 18581 3191 18615
rect 5641 18581 5675 18615
rect 7665 18581 7699 18615
rect 9413 18581 9447 18615
rect 9689 18581 9723 18615
rect 12541 18581 12575 18615
rect 3801 18377 3835 18411
rect 8401 18377 8435 18411
rect 11437 18377 11471 18411
rect 14013 18377 14047 18411
rect 2697 18309 2731 18343
rect 8953 18309 8987 18343
rect 13461 18309 13495 18343
rect 3249 18241 3283 18275
rect 7021 18241 7055 18275
rect 9413 18241 9447 18275
rect 11897 18241 11931 18275
rect 13001 18241 13035 18275
rect 14565 18241 14599 18275
rect 1409 18173 1443 18207
rect 2237 18173 2271 18207
rect 3157 18173 3191 18207
rect 4169 18173 4203 18207
rect 4261 18173 4295 18207
rect 9505 18173 9539 18207
rect 12817 18173 12851 18207
rect 2605 18105 2639 18139
rect 4506 18105 4540 18139
rect 6193 18105 6227 18139
rect 7288 18105 7322 18139
rect 9750 18105 9784 18139
rect 12265 18105 12299 18139
rect 12909 18105 12943 18139
rect 14473 18105 14507 18139
rect 1593 18037 1627 18071
rect 3065 18037 3099 18071
rect 5641 18037 5675 18071
rect 6653 18037 6687 18071
rect 10885 18037 10919 18071
rect 12449 18037 12483 18071
rect 13921 18037 13955 18071
rect 14381 18037 14415 18071
rect 2237 17833 2271 17867
rect 2789 17833 2823 17867
rect 4077 17833 4111 17867
rect 4537 17833 4571 17867
rect 5181 17833 5215 17867
rect 5641 17833 5675 17867
rect 9505 17833 9539 17867
rect 14473 17833 14507 17867
rect 3893 17765 3927 17799
rect 6193 17765 6227 17799
rect 9965 17765 9999 17799
rect 1409 17697 1443 17731
rect 4445 17697 4479 17731
rect 6920 17697 6954 17731
rect 10149 17697 10183 17731
rect 11428 17697 11462 17731
rect 2881 17629 2915 17663
rect 3065 17629 3099 17663
rect 4721 17629 4755 17663
rect 6653 17629 6687 17663
rect 11161 17629 11195 17663
rect 10333 17561 10367 17595
rect 1961 17493 1995 17527
rect 2421 17493 2455 17527
rect 3525 17493 3559 17527
rect 5549 17493 5583 17527
rect 6469 17493 6503 17527
rect 8033 17493 8067 17527
rect 12541 17493 12575 17527
rect 13277 17493 13311 17527
rect 14105 17493 14139 17527
rect 2145 17289 2179 17323
rect 4905 17289 4939 17323
rect 5273 17289 5307 17323
rect 6285 17289 6319 17323
rect 6653 17289 6687 17323
rect 8585 17289 8619 17323
rect 10517 17289 10551 17323
rect 12817 17289 12851 17323
rect 14657 17289 14691 17323
rect 5641 17221 5675 17255
rect 8309 17221 8343 17255
rect 9413 17221 9447 17255
rect 11253 17221 11287 17255
rect 13093 17221 13127 17255
rect 7297 17153 7331 17187
rect 7389 17153 7423 17187
rect 7941 17153 7975 17187
rect 9965 17153 9999 17187
rect 11345 17153 11379 17187
rect 13277 17153 13311 17187
rect 1409 17085 1443 17119
rect 2881 17085 2915 17119
rect 2973 17085 3007 17119
rect 5457 17085 5491 17119
rect 8401 17085 8435 17119
rect 9321 17085 9355 17119
rect 9781 17085 9815 17119
rect 2513 17017 2547 17051
rect 3240 17017 3274 17051
rect 7205 17017 7239 17051
rect 8953 17017 8987 17051
rect 9873 17017 9907 17051
rect 13522 17017 13556 17051
rect 1593 16949 1627 16983
rect 4353 16949 4387 16983
rect 6837 16949 6871 16983
rect 11805 16949 11839 16983
rect 1593 16745 1627 16779
rect 2421 16745 2455 16779
rect 3433 16745 3467 16779
rect 4445 16745 4479 16779
rect 5641 16745 5675 16779
rect 6745 16745 6779 16779
rect 7205 16745 7239 16779
rect 8217 16745 8251 16779
rect 8677 16745 8711 16779
rect 9505 16745 9539 16779
rect 9965 16745 9999 16779
rect 10333 16745 10367 16779
rect 13093 16745 13127 16779
rect 15761 16745 15795 16779
rect 4537 16677 4571 16711
rect 7665 16677 7699 16711
rect 1409 16609 1443 16643
rect 2513 16609 2547 16643
rect 3065 16609 3099 16643
rect 3893 16609 3927 16643
rect 5089 16609 5123 16643
rect 5549 16609 5583 16643
rect 6009 16609 6043 16643
rect 7573 16609 7607 16643
rect 11713 16609 11747 16643
rect 11980 16609 12014 16643
rect 15669 16609 15703 16643
rect 4721 16541 4755 16575
rect 6101 16541 6135 16575
rect 6285 16541 6319 16575
rect 7757 16541 7791 16575
rect 10425 16541 10459 16575
rect 10517 16541 10551 16575
rect 15945 16541 15979 16575
rect 1961 16405 1995 16439
rect 2697 16405 2731 16439
rect 4077 16405 4111 16439
rect 7021 16405 7055 16439
rect 15301 16405 15335 16439
rect 4721 16201 4755 16235
rect 5273 16201 5307 16235
rect 6193 16201 6227 16235
rect 6653 16201 6687 16235
rect 8585 16201 8619 16235
rect 9781 16201 9815 16235
rect 11805 16201 11839 16235
rect 16405 16201 16439 16235
rect 16037 16133 16071 16167
rect 2329 16065 2363 16099
rect 9321 16065 9355 16099
rect 9873 16065 9907 16099
rect 1409 15997 1443 16031
rect 2789 15997 2823 16031
rect 3045 15997 3079 16031
rect 7205 15997 7239 16031
rect 13553 15997 13587 16031
rect 13737 15997 13771 16031
rect 15669 15997 15703 16031
rect 5641 15929 5675 15963
rect 7450 15929 7484 15963
rect 10140 15929 10174 15963
rect 13982 15929 14016 15963
rect 1593 15861 1627 15895
rect 2697 15861 2731 15895
rect 4169 15861 4203 15895
rect 5733 15861 5767 15895
rect 7113 15861 7147 15895
rect 11253 15861 11287 15895
rect 12173 15861 12207 15895
rect 15117 15861 15151 15895
rect 1593 15657 1627 15691
rect 2237 15657 2271 15691
rect 2421 15657 2455 15691
rect 2881 15657 2915 15691
rect 3525 15657 3559 15691
rect 4261 15657 4295 15691
rect 4629 15657 4663 15691
rect 5273 15657 5307 15691
rect 8125 15657 8159 15691
rect 9413 15657 9447 15691
rect 10333 15657 10367 15691
rect 10793 15657 10827 15691
rect 11253 15657 11287 15691
rect 12357 15657 12391 15691
rect 12817 15657 12851 15691
rect 13829 15657 13863 15691
rect 14381 15657 14415 15691
rect 3893 15589 3927 15623
rect 6070 15589 6104 15623
rect 7849 15589 7883 15623
rect 11161 15589 11195 15623
rect 15761 15589 15795 15623
rect 1409 15521 1443 15555
rect 1961 15521 1995 15555
rect 2789 15521 2823 15555
rect 4077 15521 4111 15555
rect 5825 15521 5859 15555
rect 12725 15521 12759 15555
rect 14197 15521 14231 15555
rect 14657 15521 14691 15555
rect 15669 15521 15703 15555
rect 3065 15453 3099 15487
rect 8585 15453 8619 15487
rect 11437 15453 11471 15487
rect 13001 15453 13035 15487
rect 15853 15453 15887 15487
rect 9045 15385 9079 15419
rect 10057 15385 10091 15419
rect 5549 15317 5583 15351
rect 7205 15317 7239 15351
rect 15301 15317 15335 15351
rect 1961 15113 1995 15147
rect 3893 15113 3927 15147
rect 8585 15113 8619 15147
rect 10149 15113 10183 15147
rect 10885 15113 10919 15147
rect 11253 15113 11287 15147
rect 11529 15113 11563 15147
rect 12265 15113 12299 15147
rect 13093 15113 13127 15147
rect 1593 15045 1627 15079
rect 6285 15045 6319 15079
rect 2881 14977 2915 15011
rect 3065 14977 3099 15011
rect 4721 14977 4755 15011
rect 5733 14977 5767 15011
rect 7389 14977 7423 15011
rect 7849 14977 7883 15011
rect 8309 14977 8343 15011
rect 1409 14909 1443 14943
rect 3985 14909 4019 14943
rect 5549 14909 5583 14943
rect 5641 14909 5675 14943
rect 6653 14909 6687 14943
rect 7205 14909 7239 14943
rect 8769 14909 8803 14943
rect 9036 14909 9070 14943
rect 13829 14909 13863 14943
rect 13921 14909 13955 14943
rect 2329 14841 2363 14875
rect 2789 14841 2823 14875
rect 5089 14841 5123 14875
rect 12725 14841 12759 14875
rect 13461 14841 13495 14875
rect 14166 14841 14200 14875
rect 2421 14773 2455 14807
rect 3525 14773 3559 14807
rect 4169 14773 4203 14807
rect 5181 14773 5215 14807
rect 6837 14773 6871 14807
rect 7297 14773 7331 14807
rect 15301 14773 15335 14807
rect 15853 14773 15887 14807
rect 16221 14773 16255 14807
rect 16681 14773 16715 14807
rect 1593 14569 1627 14603
rect 3801 14569 3835 14603
rect 6009 14569 6043 14603
rect 7941 14569 7975 14603
rect 9689 14569 9723 14603
rect 14105 14569 14139 14603
rect 14933 14569 14967 14603
rect 2881 14501 2915 14535
rect 4344 14501 4378 14535
rect 15761 14501 15795 14535
rect 1409 14433 1443 14467
rect 2789 14433 2823 14467
rect 4077 14433 4111 14467
rect 6817 14433 6851 14467
rect 10057 14433 10091 14467
rect 10701 14433 10735 14467
rect 12981 14433 13015 14467
rect 15669 14433 15703 14467
rect 3065 14365 3099 14399
rect 3525 14365 3559 14399
rect 6561 14365 6595 14399
rect 9505 14365 9539 14399
rect 10149 14365 10183 14399
rect 10241 14365 10275 14399
rect 12725 14365 12759 14399
rect 15945 14365 15979 14399
rect 12265 14297 12299 14331
rect 1961 14229 1995 14263
rect 2237 14229 2271 14263
rect 2421 14229 2455 14263
rect 5457 14229 5491 14263
rect 6469 14229 6503 14263
rect 8861 14229 8895 14263
rect 11897 14229 11931 14263
rect 12541 14229 12575 14263
rect 15301 14229 15335 14263
rect 1593 14025 1627 14059
rect 4169 14025 4203 14059
rect 4537 14025 4571 14059
rect 5181 14025 5215 14059
rect 6193 14025 6227 14059
rect 6653 14025 6687 14059
rect 7205 14025 7239 14059
rect 8585 14025 8619 14059
rect 9873 14025 9907 14059
rect 10149 14025 10183 14059
rect 10333 14025 10367 14059
rect 11345 14025 11379 14059
rect 12265 14025 12299 14059
rect 12725 14025 12759 14059
rect 13277 14025 13311 14059
rect 14289 14025 14323 14059
rect 3157 13957 3191 13991
rect 14565 13957 14599 13991
rect 14657 13957 14691 13991
rect 2237 13889 2271 13923
rect 3709 13889 3743 13923
rect 5089 13889 5123 13923
rect 5733 13889 5767 13923
rect 7757 13889 7791 13923
rect 9413 13889 9447 13923
rect 10885 13889 10919 13923
rect 13185 13889 13219 13923
rect 13921 13889 13955 13923
rect 2053 13821 2087 13855
rect 2697 13821 2731 13855
rect 3065 13821 3099 13855
rect 3617 13821 3651 13855
rect 5641 13821 5675 13855
rect 7665 13821 7699 13855
rect 9137 13821 9171 13855
rect 10793 13821 10827 13855
rect 14565 13821 14599 13855
rect 14841 13821 14875 13855
rect 15108 13821 15142 13855
rect 16773 13821 16807 13855
rect 3525 13753 3559 13787
rect 5549 13753 5583 13787
rect 9229 13753 9263 13787
rect 10701 13753 10735 13787
rect 11805 13753 11839 13787
rect 13645 13753 13679 13787
rect 1961 13685 1995 13719
rect 7113 13685 7147 13719
rect 7573 13685 7607 13719
rect 8309 13685 8343 13719
rect 8769 13685 8803 13719
rect 13737 13685 13771 13719
rect 16221 13685 16255 13719
rect 2881 13481 2915 13515
rect 3525 13481 3559 13515
rect 4261 13481 4295 13515
rect 4813 13481 4847 13515
rect 5549 13481 5583 13515
rect 5917 13481 5951 13515
rect 6009 13481 6043 13515
rect 7573 13481 7607 13515
rect 9689 13481 9723 13515
rect 10149 13481 10183 13515
rect 10701 13481 10735 13515
rect 11805 13481 11839 13515
rect 13277 13481 13311 13515
rect 13829 13481 13863 13515
rect 16681 13481 16715 13515
rect 17325 13481 17359 13515
rect 7297 13413 7331 13447
rect 11069 13413 11103 13447
rect 12173 13413 12207 13447
rect 15117 13413 15151 13447
rect 17233 13413 17267 13447
rect 1409 13345 1443 13379
rect 2329 13345 2363 13379
rect 2789 13345 2823 13379
rect 4905 13345 4939 13379
rect 6377 13345 6411 13379
rect 8401 13345 8435 13379
rect 10057 13345 10091 13379
rect 13737 13345 13771 13379
rect 14381 13345 14415 13379
rect 15669 13345 15703 13379
rect 15761 13345 15795 13379
rect 3065 13277 3099 13311
rect 5089 13277 5123 13311
rect 6469 13277 6503 13311
rect 6561 13277 6595 13311
rect 8493 13277 8527 13311
rect 8677 13277 8711 13311
rect 10333 13277 10367 13311
rect 12265 13277 12299 13311
rect 12449 13277 12483 13311
rect 13921 13277 13955 13311
rect 15945 13277 15979 13311
rect 16313 13277 16347 13311
rect 17417 13277 17451 13311
rect 1593 13209 1627 13243
rect 1961 13209 1995 13243
rect 3893 13209 3927 13243
rect 13369 13209 13403 13243
rect 2421 13141 2455 13175
rect 4445 13141 4479 13175
rect 8033 13141 8067 13175
rect 9229 13141 9263 13175
rect 11437 13141 11471 13175
rect 12909 13141 12943 13175
rect 15301 13141 15335 13175
rect 16865 13141 16899 13175
rect 4353 12937 4387 12971
rect 6101 12937 6135 12971
rect 8033 12937 8067 12971
rect 8401 12937 8435 12971
rect 9045 12937 9079 12971
rect 11069 12937 11103 12971
rect 12541 12937 12575 12971
rect 13553 12937 13587 12971
rect 14013 12937 14047 12971
rect 14565 12937 14599 12971
rect 14933 12937 14967 12971
rect 17417 12937 17451 12971
rect 4077 12869 4111 12903
rect 6837 12869 6871 12903
rect 4997 12801 5031 12835
rect 5181 12801 5215 12835
rect 6653 12801 6687 12835
rect 7389 12801 7423 12835
rect 9137 12801 9171 12835
rect 13001 12801 13035 12835
rect 13185 12801 13219 12835
rect 17877 12801 17911 12835
rect 2053 12733 2087 12767
rect 4905 12733 4939 12767
rect 9404 12733 9438 12767
rect 11437 12733 11471 12767
rect 12909 12733 12943 12767
rect 15485 12733 15519 12767
rect 15741 12733 15775 12767
rect 18061 12733 18095 12767
rect 18328 12733 18362 12767
rect 2320 12665 2354 12699
rect 11897 12665 11931 12699
rect 12173 12665 12207 12699
rect 15393 12665 15427 12699
rect 1869 12597 1903 12631
rect 3433 12597 3467 12631
rect 4537 12597 4571 12631
rect 5641 12597 5675 12631
rect 7205 12597 7239 12631
rect 7297 12597 7331 12631
rect 10517 12597 10551 12631
rect 14105 12597 14139 12631
rect 16865 12597 16899 12631
rect 19441 12597 19475 12631
rect 2789 12393 2823 12427
rect 3801 12393 3835 12427
rect 5089 12393 5123 12427
rect 6745 12393 6779 12427
rect 7297 12393 7331 12427
rect 7849 12393 7883 12427
rect 9137 12393 9171 12427
rect 9689 12393 9723 12427
rect 10149 12393 10183 12427
rect 11253 12393 11287 12427
rect 12817 12393 12851 12427
rect 13645 12393 13679 12427
rect 14289 12393 14323 12427
rect 14749 12393 14783 12427
rect 15853 12393 15887 12427
rect 18061 12393 18095 12427
rect 7757 12325 7791 12359
rect 12633 12325 12667 12359
rect 1676 12257 1710 12291
rect 4077 12257 4111 12291
rect 5632 12257 5666 12291
rect 8217 12257 8251 12291
rect 10057 12257 10091 12291
rect 11621 12257 11655 12291
rect 11713 12257 11747 12291
rect 13185 12257 13219 12291
rect 1409 12189 1443 12223
rect 3433 12189 3467 12223
rect 5365 12189 5399 12223
rect 8309 12189 8343 12223
rect 8493 12189 8527 12223
rect 10333 12189 10367 12223
rect 11897 12189 11931 12223
rect 13277 12189 13311 12223
rect 13461 12189 13495 12223
rect 11161 12121 11195 12155
rect 17325 12325 17359 12359
rect 15761 12257 15795 12291
rect 16773 12257 16807 12291
rect 16037 12189 16071 12223
rect 17417 12189 17451 12223
rect 17601 12189 17635 12223
rect 4261 12053 4295 12087
rect 4721 12053 4755 12087
rect 10793 12053 10827 12087
rect 13645 12053 13679 12087
rect 13829 12053 13863 12087
rect 15025 12053 15059 12087
rect 15393 12053 15427 12087
rect 16405 12053 16439 12087
rect 16957 12053 16991 12087
rect 1593 11849 1627 11883
rect 4813 11849 4847 11883
rect 6285 11849 6319 11883
rect 9137 11849 9171 11883
rect 9781 11849 9815 11883
rect 10149 11849 10183 11883
rect 10793 11849 10827 11883
rect 11805 11849 11839 11883
rect 14473 11849 14507 11883
rect 15025 11849 15059 11883
rect 16405 11849 16439 11883
rect 1961 11781 1995 11815
rect 8861 11781 8895 11815
rect 10701 11781 10735 11815
rect 16037 11781 16071 11815
rect 11345 11713 11379 11747
rect 12449 11713 12483 11747
rect 15577 11713 15611 11747
rect 1409 11645 1443 11679
rect 2881 11645 2915 11679
rect 3148 11645 3182 11679
rect 6837 11645 6871 11679
rect 7093 11645 7127 11679
rect 11253 11645 11287 11679
rect 12265 11645 12299 11679
rect 2421 11577 2455 11611
rect 5825 11577 5859 11611
rect 11161 11577 11195 11611
rect 12541 11645 12575 11679
rect 12808 11645 12842 11679
rect 17049 11645 17083 11679
rect 15393 11577 15427 11611
rect 2789 11509 2823 11543
rect 4261 11509 4295 11543
rect 5457 11509 5491 11543
rect 6653 11509 6687 11543
rect 8217 11509 8251 11543
rect 12449 11509 12483 11543
rect 13921 11509 13955 11543
rect 14841 11509 14875 11543
rect 15485 11509 15519 11543
rect 17325 11509 17359 11543
rect 17785 11509 17819 11543
rect 1593 11305 1627 11339
rect 1961 11305 1995 11339
rect 2421 11305 2455 11339
rect 3801 11305 3835 11339
rect 4353 11305 4387 11339
rect 5273 11305 5307 11339
rect 6837 11305 6871 11339
rect 7481 11305 7515 11339
rect 7849 11305 7883 11339
rect 8953 11305 8987 11339
rect 9505 11305 9539 11339
rect 12909 11305 12943 11339
rect 13277 11305 13311 11339
rect 14289 11305 14323 11339
rect 14749 11305 14783 11339
rect 16037 11305 16071 11339
rect 17233 11305 17267 11339
rect 2881 11237 2915 11271
rect 3433 11237 3467 11271
rect 5724 11237 5758 11271
rect 13921 11237 13955 11271
rect 17141 11237 17175 11271
rect 17693 11237 17727 11271
rect 1409 11169 1443 11203
rect 2789 11169 2823 11203
rect 4169 11169 4203 11203
rect 5457 11169 5491 11203
rect 8309 11169 8343 11203
rect 10692 11169 10726 11203
rect 15025 11169 15059 11203
rect 15577 11169 15611 11203
rect 17601 11169 17635 11203
rect 2973 11101 3007 11135
rect 4629 11101 4663 11135
rect 8401 11101 8435 11135
rect 8493 11101 8527 11135
rect 10425 11101 10459 11135
rect 13369 11101 13403 11135
rect 13461 11101 13495 11135
rect 16129 11101 16163 11135
rect 16313 11101 16347 11135
rect 16773 11101 16807 11135
rect 17877 11101 17911 11135
rect 2329 11033 2363 11067
rect 7941 11033 7975 11067
rect 11805 11033 11839 11067
rect 15669 11033 15703 11067
rect 9965 10965 9999 10999
rect 10333 10965 10367 10999
rect 12541 10965 12575 10999
rect 18337 10965 18371 10999
rect 1409 10761 1443 10795
rect 3249 10761 3283 10795
rect 4353 10761 4387 10795
rect 5181 10761 5215 10795
rect 6653 10761 6687 10795
rect 7297 10761 7331 10795
rect 9689 10761 9723 10795
rect 11345 10761 11379 10795
rect 13461 10761 13495 10795
rect 14657 10761 14691 10795
rect 14933 10761 14967 10795
rect 15393 10761 15427 10795
rect 18061 10761 18095 10795
rect 10241 10693 10275 10727
rect 2053 10625 2087 10659
rect 3065 10625 3099 10659
rect 3801 10625 3835 10659
rect 4721 10625 4755 10659
rect 5089 10625 5123 10659
rect 5825 10625 5859 10659
rect 10793 10625 10827 10659
rect 13093 10625 13127 10659
rect 15485 10625 15519 10659
rect 18613 10625 18647 10659
rect 1777 10557 1811 10591
rect 3709 10557 3743 10591
rect 5641 10557 5675 10591
rect 6285 10557 6319 10591
rect 7665 10557 7699 10591
rect 7757 10557 7791 10591
rect 10701 10557 10735 10591
rect 12817 10557 12851 10591
rect 12909 10557 12943 10591
rect 13829 10557 13863 10591
rect 1869 10489 1903 10523
rect 2789 10489 2823 10523
rect 3617 10489 3651 10523
rect 8024 10489 8058 10523
rect 10057 10489 10091 10523
rect 10609 10489 10643 10523
rect 12265 10489 12299 10523
rect 15752 10489 15786 10523
rect 17877 10489 17911 10523
rect 18521 10489 18555 10523
rect 5549 10421 5583 10455
rect 9137 10421 9171 10455
rect 11621 10421 11655 10455
rect 12449 10421 12483 10455
rect 14197 10421 14231 10455
rect 16865 10421 16899 10455
rect 17417 10421 17451 10455
rect 18429 10421 18463 10455
rect 3433 10217 3467 10251
rect 3801 10217 3835 10251
rect 4905 10217 4939 10251
rect 6285 10217 6319 10251
rect 6469 10217 6503 10251
rect 8493 10217 8527 10251
rect 9413 10217 9447 10251
rect 11069 10217 11103 10251
rect 12541 10217 12575 10251
rect 13829 10217 13863 10251
rect 15117 10217 15151 10251
rect 15577 10217 15611 10251
rect 18061 10217 18095 10251
rect 18521 10217 18555 10251
rect 18981 10217 19015 10251
rect 6929 10149 6963 10183
rect 7941 10149 7975 10183
rect 9045 10149 9079 10183
rect 14197 10149 14231 10183
rect 1777 10081 1811 10115
rect 2421 10081 2455 10115
rect 5273 10081 5307 10115
rect 6837 10081 6871 10115
rect 8401 10081 8435 10115
rect 9945 10081 9979 10115
rect 13185 10081 13219 10115
rect 16293 10081 16327 10115
rect 18889 10081 18923 10115
rect 1869 10013 1903 10047
rect 1961 10013 1995 10047
rect 5365 10013 5399 10047
rect 5457 10013 5491 10047
rect 7113 10013 7147 10047
rect 8585 10013 8619 10047
rect 9689 10013 9723 10047
rect 13277 10013 13311 10047
rect 13461 10013 13495 10047
rect 16037 10013 16071 10047
rect 19073 10013 19107 10047
rect 1409 9945 1443 9979
rect 12817 9945 12851 9979
rect 3065 9877 3099 9911
rect 4353 9877 4387 9911
rect 4629 9877 4663 9911
rect 5917 9877 5951 9911
rect 7481 9877 7515 9911
rect 8033 9877 8067 9911
rect 11621 9877 11655 9911
rect 11989 9877 12023 9911
rect 14565 9877 14599 9911
rect 15945 9877 15979 9911
rect 17417 9877 17451 9911
rect 1409 9673 1443 9707
rect 5365 9673 5399 9707
rect 6285 9673 6319 9707
rect 9689 9673 9723 9707
rect 13277 9673 13311 9707
rect 19073 9673 19107 9707
rect 2421 9605 2455 9639
rect 8217 9605 8251 9639
rect 12265 9605 12299 9639
rect 15209 9605 15243 9639
rect 16313 9605 16347 9639
rect 18061 9605 18095 9639
rect 19809 9605 19843 9639
rect 1961 9537 1995 9571
rect 5549 9537 5583 9571
rect 10333 9537 10367 9571
rect 11345 9537 11379 9571
rect 16865 9537 16899 9571
rect 18613 9537 18647 9571
rect 3065 9469 3099 9503
rect 3332 9469 3366 9503
rect 6837 9469 6871 9503
rect 7104 9469 7138 9503
rect 13829 9469 13863 9503
rect 16037 9469 16071 9503
rect 16681 9469 16715 9503
rect 19441 9469 19475 9503
rect 1869 9401 1903 9435
rect 11253 9401 11287 9435
rect 12909 9401 12943 9435
rect 14074 9401 14108 9435
rect 16773 9401 16807 9435
rect 18429 9401 18463 9435
rect 1777 9333 1811 9367
rect 2789 9333 2823 9367
rect 4445 9333 4479 9367
rect 4997 9333 5031 9367
rect 6561 9333 6595 9367
rect 8769 9333 8803 9367
rect 9321 9333 9355 9367
rect 10609 9333 10643 9367
rect 10793 9333 10827 9367
rect 11161 9333 11195 9367
rect 11805 9333 11839 9367
rect 13645 9333 13679 9367
rect 17417 9333 17451 9367
rect 17785 9333 17819 9367
rect 18521 9333 18555 9367
rect 3433 9129 3467 9163
rect 5457 9129 5491 9163
rect 6561 9129 6595 9163
rect 8033 9129 8067 9163
rect 8401 9129 8435 9163
rect 9689 9129 9723 9163
rect 10149 9129 10183 9163
rect 11621 9129 11655 9163
rect 15669 9129 15703 9163
rect 18981 9129 19015 9163
rect 19349 9129 19383 9163
rect 4077 9061 4111 9095
rect 11161 9061 11195 9095
rect 14933 9061 14967 9095
rect 15577 9061 15611 9095
rect 16497 9061 16531 9095
rect 1501 8993 1535 9027
rect 1768 8993 1802 9027
rect 4997 8993 5031 9027
rect 5365 8993 5399 9027
rect 5825 8993 5859 9027
rect 5917 8993 5951 9027
rect 8493 8993 8527 9027
rect 10057 8993 10091 9027
rect 12061 8993 12095 9027
rect 16681 8993 16715 9027
rect 16948 8993 16982 9027
rect 6009 8925 6043 8959
rect 8585 8925 8619 8959
rect 10333 8925 10367 8959
rect 11805 8925 11839 8959
rect 14197 8925 14231 8959
rect 14565 8925 14599 8959
rect 16221 8925 16255 8959
rect 2881 8857 2915 8891
rect 3801 8857 3835 8891
rect 4537 8857 4571 8891
rect 9413 8857 9447 8891
rect 6929 8789 6963 8823
rect 7205 8789 7239 8823
rect 7573 8789 7607 8823
rect 9045 8789 9079 8823
rect 10885 8789 10919 8823
rect 13185 8789 13219 8823
rect 13921 8789 13955 8823
rect 18061 8789 18095 8823
rect 18613 8789 18647 8823
rect 2697 8585 2731 8619
rect 10057 8585 10091 8619
rect 10701 8585 10735 8619
rect 11805 8585 11839 8619
rect 12173 8585 12207 8619
rect 14381 8585 14415 8619
rect 17141 8585 17175 8619
rect 17877 8585 17911 8619
rect 12817 8517 12851 8551
rect 15301 8517 15335 8551
rect 16129 8517 16163 8551
rect 1409 8449 1443 8483
rect 3157 8449 3191 8483
rect 3249 8449 3283 8483
rect 6653 8449 6687 8483
rect 7389 8449 7423 8483
rect 11345 8449 11379 8483
rect 13001 8449 13035 8483
rect 16681 8449 16715 8483
rect 18521 8449 18555 8483
rect 18705 8449 18739 8483
rect 3985 8381 4019 8415
rect 4261 8381 4295 8415
rect 4528 8381 4562 8415
rect 6285 8381 6319 8415
rect 7297 8381 7331 8415
rect 8585 8381 8619 8415
rect 8677 8381 8711 8415
rect 15945 8381 15979 8415
rect 16589 8381 16623 8415
rect 2605 8313 2639 8347
rect 3065 8313 3099 8347
rect 3801 8313 3835 8347
rect 7205 8313 7239 8347
rect 8217 8313 8251 8347
rect 8944 8313 8978 8347
rect 13246 8313 13280 8347
rect 16497 8313 16531 8347
rect 18429 8313 18463 8347
rect 19073 8313 19107 8347
rect 1961 8245 1995 8279
rect 3985 8245 4019 8279
rect 4077 8245 4111 8279
rect 5641 8245 5675 8279
rect 6837 8245 6871 8279
rect 11161 8245 11195 8279
rect 15669 8245 15703 8279
rect 18061 8245 18095 8279
rect 1869 8041 1903 8075
rect 2789 8041 2823 8075
rect 4445 8041 4479 8075
rect 7481 8041 7515 8075
rect 8125 8041 8159 8075
rect 10885 8041 10919 8075
rect 11713 8041 11747 8075
rect 12081 8041 12115 8075
rect 13277 8041 13311 8075
rect 13645 8041 13679 8075
rect 16405 8041 16439 8075
rect 17049 8041 17083 8075
rect 17601 8041 17635 8075
rect 1777 7905 1811 7939
rect 3065 7905 3099 7939
rect 5181 7905 5215 7939
rect 6357 7905 6391 7939
rect 10057 7905 10091 7939
rect 13737 7905 13771 7939
rect 17969 7905 18003 7939
rect 2053 7837 2087 7871
rect 4537 7837 4571 7871
rect 4721 7837 4755 7871
rect 6101 7837 6135 7871
rect 8585 7837 8619 7871
rect 10149 7837 10183 7871
rect 10241 7837 10275 7871
rect 12173 7837 12207 7871
rect 12265 7837 12299 7871
rect 13093 7837 13127 7871
rect 13921 7837 13955 7871
rect 15117 7837 15151 7871
rect 16497 7837 16531 7871
rect 16681 7837 16715 7871
rect 18061 7837 18095 7871
rect 18245 7837 18279 7871
rect 18981 7837 19015 7871
rect 9413 7769 9447 7803
rect 9689 7769 9723 7803
rect 14749 7769 14783 7803
rect 17417 7769 17451 7803
rect 1409 7701 1443 7735
rect 3525 7701 3559 7735
rect 3801 7701 3835 7735
rect 4077 7701 4111 7735
rect 5549 7701 5583 7735
rect 5917 7701 5951 7735
rect 8401 7701 8435 7735
rect 9045 7701 9079 7735
rect 11253 7701 11287 7735
rect 11529 7701 11563 7735
rect 14289 7701 14323 7735
rect 15761 7701 15795 7735
rect 16037 7701 16071 7735
rect 18613 7701 18647 7735
rect 19717 7701 19751 7735
rect 2421 7497 2455 7531
rect 2605 7497 2639 7531
rect 2973 7497 3007 7531
rect 8217 7497 8251 7531
rect 8677 7497 8711 7531
rect 10793 7497 10827 7531
rect 11897 7497 11931 7531
rect 13645 7497 13679 7531
rect 14657 7497 14691 7531
rect 15485 7497 15519 7531
rect 15669 7497 15703 7531
rect 1869 7361 1903 7395
rect 2053 7361 2087 7395
rect 1777 7225 1811 7259
rect 5181 7429 5215 7463
rect 6653 7429 6687 7463
rect 8401 7429 8435 7463
rect 8493 7429 8527 7463
rect 10149 7429 10183 7463
rect 19625 7429 19659 7463
rect 3433 7361 3467 7395
rect 3617 7361 3651 7395
rect 5825 7361 5859 7395
rect 7297 7361 7331 7395
rect 7481 7361 7515 7395
rect 3341 7293 3375 7327
rect 7205 7293 7239 7327
rect 9321 7361 9355 7395
rect 9781 7361 9815 7395
rect 11345 7361 11379 7395
rect 12449 7361 12483 7395
rect 13185 7361 13219 7395
rect 14105 7361 14139 7395
rect 14289 7361 14323 7395
rect 15209 7361 15243 7395
rect 16313 7361 16347 7395
rect 18521 7361 18555 7395
rect 18613 7361 18647 7395
rect 19533 7361 19567 7395
rect 20177 7361 20211 7395
rect 9045 7293 9079 7327
rect 11253 7293 11287 7327
rect 16037 7293 16071 7327
rect 17601 7293 17635 7327
rect 18429 7293 18463 7327
rect 19073 7293 19107 7327
rect 2789 7225 2823 7259
rect 5089 7225 5123 7259
rect 5641 7225 5675 7259
rect 8401 7225 8435 7259
rect 9137 7225 9171 7259
rect 12173 7225 12207 7259
rect 13553 7225 13587 7259
rect 14013 7225 14047 7259
rect 17233 7225 17267 7259
rect 1409 7157 1443 7191
rect 2605 7157 2639 7191
rect 4077 7157 4111 7191
rect 4445 7157 4479 7191
rect 5549 7157 5583 7191
rect 6193 7157 6227 7191
rect 6837 7157 6871 7191
rect 10609 7157 10643 7191
rect 11161 7157 11195 7191
rect 16129 7157 16163 7191
rect 16773 7157 16807 7191
rect 18061 7157 18095 7191
rect 19993 7157 20027 7191
rect 20085 7157 20119 7191
rect 1409 6953 1443 6987
rect 3525 6953 3559 6987
rect 9045 6953 9079 6987
rect 9413 6953 9447 6987
rect 9689 6953 9723 6987
rect 10057 6953 10091 6987
rect 13921 6953 13955 6987
rect 17785 6953 17819 6987
rect 18429 6953 18463 6987
rect 19257 6953 19291 6987
rect 1869 6885 1903 6919
rect 2881 6885 2915 6919
rect 13185 6885 13219 6919
rect 2789 6817 2823 6851
rect 4445 6817 4479 6851
rect 6265 6817 6299 6851
rect 8493 6817 8527 6851
rect 11621 6817 11655 6851
rect 15393 6817 15427 6851
rect 16672 6817 16706 6851
rect 3065 6749 3099 6783
rect 4537 6749 4571 6783
rect 4721 6749 4755 6783
rect 6009 6749 6043 6783
rect 10149 6749 10183 6783
rect 10241 6749 10275 6783
rect 11713 6749 11747 6783
rect 11897 6749 11931 6783
rect 13277 6749 13311 6783
rect 13461 6749 13495 6783
rect 14565 6749 14599 6783
rect 16405 6749 16439 6783
rect 19349 6749 19383 6783
rect 19441 6749 19475 6783
rect 3893 6681 3927 6715
rect 12817 6681 12851 6715
rect 18889 6681 18923 6715
rect 20545 6681 20579 6715
rect 2237 6613 2271 6647
rect 2421 6613 2455 6647
rect 4077 6613 4111 6647
rect 5181 6613 5215 6647
rect 5641 6613 5675 6647
rect 7389 6613 7423 6647
rect 7941 6613 7975 6647
rect 8309 6613 8343 6647
rect 10793 6613 10827 6647
rect 11253 6613 11287 6647
rect 12541 6613 12575 6647
rect 14289 6613 14323 6647
rect 15025 6613 15059 6647
rect 16221 6613 16255 6647
rect 18705 6613 18739 6647
rect 19993 6613 20027 6647
rect 4997 6409 5031 6443
rect 5181 6409 5215 6443
rect 6837 6409 6871 6443
rect 8309 6409 8343 6443
rect 9045 6409 9079 6443
rect 9413 6409 9447 6443
rect 11437 6409 11471 6443
rect 11897 6409 11931 6443
rect 14197 6409 14231 6443
rect 16405 6409 16439 6443
rect 17785 6409 17819 6443
rect 20545 6409 20579 6443
rect 8585 6341 8619 6375
rect 19441 6341 19475 6375
rect 20361 6341 20395 6375
rect 5641 6273 5675 6307
rect 5825 6273 5859 6307
rect 7481 6273 7515 6307
rect 7849 6273 7883 6307
rect 9505 6273 9539 6307
rect 13001 6273 13035 6307
rect 14289 6273 14323 6307
rect 18061 6273 18095 6307
rect 21005 6273 21039 6307
rect 21189 6273 21223 6307
rect 2237 6205 2271 6239
rect 2504 6205 2538 6239
rect 5549 6205 5583 6239
rect 7297 6205 7331 6239
rect 16865 6205 16899 6239
rect 17417 6205 17451 6239
rect 18328 6205 18362 6239
rect 20913 6205 20947 6239
rect 21557 6205 21591 6239
rect 22293 6205 22327 6239
rect 22753 6205 22787 6239
rect 2145 6137 2179 6171
rect 7205 6137 7239 6171
rect 9772 6137 9806 6171
rect 12817 6137 12851 6171
rect 14556 6137 14590 6171
rect 19993 6137 20027 6171
rect 1685 6069 1719 6103
rect 3617 6069 3651 6103
rect 4261 6069 4295 6103
rect 4629 6069 4663 6103
rect 6193 6069 6227 6103
rect 6653 6069 6687 6103
rect 10885 6069 10919 6103
rect 12173 6069 12207 6103
rect 12449 6069 12483 6103
rect 12909 6069 12943 6103
rect 13461 6069 13495 6103
rect 15669 6069 15703 6103
rect 17049 6069 17083 6103
rect 22477 6069 22511 6103
rect 2789 5865 2823 5899
rect 5457 5865 5491 5899
rect 6101 5865 6135 5899
rect 6469 5865 6503 5899
rect 6561 5865 6595 5899
rect 7941 5865 7975 5899
rect 9505 5865 9539 5899
rect 11069 5865 11103 5899
rect 14381 5865 14415 5899
rect 18153 5865 18187 5899
rect 18981 5865 19015 5899
rect 19717 5865 19751 5899
rect 20913 5865 20947 5899
rect 11713 5797 11747 5831
rect 15577 5797 15611 5831
rect 17018 5797 17052 5831
rect 20545 5797 20579 5831
rect 1409 5729 1443 5763
rect 1676 5729 1710 5763
rect 4077 5729 4111 5763
rect 4344 5729 4378 5763
rect 6929 5729 6963 5763
rect 8309 5729 8343 5763
rect 9689 5729 9723 5763
rect 9956 5729 9990 5763
rect 12173 5729 12207 5763
rect 12440 5729 12474 5763
rect 15669 5729 15703 5763
rect 19625 5729 19659 5763
rect 21281 5729 21315 5763
rect 23305 5729 23339 5763
rect 7021 5661 7055 5695
rect 7205 5661 7239 5695
rect 8585 5661 8619 5695
rect 16773 5661 16807 5695
rect 19809 5661 19843 5695
rect 21373 5661 21407 5695
rect 21465 5661 21499 5695
rect 9045 5593 9079 5627
rect 14657 5593 14691 5627
rect 15853 5593 15887 5627
rect 19257 5593 19291 5627
rect 3709 5525 3743 5559
rect 7573 5525 7607 5559
rect 12081 5525 12115 5559
rect 13553 5525 13587 5559
rect 15117 5525 15151 5559
rect 16497 5525 16531 5559
rect 23489 5525 23523 5559
rect 2421 5321 2455 5355
rect 2881 5321 2915 5355
rect 4629 5321 4663 5355
rect 9137 5321 9171 5355
rect 13001 5321 13035 5355
rect 14933 5321 14967 5355
rect 17417 5321 17451 5355
rect 18061 5321 18095 5355
rect 19625 5321 19659 5355
rect 21649 5321 21683 5355
rect 22109 5321 22143 5355
rect 23305 5321 23339 5355
rect 1409 5253 1443 5287
rect 12173 5253 12207 5287
rect 16313 5253 16347 5287
rect 20637 5253 20671 5287
rect 22385 5253 22419 5287
rect 1869 5185 1903 5219
rect 2053 5185 2087 5219
rect 4261 5185 4295 5219
rect 5825 5185 5859 5219
rect 8861 5185 8895 5219
rect 17049 5185 17083 5219
rect 17785 5185 17819 5219
rect 18613 5185 18647 5219
rect 20177 5185 20211 5219
rect 21005 5185 21039 5219
rect 1777 5117 1811 5151
rect 4077 5117 4111 5151
rect 6561 5117 6595 5151
rect 6837 5117 6871 5151
rect 7104 5117 7138 5151
rect 9321 5117 9355 5151
rect 9588 5117 9622 5151
rect 12541 5117 12575 5151
rect 13553 5117 13587 5151
rect 15669 5117 15703 5151
rect 16773 5117 16807 5151
rect 18429 5117 18463 5151
rect 18521 5117 18555 5151
rect 21189 5117 21223 5151
rect 22753 5117 22787 5151
rect 3525 5049 3559 5083
rect 5089 5049 5123 5083
rect 11253 5049 11287 5083
rect 13369 5049 13403 5083
rect 13798 5049 13832 5083
rect 16865 5049 16899 5083
rect 19993 5049 20027 5083
rect 3617 4981 3651 5015
rect 3985 4981 4019 5015
rect 5181 4981 5215 5015
rect 5549 4981 5583 5015
rect 5641 4981 5675 5015
rect 6285 4981 6319 5015
rect 8217 4981 8251 5015
rect 10701 4981 10735 5015
rect 11621 4981 11655 5015
rect 12725 4981 12759 5015
rect 16405 4981 16439 5015
rect 19073 4981 19107 5015
rect 19533 4981 19567 5015
rect 20085 4981 20119 5015
rect 21373 4981 21407 5015
rect 1685 4777 1719 4811
rect 2881 4777 2915 4811
rect 3709 4777 3743 4811
rect 4353 4777 4387 4811
rect 5917 4777 5951 4811
rect 6009 4777 6043 4811
rect 7113 4777 7147 4811
rect 9321 4777 9355 4811
rect 10977 4777 11011 4811
rect 11437 4777 11471 4811
rect 11989 4777 12023 4811
rect 12909 4777 12943 4811
rect 13921 4777 13955 4811
rect 16129 4777 16163 4811
rect 16497 4777 16531 4811
rect 16957 4777 16991 4811
rect 20269 4777 20303 4811
rect 21557 4777 21591 4811
rect 21833 4777 21867 4811
rect 2789 4709 2823 4743
rect 6929 4709 6963 4743
rect 10517 4709 10551 4743
rect 13001 4709 13035 4743
rect 19349 4709 19383 4743
rect 7481 4641 7515 4675
rect 9965 4641 9999 4675
rect 10793 4641 10827 4675
rect 11345 4641 11379 4675
rect 14105 4641 14139 4675
rect 15301 4641 15335 4675
rect 16865 4641 16899 4675
rect 17509 4641 17543 4675
rect 17877 4641 17911 4675
rect 18429 4641 18463 4675
rect 19625 4641 19659 4675
rect 20913 4641 20947 4675
rect 2973 4573 3007 4607
rect 6101 4573 6135 4607
rect 7573 4573 7607 4607
rect 7665 4573 7699 4607
rect 11621 4573 11655 4607
rect 13093 4573 13127 4607
rect 13645 4573 13679 4607
rect 15025 4573 15059 4607
rect 17141 4573 17175 4607
rect 18521 4573 18555 4607
rect 18613 4573 18647 4607
rect 2421 4505 2455 4539
rect 5273 4505 5307 4539
rect 12541 4505 12575 4539
rect 14657 4505 14691 4539
rect 15485 4505 15519 4539
rect 19809 4505 19843 4539
rect 2329 4437 2363 4471
rect 4629 4437 4663 4471
rect 5549 4437 5583 4471
rect 8125 4437 8159 4471
rect 8493 4437 8527 4471
rect 8861 4437 8895 4471
rect 10149 4437 10183 4471
rect 12449 4437 12483 4471
rect 14289 4437 14323 4471
rect 18061 4437 18095 4471
rect 20545 4437 20579 4471
rect 21097 4437 21131 4471
rect 3801 4233 3835 4267
rect 6193 4233 6227 4267
rect 7573 4233 7607 4267
rect 10701 4233 10735 4267
rect 11713 4233 11747 4267
rect 14013 4233 14047 4267
rect 15301 4233 15335 4267
rect 19625 4233 19659 4267
rect 21097 4233 21131 4267
rect 12449 4165 12483 4199
rect 2973 4097 3007 4131
rect 3893 4097 3927 4131
rect 6653 4097 6687 4131
rect 8309 4097 8343 4131
rect 9873 4097 9907 4131
rect 11253 4097 11287 4131
rect 12909 4097 12943 4131
rect 13093 4097 13127 4131
rect 13921 4097 13955 4131
rect 14565 4097 14599 4131
rect 16589 4097 16623 4131
rect 16681 4097 16715 4131
rect 18705 4097 18739 4131
rect 19165 4097 19199 4131
rect 20269 4097 20303 4131
rect 3433 4029 3467 4063
rect 8125 4029 8159 4063
rect 8769 4029 8803 4063
rect 11069 4029 11103 4063
rect 13461 4029 13495 4063
rect 14381 4029 14415 4063
rect 16497 4029 16531 4063
rect 18429 4029 18463 4063
rect 20085 4029 20119 4063
rect 20637 4029 20671 4063
rect 21189 4029 21223 4063
rect 21741 4029 21775 4063
rect 22109 4029 22143 4063
rect 22293 4029 22327 4063
rect 22753 4029 22787 4063
rect 1869 3961 1903 3995
rect 2237 3961 2271 3995
rect 2789 3961 2823 3995
rect 4160 3961 4194 3995
rect 5825 3961 5859 3995
rect 9781 3961 9815 3995
rect 14473 3961 14507 3995
rect 16037 3961 16071 3995
rect 18521 3961 18555 3995
rect 2329 3893 2363 3927
rect 2697 3893 2731 3927
rect 5273 3893 5307 3927
rect 7205 3893 7239 3927
rect 7757 3893 7791 3927
rect 8217 3893 8251 3927
rect 9137 3893 9171 3927
rect 9321 3893 9355 3927
rect 9689 3893 9723 3927
rect 12173 3893 12207 3927
rect 12817 3893 12851 3927
rect 16129 3893 16163 3927
rect 17417 3893 17451 3927
rect 17785 3893 17819 3927
rect 18061 3893 18095 3927
rect 19441 3893 19475 3927
rect 19993 3893 20027 3927
rect 21373 3893 21407 3927
rect 22477 3893 22511 3927
rect 1593 3689 1627 3723
rect 2237 3689 2271 3723
rect 3157 3689 3191 3723
rect 3617 3689 3651 3723
rect 5365 3689 5399 3723
rect 6929 3689 6963 3723
rect 8033 3689 8067 3723
rect 9413 3689 9447 3723
rect 10149 3689 10183 3723
rect 11253 3689 11287 3723
rect 13093 3689 13127 3723
rect 13645 3689 13679 3723
rect 14013 3689 14047 3723
rect 14381 3689 14415 3723
rect 14657 3689 14691 3723
rect 15945 3689 15979 3723
rect 16589 3689 16623 3723
rect 18061 3689 18095 3723
rect 18705 3689 18739 3723
rect 20177 3689 20211 3723
rect 2145 3621 2179 3655
rect 2881 3621 2915 3655
rect 5816 3621 5850 3655
rect 10609 3621 10643 3655
rect 11980 3621 12014 3655
rect 5549 3553 5583 3587
rect 8401 3553 8435 3587
rect 9965 3553 9999 3587
rect 10517 3553 10551 3587
rect 11713 3553 11747 3587
rect 14197 3553 14231 3587
rect 15301 3553 15335 3587
rect 16948 3553 16982 3587
rect 19533 3553 19567 3587
rect 19625 3553 19659 3587
rect 20545 3553 20579 3587
rect 21097 3553 21131 3587
rect 22201 3553 22235 3587
rect 2421 3485 2455 3519
rect 8493 3485 8527 3519
rect 8585 3485 8619 3519
rect 10793 3485 10827 3519
rect 16681 3485 16715 3519
rect 19717 3485 19751 3519
rect 7573 3417 7607 3451
rect 15485 3417 15519 3451
rect 19165 3417 19199 3451
rect 1777 3349 1811 3383
rect 4537 3349 4571 3383
rect 4905 3349 4939 3383
rect 7849 3349 7883 3383
rect 15025 3349 15059 3383
rect 18981 3349 19015 3383
rect 21281 3349 21315 3383
rect 22385 3349 22419 3383
rect 1869 3145 1903 3179
rect 3525 3145 3559 3179
rect 4077 3145 4111 3179
rect 4905 3145 4939 3179
rect 6837 3145 6871 3179
rect 8125 3145 8159 3179
rect 9781 3145 9815 3179
rect 10793 3145 10827 3179
rect 11161 3145 11195 3179
rect 11805 3145 11839 3179
rect 12173 3145 12207 3179
rect 14013 3145 14047 3179
rect 14565 3145 14599 3179
rect 15025 3145 15059 3179
rect 16497 3145 16531 3179
rect 17417 3145 17451 3179
rect 17785 3145 17819 3179
rect 18061 3145 18095 3179
rect 19165 3145 19199 3179
rect 19625 3145 19659 3179
rect 22569 3145 22603 3179
rect 23857 3145 23891 3179
rect 17049 3077 17083 3111
rect 5365 3009 5399 3043
rect 5457 3009 5491 3043
rect 7481 3009 7515 3043
rect 8401 3009 8435 3043
rect 12633 3009 12667 3043
rect 18705 3009 18739 3043
rect 20269 3009 20303 3043
rect 20637 3009 20671 3043
rect 2145 2941 2179 2975
rect 2412 2941 2446 2975
rect 11253 2941 11287 2975
rect 15117 2941 15151 2975
rect 15373 2941 15407 2975
rect 18429 2941 18463 2975
rect 19993 2941 20027 2975
rect 21373 2941 21407 2975
rect 21649 2941 21683 2975
rect 22201 2941 22235 2975
rect 23673 2941 23707 2975
rect 24225 2941 24259 2975
rect 4813 2873 4847 2907
rect 5273 2873 5307 2907
rect 6653 2873 6687 2907
rect 7297 2873 7331 2907
rect 8668 2873 8702 2907
rect 10333 2873 10367 2907
rect 12900 2873 12934 2907
rect 18521 2873 18555 2907
rect 6193 2805 6227 2839
rect 7205 2805 7239 2839
rect 11437 2805 11471 2839
rect 20085 2805 20119 2839
rect 21005 2805 21039 2839
rect 21833 2805 21867 2839
rect 2421 2601 2455 2635
rect 3525 2601 3559 2635
rect 3893 2601 3927 2635
rect 5457 2601 5491 2635
rect 6377 2601 6411 2635
rect 7941 2601 7975 2635
rect 8125 2601 8159 2635
rect 9597 2601 9631 2635
rect 10149 2601 10183 2635
rect 10793 2601 10827 2635
rect 11345 2601 11379 2635
rect 12449 2601 12483 2635
rect 13001 2601 13035 2635
rect 14197 2601 14231 2635
rect 15485 2601 15519 2635
rect 16681 2601 16715 2635
rect 18061 2601 18095 2635
rect 18337 2601 18371 2635
rect 20821 2601 20855 2635
rect 21465 2601 21499 2635
rect 1961 2533 1995 2567
rect 2789 2533 2823 2567
rect 4322 2533 4356 2567
rect 10241 2533 10275 2567
rect 15945 2533 15979 2567
rect 18797 2533 18831 2567
rect 19441 2533 19475 2567
rect 4077 2465 4111 2499
rect 6009 2465 6043 2499
rect 7113 2465 7147 2499
rect 8493 2465 8527 2499
rect 9137 2465 9171 2499
rect 11437 2465 11471 2499
rect 13093 2465 13127 2499
rect 14289 2465 14323 2499
rect 14841 2465 14875 2499
rect 15853 2465 15887 2499
rect 17141 2465 17175 2499
rect 17693 2465 17727 2499
rect 18705 2465 18739 2499
rect 19901 2465 19935 2499
rect 20453 2465 20487 2499
rect 22201 2465 22235 2499
rect 22753 2465 22787 2499
rect 24041 2465 24075 2499
rect 24593 2465 24627 2499
rect 1409 2397 1443 2431
rect 2329 2397 2363 2431
rect 2881 2397 2915 2431
rect 3065 2397 3099 2431
rect 7665 2397 7699 2431
rect 8585 2397 8619 2431
rect 8769 2397 8803 2431
rect 10425 2397 10459 2431
rect 11989 2397 12023 2431
rect 13277 2397 13311 2431
rect 13645 2397 13679 2431
rect 16037 2397 16071 2431
rect 18889 2397 18923 2431
rect 19717 2397 19751 2431
rect 9781 2329 9815 2363
rect 11621 2329 11655 2363
rect 12633 2329 12667 2363
rect 14473 2329 14507 2363
rect 7297 2261 7331 2295
rect 15301 2261 15335 2295
rect 17325 2261 17359 2295
rect 20085 2261 20119 2295
rect 22385 2261 22419 2295
rect 24225 2261 24259 2295
<< metal1 >>
rect 7558 27412 7564 27464
rect 7616 27452 7622 27464
rect 7650 27452 7656 27464
rect 7616 27424 7656 27452
rect 7616 27412 7622 27424
rect 7650 27412 7656 27424
rect 7708 27412 7714 27464
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1397 25347 1455 25353
rect 1397 25313 1409 25347
rect 1443 25344 1455 25347
rect 1946 25344 1952 25356
rect 1443 25316 1952 25344
rect 1443 25313 1455 25316
rect 1397 25307 1455 25313
rect 1946 25304 1952 25316
rect 2004 25304 2010 25356
rect 2406 25304 2412 25356
rect 2464 25344 2470 25356
rect 2501 25347 2559 25353
rect 2501 25344 2513 25347
rect 2464 25316 2513 25344
rect 2464 25304 2470 25316
rect 2501 25313 2513 25316
rect 2547 25344 2559 25347
rect 5350 25344 5356 25356
rect 2547 25316 5356 25344
rect 2547 25313 2559 25316
rect 2501 25307 2559 25313
rect 5350 25304 5356 25316
rect 5408 25304 5414 25356
rect 1581 25211 1639 25217
rect 1581 25177 1593 25211
rect 1627 25208 1639 25211
rect 2958 25208 2964 25220
rect 1627 25180 2964 25208
rect 1627 25177 1639 25180
rect 1581 25171 1639 25177
rect 2958 25168 2964 25180
rect 3016 25168 3022 25220
rect 2041 25143 2099 25149
rect 2041 25109 2053 25143
rect 2087 25140 2099 25143
rect 2130 25140 2136 25152
rect 2087 25112 2136 25140
rect 2087 25109 2099 25112
rect 2041 25103 2099 25109
rect 2130 25100 2136 25112
rect 2188 25100 2194 25152
rect 2314 25140 2320 25152
rect 2275 25112 2320 25140
rect 2314 25100 2320 25112
rect 2372 25100 2378 25152
rect 2685 25143 2743 25149
rect 2685 25109 2697 25143
rect 2731 25140 2743 25143
rect 2866 25140 2872 25152
rect 2731 25112 2872 25140
rect 2731 25109 2743 25112
rect 2685 25103 2743 25109
rect 2866 25100 2872 25112
rect 2924 25100 2930 25152
rect 3050 25140 3056 25152
rect 3011 25112 3056 25140
rect 3050 25100 3056 25112
rect 3108 25100 3114 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 2406 24936 2412 24948
rect 2367 24908 2412 24936
rect 2406 24896 2412 24908
rect 2464 24896 2470 24948
rect 4062 24828 4068 24880
rect 4120 24868 4126 24880
rect 6178 24868 6184 24880
rect 4120 24840 6184 24868
rect 4120 24828 4126 24840
rect 6178 24828 6184 24840
rect 6236 24828 6242 24880
rect 2038 24800 2044 24812
rect 1412 24772 2044 24800
rect 1412 24741 1440 24772
rect 2038 24760 2044 24772
rect 2096 24760 2102 24812
rect 3237 24803 3295 24809
rect 3237 24769 3249 24803
rect 3283 24800 3295 24803
rect 3283 24772 3372 24800
rect 3283 24769 3295 24772
rect 3237 24763 3295 24769
rect 3344 24744 3372 24772
rect 1397 24735 1455 24741
rect 1397 24701 1409 24735
rect 1443 24701 1455 24735
rect 3050 24732 3056 24744
rect 3011 24704 3056 24732
rect 1397 24695 1455 24701
rect 3050 24692 3056 24704
rect 3108 24692 3114 24744
rect 3326 24692 3332 24744
rect 3384 24692 3390 24744
rect 3602 24732 3608 24744
rect 3563 24704 3608 24732
rect 3602 24692 3608 24704
rect 3660 24692 3666 24744
rect 12342 24692 12348 24744
rect 12400 24732 12406 24744
rect 15933 24735 15991 24741
rect 15933 24732 15945 24735
rect 12400 24704 15945 24732
rect 12400 24692 12406 24704
rect 15933 24701 15945 24704
rect 15979 24732 15991 24735
rect 16485 24735 16543 24741
rect 16485 24732 16497 24735
rect 15979 24704 16497 24732
rect 15979 24701 15991 24704
rect 15933 24695 15991 24701
rect 16485 24701 16497 24704
rect 16531 24701 16543 24735
rect 16485 24695 16543 24701
rect 2961 24667 3019 24673
rect 2961 24633 2973 24667
rect 3007 24664 3019 24667
rect 3007 24636 3188 24664
rect 3007 24633 3019 24636
rect 2961 24627 3019 24633
rect 1394 24556 1400 24608
rect 1452 24596 1458 24608
rect 1581 24599 1639 24605
rect 1581 24596 1593 24599
rect 1452 24568 1593 24596
rect 1452 24556 1458 24568
rect 1581 24565 1593 24568
rect 1627 24565 1639 24599
rect 2590 24596 2596 24608
rect 2551 24568 2596 24596
rect 1581 24559 1639 24565
rect 2590 24556 2596 24568
rect 2648 24556 2654 24608
rect 3160 24596 3188 24636
rect 3418 24596 3424 24608
rect 3160 24568 3424 24596
rect 3418 24556 3424 24568
rect 3476 24596 3482 24608
rect 3620 24596 3648 24692
rect 3476 24568 3648 24596
rect 3476 24556 3482 24568
rect 6914 24556 6920 24608
rect 6972 24596 6978 24608
rect 7469 24599 7527 24605
rect 7469 24596 7481 24599
rect 6972 24568 7481 24596
rect 6972 24556 6978 24568
rect 7469 24565 7481 24568
rect 7515 24596 7527 24599
rect 7834 24596 7840 24608
rect 7515 24568 7840 24596
rect 7515 24565 7527 24568
rect 7469 24559 7527 24565
rect 7834 24556 7840 24568
rect 7892 24556 7898 24608
rect 16114 24596 16120 24608
rect 16075 24568 16120 24596
rect 16114 24556 16120 24568
rect 16172 24556 16178 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1946 24392 1952 24404
rect 1907 24364 1952 24392
rect 1946 24352 1952 24364
rect 2004 24352 2010 24404
rect 2774 24352 2780 24404
rect 2832 24392 2838 24404
rect 2869 24395 2927 24401
rect 2869 24392 2881 24395
rect 2832 24364 2881 24392
rect 2832 24352 2838 24364
rect 2869 24361 2881 24364
rect 2915 24361 2927 24395
rect 2869 24355 2927 24361
rect 4798 24352 4804 24404
rect 4856 24392 4862 24404
rect 5994 24392 6000 24404
rect 4856 24364 6000 24392
rect 4856 24352 4862 24364
rect 5994 24352 6000 24364
rect 6052 24392 6058 24404
rect 6365 24395 6423 24401
rect 6365 24392 6377 24395
rect 6052 24364 6377 24392
rect 6052 24352 6058 24364
rect 6365 24361 6377 24364
rect 6411 24361 6423 24395
rect 7834 24392 7840 24404
rect 7795 24364 7840 24392
rect 6365 24355 6423 24361
rect 7834 24352 7840 24364
rect 7892 24352 7898 24404
rect 14274 24392 14280 24404
rect 14235 24364 14280 24392
rect 14274 24352 14280 24364
rect 14332 24352 14338 24404
rect 15470 24392 15476 24404
rect 15431 24364 15476 24392
rect 15470 24352 15476 24364
rect 15528 24352 15534 24404
rect 16669 24395 16727 24401
rect 16669 24361 16681 24395
rect 16715 24392 16727 24395
rect 18506 24392 18512 24404
rect 16715 24364 18512 24392
rect 16715 24361 16727 24364
rect 16669 24355 16727 24361
rect 18506 24352 18512 24364
rect 18564 24352 18570 24404
rect 18874 24392 18880 24404
rect 18835 24364 18880 24392
rect 18874 24352 18880 24364
rect 18932 24352 18938 24404
rect 21085 24395 21143 24401
rect 21085 24361 21097 24395
rect 21131 24392 21143 24395
rect 22462 24392 22468 24404
rect 21131 24364 22468 24392
rect 21131 24361 21143 24364
rect 21085 24355 21143 24361
rect 22462 24352 22468 24364
rect 22520 24352 22526 24404
rect 6086 24284 6092 24336
rect 6144 24324 6150 24336
rect 6273 24327 6331 24333
rect 6273 24324 6285 24327
rect 6144 24296 6285 24324
rect 6144 24284 6150 24296
rect 6273 24293 6285 24296
rect 6319 24293 6331 24327
rect 6273 24287 6331 24293
rect 1397 24259 1455 24265
rect 1397 24225 1409 24259
rect 1443 24256 1455 24259
rect 2038 24256 2044 24268
rect 1443 24228 2044 24256
rect 1443 24225 1455 24228
rect 1397 24219 1455 24225
rect 2038 24216 2044 24228
rect 2096 24256 2102 24268
rect 2777 24259 2835 24265
rect 2777 24256 2789 24259
rect 2096 24228 2789 24256
rect 2096 24216 2102 24228
rect 2777 24225 2789 24228
rect 2823 24225 2835 24259
rect 2777 24219 2835 24225
rect 3602 24216 3608 24268
rect 3660 24256 3666 24268
rect 4433 24259 4491 24265
rect 4433 24256 4445 24259
rect 3660 24228 4445 24256
rect 3660 24216 3666 24228
rect 4433 24225 4445 24228
rect 4479 24225 4491 24259
rect 4433 24219 4491 24225
rect 11790 24216 11796 24268
rect 11848 24256 11854 24268
rect 12069 24259 12127 24265
rect 12069 24256 12081 24259
rect 11848 24228 12081 24256
rect 11848 24216 11854 24228
rect 12069 24225 12081 24228
rect 12115 24225 12127 24259
rect 12069 24219 12127 24225
rect 13630 24216 13636 24268
rect 13688 24256 13694 24268
rect 14093 24259 14151 24265
rect 14093 24256 14105 24259
rect 13688 24228 14105 24256
rect 13688 24216 13694 24228
rect 14093 24225 14105 24228
rect 14139 24225 14151 24259
rect 15286 24256 15292 24268
rect 15247 24228 15292 24256
rect 14093 24219 14151 24225
rect 15286 24216 15292 24228
rect 15344 24216 15350 24268
rect 16485 24259 16543 24265
rect 16485 24225 16497 24259
rect 16531 24256 16543 24259
rect 16850 24256 16856 24268
rect 16531 24228 16856 24256
rect 16531 24225 16543 24228
rect 16485 24219 16543 24225
rect 16850 24216 16856 24228
rect 16908 24216 16914 24268
rect 17402 24216 17408 24268
rect 17460 24256 17466 24268
rect 17589 24259 17647 24265
rect 17589 24256 17601 24259
rect 17460 24228 17601 24256
rect 17460 24216 17466 24228
rect 17589 24225 17601 24228
rect 17635 24225 17647 24259
rect 17589 24219 17647 24225
rect 18693 24259 18751 24265
rect 18693 24225 18705 24259
rect 18739 24256 18751 24259
rect 18966 24256 18972 24268
rect 18739 24228 18972 24256
rect 18739 24225 18751 24228
rect 18693 24219 18751 24225
rect 18966 24216 18972 24228
rect 19024 24216 19030 24268
rect 20806 24216 20812 24268
rect 20864 24256 20870 24268
rect 20901 24259 20959 24265
rect 20901 24256 20913 24259
rect 20864 24228 20913 24256
rect 20864 24216 20870 24228
rect 20901 24225 20913 24228
rect 20947 24225 20959 24259
rect 20901 24219 20959 24225
rect 3053 24191 3111 24197
rect 3053 24157 3065 24191
rect 3099 24188 3111 24191
rect 3326 24188 3332 24200
rect 3099 24160 3332 24188
rect 3099 24157 3111 24160
rect 3053 24151 3111 24157
rect 3326 24148 3332 24160
rect 3384 24148 3390 24200
rect 4522 24148 4528 24200
rect 4580 24188 4586 24200
rect 4709 24191 4767 24197
rect 4580 24160 4625 24188
rect 4580 24148 4586 24160
rect 4709 24157 4721 24191
rect 4755 24157 4767 24191
rect 4709 24151 4767 24157
rect 6549 24191 6607 24197
rect 6549 24157 6561 24191
rect 6595 24188 6607 24191
rect 7374 24188 7380 24200
rect 6595 24160 7380 24188
rect 6595 24157 6607 24160
rect 6549 24151 6607 24157
rect 2409 24123 2467 24129
rect 2409 24089 2421 24123
rect 2455 24120 2467 24123
rect 2498 24120 2504 24132
rect 2455 24092 2504 24120
rect 2455 24089 2467 24092
rect 2409 24083 2467 24089
rect 2498 24080 2504 24092
rect 2556 24120 2562 24132
rect 3789 24123 3847 24129
rect 3789 24120 3801 24123
rect 2556 24092 3801 24120
rect 2556 24080 2562 24092
rect 3789 24089 3801 24092
rect 3835 24089 3847 24123
rect 4724 24120 4752 24151
rect 7374 24148 7380 24160
rect 7432 24148 7438 24200
rect 7929 24191 7987 24197
rect 7929 24157 7941 24191
rect 7975 24157 7987 24191
rect 8110 24188 8116 24200
rect 8071 24160 8116 24188
rect 7929 24151 7987 24157
rect 5350 24120 5356 24132
rect 3789 24083 3847 24089
rect 3896 24092 5356 24120
rect 1670 24012 1676 24064
rect 1728 24052 1734 24064
rect 2225 24055 2283 24061
rect 2225 24052 2237 24055
rect 1728 24024 2237 24052
rect 1728 24012 1734 24024
rect 2225 24021 2237 24024
rect 2271 24052 2283 24055
rect 2682 24052 2688 24064
rect 2271 24024 2688 24052
rect 2271 24021 2283 24024
rect 2225 24015 2283 24021
rect 2682 24012 2688 24024
rect 2740 24012 2746 24064
rect 3326 24012 3332 24064
rect 3384 24052 3390 24064
rect 3421 24055 3479 24061
rect 3421 24052 3433 24055
rect 3384 24024 3433 24052
rect 3384 24012 3390 24024
rect 3421 24021 3433 24024
rect 3467 24052 3479 24055
rect 3896 24052 3924 24092
rect 5350 24080 5356 24092
rect 5408 24080 5414 24132
rect 5905 24123 5963 24129
rect 5905 24089 5917 24123
rect 5951 24120 5963 24123
rect 7944 24120 7972 24151
rect 8110 24148 8116 24160
rect 8168 24148 8174 24200
rect 9030 24120 9036 24132
rect 5951 24092 9036 24120
rect 5951 24089 5963 24092
rect 5905 24083 5963 24089
rect 9030 24080 9036 24092
rect 9088 24080 9094 24132
rect 12250 24120 12256 24132
rect 12211 24092 12256 24120
rect 12250 24080 12256 24092
rect 12308 24080 12314 24132
rect 17770 24120 17776 24132
rect 17731 24092 17776 24120
rect 17770 24080 17776 24092
rect 17828 24080 17834 24132
rect 4062 24052 4068 24064
rect 3467 24024 3924 24052
rect 4023 24024 4068 24052
rect 3467 24021 3479 24024
rect 3421 24015 3479 24021
rect 4062 24012 4068 24024
rect 4120 24012 4126 24064
rect 5261 24055 5319 24061
rect 5261 24021 5273 24055
rect 5307 24052 5319 24055
rect 5442 24052 5448 24064
rect 5307 24024 5448 24052
rect 5307 24021 5319 24024
rect 5261 24015 5319 24021
rect 5442 24012 5448 24024
rect 5500 24012 5506 24064
rect 6914 24052 6920 24064
rect 6875 24024 6920 24052
rect 6914 24012 6920 24024
rect 6972 24012 6978 24064
rect 7374 24052 7380 24064
rect 7335 24024 7380 24052
rect 7374 24012 7380 24024
rect 7432 24012 7438 24064
rect 7466 24012 7472 24064
rect 7524 24052 7530 24064
rect 7524 24024 7569 24052
rect 7524 24012 7530 24024
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 2038 23848 2044 23860
rect 1999 23820 2044 23848
rect 2038 23808 2044 23820
rect 2096 23808 2102 23860
rect 2133 23851 2191 23857
rect 2133 23817 2145 23851
rect 2179 23848 2191 23851
rect 2314 23848 2320 23860
rect 2179 23820 2320 23848
rect 2179 23817 2191 23820
rect 2133 23811 2191 23817
rect 2314 23808 2320 23820
rect 2372 23808 2378 23860
rect 2774 23808 2780 23860
rect 2832 23848 2838 23860
rect 3142 23848 3148 23860
rect 2832 23820 3148 23848
rect 2832 23808 2838 23820
rect 3142 23808 3148 23820
rect 3200 23808 3206 23860
rect 3234 23808 3240 23860
rect 3292 23848 3298 23860
rect 3602 23848 3608 23860
rect 3292 23820 3608 23848
rect 3292 23808 3298 23820
rect 3602 23808 3608 23820
rect 3660 23808 3666 23860
rect 5350 23808 5356 23860
rect 5408 23848 5414 23860
rect 5445 23851 5503 23857
rect 5445 23848 5457 23851
rect 5408 23820 5457 23848
rect 5408 23808 5414 23820
rect 5445 23817 5457 23820
rect 5491 23817 5503 23851
rect 5994 23848 6000 23860
rect 5955 23820 6000 23848
rect 5445 23811 5503 23817
rect 5994 23808 6000 23820
rect 6052 23808 6058 23860
rect 6086 23808 6092 23860
rect 6144 23848 6150 23860
rect 6270 23848 6276 23860
rect 6144 23820 6276 23848
rect 6144 23808 6150 23820
rect 6270 23808 6276 23820
rect 6328 23848 6334 23860
rect 6365 23851 6423 23857
rect 6365 23848 6377 23851
rect 6328 23820 6377 23848
rect 6328 23808 6334 23820
rect 6365 23817 6377 23820
rect 6411 23817 6423 23851
rect 6365 23811 6423 23817
rect 9030 23808 9036 23860
rect 9088 23848 9094 23860
rect 9125 23851 9183 23857
rect 9125 23848 9137 23851
rect 9088 23820 9137 23848
rect 9088 23808 9094 23820
rect 9125 23817 9137 23820
rect 9171 23817 9183 23851
rect 9125 23811 9183 23817
rect 10321 23851 10379 23857
rect 10321 23817 10333 23851
rect 10367 23848 10379 23851
rect 10778 23848 10784 23860
rect 10367 23820 10784 23848
rect 10367 23817 10379 23820
rect 10321 23811 10379 23817
rect 10778 23808 10784 23820
rect 10836 23808 10842 23860
rect 12618 23848 12624 23860
rect 12579 23820 12624 23848
rect 12618 23808 12624 23820
rect 12676 23808 12682 23860
rect 13081 23851 13139 23857
rect 13081 23817 13093 23851
rect 13127 23848 13139 23851
rect 13354 23848 13360 23860
rect 13127 23820 13360 23848
rect 13127 23817 13139 23820
rect 13081 23811 13139 23817
rect 2682 23712 2688 23724
rect 2643 23684 2688 23712
rect 2682 23672 2688 23684
rect 2740 23672 2746 23724
rect 2498 23644 2504 23656
rect 2459 23616 2504 23644
rect 2498 23604 2504 23616
rect 2556 23604 2562 23656
rect 2590 23604 2596 23656
rect 2648 23644 2654 23656
rect 4065 23647 4123 23653
rect 2648 23616 2693 23644
rect 2648 23604 2654 23616
rect 4065 23613 4077 23647
rect 4111 23644 4123 23647
rect 4154 23644 4160 23656
rect 4111 23616 4160 23644
rect 4111 23613 4123 23616
rect 4065 23607 4123 23613
rect 4154 23604 4160 23616
rect 4212 23604 4218 23656
rect 6362 23604 6368 23656
rect 6420 23644 6426 23656
rect 6825 23647 6883 23653
rect 6825 23644 6837 23647
rect 6420 23616 6837 23644
rect 6420 23604 6426 23616
rect 6825 23613 6837 23616
rect 6871 23644 6883 23647
rect 6914 23644 6920 23656
rect 6871 23616 6920 23644
rect 6871 23613 6883 23616
rect 6825 23607 6883 23613
rect 6914 23604 6920 23616
rect 6972 23604 6978 23656
rect 9858 23604 9864 23656
rect 9916 23644 9922 23656
rect 10137 23647 10195 23653
rect 10137 23644 10149 23647
rect 9916 23616 10149 23644
rect 9916 23604 9922 23616
rect 10137 23613 10149 23616
rect 10183 23644 10195 23647
rect 10689 23647 10747 23653
rect 10689 23644 10701 23647
rect 10183 23616 10701 23644
rect 10183 23613 10195 23616
rect 10137 23607 10195 23613
rect 10689 23613 10701 23616
rect 10735 23613 10747 23647
rect 10689 23607 10747 23613
rect 10778 23604 10784 23656
rect 10836 23644 10842 23656
rect 11241 23647 11299 23653
rect 11241 23644 11253 23647
rect 10836 23616 11253 23644
rect 10836 23604 10842 23616
rect 11241 23613 11253 23616
rect 11287 23644 11299 23647
rect 11793 23647 11851 23653
rect 11793 23644 11805 23647
rect 11287 23616 11805 23644
rect 11287 23613 11299 23616
rect 11241 23607 11299 23613
rect 11793 23613 11805 23616
rect 11839 23613 11851 23647
rect 11793 23607 11851 23613
rect 12437 23647 12495 23653
rect 12437 23613 12449 23647
rect 12483 23644 12495 23647
rect 13096 23644 13124 23811
rect 13354 23808 13360 23820
rect 13412 23808 13418 23860
rect 14461 23851 14519 23857
rect 14461 23817 14473 23851
rect 14507 23848 14519 23851
rect 15654 23848 15660 23860
rect 14507 23820 15660 23848
rect 14507 23817 14519 23820
rect 14461 23811 14519 23817
rect 13998 23780 14004 23792
rect 13959 23752 14004 23780
rect 13998 23740 14004 23752
rect 14056 23740 14062 23792
rect 12483 23616 13124 23644
rect 13817 23647 13875 23653
rect 12483 23613 12495 23616
rect 12437 23607 12495 23613
rect 13817 23613 13829 23647
rect 13863 23644 13875 23647
rect 14476 23644 14504 23811
rect 15654 23808 15660 23820
rect 15712 23808 15718 23860
rect 17034 23848 17040 23860
rect 16995 23820 17040 23848
rect 17034 23808 17040 23820
rect 17092 23808 17098 23860
rect 18230 23848 18236 23860
rect 18191 23820 18236 23848
rect 18230 23808 18236 23820
rect 18288 23808 18294 23860
rect 19613 23851 19671 23857
rect 19613 23817 19625 23851
rect 19659 23848 19671 23851
rect 19702 23848 19708 23860
rect 19659 23820 19708 23848
rect 19659 23817 19671 23820
rect 19613 23811 19671 23817
rect 19702 23808 19708 23820
rect 19760 23808 19766 23860
rect 21358 23848 21364 23860
rect 21319 23820 21364 23848
rect 21358 23808 21364 23820
rect 21416 23808 21422 23860
rect 23845 23851 23903 23857
rect 23845 23817 23857 23851
rect 23891 23848 23903 23851
rect 25314 23848 25320 23860
rect 23891 23820 25320 23848
rect 23891 23817 23903 23820
rect 23845 23811 23903 23817
rect 25314 23808 25320 23820
rect 25372 23808 25378 23860
rect 15102 23780 15108 23792
rect 15063 23752 15108 23780
rect 15102 23740 15108 23752
rect 15160 23740 15166 23792
rect 14921 23647 14979 23653
rect 14921 23644 14933 23647
rect 13863 23616 14504 23644
rect 14752 23616 14933 23644
rect 13863 23613 13875 23616
rect 13817 23607 13875 23613
rect 3970 23576 3976 23588
rect 3931 23548 3976 23576
rect 3970 23536 3976 23548
rect 4028 23536 4034 23588
rect 4332 23579 4390 23585
rect 4332 23545 4344 23579
rect 4378 23576 4390 23579
rect 4890 23576 4896 23588
rect 4378 23548 4896 23576
rect 4378 23545 4390 23548
rect 4332 23539 4390 23545
rect 4890 23536 4896 23548
rect 4948 23536 4954 23588
rect 7092 23579 7150 23585
rect 7092 23545 7104 23579
rect 7138 23576 7150 23579
rect 7374 23576 7380 23588
rect 7138 23548 7380 23576
rect 7138 23545 7150 23548
rect 7092 23539 7150 23545
rect 7374 23536 7380 23548
rect 7432 23536 7438 23588
rect 7558 23536 7564 23588
rect 7616 23576 7622 23588
rect 7926 23576 7932 23588
rect 7616 23548 7932 23576
rect 7616 23536 7622 23548
rect 7926 23536 7932 23548
rect 7984 23536 7990 23588
rect 1673 23511 1731 23517
rect 1673 23477 1685 23511
rect 1719 23508 1731 23511
rect 3326 23508 3332 23520
rect 1719 23480 3332 23508
rect 1719 23477 1731 23480
rect 1673 23471 1731 23477
rect 3326 23468 3332 23480
rect 3384 23468 3390 23520
rect 6822 23468 6828 23520
rect 6880 23508 6886 23520
rect 8110 23508 8116 23520
rect 6880 23480 8116 23508
rect 6880 23468 6886 23480
rect 8110 23468 8116 23480
rect 8168 23508 8174 23520
rect 8205 23511 8263 23517
rect 8205 23508 8217 23511
rect 8168 23480 8217 23508
rect 8168 23468 8174 23480
rect 8205 23477 8217 23480
rect 8251 23508 8263 23511
rect 8757 23511 8815 23517
rect 8757 23508 8769 23511
rect 8251 23480 8769 23508
rect 8251 23477 8263 23480
rect 8205 23471 8263 23477
rect 8757 23477 8769 23480
rect 8803 23477 8815 23511
rect 11422 23508 11428 23520
rect 11383 23480 11428 23508
rect 8757 23471 8815 23477
rect 11422 23468 11428 23480
rect 11480 23468 11486 23520
rect 11790 23468 11796 23520
rect 11848 23508 11854 23520
rect 12161 23511 12219 23517
rect 12161 23508 12173 23511
rect 11848 23480 12173 23508
rect 11848 23468 11854 23480
rect 12161 23477 12173 23480
rect 12207 23477 12219 23511
rect 13630 23508 13636 23520
rect 13591 23480 13636 23508
rect 12161 23471 12219 23477
rect 13630 23468 13636 23480
rect 13688 23468 13694 23520
rect 14550 23468 14556 23520
rect 14608 23508 14614 23520
rect 14752 23517 14780 23616
rect 14921 23613 14933 23616
rect 14967 23613 14979 23647
rect 14921 23607 14979 23613
rect 16853 23647 16911 23653
rect 16853 23613 16865 23647
rect 16899 23613 16911 23647
rect 16853 23607 16911 23613
rect 16868 23576 16896 23607
rect 17402 23604 17408 23656
rect 17460 23644 17466 23656
rect 17773 23647 17831 23653
rect 17773 23644 17785 23647
rect 17460 23616 17785 23644
rect 17460 23604 17466 23616
rect 17773 23613 17785 23616
rect 17819 23613 17831 23647
rect 17773 23607 17831 23613
rect 18049 23647 18107 23653
rect 18049 23613 18061 23647
rect 18095 23644 18107 23647
rect 19426 23644 19432 23656
rect 18095 23616 18644 23644
rect 19387 23616 19432 23644
rect 18095 23613 18107 23616
rect 18049 23607 18107 23613
rect 16868 23548 17540 23576
rect 14737 23511 14795 23517
rect 14737 23508 14749 23511
rect 14608 23480 14749 23508
rect 14608 23468 14614 23480
rect 14737 23477 14749 23480
rect 14783 23477 14795 23511
rect 14737 23471 14795 23477
rect 15286 23468 15292 23520
rect 15344 23508 15350 23520
rect 15473 23511 15531 23517
rect 15473 23508 15485 23511
rect 15344 23480 15485 23508
rect 15344 23468 15350 23480
rect 15473 23477 15485 23480
rect 15519 23477 15531 23511
rect 15473 23471 15531 23477
rect 16577 23511 16635 23517
rect 16577 23477 16589 23511
rect 16623 23508 16635 23511
rect 16850 23508 16856 23520
rect 16623 23480 16856 23508
rect 16623 23477 16635 23480
rect 16577 23471 16635 23477
rect 16850 23468 16856 23480
rect 16908 23468 16914 23520
rect 17512 23517 17540 23548
rect 18616 23520 18644 23616
rect 19426 23604 19432 23616
rect 19484 23644 19490 23656
rect 19981 23647 20039 23653
rect 19981 23644 19993 23647
rect 19484 23616 19993 23644
rect 19484 23604 19490 23616
rect 19981 23613 19993 23616
rect 20027 23613 20039 23647
rect 19981 23607 20039 23613
rect 21082 23604 21088 23656
rect 21140 23644 21146 23656
rect 21177 23647 21235 23653
rect 21177 23644 21189 23647
rect 21140 23616 21189 23644
rect 21140 23604 21146 23616
rect 21177 23613 21189 23616
rect 21223 23644 21235 23647
rect 21729 23647 21787 23653
rect 21729 23644 21741 23647
rect 21223 23616 21741 23644
rect 21223 23613 21235 23616
rect 21177 23607 21235 23613
rect 21729 23613 21741 23616
rect 21775 23613 21787 23647
rect 21729 23607 21787 23613
rect 23474 23604 23480 23656
rect 23532 23644 23538 23656
rect 23661 23647 23719 23653
rect 23661 23644 23673 23647
rect 23532 23616 23673 23644
rect 23532 23604 23538 23616
rect 23661 23613 23673 23616
rect 23707 23644 23719 23647
rect 24213 23647 24271 23653
rect 24213 23644 24225 23647
rect 23707 23616 24225 23644
rect 23707 23613 23719 23616
rect 23661 23607 23719 23613
rect 24213 23613 24225 23616
rect 24259 23613 24271 23647
rect 24213 23607 24271 23613
rect 17497 23511 17555 23517
rect 17497 23477 17509 23511
rect 17543 23508 17555 23511
rect 17586 23508 17592 23520
rect 17543 23480 17592 23508
rect 17543 23477 17555 23480
rect 17497 23471 17555 23477
rect 17586 23468 17592 23480
rect 17644 23468 17650 23520
rect 18598 23508 18604 23520
rect 18559 23480 18604 23508
rect 18598 23468 18604 23480
rect 18656 23468 18662 23520
rect 18966 23508 18972 23520
rect 18927 23480 18972 23508
rect 18966 23468 18972 23480
rect 19024 23468 19030 23520
rect 20806 23468 20812 23520
rect 20864 23508 20870 23520
rect 20901 23511 20959 23517
rect 20901 23508 20913 23511
rect 20864 23480 20913 23508
rect 20864 23468 20870 23480
rect 20901 23477 20913 23480
rect 20947 23477 20959 23511
rect 20901 23471 20959 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 2133 23307 2191 23313
rect 2133 23273 2145 23307
rect 2179 23304 2191 23307
rect 2314 23304 2320 23316
rect 2179 23276 2320 23304
rect 2179 23273 2191 23276
rect 2133 23267 2191 23273
rect 2314 23264 2320 23276
rect 2372 23264 2378 23316
rect 2774 23264 2780 23316
rect 2832 23304 2838 23316
rect 3145 23307 3203 23313
rect 3145 23304 3157 23307
rect 2832 23276 3157 23304
rect 2832 23264 2838 23276
rect 3145 23273 3157 23276
rect 3191 23273 3203 23307
rect 3145 23267 3203 23273
rect 3970 23264 3976 23316
rect 4028 23304 4034 23316
rect 5258 23304 5264 23316
rect 4028 23276 5264 23304
rect 4028 23264 4034 23276
rect 5258 23264 5264 23276
rect 5316 23264 5322 23316
rect 9858 23304 9864 23316
rect 9819 23276 9864 23304
rect 9858 23264 9864 23276
rect 9916 23264 9922 23316
rect 12713 23307 12771 23313
rect 12713 23273 12725 23307
rect 12759 23304 12771 23307
rect 13630 23304 13636 23316
rect 12759 23276 13636 23304
rect 12759 23273 12771 23276
rect 12713 23267 12771 23273
rect 13630 23264 13636 23276
rect 13688 23264 13694 23316
rect 14093 23307 14151 23313
rect 14093 23273 14105 23307
rect 14139 23304 14151 23307
rect 14826 23304 14832 23316
rect 14139 23276 14832 23304
rect 14139 23273 14151 23276
rect 14093 23267 14151 23273
rect 14826 23264 14832 23276
rect 14884 23264 14890 23316
rect 17218 23304 17224 23316
rect 17179 23276 17224 23304
rect 17218 23264 17224 23276
rect 17276 23264 17282 23316
rect 18325 23307 18383 23313
rect 18325 23273 18337 23307
rect 18371 23304 18383 23307
rect 18966 23304 18972 23316
rect 18371 23276 18972 23304
rect 18371 23273 18383 23276
rect 18325 23267 18383 23273
rect 18966 23264 18972 23276
rect 19024 23264 19030 23316
rect 21082 23304 21088 23316
rect 21043 23276 21088 23304
rect 21082 23264 21088 23276
rect 21140 23264 21146 23316
rect 22373 23307 22431 23313
rect 22373 23273 22385 23307
rect 22419 23304 22431 23307
rect 23474 23304 23480 23316
rect 22419 23276 23480 23304
rect 22419 23273 22431 23276
rect 22373 23267 22431 23273
rect 23474 23264 23480 23276
rect 23532 23264 23538 23316
rect 2222 23196 2228 23248
rect 2280 23236 2286 23248
rect 2590 23236 2596 23248
rect 2280 23208 2596 23236
rect 2280 23196 2286 23208
rect 2590 23196 2596 23208
rect 2648 23196 2654 23248
rect 3602 23196 3608 23248
rect 3660 23236 3666 23248
rect 4154 23236 4160 23248
rect 3660 23208 4160 23236
rect 3660 23196 3666 23208
rect 4154 23196 4160 23208
rect 4212 23236 4218 23248
rect 4341 23239 4399 23245
rect 4341 23236 4353 23239
rect 4212 23208 4353 23236
rect 4212 23196 4218 23208
rect 4341 23205 4353 23208
rect 4387 23236 4399 23239
rect 6362 23236 6368 23248
rect 4387 23208 6368 23236
rect 4387 23205 4399 23208
rect 4341 23199 4399 23205
rect 6362 23196 6368 23208
rect 6420 23196 6426 23248
rect 6632 23239 6690 23245
rect 6632 23205 6644 23239
rect 6678 23236 6690 23239
rect 6822 23236 6828 23248
rect 6678 23208 6828 23236
rect 6678 23205 6690 23208
rect 6632 23199 6690 23205
rect 6822 23196 6828 23208
rect 6880 23196 6886 23248
rect 5166 23168 5172 23180
rect 5127 23140 5172 23168
rect 5166 23128 5172 23140
rect 5224 23128 5230 23180
rect 5997 23171 6055 23177
rect 5997 23137 6009 23171
rect 6043 23168 6055 23171
rect 7374 23168 7380 23180
rect 6043 23140 7380 23168
rect 6043 23137 6055 23140
rect 5997 23131 6055 23137
rect 7374 23128 7380 23140
rect 7432 23128 7438 23180
rect 9677 23171 9735 23177
rect 9677 23137 9689 23171
rect 9723 23168 9735 23171
rect 9766 23168 9772 23180
rect 9723 23140 9772 23168
rect 9723 23137 9735 23140
rect 9677 23131 9735 23137
rect 9766 23128 9772 23140
rect 9824 23128 9830 23180
rect 12158 23128 12164 23180
rect 12216 23168 12222 23180
rect 12529 23171 12587 23177
rect 12529 23168 12541 23171
rect 12216 23140 12541 23168
rect 12216 23128 12222 23140
rect 12529 23137 12541 23140
rect 12575 23137 12587 23171
rect 12529 23131 12587 23137
rect 15289 23171 15347 23177
rect 15289 23137 15301 23171
rect 15335 23168 15347 23171
rect 15378 23168 15384 23180
rect 15335 23140 15384 23168
rect 15335 23137 15347 23140
rect 15289 23131 15347 23137
rect 15378 23128 15384 23140
rect 15436 23128 15442 23180
rect 17034 23168 17040 23180
rect 16995 23140 17040 23168
rect 17034 23128 17040 23140
rect 17092 23128 17098 23180
rect 18141 23171 18199 23177
rect 18141 23137 18153 23171
rect 18187 23168 18199 23171
rect 18230 23168 18236 23180
rect 18187 23140 18236 23168
rect 18187 23137 18199 23140
rect 18141 23131 18199 23137
rect 18230 23128 18236 23140
rect 18288 23128 18294 23180
rect 20898 23168 20904 23180
rect 20859 23140 20904 23168
rect 20898 23128 20904 23140
rect 20956 23128 20962 23180
rect 22186 23168 22192 23180
rect 22147 23140 22192 23168
rect 22186 23128 22192 23140
rect 22244 23128 22250 23180
rect 2038 23060 2044 23112
rect 2096 23100 2102 23112
rect 2225 23103 2283 23109
rect 2225 23100 2237 23103
rect 2096 23072 2237 23100
rect 2096 23060 2102 23072
rect 2225 23069 2237 23072
rect 2271 23069 2283 23103
rect 2225 23063 2283 23069
rect 2409 23103 2467 23109
rect 2409 23069 2421 23103
rect 2455 23100 2467 23103
rect 2682 23100 2688 23112
rect 2455 23072 2688 23100
rect 2455 23069 2467 23072
rect 2409 23063 2467 23069
rect 1673 23035 1731 23041
rect 1673 23001 1685 23035
rect 1719 23032 1731 23035
rect 2424 23032 2452 23063
rect 2682 23060 2688 23072
rect 2740 23060 2746 23112
rect 4154 23060 4160 23112
rect 4212 23100 4218 23112
rect 4430 23100 4436 23112
rect 4212 23072 4436 23100
rect 4212 23060 4218 23072
rect 4430 23060 4436 23072
rect 4488 23060 4494 23112
rect 5445 23103 5503 23109
rect 5445 23069 5457 23103
rect 5491 23069 5503 23103
rect 6362 23100 6368 23112
rect 6323 23072 6368 23100
rect 5445 23063 5503 23069
rect 1719 23004 2452 23032
rect 4709 23035 4767 23041
rect 1719 23001 1731 23004
rect 1673 22995 1731 23001
rect 4709 23001 4721 23035
rect 4755 23032 4767 23035
rect 4890 23032 4896 23044
rect 4755 23004 4896 23032
rect 4755 23001 4767 23004
rect 4709 22995 4767 23001
rect 4890 22992 4896 23004
rect 4948 23032 4954 23044
rect 5460 23032 5488 23063
rect 6362 23060 6368 23072
rect 6420 23060 6426 23112
rect 13538 23100 13544 23112
rect 13499 23072 13544 23100
rect 13538 23060 13544 23072
rect 13596 23060 13602 23112
rect 4948 23004 6040 23032
rect 4948 22992 4954 23004
rect 1765 22967 1823 22973
rect 1765 22933 1777 22967
rect 1811 22964 1823 22967
rect 1854 22964 1860 22976
rect 1811 22936 1860 22964
rect 1811 22933 1823 22936
rect 1765 22927 1823 22933
rect 1854 22924 1860 22936
rect 1912 22924 1918 22976
rect 2866 22964 2872 22976
rect 2827 22936 2872 22964
rect 2866 22924 2872 22936
rect 2924 22964 2930 22976
rect 3326 22964 3332 22976
rect 2924 22936 3332 22964
rect 2924 22924 2930 22936
rect 3326 22924 3332 22936
rect 3384 22964 3390 22976
rect 3789 22967 3847 22973
rect 3789 22964 3801 22967
rect 3384 22936 3801 22964
rect 3384 22924 3390 22936
rect 3789 22933 3801 22936
rect 3835 22933 3847 22967
rect 4798 22964 4804 22976
rect 4759 22936 4804 22964
rect 3789 22927 3847 22933
rect 4798 22924 4804 22936
rect 4856 22924 4862 22976
rect 6012 22964 6040 23004
rect 7745 22967 7803 22973
rect 7745 22964 7757 22967
rect 6012 22936 7757 22964
rect 7745 22933 7757 22936
rect 7791 22933 7803 22967
rect 8478 22964 8484 22976
rect 8439 22936 8484 22964
rect 7745 22927 7803 22933
rect 8478 22924 8484 22936
rect 8536 22924 8542 22976
rect 14458 22964 14464 22976
rect 14419 22936 14464 22964
rect 14458 22924 14464 22936
rect 14516 22924 14522 22976
rect 15470 22964 15476 22976
rect 15431 22936 15476 22964
rect 15470 22924 15476 22936
rect 15528 22924 15534 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 2041 22763 2099 22769
rect 2041 22729 2053 22763
rect 2087 22760 2099 22763
rect 2130 22760 2136 22772
rect 2087 22732 2136 22760
rect 2087 22729 2099 22732
rect 2041 22723 2099 22729
rect 1397 22559 1455 22565
rect 1397 22525 1409 22559
rect 1443 22556 1455 22559
rect 2056 22556 2084 22723
rect 2130 22720 2136 22732
rect 2188 22720 2194 22772
rect 2593 22763 2651 22769
rect 2593 22729 2605 22763
rect 2639 22760 2651 22763
rect 3602 22760 3608 22772
rect 2639 22732 3608 22760
rect 2639 22729 2651 22732
rect 2593 22723 2651 22729
rect 2222 22584 2228 22636
rect 2280 22624 2286 22636
rect 2700 22633 2728 22732
rect 3602 22720 3608 22732
rect 3660 22720 3666 22772
rect 4890 22760 4896 22772
rect 4851 22732 4896 22760
rect 4890 22720 4896 22732
rect 4948 22720 4954 22772
rect 6178 22760 6184 22772
rect 6139 22732 6184 22760
rect 6178 22720 6184 22732
rect 6236 22720 6242 22772
rect 6362 22720 6368 22772
rect 6420 22760 6426 22772
rect 7466 22760 7472 22772
rect 6420 22732 7472 22760
rect 6420 22720 6426 22732
rect 7466 22720 7472 22732
rect 7524 22720 7530 22772
rect 15749 22763 15807 22769
rect 15749 22729 15761 22763
rect 15795 22760 15807 22763
rect 16390 22760 16396 22772
rect 15795 22732 16396 22760
rect 15795 22729 15807 22732
rect 15749 22723 15807 22729
rect 16390 22720 16396 22732
rect 16448 22720 16454 22772
rect 16850 22760 16856 22772
rect 16811 22732 16856 22760
rect 16850 22720 16856 22732
rect 16908 22720 16914 22772
rect 17034 22720 17040 22772
rect 17092 22760 17098 22772
rect 17129 22763 17187 22769
rect 17129 22760 17141 22763
rect 17092 22732 17141 22760
rect 17092 22720 17098 22732
rect 17129 22729 17141 22732
rect 17175 22729 17187 22763
rect 20898 22760 20904 22772
rect 20859 22732 20904 22760
rect 17129 22723 17187 22729
rect 20898 22720 20904 22732
rect 20956 22720 20962 22772
rect 6825 22695 6883 22701
rect 6825 22692 6837 22695
rect 5644 22664 6837 22692
rect 5644 22636 5672 22664
rect 6825 22661 6837 22664
rect 6871 22661 6883 22695
rect 8386 22692 8392 22704
rect 8347 22664 8392 22692
rect 6825 22655 6883 22661
rect 8386 22652 8392 22664
rect 8444 22652 8450 22704
rect 12894 22692 12900 22704
rect 12855 22664 12900 22692
rect 12894 22652 12900 22664
rect 12952 22652 12958 22704
rect 2685 22627 2743 22633
rect 2685 22624 2697 22627
rect 2280 22596 2697 22624
rect 2280 22584 2286 22596
rect 2685 22593 2697 22596
rect 2731 22593 2743 22627
rect 5626 22624 5632 22636
rect 5539 22596 5632 22624
rect 2685 22587 2743 22593
rect 5626 22584 5632 22596
rect 5684 22584 5690 22636
rect 5813 22627 5871 22633
rect 5813 22593 5825 22627
rect 5859 22593 5871 22627
rect 5813 22587 5871 22593
rect 1443 22528 2084 22556
rect 2952 22559 3010 22565
rect 1443 22525 1455 22528
rect 1397 22519 1455 22525
rect 2952 22525 2964 22559
rect 2998 22525 3010 22559
rect 5534 22556 5540 22568
rect 5495 22528 5540 22556
rect 2952 22519 3010 22525
rect 1578 22420 1584 22432
rect 1539 22392 1584 22420
rect 1578 22380 1584 22392
rect 1636 22380 1642 22432
rect 2866 22380 2872 22432
rect 2924 22420 2930 22432
rect 2967 22420 2995 22519
rect 5534 22516 5540 22528
rect 5592 22516 5598 22568
rect 5828 22556 5856 22587
rect 7374 22584 7380 22636
rect 7432 22624 7438 22636
rect 7469 22627 7527 22633
rect 7469 22624 7481 22627
rect 7432 22596 7481 22624
rect 7432 22584 7438 22596
rect 7469 22593 7481 22596
rect 7515 22624 7527 22627
rect 8478 22624 8484 22636
rect 7515 22596 8484 22624
rect 7515 22593 7527 22596
rect 7469 22587 7527 22593
rect 8478 22584 8484 22596
rect 8536 22624 8542 22636
rect 8941 22627 8999 22633
rect 8941 22624 8953 22627
rect 8536 22596 8953 22624
rect 8536 22584 8542 22596
rect 8941 22593 8953 22596
rect 8987 22593 8999 22627
rect 8941 22587 8999 22593
rect 14458 22584 14464 22636
rect 14516 22624 14522 22636
rect 14553 22627 14611 22633
rect 14553 22624 14565 22627
rect 14516 22596 14565 22624
rect 14516 22584 14522 22596
rect 14553 22593 14565 22596
rect 14599 22593 14611 22627
rect 14553 22587 14611 22593
rect 6822 22556 6828 22568
rect 5828 22528 6828 22556
rect 6822 22516 6828 22528
rect 6880 22516 6886 22568
rect 12158 22556 12164 22568
rect 12119 22528 12164 22556
rect 12158 22516 12164 22528
rect 12216 22516 12222 22568
rect 12713 22559 12771 22565
rect 12713 22525 12725 22559
rect 12759 22556 12771 22559
rect 12894 22556 12900 22568
rect 12759 22528 12900 22556
rect 12759 22525 12771 22528
rect 12713 22519 12771 22525
rect 12894 22516 12900 22528
rect 12952 22556 12958 22568
rect 13265 22559 13323 22565
rect 13265 22556 13277 22559
rect 12952 22528 13277 22556
rect 12952 22516 12958 22528
rect 13265 22525 13277 22528
rect 13311 22525 13323 22559
rect 13265 22519 13323 22525
rect 15470 22516 15476 22568
rect 15528 22556 15534 22568
rect 15565 22559 15623 22565
rect 15565 22556 15577 22559
rect 15528 22528 15577 22556
rect 15528 22516 15534 22528
rect 15565 22525 15577 22528
rect 15611 22556 15623 22559
rect 16117 22559 16175 22565
rect 16117 22556 16129 22559
rect 15611 22528 16129 22556
rect 15611 22525 15623 22528
rect 15565 22519 15623 22525
rect 16117 22525 16129 22528
rect 16163 22525 16175 22559
rect 16117 22519 16175 22525
rect 16669 22559 16727 22565
rect 16669 22525 16681 22559
rect 16715 22556 16727 22559
rect 16715 22528 17632 22556
rect 16715 22525 16727 22528
rect 16669 22519 16727 22525
rect 6362 22448 6368 22500
rect 6420 22488 6426 22500
rect 6549 22491 6607 22497
rect 6549 22488 6561 22491
rect 6420 22460 6561 22488
rect 6420 22448 6426 22460
rect 6549 22457 6561 22460
rect 6595 22488 6607 22491
rect 7285 22491 7343 22497
rect 7285 22488 7297 22491
rect 6595 22460 7297 22488
rect 6595 22457 6607 22460
rect 6549 22451 6607 22457
rect 7285 22457 7297 22460
rect 7331 22457 7343 22491
rect 8849 22491 8907 22497
rect 8849 22488 8861 22491
rect 7285 22451 7343 22457
rect 8220 22460 8861 22488
rect 2924 22392 2995 22420
rect 2924 22380 2930 22392
rect 3786 22380 3792 22432
rect 3844 22420 3850 22432
rect 4065 22423 4123 22429
rect 4065 22420 4077 22423
rect 3844 22392 4077 22420
rect 3844 22380 3850 22392
rect 4065 22389 4077 22392
rect 4111 22389 4123 22423
rect 5166 22420 5172 22432
rect 5127 22392 5172 22420
rect 4065 22383 4123 22389
rect 5166 22380 5172 22392
rect 5224 22380 5230 22432
rect 6178 22380 6184 22432
rect 6236 22420 6242 22432
rect 7193 22423 7251 22429
rect 7193 22420 7205 22423
rect 6236 22392 7205 22420
rect 6236 22380 6242 22392
rect 7193 22389 7205 22392
rect 7239 22389 7251 22423
rect 7193 22383 7251 22389
rect 7466 22380 7472 22432
rect 7524 22420 7530 22432
rect 7837 22423 7895 22429
rect 7837 22420 7849 22423
rect 7524 22392 7849 22420
rect 7524 22380 7530 22392
rect 7837 22389 7849 22392
rect 7883 22389 7895 22423
rect 7837 22383 7895 22389
rect 8110 22380 8116 22432
rect 8168 22420 8174 22432
rect 8220 22429 8248 22460
rect 8849 22457 8861 22460
rect 8895 22457 8907 22491
rect 8849 22451 8907 22457
rect 13909 22491 13967 22497
rect 13909 22457 13921 22491
rect 13955 22488 13967 22491
rect 14369 22491 14427 22497
rect 14369 22488 14381 22491
rect 13955 22460 14381 22488
rect 13955 22457 13967 22460
rect 13909 22451 13967 22457
rect 14369 22457 14381 22460
rect 14415 22488 14427 22491
rect 14550 22488 14556 22500
rect 14415 22460 14556 22488
rect 14415 22457 14427 22460
rect 14369 22451 14427 22457
rect 14550 22448 14556 22460
rect 14608 22488 14614 22500
rect 14826 22488 14832 22500
rect 14608 22460 14832 22488
rect 14608 22448 14614 22460
rect 14826 22448 14832 22460
rect 14884 22448 14890 22500
rect 17604 22497 17632 22528
rect 19334 22516 19340 22568
rect 19392 22556 19398 22568
rect 22186 22556 22192 22568
rect 19392 22528 22192 22556
rect 19392 22516 19398 22528
rect 22186 22516 22192 22528
rect 22244 22516 22250 22568
rect 17589 22491 17647 22497
rect 17589 22457 17601 22491
rect 17635 22488 17647 22491
rect 18506 22488 18512 22500
rect 17635 22460 18512 22488
rect 17635 22457 17647 22460
rect 17589 22451 17647 22457
rect 18506 22448 18512 22460
rect 18564 22448 18570 22500
rect 8205 22423 8263 22429
rect 8205 22420 8217 22423
rect 8168 22392 8217 22420
rect 8168 22380 8174 22392
rect 8205 22389 8217 22392
rect 8251 22389 8263 22423
rect 8205 22383 8263 22389
rect 8478 22380 8484 22432
rect 8536 22420 8542 22432
rect 8757 22423 8815 22429
rect 8757 22420 8769 22423
rect 8536 22392 8769 22420
rect 8536 22380 8542 22392
rect 8757 22389 8769 22392
rect 8803 22389 8815 22423
rect 9766 22420 9772 22432
rect 9727 22392 9772 22420
rect 8757 22383 8815 22389
rect 9766 22380 9772 22392
rect 9824 22380 9830 22432
rect 9858 22380 9864 22432
rect 9916 22420 9922 22432
rect 9953 22423 10011 22429
rect 9953 22420 9965 22423
rect 9916 22392 9965 22420
rect 9916 22380 9922 22392
rect 9953 22389 9965 22392
rect 9999 22389 10011 22423
rect 13998 22420 14004 22432
rect 13959 22392 14004 22420
rect 9953 22383 10011 22389
rect 13998 22380 14004 22392
rect 14056 22380 14062 22432
rect 14461 22423 14519 22429
rect 14461 22389 14473 22423
rect 14507 22420 14519 22423
rect 14734 22420 14740 22432
rect 14507 22392 14740 22420
rect 14507 22389 14519 22392
rect 14461 22383 14519 22389
rect 14734 22380 14740 22392
rect 14792 22380 14798 22432
rect 15378 22420 15384 22432
rect 15339 22392 15384 22420
rect 15378 22380 15384 22392
rect 15436 22380 15442 22432
rect 18230 22420 18236 22432
rect 18191 22392 18236 22420
rect 18230 22380 18236 22392
rect 18288 22380 18294 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1946 22176 1952 22228
rect 2004 22216 2010 22228
rect 4065 22219 4123 22225
rect 4065 22216 4077 22219
rect 2004 22188 4077 22216
rect 2004 22176 2010 22188
rect 4065 22185 4077 22188
rect 4111 22185 4123 22219
rect 5166 22216 5172 22228
rect 4065 22179 4123 22185
rect 4264 22188 5172 22216
rect 2222 22148 2228 22160
rect 1412 22120 2228 22148
rect 1412 22089 1440 22120
rect 2222 22108 2228 22120
rect 2280 22108 2286 22160
rect 4264 22148 4292 22188
rect 5166 22176 5172 22188
rect 5224 22176 5230 22228
rect 5626 22216 5632 22228
rect 5587 22188 5632 22216
rect 5626 22176 5632 22188
rect 5684 22176 5690 22228
rect 6273 22219 6331 22225
rect 6273 22185 6285 22219
rect 6319 22216 6331 22219
rect 6822 22216 6828 22228
rect 6319 22188 6828 22216
rect 6319 22185 6331 22188
rect 6273 22179 6331 22185
rect 4430 22148 4436 22160
rect 4080 22120 4292 22148
rect 4391 22120 4436 22148
rect 1670 22089 1676 22092
rect 1397 22083 1455 22089
rect 1397 22049 1409 22083
rect 1443 22049 1455 22083
rect 1664 22080 1676 22089
rect 1631 22052 1676 22080
rect 1397 22043 1455 22049
rect 1664 22043 1676 22052
rect 1670 22040 1676 22043
rect 1728 22040 1734 22092
rect 2406 22040 2412 22092
rect 2464 22040 2470 22092
rect 3881 22083 3939 22089
rect 3881 22049 3893 22083
rect 3927 22080 3939 22083
rect 3970 22080 3976 22092
rect 3927 22052 3976 22080
rect 3927 22049 3939 22052
rect 3881 22043 3939 22049
rect 3970 22040 3976 22052
rect 4028 22040 4034 22092
rect 4080 22080 4108 22120
rect 4430 22108 4436 22120
rect 4488 22148 4494 22160
rect 5534 22148 5540 22160
rect 4488 22120 5540 22148
rect 4488 22108 4494 22120
rect 5534 22108 5540 22120
rect 5592 22108 5598 22160
rect 4522 22080 4528 22092
rect 4080 22052 4200 22080
rect 4483 22052 4528 22080
rect 1762 21836 1768 21888
rect 1820 21876 1826 21888
rect 2424 21876 2452 22040
rect 2682 21904 2688 21956
rect 2740 21944 2746 21956
rect 2777 21947 2835 21953
rect 2777 21944 2789 21947
rect 2740 21916 2789 21944
rect 2740 21904 2746 21916
rect 2777 21913 2789 21916
rect 2823 21913 2835 21947
rect 2777 21907 2835 21913
rect 1820 21848 2452 21876
rect 3513 21879 3571 21885
rect 1820 21836 1826 21848
rect 3513 21845 3525 21879
rect 3559 21876 3571 21879
rect 4172 21876 4200 22052
rect 4522 22040 4528 22052
rect 4580 22040 4586 22092
rect 5261 22083 5319 22089
rect 5261 22049 5273 22083
rect 5307 22080 5319 22083
rect 6288 22080 6316 22179
rect 6822 22176 6828 22188
rect 6880 22176 6886 22228
rect 7929 22219 7987 22225
rect 7929 22185 7941 22219
rect 7975 22216 7987 22219
rect 8478 22216 8484 22228
rect 7975 22188 8484 22216
rect 7975 22185 7987 22188
rect 7929 22179 7987 22185
rect 8478 22176 8484 22188
rect 8536 22176 8542 22228
rect 13814 22216 13820 22228
rect 13727 22188 13820 22216
rect 13814 22176 13820 22188
rect 13872 22216 13878 22228
rect 13998 22216 14004 22228
rect 13872 22188 14004 22216
rect 13872 22176 13878 22188
rect 13998 22176 14004 22188
rect 14056 22176 14062 22228
rect 14366 22176 14372 22228
rect 14424 22216 14430 22228
rect 14734 22216 14740 22228
rect 14424 22188 14740 22216
rect 14424 22176 14430 22188
rect 14734 22176 14740 22188
rect 14792 22176 14798 22228
rect 5307 22052 6316 22080
rect 5307 22049 5319 22052
rect 5261 22043 5319 22049
rect 6638 22040 6644 22092
rect 6696 22080 6702 22092
rect 6733 22083 6791 22089
rect 6733 22080 6745 22083
rect 6696 22052 6745 22080
rect 6696 22040 6702 22052
rect 6733 22049 6745 22052
rect 6779 22049 6791 22083
rect 6733 22043 6791 22049
rect 6822 22040 6828 22092
rect 6880 22080 6886 22092
rect 8754 22080 8760 22092
rect 6880 22052 8760 22080
rect 6880 22040 6886 22052
rect 8754 22040 8760 22052
rect 8812 22040 8818 22092
rect 10870 22080 10876 22092
rect 10831 22052 10876 22080
rect 10870 22040 10876 22052
rect 10928 22040 10934 22092
rect 13262 22040 13268 22092
rect 13320 22080 13326 22092
rect 13725 22083 13783 22089
rect 13725 22080 13737 22083
rect 13320 22052 13737 22080
rect 13320 22040 13326 22052
rect 13725 22049 13737 22052
rect 13771 22049 13783 22083
rect 13725 22043 13783 22049
rect 14458 22040 14464 22092
rect 14516 22080 14522 22092
rect 15562 22089 15568 22092
rect 15545 22083 15568 22089
rect 15545 22080 15557 22083
rect 14516 22052 15557 22080
rect 14516 22040 14522 22052
rect 15545 22049 15557 22052
rect 15620 22080 15626 22092
rect 15620 22052 15693 22080
rect 15545 22043 15568 22049
rect 15562 22040 15568 22043
rect 15620 22040 15626 22052
rect 4614 22012 4620 22024
rect 4575 21984 4620 22012
rect 4614 21972 4620 21984
rect 4672 21972 4678 22024
rect 7009 22015 7067 22021
rect 7009 21981 7021 22015
rect 7055 22012 7067 22015
rect 10962 22012 10968 22024
rect 7055 21984 7420 22012
rect 10923 21984 10968 22012
rect 7055 21981 7067 21984
rect 7009 21975 7067 21981
rect 6365 21947 6423 21953
rect 6365 21913 6377 21947
rect 6411 21944 6423 21947
rect 6730 21944 6736 21956
rect 6411 21916 6736 21944
rect 6411 21913 6423 21916
rect 6365 21907 6423 21913
rect 6730 21904 6736 21916
rect 6788 21904 6794 21956
rect 7392 21888 7420 21984
rect 10962 21972 10968 21984
rect 11020 21972 11026 22024
rect 11054 21972 11060 22024
rect 11112 22012 11118 22024
rect 11149 22015 11207 22021
rect 11149 22012 11161 22015
rect 11112 21984 11161 22012
rect 11112 21972 11118 21984
rect 11149 21981 11161 21984
rect 11195 21981 11207 22015
rect 11149 21975 11207 21981
rect 13630 21972 13636 22024
rect 13688 22012 13694 22024
rect 13909 22015 13967 22021
rect 13909 22012 13921 22015
rect 13688 21984 13921 22012
rect 13688 21972 13694 21984
rect 13909 21981 13921 21984
rect 13955 21981 13967 22015
rect 13909 21975 13967 21981
rect 14090 21972 14096 22024
rect 14148 22012 14154 22024
rect 15289 22015 15347 22021
rect 15289 22012 15301 22015
rect 14148 21984 15301 22012
rect 14148 21972 14154 21984
rect 15289 21981 15301 21984
rect 15335 21981 15347 22015
rect 15289 21975 15347 21981
rect 9674 21904 9680 21956
rect 9732 21944 9738 21956
rect 10505 21947 10563 21953
rect 10505 21944 10517 21947
rect 9732 21916 10517 21944
rect 9732 21904 9738 21916
rect 10505 21913 10517 21916
rect 10551 21913 10563 21947
rect 10505 21907 10563 21913
rect 12529 21947 12587 21953
rect 12529 21913 12541 21947
rect 12575 21944 12587 21947
rect 13722 21944 13728 21956
rect 12575 21916 13728 21944
rect 12575 21913 12587 21916
rect 12529 21907 12587 21913
rect 13722 21904 13728 21916
rect 13780 21904 13786 21956
rect 16666 21944 16672 21956
rect 16627 21916 16672 21944
rect 16666 21904 16672 21916
rect 16724 21904 16730 21956
rect 7374 21876 7380 21888
rect 3559 21848 4200 21876
rect 7335 21848 7380 21876
rect 3559 21845 3571 21848
rect 3513 21839 3571 21845
rect 7374 21836 7380 21848
rect 7432 21836 7438 21888
rect 7650 21836 7656 21888
rect 7708 21876 7714 21888
rect 7745 21879 7803 21885
rect 7745 21876 7757 21879
rect 7708 21848 7757 21876
rect 7708 21836 7714 21848
rect 7745 21845 7757 21848
rect 7791 21845 7803 21879
rect 7745 21839 7803 21845
rect 9033 21879 9091 21885
rect 9033 21845 9045 21879
rect 9079 21876 9091 21879
rect 9490 21876 9496 21888
rect 9079 21848 9496 21876
rect 9079 21845 9091 21848
rect 9033 21839 9091 21845
rect 9490 21836 9496 21848
rect 9548 21876 9554 21888
rect 10321 21879 10379 21885
rect 10321 21876 10333 21879
rect 9548 21848 10333 21876
rect 9548 21836 9554 21848
rect 10321 21845 10333 21848
rect 10367 21876 10379 21879
rect 11054 21876 11060 21888
rect 10367 21848 11060 21876
rect 10367 21845 10379 21848
rect 10321 21839 10379 21845
rect 11054 21836 11060 21848
rect 11112 21836 11118 21888
rect 11146 21836 11152 21888
rect 11204 21876 11210 21888
rect 11517 21879 11575 21885
rect 11517 21876 11529 21879
rect 11204 21848 11529 21876
rect 11204 21836 11210 21848
rect 11517 21845 11529 21848
rect 11563 21845 11575 21879
rect 13262 21876 13268 21888
rect 13223 21848 13268 21876
rect 11517 21839 11575 21845
rect 13262 21836 13268 21848
rect 13320 21836 13326 21888
rect 13354 21836 13360 21888
rect 13412 21876 13418 21888
rect 14461 21879 14519 21885
rect 13412 21848 13457 21876
rect 13412 21836 13418 21848
rect 14461 21845 14473 21879
rect 14507 21876 14519 21879
rect 14550 21876 14556 21888
rect 14507 21848 14556 21876
rect 14507 21845 14519 21848
rect 14461 21839 14519 21845
rect 14550 21836 14556 21848
rect 14608 21836 14614 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 4706 21672 4712 21684
rect 4667 21644 4712 21672
rect 4706 21632 4712 21644
rect 4764 21632 4770 21684
rect 6457 21675 6515 21681
rect 6457 21641 6469 21675
rect 6503 21672 6515 21675
rect 6822 21672 6828 21684
rect 6503 21644 6828 21672
rect 6503 21641 6515 21644
rect 6457 21635 6515 21641
rect 6822 21632 6828 21644
rect 6880 21632 6886 21684
rect 10597 21675 10655 21681
rect 10597 21641 10609 21675
rect 10643 21672 10655 21675
rect 10870 21672 10876 21684
rect 10643 21644 10876 21672
rect 10643 21641 10655 21644
rect 10597 21635 10655 21641
rect 10870 21632 10876 21644
rect 10928 21632 10934 21684
rect 13541 21675 13599 21681
rect 13541 21641 13553 21675
rect 13587 21672 13599 21675
rect 13630 21672 13636 21684
rect 13587 21644 13636 21672
rect 13587 21641 13599 21644
rect 13541 21635 13599 21641
rect 13630 21632 13636 21644
rect 13688 21632 13694 21684
rect 15562 21672 15568 21684
rect 15523 21644 15568 21672
rect 15562 21632 15568 21644
rect 15620 21632 15626 21684
rect 10229 21607 10287 21613
rect 10229 21573 10241 21607
rect 10275 21604 10287 21607
rect 10962 21604 10968 21616
rect 10275 21576 10968 21604
rect 10275 21573 10287 21576
rect 10229 21567 10287 21573
rect 10962 21564 10968 21576
rect 11020 21564 11026 21616
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21536 1731 21539
rect 2133 21539 2191 21545
rect 2133 21536 2145 21539
rect 1719 21508 2145 21536
rect 1719 21505 1731 21508
rect 1673 21499 1731 21505
rect 2133 21505 2145 21508
rect 2179 21536 2191 21539
rect 2222 21536 2228 21548
rect 2179 21508 2228 21536
rect 2179 21505 2191 21508
rect 2133 21499 2191 21505
rect 2222 21496 2228 21508
rect 2280 21496 2286 21548
rect 5166 21496 5172 21548
rect 5224 21536 5230 21548
rect 5445 21539 5503 21545
rect 5445 21536 5457 21539
rect 5224 21508 5457 21536
rect 5224 21496 5230 21508
rect 5445 21505 5457 21508
rect 5491 21505 5503 21539
rect 5445 21499 5503 21505
rect 7653 21539 7711 21545
rect 7653 21505 7665 21539
rect 7699 21536 7711 21539
rect 8021 21539 8079 21545
rect 8021 21536 8033 21539
rect 7699 21508 8033 21536
rect 7699 21505 7711 21508
rect 7653 21499 7711 21505
rect 8021 21505 8033 21508
rect 8067 21536 8079 21539
rect 8202 21536 8208 21548
rect 8067 21508 8208 21536
rect 8067 21505 8079 21508
rect 8021 21499 8079 21505
rect 8202 21496 8208 21508
rect 8260 21496 8266 21548
rect 9490 21536 9496 21548
rect 9451 21508 9496 21536
rect 9490 21496 9496 21508
rect 9548 21496 9554 21548
rect 11422 21536 11428 21548
rect 11383 21508 11428 21536
rect 11422 21496 11428 21508
rect 11480 21496 11486 21548
rect 12986 21536 12992 21548
rect 12947 21508 12992 21536
rect 12986 21496 12992 21508
rect 13044 21496 13050 21548
rect 4433 21471 4491 21477
rect 4433 21437 4445 21471
rect 4479 21468 4491 21471
rect 5261 21471 5319 21477
rect 5261 21468 5273 21471
rect 4479 21440 5273 21468
rect 4479 21437 4491 21440
rect 4433 21431 4491 21437
rect 5261 21437 5273 21440
rect 5307 21468 5319 21471
rect 5350 21468 5356 21480
rect 5307 21440 5356 21468
rect 5307 21437 5319 21440
rect 5261 21431 5319 21437
rect 5350 21428 5356 21440
rect 5408 21428 5414 21480
rect 8110 21468 8116 21480
rect 5920 21440 8116 21468
rect 2314 21360 2320 21412
rect 2372 21400 2378 21412
rect 2470 21403 2528 21409
rect 2470 21400 2482 21403
rect 2372 21372 2482 21400
rect 2372 21360 2378 21372
rect 2470 21369 2482 21372
rect 2516 21400 2528 21403
rect 2682 21400 2688 21412
rect 2516 21372 2688 21400
rect 2516 21369 2528 21372
rect 2470 21363 2528 21369
rect 2682 21360 2688 21372
rect 2740 21360 2746 21412
rect 4706 21360 4712 21412
rect 4764 21400 4770 21412
rect 5920 21400 5948 21440
rect 8110 21428 8116 21440
rect 8168 21428 8174 21480
rect 11238 21468 11244 21480
rect 11151 21440 11244 21468
rect 11238 21428 11244 21440
rect 11296 21468 11302 21480
rect 11793 21471 11851 21477
rect 11793 21468 11805 21471
rect 11296 21440 11805 21468
rect 11296 21428 11302 21440
rect 11793 21437 11805 21440
rect 11839 21437 11851 21471
rect 14185 21471 14243 21477
rect 14185 21468 14197 21471
rect 11793 21431 11851 21437
rect 14108 21440 14197 21468
rect 4764 21372 5948 21400
rect 4764 21360 4770 21372
rect 3602 21332 3608 21344
rect 3563 21304 3608 21332
rect 3602 21292 3608 21304
rect 3660 21292 3666 21344
rect 4893 21335 4951 21341
rect 4893 21301 4905 21335
rect 4939 21332 4951 21335
rect 4982 21332 4988 21344
rect 4939 21304 4988 21332
rect 4939 21301 4951 21304
rect 4893 21295 4951 21301
rect 4982 21292 4988 21304
rect 5040 21292 5046 21344
rect 5368 21341 5396 21372
rect 5994 21360 6000 21412
rect 6052 21400 6058 21412
rect 6089 21403 6147 21409
rect 6089 21400 6101 21403
rect 6052 21372 6101 21400
rect 6052 21360 6058 21372
rect 6089 21369 6101 21372
rect 6135 21400 6147 21403
rect 6638 21400 6644 21412
rect 6135 21372 6644 21400
rect 6135 21369 6147 21372
rect 6089 21363 6147 21369
rect 6638 21360 6644 21372
rect 6696 21400 6702 21412
rect 6822 21400 6828 21412
rect 6696 21372 6828 21400
rect 6696 21360 6702 21372
rect 6822 21360 6828 21372
rect 6880 21360 6886 21412
rect 7377 21403 7435 21409
rect 7377 21369 7389 21403
rect 7423 21400 7435 21403
rect 7558 21400 7564 21412
rect 7423 21372 7564 21400
rect 7423 21369 7435 21372
rect 7377 21363 7435 21369
rect 7558 21360 7564 21372
rect 7616 21400 7622 21412
rect 8389 21403 8447 21409
rect 8389 21400 8401 21403
rect 7616 21372 8401 21400
rect 7616 21360 7622 21372
rect 8389 21369 8401 21372
rect 8435 21369 8447 21403
rect 8846 21400 8852 21412
rect 8759 21372 8852 21400
rect 8389 21363 8447 21369
rect 8846 21360 8852 21372
rect 8904 21400 8910 21412
rect 9401 21403 9459 21409
rect 9401 21400 9413 21403
rect 8904 21372 9413 21400
rect 8904 21360 8910 21372
rect 9401 21369 9413 21372
rect 9447 21369 9459 21403
rect 9401 21363 9459 21369
rect 12253 21403 12311 21409
rect 12253 21369 12265 21403
rect 12299 21400 12311 21403
rect 12805 21403 12863 21409
rect 12805 21400 12817 21403
rect 12299 21372 12817 21400
rect 12299 21369 12311 21372
rect 12253 21363 12311 21369
rect 12805 21369 12817 21372
rect 12851 21400 12863 21403
rect 13078 21400 13084 21412
rect 12851 21372 13084 21400
rect 12851 21369 12863 21372
rect 12805 21363 12863 21369
rect 13078 21360 13084 21372
rect 13136 21360 13142 21412
rect 14108 21344 14136 21440
rect 14185 21437 14197 21440
rect 14231 21468 14243 21471
rect 16117 21471 16175 21477
rect 16117 21468 16129 21471
rect 14231 21440 16129 21468
rect 14231 21437 14243 21440
rect 14185 21431 14243 21437
rect 16117 21437 16129 21440
rect 16163 21437 16175 21471
rect 16117 21431 16175 21437
rect 14452 21403 14510 21409
rect 14452 21369 14464 21403
rect 14498 21400 14510 21403
rect 14550 21400 14556 21412
rect 14498 21372 14556 21400
rect 14498 21369 14510 21372
rect 14452 21363 14510 21369
rect 14550 21360 14556 21372
rect 14608 21360 14614 21412
rect 5353 21335 5411 21341
rect 5353 21301 5365 21335
rect 5399 21301 5411 21335
rect 7006 21332 7012 21344
rect 6967 21304 7012 21332
rect 5353 21295 5411 21301
rect 7006 21292 7012 21304
rect 7064 21292 7070 21344
rect 7469 21335 7527 21341
rect 7469 21301 7481 21335
rect 7515 21332 7527 21335
rect 7650 21332 7656 21344
rect 7515 21304 7656 21332
rect 7515 21301 7527 21304
rect 7469 21295 7527 21301
rect 7650 21292 7656 21304
rect 7708 21292 7714 21344
rect 8938 21332 8944 21344
rect 8899 21304 8944 21332
rect 8938 21292 8944 21304
rect 8996 21292 9002 21344
rect 9030 21292 9036 21344
rect 9088 21332 9094 21344
rect 9309 21335 9367 21341
rect 9309 21332 9321 21335
rect 9088 21304 9321 21332
rect 9088 21292 9094 21304
rect 9309 21301 9321 21304
rect 9355 21301 9367 21335
rect 9309 21295 9367 21301
rect 10781 21335 10839 21341
rect 10781 21301 10793 21335
rect 10827 21332 10839 21335
rect 10962 21332 10968 21344
rect 10827 21304 10968 21332
rect 10827 21301 10839 21304
rect 10781 21295 10839 21301
rect 10962 21292 10968 21304
rect 11020 21292 11026 21344
rect 11146 21332 11152 21344
rect 11107 21304 11152 21332
rect 11146 21292 11152 21304
rect 11204 21292 11210 21344
rect 12158 21292 12164 21344
rect 12216 21332 12222 21344
rect 12437 21335 12495 21341
rect 12437 21332 12449 21335
rect 12216 21304 12449 21332
rect 12216 21292 12222 21304
rect 12437 21301 12449 21304
rect 12483 21301 12495 21335
rect 12437 21295 12495 21301
rect 12897 21335 12955 21341
rect 12897 21301 12909 21335
rect 12943 21332 12955 21335
rect 13630 21332 13636 21344
rect 12943 21304 13636 21332
rect 12943 21301 12955 21304
rect 12897 21295 12955 21301
rect 13630 21292 13636 21304
rect 13688 21292 13694 21344
rect 14090 21332 14096 21344
rect 14051 21304 14096 21332
rect 14090 21292 14096 21304
rect 14148 21292 14154 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 2314 21128 2320 21140
rect 2275 21100 2320 21128
rect 2314 21088 2320 21100
rect 2372 21088 2378 21140
rect 2409 21131 2467 21137
rect 2409 21097 2421 21131
rect 2455 21128 2467 21131
rect 3513 21131 3571 21137
rect 3513 21128 3525 21131
rect 2455 21100 3525 21128
rect 2455 21097 2467 21100
rect 2409 21091 2467 21097
rect 3513 21097 3525 21100
rect 3559 21128 3571 21131
rect 4522 21128 4528 21140
rect 3559 21100 4528 21128
rect 3559 21097 3571 21100
rect 3513 21091 3571 21097
rect 4522 21088 4528 21100
rect 4580 21088 4586 21140
rect 5534 21088 5540 21140
rect 5592 21128 5598 21140
rect 5721 21131 5779 21137
rect 5721 21128 5733 21131
rect 5592 21100 5733 21128
rect 5592 21088 5598 21100
rect 5721 21097 5733 21100
rect 5767 21097 5779 21131
rect 5721 21091 5779 21097
rect 5905 21131 5963 21137
rect 5905 21097 5917 21131
rect 5951 21097 5963 21131
rect 5905 21091 5963 21097
rect 2866 21060 2872 21072
rect 2827 21032 2872 21060
rect 2866 21020 2872 21032
rect 2924 21020 2930 21072
rect 3786 21060 3792 21072
rect 3747 21032 3792 21060
rect 3786 21020 3792 21032
rect 3844 21020 3850 21072
rect 4801 21063 4859 21069
rect 4801 21029 4813 21063
rect 4847 21060 4859 21063
rect 5920 21060 5948 21091
rect 6178 21088 6184 21140
rect 6236 21128 6242 21140
rect 6273 21131 6331 21137
rect 6273 21128 6285 21131
rect 6236 21100 6285 21128
rect 6236 21088 6242 21100
rect 6273 21097 6285 21100
rect 6319 21097 6331 21131
rect 6273 21091 6331 21097
rect 7469 21131 7527 21137
rect 7469 21097 7481 21131
rect 7515 21128 7527 21131
rect 7558 21128 7564 21140
rect 7515 21100 7564 21128
rect 7515 21097 7527 21100
rect 7469 21091 7527 21097
rect 7558 21088 7564 21100
rect 7616 21088 7622 21140
rect 7834 21128 7840 21140
rect 7795 21100 7840 21128
rect 7834 21088 7840 21100
rect 7892 21088 7898 21140
rect 9030 21128 9036 21140
rect 8991 21100 9036 21128
rect 9030 21088 9036 21100
rect 9088 21088 9094 21140
rect 11422 21088 11428 21140
rect 11480 21128 11486 21140
rect 11609 21131 11667 21137
rect 11609 21128 11621 21131
rect 11480 21100 11621 21128
rect 11480 21088 11486 21100
rect 11609 21097 11621 21100
rect 11655 21128 11667 21131
rect 12713 21131 12771 21137
rect 12713 21128 12725 21131
rect 11655 21100 12725 21128
rect 11655 21097 11667 21100
rect 11609 21091 11667 21097
rect 12713 21097 12725 21100
rect 12759 21128 12771 21131
rect 12986 21128 12992 21140
rect 12759 21100 12992 21128
rect 12759 21097 12771 21100
rect 12713 21091 12771 21097
rect 12986 21088 12992 21100
rect 13044 21088 13050 21140
rect 13262 21088 13268 21140
rect 13320 21128 13326 21140
rect 13541 21131 13599 21137
rect 13541 21128 13553 21131
rect 13320 21100 13553 21128
rect 13320 21088 13326 21100
rect 13541 21097 13553 21100
rect 13587 21097 13599 21131
rect 15562 21128 15568 21140
rect 15523 21100 15568 21128
rect 13541 21091 13599 21097
rect 15562 21088 15568 21100
rect 15620 21088 15626 21140
rect 5994 21060 6000 21072
rect 4847 21032 6000 21060
rect 4847 21029 4859 21032
rect 4801 21023 4859 21029
rect 5994 21020 6000 21032
rect 6052 21020 6058 21072
rect 7377 21063 7435 21069
rect 7377 21029 7389 21063
rect 7423 21060 7435 21063
rect 7852 21060 7880 21088
rect 7423 21032 7880 21060
rect 7423 21029 7435 21032
rect 7377 21023 7435 21029
rect 9490 21020 9496 21072
rect 9548 21060 9554 21072
rect 9922 21063 9980 21069
rect 9922 21060 9934 21063
rect 9548 21032 9934 21060
rect 9548 21020 9554 21032
rect 9922 21029 9934 21032
rect 9968 21029 9980 21063
rect 9922 21023 9980 21029
rect 13449 21063 13507 21069
rect 13449 21029 13461 21063
rect 13495 21060 13507 21063
rect 13722 21060 13728 21072
rect 13495 21032 13728 21060
rect 13495 21029 13507 21032
rect 13449 21023 13507 21029
rect 13722 21020 13728 21032
rect 13780 21020 13786 21072
rect 13998 21020 14004 21072
rect 14056 21020 14062 21072
rect 1394 20992 1400 21004
rect 1355 20964 1400 20992
rect 1394 20952 1400 20964
rect 1452 20952 1458 21004
rect 2774 20952 2780 21004
rect 2832 20992 2838 21004
rect 4709 20995 4767 21001
rect 2832 20964 2877 20992
rect 2832 20952 2838 20964
rect 4709 20961 4721 20995
rect 4755 20992 4767 20995
rect 4982 20992 4988 21004
rect 4755 20964 4988 20992
rect 4755 20961 4767 20964
rect 4709 20955 4767 20961
rect 4982 20952 4988 20964
rect 5040 20992 5046 21004
rect 5442 20992 5448 21004
rect 5040 20964 5448 20992
rect 5040 20952 5046 20964
rect 5442 20952 5448 20964
rect 5500 20952 5506 21004
rect 12153 20995 12211 21001
rect 12153 20992 12165 20995
rect 12084 20964 12165 20992
rect 2958 20924 2964 20936
rect 2919 20896 2964 20924
rect 2958 20884 2964 20896
rect 3016 20884 3022 20936
rect 3602 20884 3608 20936
rect 3660 20924 3666 20936
rect 4890 20924 4896 20936
rect 3660 20896 4660 20924
rect 4851 20896 4896 20924
rect 3660 20884 3666 20896
rect 1670 20816 1676 20868
rect 1728 20856 1734 20868
rect 1949 20859 2007 20865
rect 1949 20856 1961 20859
rect 1728 20828 1961 20856
rect 1728 20816 1734 20828
rect 1949 20825 1961 20828
rect 1995 20856 2007 20859
rect 3786 20856 3792 20868
rect 1995 20828 3792 20856
rect 1995 20825 2007 20828
rect 1949 20819 2007 20825
rect 3786 20816 3792 20828
rect 3844 20816 3850 20868
rect 1578 20788 1584 20800
rect 1539 20760 1584 20788
rect 1578 20748 1584 20760
rect 1636 20748 1642 20800
rect 4154 20748 4160 20800
rect 4212 20788 4218 20800
rect 4341 20791 4399 20797
rect 4341 20788 4353 20791
rect 4212 20760 4353 20788
rect 4212 20748 4218 20760
rect 4341 20757 4353 20760
rect 4387 20757 4399 20791
rect 4632 20788 4660 20896
rect 4890 20884 4896 20896
rect 4948 20884 4954 20936
rect 6362 20924 6368 20936
rect 6323 20896 6368 20924
rect 6362 20884 6368 20896
rect 6420 20884 6426 20936
rect 6457 20927 6515 20933
rect 6457 20893 6469 20927
rect 6503 20893 6515 20927
rect 6457 20887 6515 20893
rect 6086 20856 6092 20868
rect 5552 20828 6092 20856
rect 5552 20800 5580 20828
rect 6086 20816 6092 20828
rect 6144 20856 6150 20868
rect 6472 20856 6500 20887
rect 7190 20884 7196 20936
rect 7248 20924 7254 20936
rect 7929 20927 7987 20933
rect 7929 20924 7941 20927
rect 7248 20896 7941 20924
rect 7248 20884 7254 20896
rect 7929 20893 7941 20896
rect 7975 20893 7987 20927
rect 7929 20887 7987 20893
rect 8113 20927 8171 20933
rect 8113 20893 8125 20927
rect 8159 20924 8171 20927
rect 9677 20927 9735 20933
rect 8159 20896 8432 20924
rect 8159 20893 8171 20896
rect 8113 20887 8171 20893
rect 6144 20828 6500 20856
rect 6144 20816 6150 20828
rect 8404 20800 8432 20896
rect 9677 20893 9689 20927
rect 9723 20893 9735 20927
rect 12084 20924 12112 20964
rect 12153 20961 12165 20964
rect 12199 20961 12211 20995
rect 12153 20955 12211 20961
rect 13081 20995 13139 21001
rect 13081 20961 13093 20995
rect 13127 20992 13139 20995
rect 13354 20992 13360 21004
rect 13127 20964 13360 20992
rect 13127 20961 13139 20964
rect 13081 20955 13139 20961
rect 13096 20924 13124 20955
rect 13354 20952 13360 20964
rect 13412 20952 13418 21004
rect 13909 20995 13967 21001
rect 13909 20961 13921 20995
rect 13955 20992 13967 20995
rect 14016 20992 14044 21020
rect 14734 20992 14740 21004
rect 13955 20964 14740 20992
rect 13955 20961 13967 20964
rect 13909 20955 13967 20961
rect 14734 20952 14740 20964
rect 14792 20952 14798 21004
rect 13998 20924 14004 20936
rect 12084 20896 13124 20924
rect 13959 20896 14004 20924
rect 9677 20887 9735 20893
rect 5166 20788 5172 20800
rect 4632 20760 5172 20788
rect 4341 20751 4399 20757
rect 5166 20748 5172 20760
rect 5224 20788 5230 20800
rect 5353 20791 5411 20797
rect 5353 20788 5365 20791
rect 5224 20760 5365 20788
rect 5224 20748 5230 20760
rect 5353 20757 5365 20760
rect 5399 20788 5411 20791
rect 5534 20788 5540 20800
rect 5399 20760 5540 20788
rect 5399 20757 5411 20760
rect 5353 20751 5411 20757
rect 5534 20748 5540 20760
rect 5592 20748 5598 20800
rect 7009 20791 7067 20797
rect 7009 20757 7021 20791
rect 7055 20788 7067 20791
rect 7374 20788 7380 20800
rect 7055 20760 7380 20788
rect 7055 20757 7067 20760
rect 7009 20751 7067 20757
rect 7374 20748 7380 20760
rect 7432 20788 7438 20800
rect 8110 20788 8116 20800
rect 7432 20760 8116 20788
rect 7432 20748 7438 20760
rect 8110 20748 8116 20760
rect 8168 20748 8174 20800
rect 8386 20748 8392 20800
rect 8444 20788 8450 20800
rect 8481 20791 8539 20797
rect 8481 20788 8493 20791
rect 8444 20760 8493 20788
rect 8444 20748 8450 20760
rect 8481 20757 8493 20760
rect 8527 20757 8539 20791
rect 9692 20788 9720 20887
rect 13998 20884 14004 20896
rect 14056 20884 14062 20936
rect 14185 20927 14243 20933
rect 14185 20893 14197 20927
rect 14231 20924 14243 20927
rect 14458 20924 14464 20936
rect 14231 20896 14464 20924
rect 14231 20893 14243 20896
rect 14185 20887 14243 20893
rect 14458 20884 14464 20896
rect 14516 20884 14522 20936
rect 9858 20788 9864 20800
rect 9692 20760 9864 20788
rect 8481 20751 8539 20757
rect 9858 20748 9864 20760
rect 9916 20748 9922 20800
rect 10870 20748 10876 20800
rect 10928 20788 10934 20800
rect 11057 20791 11115 20797
rect 11057 20788 11069 20791
rect 10928 20760 11069 20788
rect 10928 20748 10934 20760
rect 11057 20757 11069 20760
rect 11103 20757 11115 20791
rect 12342 20788 12348 20800
rect 12303 20760 12348 20788
rect 11057 20751 11115 20757
rect 12342 20748 12348 20760
rect 12400 20748 12406 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 2133 20587 2191 20593
rect 2133 20553 2145 20587
rect 2179 20584 2191 20587
rect 2958 20584 2964 20596
rect 2179 20556 2964 20584
rect 2179 20553 2191 20556
rect 2133 20547 2191 20553
rect 2958 20544 2964 20556
rect 3016 20544 3022 20596
rect 5534 20584 5540 20596
rect 5495 20556 5540 20584
rect 5534 20544 5540 20556
rect 5592 20544 5598 20596
rect 6178 20544 6184 20596
rect 6236 20584 6242 20596
rect 6273 20587 6331 20593
rect 6273 20584 6285 20587
rect 6236 20556 6285 20584
rect 6236 20544 6242 20556
rect 6273 20553 6285 20556
rect 6319 20584 6331 20587
rect 7190 20584 7196 20596
rect 6319 20556 7196 20584
rect 6319 20553 6331 20556
rect 6273 20547 6331 20553
rect 7190 20544 7196 20556
rect 7248 20544 7254 20596
rect 8294 20544 8300 20596
rect 8352 20584 8358 20596
rect 8757 20587 8815 20593
rect 8757 20584 8769 20587
rect 8352 20556 8769 20584
rect 8352 20544 8358 20556
rect 8757 20553 8769 20556
rect 8803 20584 8815 20587
rect 9309 20587 9367 20593
rect 9309 20584 9321 20587
rect 8803 20556 9321 20584
rect 8803 20553 8815 20556
rect 8757 20547 8815 20553
rect 9309 20553 9321 20556
rect 9355 20553 9367 20587
rect 9309 20547 9367 20553
rect 9324 20448 9352 20547
rect 11054 20544 11060 20596
rect 11112 20584 11118 20596
rect 11241 20587 11299 20593
rect 11241 20584 11253 20587
rect 11112 20556 11253 20584
rect 11112 20544 11118 20556
rect 11241 20553 11253 20556
rect 11287 20553 11299 20587
rect 11241 20547 11299 20553
rect 13998 20544 14004 20596
rect 14056 20584 14062 20596
rect 14369 20587 14427 20593
rect 14369 20584 14381 20587
rect 14056 20556 14381 20584
rect 14056 20544 14062 20556
rect 14369 20553 14381 20556
rect 14415 20553 14427 20587
rect 14734 20584 14740 20596
rect 14695 20556 14740 20584
rect 14369 20547 14427 20553
rect 14734 20544 14740 20556
rect 14792 20544 14798 20596
rect 15197 20587 15255 20593
rect 15197 20553 15209 20587
rect 15243 20584 15255 20587
rect 15562 20584 15568 20596
rect 15243 20556 15568 20584
rect 15243 20553 15255 20556
rect 15197 20547 15255 20553
rect 15562 20544 15568 20556
rect 15620 20544 15626 20596
rect 9324 20420 9996 20448
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20380 1455 20383
rect 2406 20380 2412 20392
rect 1443 20352 2412 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 2406 20340 2412 20352
rect 2464 20340 2470 20392
rect 2501 20383 2559 20389
rect 2501 20349 2513 20383
rect 2547 20380 2559 20383
rect 2682 20380 2688 20392
rect 2547 20352 2688 20380
rect 2547 20349 2559 20352
rect 2501 20343 2559 20349
rect 2682 20340 2688 20352
rect 2740 20340 2746 20392
rect 3329 20383 3387 20389
rect 3329 20349 3341 20383
rect 3375 20380 3387 20383
rect 3421 20383 3479 20389
rect 3421 20380 3433 20383
rect 3375 20352 3433 20380
rect 3375 20349 3387 20352
rect 3329 20343 3387 20349
rect 3421 20349 3433 20352
rect 3467 20380 3479 20383
rect 4062 20380 4068 20392
rect 3467 20352 4068 20380
rect 3467 20349 3479 20352
rect 3421 20343 3479 20349
rect 4062 20340 4068 20352
rect 4120 20380 4126 20392
rect 7374 20380 7380 20392
rect 4120 20352 7380 20380
rect 4120 20340 4126 20352
rect 7374 20340 7380 20352
rect 7432 20340 7438 20392
rect 9861 20383 9919 20389
rect 9861 20349 9873 20383
rect 9907 20349 9919 20383
rect 9968 20380 9996 20420
rect 10117 20383 10175 20389
rect 10117 20380 10129 20383
rect 9968 20352 10129 20380
rect 9861 20343 9919 20349
rect 10117 20349 10129 20352
rect 10163 20349 10175 20383
rect 10117 20343 10175 20349
rect 12437 20383 12495 20389
rect 12437 20349 12449 20383
rect 12483 20349 12495 20383
rect 12437 20343 12495 20349
rect 2866 20312 2872 20324
rect 2827 20284 2872 20312
rect 2866 20272 2872 20284
rect 2924 20272 2930 20324
rect 3602 20272 3608 20324
rect 3660 20321 3666 20324
rect 3660 20315 3724 20321
rect 3660 20281 3678 20315
rect 3712 20281 3724 20315
rect 3660 20275 3724 20281
rect 7644 20315 7702 20321
rect 7644 20281 7656 20315
rect 7690 20312 7702 20315
rect 8386 20312 8392 20324
rect 7690 20284 8392 20312
rect 7690 20281 7702 20284
rect 7644 20275 7702 20281
rect 3660 20272 3666 20275
rect 8386 20272 8392 20284
rect 8444 20272 8450 20324
rect 9876 20256 9904 20343
rect 12253 20315 12311 20321
rect 12253 20281 12265 20315
rect 12299 20312 12311 20315
rect 12452 20312 12480 20343
rect 12526 20340 12532 20392
rect 12584 20380 12590 20392
rect 12704 20383 12762 20389
rect 12704 20380 12716 20383
rect 12584 20352 12716 20380
rect 12584 20340 12590 20352
rect 12704 20349 12716 20352
rect 12750 20380 12762 20383
rect 12986 20380 12992 20392
rect 12750 20352 12992 20380
rect 12750 20349 12762 20352
rect 12704 20343 12762 20349
rect 12986 20340 12992 20352
rect 13044 20340 13050 20392
rect 12299 20284 12756 20312
rect 12299 20281 12311 20284
rect 12253 20275 12311 20281
rect 12728 20256 12756 20284
rect 1394 20204 1400 20256
rect 1452 20244 1458 20256
rect 1581 20247 1639 20253
rect 1581 20244 1593 20247
rect 1452 20216 1593 20244
rect 1452 20204 1458 20216
rect 1581 20213 1593 20216
rect 1627 20213 1639 20247
rect 1581 20207 1639 20213
rect 2958 20204 2964 20256
rect 3016 20244 3022 20256
rect 3234 20244 3240 20256
rect 3016 20216 3240 20244
rect 3016 20204 3022 20216
rect 3234 20204 3240 20216
rect 3292 20204 3298 20256
rect 3786 20204 3792 20256
rect 3844 20244 3850 20256
rect 4430 20244 4436 20256
rect 3844 20216 4436 20244
rect 3844 20204 3850 20216
rect 4430 20204 4436 20216
rect 4488 20244 4494 20256
rect 4801 20247 4859 20253
rect 4801 20244 4813 20247
rect 4488 20216 4813 20244
rect 4488 20204 4494 20216
rect 4801 20213 4813 20216
rect 4847 20244 4859 20247
rect 4890 20244 4896 20256
rect 4847 20216 4896 20244
rect 4847 20213 4859 20216
rect 4801 20207 4859 20213
rect 4890 20204 4896 20216
rect 4948 20204 4954 20256
rect 5997 20247 6055 20253
rect 5997 20213 6009 20247
rect 6043 20244 6055 20247
rect 6178 20244 6184 20256
rect 6043 20216 6184 20244
rect 6043 20213 6055 20216
rect 5997 20207 6055 20213
rect 6178 20204 6184 20216
rect 6236 20244 6242 20256
rect 6362 20244 6368 20256
rect 6236 20216 6368 20244
rect 6236 20204 6242 20216
rect 6362 20204 6368 20216
rect 6420 20204 6426 20256
rect 9769 20247 9827 20253
rect 9769 20213 9781 20247
rect 9815 20244 9827 20247
rect 9858 20244 9864 20256
rect 9815 20216 9864 20244
rect 9815 20213 9827 20216
rect 9769 20207 9827 20213
rect 9858 20204 9864 20216
rect 9916 20204 9922 20256
rect 11882 20244 11888 20256
rect 11843 20216 11888 20244
rect 11882 20204 11888 20216
rect 11940 20204 11946 20256
rect 12710 20204 12716 20256
rect 12768 20204 12774 20256
rect 13538 20204 13544 20256
rect 13596 20244 13602 20256
rect 13817 20247 13875 20253
rect 13817 20244 13829 20247
rect 13596 20216 13829 20244
rect 13596 20204 13602 20216
rect 13817 20213 13829 20216
rect 13863 20213 13875 20247
rect 13817 20207 13875 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1946 20040 1952 20052
rect 1907 20012 1952 20040
rect 1946 20000 1952 20012
rect 2004 20000 2010 20052
rect 2406 20040 2412 20052
rect 2367 20012 2412 20040
rect 2406 20000 2412 20012
rect 2464 20000 2470 20052
rect 3513 20043 3571 20049
rect 3513 20009 3525 20043
rect 3559 20040 3571 20043
rect 3602 20040 3608 20052
rect 3559 20012 3608 20040
rect 3559 20009 3571 20012
rect 3513 20003 3571 20009
rect 3602 20000 3608 20012
rect 3660 20000 3666 20052
rect 5994 20040 6000 20052
rect 5955 20012 6000 20040
rect 5994 20000 6000 20012
rect 6052 20000 6058 20052
rect 6914 20040 6920 20052
rect 6875 20012 6920 20040
rect 6914 20000 6920 20012
rect 6972 20000 6978 20052
rect 8573 20043 8631 20049
rect 8573 20009 8585 20043
rect 8619 20040 8631 20043
rect 9030 20040 9036 20052
rect 8619 20012 9036 20040
rect 8619 20009 8631 20012
rect 8573 20003 8631 20009
rect 9030 20000 9036 20012
rect 9088 20000 9094 20052
rect 9309 20043 9367 20049
rect 9309 20009 9321 20043
rect 9355 20040 9367 20043
rect 9674 20040 9680 20052
rect 9355 20012 9680 20040
rect 9355 20009 9367 20012
rect 9309 20003 9367 20009
rect 9674 20000 9680 20012
rect 9732 20000 9738 20052
rect 10321 20043 10379 20049
rect 10321 20009 10333 20043
rect 10367 20040 10379 20043
rect 11054 20040 11060 20052
rect 10367 20012 11060 20040
rect 10367 20009 10379 20012
rect 10321 20003 10379 20009
rect 11054 20000 11060 20012
rect 11112 20000 11118 20052
rect 11882 20000 11888 20052
rect 11940 20040 11946 20052
rect 12986 20040 12992 20052
rect 11940 20012 12992 20040
rect 11940 20000 11946 20012
rect 12986 20000 12992 20012
rect 13044 20040 13050 20052
rect 13541 20043 13599 20049
rect 13541 20040 13553 20043
rect 13044 20012 13553 20040
rect 13044 20000 13050 20012
rect 13541 20009 13553 20012
rect 13587 20009 13599 20043
rect 13541 20003 13599 20009
rect 4332 19975 4390 19981
rect 4332 19941 4344 19975
rect 4378 19972 4390 19975
rect 4430 19972 4436 19984
rect 4378 19944 4436 19972
rect 4378 19941 4390 19944
rect 4332 19935 4390 19941
rect 4430 19932 4436 19944
rect 4488 19932 4494 19984
rect 10772 19975 10830 19981
rect 10772 19941 10784 19975
rect 10818 19972 10830 19975
rect 10870 19972 10876 19984
rect 10818 19944 10876 19972
rect 10818 19941 10830 19944
rect 10772 19935 10830 19941
rect 10870 19932 10876 19944
rect 10928 19932 10934 19984
rect 12526 19972 12532 19984
rect 12487 19944 12532 19972
rect 12526 19932 12532 19944
rect 12584 19932 12590 19984
rect 14734 19932 14740 19984
rect 14792 19972 14798 19984
rect 15286 19972 15292 19984
rect 14792 19944 15292 19972
rect 14792 19932 14798 19944
rect 15286 19932 15292 19944
rect 15344 19932 15350 19984
rect 1397 19907 1455 19913
rect 1397 19873 1409 19907
rect 1443 19904 1455 19907
rect 2314 19904 2320 19916
rect 1443 19876 2320 19904
rect 1443 19873 1455 19876
rect 1397 19867 1455 19873
rect 2314 19864 2320 19876
rect 2372 19864 2378 19916
rect 2501 19907 2559 19913
rect 2501 19873 2513 19907
rect 2547 19904 2559 19907
rect 2547 19876 3096 19904
rect 2547 19873 2559 19876
rect 2501 19867 2559 19873
rect 2332 19768 2360 19864
rect 3068 19780 3096 19876
rect 4062 19864 4068 19916
rect 4120 19913 4126 19916
rect 4120 19904 4130 19913
rect 13449 19907 13507 19913
rect 4120 19876 4165 19904
rect 4120 19867 4130 19876
rect 13449 19873 13461 19907
rect 13495 19904 13507 19907
rect 13909 19907 13967 19913
rect 13909 19904 13921 19907
rect 13495 19876 13921 19904
rect 13495 19873 13507 19876
rect 13449 19867 13507 19873
rect 13909 19873 13921 19876
rect 13955 19904 13967 19907
rect 15102 19904 15108 19916
rect 13955 19876 15108 19904
rect 13955 19873 13967 19876
rect 13909 19867 13967 19873
rect 4120 19864 4126 19867
rect 15102 19864 15108 19876
rect 15160 19864 15166 19916
rect 7006 19836 7012 19848
rect 6967 19808 7012 19836
rect 7006 19796 7012 19808
rect 7064 19796 7070 19848
rect 7101 19839 7159 19845
rect 7101 19805 7113 19839
rect 7147 19805 7159 19839
rect 7101 19799 7159 19805
rect 2685 19771 2743 19777
rect 2685 19768 2697 19771
rect 2332 19740 2697 19768
rect 2685 19737 2697 19740
rect 2731 19737 2743 19771
rect 3050 19768 3056 19780
rect 3011 19740 3056 19768
rect 2685 19731 2743 19737
rect 3050 19728 3056 19740
rect 3108 19728 3114 19780
rect 6086 19728 6092 19780
rect 6144 19768 6150 19780
rect 6638 19768 6644 19780
rect 6144 19740 6644 19768
rect 6144 19728 6150 19740
rect 6638 19728 6644 19740
rect 6696 19768 6702 19780
rect 7116 19768 7144 19799
rect 7374 19796 7380 19848
rect 7432 19836 7438 19848
rect 8113 19839 8171 19845
rect 8113 19836 8125 19839
rect 7432 19808 8125 19836
rect 7432 19796 7438 19808
rect 8113 19805 8125 19808
rect 8159 19836 8171 19839
rect 9858 19836 9864 19848
rect 8159 19808 9864 19836
rect 8159 19805 8171 19808
rect 8113 19799 8171 19805
rect 9858 19796 9864 19808
rect 9916 19836 9922 19848
rect 9953 19839 10011 19845
rect 9953 19836 9965 19839
rect 9916 19808 9965 19836
rect 9916 19796 9922 19808
rect 9953 19805 9965 19808
rect 9999 19836 10011 19839
rect 10502 19836 10508 19848
rect 9999 19808 10508 19836
rect 9999 19805 10011 19808
rect 9953 19799 10011 19805
rect 10502 19796 10508 19808
rect 10560 19796 10566 19848
rect 13814 19796 13820 19848
rect 13872 19836 13878 19848
rect 14001 19839 14059 19845
rect 14001 19836 14013 19839
rect 13872 19808 14013 19836
rect 13872 19796 13878 19808
rect 14001 19805 14013 19808
rect 14047 19805 14059 19839
rect 14001 19799 14059 19805
rect 14093 19839 14151 19845
rect 14093 19805 14105 19839
rect 14139 19805 14151 19839
rect 14093 19799 14151 19805
rect 6696 19740 7144 19768
rect 11885 19771 11943 19777
rect 6696 19728 6702 19740
rect 11885 19737 11897 19771
rect 11931 19768 11943 19771
rect 12526 19768 12532 19780
rect 11931 19740 12532 19768
rect 11931 19737 11943 19740
rect 11885 19731 11943 19737
rect 12526 19728 12532 19740
rect 12584 19728 12590 19780
rect 13081 19771 13139 19777
rect 13081 19737 13093 19771
rect 13127 19768 13139 19771
rect 14108 19768 14136 19799
rect 14458 19768 14464 19780
rect 13127 19740 14464 19768
rect 13127 19737 13139 19740
rect 13081 19731 13139 19737
rect 14458 19728 14464 19740
rect 14516 19768 14522 19780
rect 14553 19771 14611 19777
rect 14553 19768 14565 19771
rect 14516 19740 14565 19768
rect 14516 19728 14522 19740
rect 14553 19737 14565 19740
rect 14599 19737 14611 19771
rect 14553 19731 14611 19737
rect 1578 19700 1584 19712
rect 1539 19672 1584 19700
rect 1578 19660 1584 19672
rect 1636 19660 1642 19712
rect 3786 19700 3792 19712
rect 3747 19672 3792 19700
rect 3786 19660 3792 19672
rect 3844 19660 3850 19712
rect 4430 19660 4436 19712
rect 4488 19700 4494 19712
rect 5445 19703 5503 19709
rect 5445 19700 5457 19703
rect 4488 19672 5457 19700
rect 4488 19660 4494 19672
rect 5445 19669 5457 19672
rect 5491 19669 5503 19703
rect 5445 19663 5503 19669
rect 5534 19660 5540 19712
rect 5592 19700 5598 19712
rect 6549 19703 6607 19709
rect 6549 19700 6561 19703
rect 5592 19672 6561 19700
rect 5592 19660 5598 19672
rect 6549 19669 6561 19672
rect 6595 19669 6607 19703
rect 6549 19663 6607 19669
rect 7745 19703 7803 19709
rect 7745 19669 7757 19703
rect 7791 19700 7803 19703
rect 7926 19700 7932 19712
rect 7791 19672 7932 19700
rect 7791 19669 7803 19672
rect 7745 19663 7803 19669
rect 7926 19660 7932 19672
rect 7984 19660 7990 19712
rect 8386 19700 8392 19712
rect 8347 19672 8392 19700
rect 8386 19660 8392 19672
rect 8444 19660 8450 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 2314 19496 2320 19508
rect 2275 19468 2320 19496
rect 2314 19456 2320 19468
rect 2372 19456 2378 19508
rect 6086 19456 6092 19508
rect 6144 19496 6150 19508
rect 6181 19499 6239 19505
rect 6181 19496 6193 19499
rect 6144 19468 6193 19496
rect 6144 19456 6150 19468
rect 6181 19465 6193 19468
rect 6227 19465 6239 19499
rect 6181 19459 6239 19465
rect 6914 19456 6920 19508
rect 6972 19496 6978 19508
rect 7009 19499 7067 19505
rect 7009 19496 7021 19499
rect 6972 19468 7021 19496
rect 6972 19456 6978 19468
rect 7009 19465 7021 19468
rect 7055 19496 7067 19499
rect 7190 19496 7196 19508
rect 7055 19468 7196 19496
rect 7055 19465 7067 19468
rect 7009 19459 7067 19465
rect 7190 19456 7196 19468
rect 7248 19456 7254 19508
rect 7650 19496 7656 19508
rect 7611 19468 7656 19496
rect 7650 19456 7656 19468
rect 7708 19456 7714 19508
rect 9950 19456 9956 19508
rect 10008 19496 10014 19508
rect 10502 19496 10508 19508
rect 10008 19468 10508 19496
rect 10008 19456 10014 19468
rect 10502 19456 10508 19468
rect 10560 19496 10566 19508
rect 10597 19499 10655 19505
rect 10597 19496 10609 19499
rect 10560 19468 10609 19496
rect 10560 19456 10566 19468
rect 10597 19465 10609 19468
rect 10643 19496 10655 19499
rect 12618 19496 12624 19508
rect 10643 19468 12388 19496
rect 12579 19468 12624 19496
rect 10643 19465 10655 19468
rect 10597 19459 10655 19465
rect 7466 19388 7472 19440
rect 7524 19428 7530 19440
rect 7834 19428 7840 19440
rect 7524 19400 7840 19428
rect 7524 19388 7530 19400
rect 7834 19388 7840 19400
rect 7892 19388 7898 19440
rect 12360 19428 12388 19468
rect 12618 19456 12624 19468
rect 12676 19456 12682 19508
rect 14550 19496 14556 19508
rect 13188 19468 14556 19496
rect 12710 19428 12716 19440
rect 12360 19400 12716 19428
rect 12710 19388 12716 19400
rect 12768 19388 12774 19440
rect 1302 19320 1308 19372
rect 1360 19360 1366 19372
rect 2314 19360 2320 19372
rect 1360 19332 2320 19360
rect 1360 19320 1366 19332
rect 2314 19320 2320 19332
rect 2372 19320 2378 19372
rect 4430 19360 4436 19372
rect 3988 19332 4436 19360
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19292 1455 19295
rect 2501 19295 2559 19301
rect 1443 19264 2084 19292
rect 1443 19261 1455 19264
rect 1397 19255 1455 19261
rect 2056 19168 2084 19264
rect 2501 19261 2513 19295
rect 2547 19292 2559 19295
rect 2958 19292 2964 19304
rect 2547 19264 2964 19292
rect 2547 19261 2559 19264
rect 2501 19255 2559 19261
rect 2958 19252 2964 19264
rect 3016 19292 3022 19304
rect 3697 19295 3755 19301
rect 3016 19264 3188 19292
rect 3016 19252 3022 19264
rect 1486 19116 1492 19168
rect 1544 19156 1550 19168
rect 1581 19159 1639 19165
rect 1581 19156 1593 19159
rect 1544 19128 1593 19156
rect 1544 19116 1550 19128
rect 1581 19125 1593 19128
rect 1627 19125 1639 19159
rect 2038 19156 2044 19168
rect 1999 19128 2044 19156
rect 1581 19119 1639 19125
rect 2038 19116 2044 19128
rect 2096 19116 2102 19168
rect 2682 19156 2688 19168
rect 2643 19128 2688 19156
rect 2682 19116 2688 19128
rect 2740 19116 2746 19168
rect 3160 19165 3188 19264
rect 3697 19261 3709 19295
rect 3743 19292 3755 19295
rect 3988 19292 4016 19332
rect 4430 19320 4436 19332
rect 4488 19320 4494 19372
rect 7006 19360 7012 19372
rect 6840 19332 7012 19360
rect 4154 19292 4160 19304
rect 3743 19264 4016 19292
rect 4115 19264 4160 19292
rect 3743 19261 3755 19264
rect 3697 19255 3755 19261
rect 4154 19252 4160 19264
rect 4212 19252 4218 19304
rect 5350 19292 5356 19304
rect 5311 19264 5356 19292
rect 5350 19252 5356 19264
rect 5408 19252 5414 19304
rect 5442 19252 5448 19304
rect 5500 19292 5506 19304
rect 5813 19295 5871 19301
rect 5813 19292 5825 19295
rect 5500 19264 5825 19292
rect 5500 19252 5506 19264
rect 5813 19261 5825 19264
rect 5859 19261 5871 19295
rect 5813 19255 5871 19261
rect 6641 19295 6699 19301
rect 6641 19261 6653 19295
rect 6687 19292 6699 19295
rect 6840 19292 6868 19332
rect 7006 19320 7012 19332
rect 7064 19360 7070 19372
rect 7558 19360 7564 19372
rect 7064 19332 7564 19360
rect 7064 19320 7070 19332
rect 7558 19320 7564 19332
rect 7616 19320 7622 19372
rect 8297 19363 8355 19369
rect 8297 19329 8309 19363
rect 8343 19360 8355 19363
rect 8386 19360 8392 19372
rect 8343 19332 8392 19360
rect 8343 19329 8355 19332
rect 8297 19323 8355 19329
rect 8386 19320 8392 19332
rect 8444 19320 8450 19372
rect 9861 19363 9919 19369
rect 9861 19329 9873 19363
rect 9907 19360 9919 19363
rect 10870 19360 10876 19372
rect 9907 19332 10876 19360
rect 9907 19329 9919 19332
rect 9861 19323 9919 19329
rect 6687 19264 6868 19292
rect 6687 19261 6699 19264
rect 6641 19255 6699 19261
rect 8938 19252 8944 19304
rect 8996 19292 9002 19304
rect 9585 19295 9643 19301
rect 9585 19292 9597 19295
rect 8996 19264 9597 19292
rect 8996 19252 9002 19264
rect 9585 19261 9597 19264
rect 9631 19261 9643 19295
rect 9585 19255 9643 19261
rect 9674 19252 9680 19304
rect 9732 19292 9738 19304
rect 9732 19264 9777 19292
rect 9732 19252 9738 19264
rect 4890 19224 4896 19236
rect 4803 19196 4896 19224
rect 4890 19184 4896 19196
rect 4948 19224 4954 19236
rect 7006 19224 7012 19236
rect 4948 19196 7012 19224
rect 4948 19184 4954 19196
rect 7006 19184 7012 19196
rect 7064 19184 7070 19236
rect 7926 19184 7932 19236
rect 7984 19224 7990 19236
rect 8113 19227 8171 19233
rect 8113 19224 8125 19227
rect 7984 19196 8125 19224
rect 7984 19184 7990 19196
rect 8113 19193 8125 19196
rect 8159 19193 8171 19227
rect 8113 19187 8171 19193
rect 9125 19227 9183 19233
rect 9125 19193 9137 19227
rect 9171 19224 9183 19227
rect 9876 19224 9904 19323
rect 10870 19320 10876 19332
rect 10928 19320 10934 19372
rect 11422 19360 11428 19372
rect 11383 19332 11428 19360
rect 11422 19320 11428 19332
rect 11480 19320 11486 19372
rect 13188 19369 13216 19468
rect 14550 19456 14556 19468
rect 14608 19496 14614 19508
rect 15565 19499 15623 19505
rect 15565 19496 15577 19499
rect 14608 19468 15577 19496
rect 14608 19456 14614 19468
rect 15565 19465 15577 19468
rect 15611 19465 15623 19499
rect 15565 19459 15623 19465
rect 12437 19363 12495 19369
rect 12437 19329 12449 19363
rect 12483 19360 12495 19363
rect 13173 19363 13231 19369
rect 13173 19360 13185 19363
rect 12483 19332 13185 19360
rect 12483 19329 12495 19332
rect 12437 19323 12495 19329
rect 13173 19329 13185 19332
rect 13219 19329 13231 19363
rect 13173 19323 13231 19329
rect 11054 19252 11060 19304
rect 11112 19292 11118 19304
rect 11149 19295 11207 19301
rect 11149 19292 11161 19295
rect 11112 19264 11161 19292
rect 11112 19252 11118 19264
rect 11149 19261 11161 19264
rect 11195 19261 11207 19295
rect 11149 19255 11207 19261
rect 11241 19295 11299 19301
rect 11241 19261 11253 19295
rect 11287 19292 11299 19295
rect 11885 19295 11943 19301
rect 11885 19292 11897 19295
rect 11287 19264 11897 19292
rect 11287 19261 11299 19264
rect 11241 19255 11299 19261
rect 11885 19261 11897 19264
rect 11931 19292 11943 19295
rect 12158 19292 12164 19304
rect 11931 19264 12164 19292
rect 11931 19261 11943 19264
rect 11885 19255 11943 19261
rect 12158 19252 12164 19264
rect 12216 19252 12222 19304
rect 12253 19295 12311 19301
rect 12253 19261 12265 19295
rect 12299 19292 12311 19295
rect 12345 19295 12403 19301
rect 12345 19292 12357 19295
rect 12299 19264 12357 19292
rect 12299 19261 12311 19264
rect 12253 19255 12311 19261
rect 12345 19261 12357 19264
rect 12391 19261 12403 19295
rect 12986 19292 12992 19304
rect 12947 19264 12992 19292
rect 12345 19255 12403 19261
rect 12986 19252 12992 19264
rect 13044 19252 13050 19304
rect 14090 19292 14096 19304
rect 13096 19264 14096 19292
rect 9171 19196 9904 19224
rect 9171 19193 9183 19196
rect 9125 19187 9183 19193
rect 12710 19184 12716 19236
rect 12768 19224 12774 19236
rect 13096 19224 13124 19264
rect 14090 19252 14096 19264
rect 14148 19292 14154 19304
rect 14458 19301 14464 19304
rect 14185 19295 14243 19301
rect 14185 19292 14197 19295
rect 14148 19264 14197 19292
rect 14148 19252 14154 19264
rect 14185 19261 14197 19264
rect 14231 19261 14243 19295
rect 14452 19292 14464 19301
rect 14419 19264 14464 19292
rect 14185 19255 14243 19261
rect 14452 19255 14464 19264
rect 14458 19252 14464 19255
rect 14516 19252 14522 19304
rect 12768 19196 13124 19224
rect 12768 19184 12774 19196
rect 3145 19159 3203 19165
rect 3145 19125 3157 19159
rect 3191 19156 3203 19159
rect 3234 19156 3240 19168
rect 3191 19128 3240 19156
rect 3191 19125 3203 19128
rect 3145 19119 3203 19125
rect 3234 19116 3240 19128
rect 3292 19116 3298 19168
rect 3789 19159 3847 19165
rect 3789 19125 3801 19159
rect 3835 19156 3847 19159
rect 3878 19156 3884 19168
rect 3835 19128 3884 19156
rect 3835 19125 3847 19128
rect 3789 19119 3847 19125
rect 3878 19116 3884 19128
rect 3936 19116 3942 19168
rect 4246 19156 4252 19168
rect 4207 19128 4252 19156
rect 4246 19116 4252 19128
rect 4304 19116 4310 19168
rect 5074 19116 5080 19168
rect 5132 19156 5138 19168
rect 5169 19159 5227 19165
rect 5169 19156 5181 19159
rect 5132 19128 5181 19156
rect 5132 19116 5138 19128
rect 5169 19125 5181 19128
rect 5215 19125 5227 19159
rect 5169 19119 5227 19125
rect 7561 19159 7619 19165
rect 7561 19125 7573 19159
rect 7607 19156 7619 19159
rect 8021 19159 8079 19165
rect 8021 19156 8033 19159
rect 7607 19128 8033 19156
rect 7607 19125 7619 19128
rect 7561 19119 7619 19125
rect 8021 19125 8033 19128
rect 8067 19156 8079 19159
rect 8202 19156 8208 19168
rect 8067 19128 8208 19156
rect 8067 19125 8079 19128
rect 8021 19119 8079 19125
rect 8202 19116 8208 19128
rect 8260 19116 8266 19168
rect 8386 19116 8392 19168
rect 8444 19156 8450 19168
rect 8665 19159 8723 19165
rect 8665 19156 8677 19159
rect 8444 19128 8677 19156
rect 8444 19116 8450 19128
rect 8665 19125 8677 19128
rect 8711 19125 8723 19159
rect 9214 19156 9220 19168
rect 9175 19128 9220 19156
rect 8665 19119 8723 19125
rect 9214 19116 9220 19128
rect 9272 19116 9278 19168
rect 10778 19156 10784 19168
rect 10739 19128 10784 19156
rect 10778 19116 10784 19128
rect 10836 19116 10842 19168
rect 13078 19156 13084 19168
rect 13039 19128 13084 19156
rect 13078 19116 13084 19128
rect 13136 19116 13142 19168
rect 13725 19159 13783 19165
rect 13725 19125 13737 19159
rect 13771 19156 13783 19159
rect 13814 19156 13820 19168
rect 13771 19128 13820 19156
rect 13771 19125 13783 19128
rect 13725 19119 13783 19125
rect 13814 19116 13820 19128
rect 13872 19116 13878 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 3881 18955 3939 18961
rect 3881 18921 3893 18955
rect 3927 18952 3939 18955
rect 4246 18952 4252 18964
rect 3927 18924 4252 18952
rect 3927 18921 3939 18924
rect 3881 18915 3939 18921
rect 4246 18912 4252 18924
rect 4304 18952 4310 18964
rect 4525 18955 4583 18961
rect 4525 18952 4537 18955
rect 4304 18924 4537 18952
rect 4304 18912 4310 18924
rect 4525 18921 4537 18924
rect 4571 18921 4583 18955
rect 4525 18915 4583 18921
rect 4985 18955 5043 18961
rect 4985 18921 4997 18955
rect 5031 18952 5043 18955
rect 5166 18952 5172 18964
rect 5031 18924 5172 18952
rect 5031 18921 5043 18924
rect 4985 18915 5043 18921
rect 5166 18912 5172 18924
rect 5224 18952 5230 18964
rect 6089 18955 6147 18961
rect 6089 18952 6101 18955
rect 5224 18924 6101 18952
rect 5224 18912 5230 18924
rect 6089 18921 6101 18924
rect 6135 18921 6147 18955
rect 6089 18915 6147 18921
rect 7006 18912 7012 18964
rect 7064 18952 7070 18964
rect 7193 18955 7251 18961
rect 7193 18952 7205 18955
rect 7064 18924 7205 18952
rect 7064 18912 7070 18924
rect 7193 18921 7205 18924
rect 7239 18952 7251 18955
rect 7374 18952 7380 18964
rect 7239 18924 7380 18952
rect 7239 18921 7251 18924
rect 7193 18915 7251 18921
rect 7374 18912 7380 18924
rect 7432 18912 7438 18964
rect 8018 18912 8024 18964
rect 8076 18952 8082 18964
rect 8113 18955 8171 18961
rect 8113 18952 8125 18955
rect 8076 18924 8125 18952
rect 8076 18912 8082 18924
rect 8113 18921 8125 18924
rect 8159 18921 8171 18955
rect 8113 18915 8171 18921
rect 8938 18912 8944 18964
rect 8996 18952 9002 18964
rect 9033 18955 9091 18961
rect 9033 18952 9045 18955
rect 8996 18924 9045 18952
rect 8996 18912 9002 18924
rect 9033 18921 9045 18924
rect 9079 18921 9091 18955
rect 9033 18915 9091 18921
rect 10781 18955 10839 18961
rect 10781 18921 10793 18955
rect 10827 18952 10839 18955
rect 10870 18952 10876 18964
rect 10827 18924 10876 18952
rect 10827 18921 10839 18924
rect 10781 18915 10839 18921
rect 10870 18912 10876 18924
rect 10928 18912 10934 18964
rect 11146 18912 11152 18964
rect 11204 18952 11210 18964
rect 11241 18955 11299 18961
rect 11241 18952 11253 18955
rect 11204 18924 11253 18952
rect 11204 18912 11210 18924
rect 11241 18921 11253 18924
rect 11287 18921 11299 18955
rect 11241 18915 11299 18921
rect 14093 18955 14151 18961
rect 14093 18921 14105 18955
rect 14139 18952 14151 18955
rect 14458 18952 14464 18964
rect 14139 18924 14464 18952
rect 14139 18921 14151 18924
rect 14093 18915 14151 18921
rect 14458 18912 14464 18924
rect 14516 18912 14522 18964
rect 15286 18952 15292 18964
rect 15247 18924 15292 18952
rect 15286 18912 15292 18924
rect 15344 18912 15350 18964
rect 3513 18887 3571 18893
rect 3513 18853 3525 18887
rect 3559 18884 3571 18887
rect 4154 18884 4160 18896
rect 3559 18856 4160 18884
rect 3559 18853 3571 18856
rect 3513 18847 3571 18853
rect 4154 18844 4160 18856
rect 4212 18844 4218 18896
rect 4341 18887 4399 18893
rect 4341 18853 4353 18887
rect 4387 18884 4399 18887
rect 4430 18884 4436 18896
rect 4387 18856 4436 18884
rect 4387 18853 4399 18856
rect 4341 18847 4399 18853
rect 4430 18844 4436 18856
rect 4488 18844 4494 18896
rect 4893 18887 4951 18893
rect 4893 18853 4905 18887
rect 4939 18884 4951 18887
rect 5442 18884 5448 18896
rect 4939 18856 5448 18884
rect 4939 18853 4951 18856
rect 4893 18847 4951 18853
rect 1397 18819 1455 18825
rect 1397 18785 1409 18819
rect 1443 18816 1455 18819
rect 1670 18816 1676 18828
rect 1443 18788 1676 18816
rect 1443 18785 1455 18788
rect 1397 18779 1455 18785
rect 1670 18776 1676 18788
rect 1728 18776 1734 18828
rect 2501 18819 2559 18825
rect 2501 18785 2513 18819
rect 2547 18785 2559 18819
rect 2501 18779 2559 18785
rect 2409 18683 2467 18689
rect 2409 18649 2421 18683
rect 2455 18680 2467 18683
rect 2516 18680 2544 18779
rect 3970 18776 3976 18828
rect 4028 18816 4034 18828
rect 4908 18816 4936 18847
rect 5442 18844 5448 18856
rect 5500 18844 5506 18896
rect 9490 18844 9496 18896
rect 9548 18884 9554 18896
rect 9950 18884 9956 18896
rect 9548 18856 9956 18884
rect 9548 18844 9554 18856
rect 9950 18844 9956 18856
rect 10008 18844 10014 18896
rect 11054 18844 11060 18896
rect 11112 18884 11118 18896
rect 11701 18887 11759 18893
rect 11701 18884 11713 18887
rect 11112 18856 11713 18884
rect 11112 18844 11118 18856
rect 11701 18853 11713 18856
rect 11747 18853 11759 18887
rect 11701 18847 11759 18853
rect 12161 18887 12219 18893
rect 12161 18853 12173 18887
rect 12207 18884 12219 18887
rect 13078 18884 13084 18896
rect 12207 18856 13084 18884
rect 12207 18853 12219 18856
rect 12161 18847 12219 18853
rect 13078 18844 13084 18856
rect 13136 18844 13142 18896
rect 6454 18816 6460 18828
rect 4028 18788 4936 18816
rect 6415 18788 6460 18816
rect 4028 18776 4034 18788
rect 6454 18776 6460 18788
rect 6512 18776 6518 18828
rect 6549 18819 6607 18825
rect 6549 18785 6561 18819
rect 6595 18816 6607 18819
rect 6730 18816 6736 18828
rect 6595 18788 6736 18816
rect 6595 18785 6607 18788
rect 6549 18779 6607 18785
rect 6730 18776 6736 18788
rect 6788 18816 6794 18828
rect 7466 18816 7472 18828
rect 6788 18788 7472 18816
rect 6788 18776 6794 18788
rect 7466 18776 7472 18788
rect 7524 18776 7530 18828
rect 8021 18819 8079 18825
rect 8021 18785 8033 18819
rect 8067 18785 8079 18819
rect 10042 18816 10048 18828
rect 10003 18788 10048 18816
rect 8021 18779 8079 18785
rect 3786 18708 3792 18760
rect 3844 18748 3850 18760
rect 5074 18748 5080 18760
rect 3844 18720 5080 18748
rect 3844 18708 3850 18720
rect 5074 18708 5080 18720
rect 5132 18708 5138 18760
rect 6638 18708 6644 18760
rect 6696 18748 6702 18760
rect 7834 18748 7840 18760
rect 6696 18720 6741 18748
rect 6820 18720 7840 18748
rect 6696 18708 6702 18720
rect 6820 18680 6848 18720
rect 7834 18708 7840 18720
rect 7892 18708 7898 18760
rect 2455 18652 6848 18680
rect 2455 18649 2467 18652
rect 2409 18643 2467 18649
rect 6914 18640 6920 18692
rect 6972 18680 6978 18692
rect 7469 18683 7527 18689
rect 7469 18680 7481 18683
rect 6972 18652 7481 18680
rect 6972 18640 6978 18652
rect 7469 18649 7481 18652
rect 7515 18680 7527 18683
rect 8036 18680 8064 18779
rect 10042 18776 10048 18788
rect 10100 18776 10106 18828
rect 11149 18819 11207 18825
rect 11149 18785 11161 18819
rect 11195 18816 11207 18819
rect 11422 18816 11428 18828
rect 11195 18788 11428 18816
rect 11195 18785 11207 18788
rect 11149 18779 11207 18785
rect 11422 18776 11428 18788
rect 11480 18816 11486 18828
rect 12802 18816 12808 18828
rect 11480 18788 12808 18816
rect 11480 18776 11486 18788
rect 12802 18776 12808 18788
rect 12860 18816 12866 18828
rect 12980 18819 13038 18825
rect 12980 18816 12992 18819
rect 12860 18788 12992 18816
rect 12860 18776 12866 18788
rect 12980 18785 12992 18788
rect 13026 18816 13038 18819
rect 13538 18816 13544 18828
rect 13026 18788 13544 18816
rect 13026 18785 13038 18788
rect 12980 18779 13038 18785
rect 13538 18776 13544 18788
rect 13596 18776 13602 18828
rect 8202 18708 8208 18760
rect 8260 18748 8266 18760
rect 8260 18720 8305 18748
rect 8260 18708 8266 18720
rect 9950 18708 9956 18760
rect 10008 18748 10014 18760
rect 10134 18748 10140 18760
rect 10008 18720 10140 18748
rect 10008 18708 10014 18720
rect 10134 18708 10140 18720
rect 10192 18708 10198 18760
rect 10321 18751 10379 18757
rect 10321 18717 10333 18751
rect 10367 18748 10379 18751
rect 10410 18748 10416 18760
rect 10367 18720 10416 18748
rect 10367 18717 10379 18720
rect 10321 18711 10379 18717
rect 10410 18708 10416 18720
rect 10468 18708 10474 18760
rect 12710 18748 12716 18760
rect 12671 18720 12716 18748
rect 12710 18708 12716 18720
rect 12768 18708 12774 18760
rect 7515 18652 8064 18680
rect 7515 18649 7527 18652
rect 7469 18643 7527 18649
rect 11054 18640 11060 18692
rect 11112 18680 11118 18692
rect 11112 18652 12756 18680
rect 11112 18640 11118 18652
rect 1394 18572 1400 18624
rect 1452 18612 1458 18624
rect 1581 18615 1639 18621
rect 1581 18612 1593 18615
rect 1452 18584 1593 18612
rect 1452 18572 1458 18584
rect 1581 18581 1593 18584
rect 1627 18581 1639 18615
rect 2038 18612 2044 18624
rect 1999 18584 2044 18612
rect 1581 18575 1639 18581
rect 2038 18572 2044 18584
rect 2096 18572 2102 18624
rect 2682 18612 2688 18624
rect 2643 18584 2688 18612
rect 2682 18572 2688 18584
rect 2740 18572 2746 18624
rect 3145 18615 3203 18621
rect 3145 18581 3157 18615
rect 3191 18612 3203 18615
rect 3234 18612 3240 18624
rect 3191 18584 3240 18612
rect 3191 18581 3203 18584
rect 3145 18575 3203 18581
rect 3234 18572 3240 18584
rect 3292 18572 3298 18624
rect 5629 18615 5687 18621
rect 5629 18581 5641 18615
rect 5675 18612 5687 18615
rect 6362 18612 6368 18624
rect 5675 18584 6368 18612
rect 5675 18581 5687 18584
rect 5629 18575 5687 18581
rect 6362 18572 6368 18584
rect 6420 18572 6426 18624
rect 7650 18612 7656 18624
rect 7611 18584 7656 18612
rect 7650 18572 7656 18584
rect 7708 18572 7714 18624
rect 9398 18612 9404 18624
rect 9359 18584 9404 18612
rect 9398 18572 9404 18584
rect 9456 18572 9462 18624
rect 9677 18615 9735 18621
rect 9677 18581 9689 18615
rect 9723 18612 9735 18615
rect 9858 18612 9864 18624
rect 9723 18584 9864 18612
rect 9723 18581 9735 18584
rect 9677 18575 9735 18581
rect 9858 18572 9864 18584
rect 9916 18572 9922 18624
rect 12526 18612 12532 18624
rect 12487 18584 12532 18612
rect 12526 18572 12532 18584
rect 12584 18572 12590 18624
rect 12728 18612 12756 18652
rect 15378 18612 15384 18624
rect 12728 18584 15384 18612
rect 15378 18572 15384 18584
rect 15436 18572 15442 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 3786 18408 3792 18420
rect 3747 18380 3792 18408
rect 3786 18368 3792 18380
rect 3844 18368 3850 18420
rect 8386 18408 8392 18420
rect 8347 18380 8392 18408
rect 8386 18368 8392 18380
rect 8444 18368 8450 18420
rect 9306 18368 9312 18420
rect 9364 18408 9370 18420
rect 10410 18408 10416 18420
rect 9364 18380 10416 18408
rect 9364 18368 9370 18380
rect 10410 18368 10416 18380
rect 10468 18408 10474 18420
rect 11425 18411 11483 18417
rect 11425 18408 11437 18411
rect 10468 18380 11437 18408
rect 10468 18368 10474 18380
rect 11425 18377 11437 18380
rect 11471 18377 11483 18411
rect 11425 18371 11483 18377
rect 13078 18368 13084 18420
rect 13136 18408 13142 18420
rect 14001 18411 14059 18417
rect 14001 18408 14013 18411
rect 13136 18380 14013 18408
rect 13136 18368 13142 18380
rect 14001 18377 14013 18380
rect 14047 18377 14059 18411
rect 14001 18371 14059 18377
rect 2590 18300 2596 18352
rect 2648 18340 2654 18352
rect 2685 18343 2743 18349
rect 2685 18340 2697 18343
rect 2648 18312 2697 18340
rect 2648 18300 2654 18312
rect 2685 18309 2697 18312
rect 2731 18309 2743 18343
rect 2685 18303 2743 18309
rect 8018 18300 8024 18352
rect 8076 18340 8082 18352
rect 8941 18343 8999 18349
rect 8941 18340 8953 18343
rect 8076 18312 8953 18340
rect 8076 18300 8082 18312
rect 8941 18309 8953 18312
rect 8987 18309 8999 18343
rect 8941 18303 8999 18309
rect 12710 18300 12716 18352
rect 12768 18340 12774 18352
rect 13449 18343 13507 18349
rect 13449 18340 13461 18343
rect 12768 18312 13461 18340
rect 12768 18300 12774 18312
rect 13449 18309 13461 18312
rect 13495 18309 13507 18343
rect 13449 18303 13507 18309
rect 3234 18272 3240 18284
rect 3195 18244 3240 18272
rect 3234 18232 3240 18244
rect 3292 18232 3298 18284
rect 7006 18272 7012 18284
rect 6967 18244 7012 18272
rect 7006 18232 7012 18244
rect 7064 18232 7070 18284
rect 9401 18275 9459 18281
rect 9401 18241 9413 18275
rect 9447 18272 9459 18275
rect 11885 18275 11943 18281
rect 9447 18244 9628 18272
rect 9447 18241 9459 18244
rect 9401 18235 9459 18241
rect 1397 18207 1455 18213
rect 1397 18173 1409 18207
rect 1443 18204 1455 18207
rect 2038 18204 2044 18216
rect 1443 18176 2044 18204
rect 1443 18173 1455 18176
rect 1397 18167 1455 18173
rect 2038 18164 2044 18176
rect 2096 18164 2102 18216
rect 2225 18207 2283 18213
rect 2225 18173 2237 18207
rect 2271 18204 2283 18207
rect 2958 18204 2964 18216
rect 2271 18176 2964 18204
rect 2271 18173 2283 18176
rect 2225 18167 2283 18173
rect 2958 18164 2964 18176
rect 3016 18164 3022 18216
rect 3142 18204 3148 18216
rect 3103 18176 3148 18204
rect 3142 18164 3148 18176
rect 3200 18164 3206 18216
rect 4062 18164 4068 18216
rect 4120 18204 4126 18216
rect 4157 18207 4215 18213
rect 4157 18204 4169 18207
rect 4120 18176 4169 18204
rect 4120 18164 4126 18176
rect 4157 18173 4169 18176
rect 4203 18204 4215 18207
rect 4249 18207 4307 18213
rect 4249 18204 4261 18207
rect 4203 18176 4261 18204
rect 4203 18173 4215 18176
rect 4157 18167 4215 18173
rect 4249 18173 4261 18176
rect 4295 18204 4307 18207
rect 4890 18204 4896 18216
rect 4295 18176 4896 18204
rect 4295 18173 4307 18176
rect 4249 18167 4307 18173
rect 4890 18164 4896 18176
rect 4948 18164 4954 18216
rect 9490 18204 9496 18216
rect 9451 18176 9496 18204
rect 9490 18164 9496 18176
rect 9548 18164 9554 18216
rect 9600 18204 9628 18244
rect 11885 18241 11897 18275
rect 11931 18272 11943 18275
rect 12989 18275 13047 18281
rect 12989 18272 13001 18275
rect 11931 18244 13001 18272
rect 11931 18241 11943 18244
rect 11885 18235 11943 18241
rect 12989 18241 13001 18244
rect 13035 18272 13047 18275
rect 13722 18272 13728 18284
rect 13035 18244 13728 18272
rect 13035 18241 13047 18244
rect 12989 18235 13047 18241
rect 13722 18232 13728 18244
rect 13780 18232 13786 18284
rect 14458 18232 14464 18284
rect 14516 18272 14522 18284
rect 14553 18275 14611 18281
rect 14553 18272 14565 18275
rect 14516 18244 14565 18272
rect 14516 18232 14522 18244
rect 14553 18241 14565 18244
rect 14599 18241 14611 18275
rect 14553 18235 14611 18241
rect 10042 18204 10048 18216
rect 9600 18176 10048 18204
rect 10042 18164 10048 18176
rect 10100 18204 10106 18216
rect 11054 18204 11060 18216
rect 10100 18176 11060 18204
rect 10100 18164 10106 18176
rect 11054 18164 11060 18176
rect 11112 18164 11118 18216
rect 12526 18164 12532 18216
rect 12584 18204 12590 18216
rect 12805 18207 12863 18213
rect 12805 18204 12817 18207
rect 12584 18176 12817 18204
rect 12584 18164 12590 18176
rect 12805 18173 12817 18176
rect 12851 18173 12863 18207
rect 12805 18167 12863 18173
rect 2593 18139 2651 18145
rect 2593 18105 2605 18139
rect 2639 18136 2651 18139
rect 3160 18136 3188 18164
rect 2639 18108 3188 18136
rect 2639 18105 2651 18108
rect 2593 18099 2651 18105
rect 4430 18096 4436 18148
rect 4488 18145 4494 18148
rect 4488 18139 4552 18145
rect 4488 18105 4506 18139
rect 4540 18105 4552 18139
rect 4488 18099 4552 18105
rect 4488 18096 4494 18099
rect 5074 18096 5080 18148
rect 5132 18136 5138 18148
rect 6181 18139 6239 18145
rect 6181 18136 6193 18139
rect 5132 18108 6193 18136
rect 5132 18096 5138 18108
rect 6181 18105 6193 18108
rect 6227 18136 6239 18139
rect 6454 18136 6460 18148
rect 6227 18108 6460 18136
rect 6227 18105 6239 18108
rect 6181 18099 6239 18105
rect 6454 18096 6460 18108
rect 6512 18096 6518 18148
rect 7276 18139 7334 18145
rect 7276 18105 7288 18139
rect 7322 18136 7334 18139
rect 7374 18136 7380 18148
rect 7322 18108 7380 18136
rect 7322 18105 7334 18108
rect 7276 18099 7334 18105
rect 7374 18096 7380 18108
rect 7432 18096 7438 18148
rect 9398 18096 9404 18148
rect 9456 18136 9462 18148
rect 9738 18139 9796 18145
rect 9738 18136 9750 18139
rect 9456 18108 9750 18136
rect 9456 18096 9462 18108
rect 9738 18105 9750 18108
rect 9784 18105 9796 18139
rect 12250 18136 12256 18148
rect 12163 18108 12256 18136
rect 9738 18099 9796 18105
rect 12250 18096 12256 18108
rect 12308 18136 12314 18148
rect 12897 18139 12955 18145
rect 12897 18136 12909 18139
rect 12308 18108 12909 18136
rect 12308 18096 12314 18108
rect 12897 18105 12909 18108
rect 12943 18105 12955 18139
rect 12897 18099 12955 18105
rect 14182 18096 14188 18148
rect 14240 18136 14246 18148
rect 14461 18139 14519 18145
rect 14461 18136 14473 18139
rect 14240 18108 14473 18136
rect 14240 18096 14246 18108
rect 14461 18105 14473 18108
rect 14507 18136 14519 18139
rect 14642 18136 14648 18148
rect 14507 18108 14648 18136
rect 14507 18105 14519 18108
rect 14461 18099 14519 18105
rect 14642 18096 14648 18108
rect 14700 18096 14706 18148
rect 1578 18068 1584 18080
rect 1539 18040 1584 18068
rect 1578 18028 1584 18040
rect 1636 18028 1642 18080
rect 2958 18028 2964 18080
rect 3016 18068 3022 18080
rect 3053 18071 3111 18077
rect 3053 18068 3065 18071
rect 3016 18040 3065 18068
rect 3016 18028 3022 18040
rect 3053 18037 3065 18040
rect 3099 18068 3111 18071
rect 3418 18068 3424 18080
rect 3099 18040 3424 18068
rect 3099 18037 3111 18040
rect 3053 18031 3111 18037
rect 3418 18028 3424 18040
rect 3476 18028 3482 18080
rect 5534 18028 5540 18080
rect 5592 18068 5598 18080
rect 5629 18071 5687 18077
rect 5629 18068 5641 18071
rect 5592 18040 5641 18068
rect 5592 18028 5598 18040
rect 5629 18037 5641 18040
rect 5675 18037 5687 18071
rect 5629 18031 5687 18037
rect 6641 18071 6699 18077
rect 6641 18037 6653 18071
rect 6687 18068 6699 18071
rect 6730 18068 6736 18080
rect 6687 18040 6736 18068
rect 6687 18037 6699 18040
rect 6641 18031 6699 18037
rect 6730 18028 6736 18040
rect 6788 18068 6794 18080
rect 7098 18068 7104 18080
rect 6788 18040 7104 18068
rect 6788 18028 6794 18040
rect 7098 18028 7104 18040
rect 7156 18028 7162 18080
rect 10870 18068 10876 18080
rect 10831 18040 10876 18068
rect 10870 18028 10876 18040
rect 10928 18028 10934 18080
rect 11514 18028 11520 18080
rect 11572 18068 11578 18080
rect 12437 18071 12495 18077
rect 12437 18068 12449 18071
rect 11572 18040 12449 18068
rect 11572 18028 11578 18040
rect 12437 18037 12449 18040
rect 12483 18037 12495 18071
rect 12437 18031 12495 18037
rect 13909 18071 13967 18077
rect 13909 18037 13921 18071
rect 13955 18068 13967 18071
rect 13998 18068 14004 18080
rect 13955 18040 14004 18068
rect 13955 18037 13967 18040
rect 13909 18031 13967 18037
rect 13998 18028 14004 18040
rect 14056 18068 14062 18080
rect 14369 18071 14427 18077
rect 14369 18068 14381 18071
rect 14056 18040 14381 18068
rect 14056 18028 14062 18040
rect 14369 18037 14381 18040
rect 14415 18068 14427 18071
rect 14734 18068 14740 18080
rect 14415 18040 14740 18068
rect 14415 18037 14427 18040
rect 14369 18031 14427 18037
rect 14734 18028 14740 18040
rect 14792 18028 14798 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1670 17824 1676 17876
rect 1728 17864 1734 17876
rect 2225 17867 2283 17873
rect 2225 17864 2237 17867
rect 1728 17836 2237 17864
rect 1728 17824 1734 17836
rect 2225 17833 2237 17836
rect 2271 17833 2283 17867
rect 2225 17827 2283 17833
rect 2777 17867 2835 17873
rect 2777 17833 2789 17867
rect 2823 17864 2835 17867
rect 3418 17864 3424 17876
rect 2823 17836 3424 17864
rect 2823 17833 2835 17836
rect 2777 17827 2835 17833
rect 3418 17824 3424 17836
rect 3476 17864 3482 17876
rect 4065 17867 4123 17873
rect 4065 17864 4077 17867
rect 3476 17836 4077 17864
rect 3476 17824 3482 17836
rect 4065 17833 4077 17836
rect 4111 17833 4123 17867
rect 4065 17827 4123 17833
rect 4525 17867 4583 17873
rect 4525 17833 4537 17867
rect 4571 17864 4583 17867
rect 4614 17864 4620 17876
rect 4571 17836 4620 17864
rect 4571 17833 4583 17836
rect 4525 17827 4583 17833
rect 4614 17824 4620 17836
rect 4672 17824 4678 17876
rect 5166 17864 5172 17876
rect 5127 17836 5172 17864
rect 5166 17824 5172 17836
rect 5224 17824 5230 17876
rect 5629 17867 5687 17873
rect 5629 17833 5641 17867
rect 5675 17864 5687 17867
rect 6822 17864 6828 17876
rect 5675 17836 6828 17864
rect 5675 17833 5687 17836
rect 5629 17827 5687 17833
rect 6822 17824 6828 17836
rect 6880 17824 6886 17876
rect 9030 17824 9036 17876
rect 9088 17864 9094 17876
rect 9490 17864 9496 17876
rect 9088 17836 9496 17864
rect 9088 17824 9094 17836
rect 9490 17824 9496 17836
rect 9548 17824 9554 17876
rect 14458 17864 14464 17876
rect 14419 17836 14464 17864
rect 14458 17824 14464 17836
rect 14516 17824 14522 17876
rect 3881 17799 3939 17805
rect 3881 17765 3893 17799
rect 3927 17796 3939 17799
rect 3970 17796 3976 17808
rect 3927 17768 3976 17796
rect 3927 17765 3939 17768
rect 3881 17759 3939 17765
rect 3970 17756 3976 17768
rect 4028 17756 4034 17808
rect 6181 17799 6239 17805
rect 6181 17765 6193 17799
rect 6227 17796 6239 17799
rect 6638 17796 6644 17808
rect 6227 17768 6644 17796
rect 6227 17765 6239 17768
rect 6181 17759 6239 17765
rect 6638 17756 6644 17768
rect 6696 17756 6702 17808
rect 9950 17796 9956 17808
rect 9911 17768 9956 17796
rect 9950 17756 9956 17768
rect 10008 17756 10014 17808
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17728 1455 17731
rect 4433 17731 4491 17737
rect 4433 17728 4445 17731
rect 1443 17700 4445 17728
rect 1443 17697 1455 17700
rect 1397 17691 1455 17697
rect 4433 17697 4445 17700
rect 4479 17728 4491 17731
rect 5166 17728 5172 17740
rect 4479 17700 5172 17728
rect 4479 17697 4491 17700
rect 4433 17691 4491 17697
rect 5166 17688 5172 17700
rect 5224 17688 5230 17740
rect 6730 17688 6736 17740
rect 6788 17728 6794 17740
rect 6908 17731 6966 17737
rect 6908 17728 6920 17731
rect 6788 17700 6920 17728
rect 6788 17688 6794 17700
rect 6908 17697 6920 17700
rect 6954 17728 6966 17731
rect 8202 17728 8208 17740
rect 6954 17700 8208 17728
rect 6954 17697 6966 17700
rect 6908 17691 6966 17697
rect 8202 17688 8208 17700
rect 8260 17688 8266 17740
rect 10137 17731 10195 17737
rect 10137 17697 10149 17731
rect 10183 17728 10195 17731
rect 10778 17728 10784 17740
rect 10183 17700 10784 17728
rect 10183 17697 10195 17700
rect 10137 17691 10195 17697
rect 10778 17688 10784 17700
rect 10836 17688 10842 17740
rect 11422 17737 11428 17740
rect 11416 17728 11428 17737
rect 11383 17700 11428 17728
rect 11416 17691 11428 17700
rect 11422 17688 11428 17691
rect 11480 17688 11486 17740
rect 2590 17620 2596 17672
rect 2648 17660 2654 17672
rect 2869 17663 2927 17669
rect 2869 17660 2881 17663
rect 2648 17632 2881 17660
rect 2648 17620 2654 17632
rect 2869 17629 2881 17632
rect 2915 17629 2927 17663
rect 3050 17660 3056 17672
rect 3011 17632 3056 17660
rect 2869 17623 2927 17629
rect 3050 17620 3056 17632
rect 3108 17620 3114 17672
rect 4709 17663 4767 17669
rect 4709 17629 4721 17663
rect 4755 17660 4767 17663
rect 4890 17660 4896 17672
rect 4755 17632 4896 17660
rect 4755 17629 4767 17632
rect 4709 17623 4767 17629
rect 4890 17620 4896 17632
rect 4948 17660 4954 17672
rect 5534 17660 5540 17672
rect 4948 17632 5540 17660
rect 4948 17620 4954 17632
rect 5534 17620 5540 17632
rect 5592 17620 5598 17672
rect 6641 17663 6699 17669
rect 6641 17629 6653 17663
rect 6687 17629 6699 17663
rect 6641 17623 6699 17629
rect 2222 17552 2228 17604
rect 2280 17592 2286 17604
rect 3068 17592 3096 17620
rect 2280 17564 3096 17592
rect 2280 17552 2286 17564
rect 1946 17524 1952 17536
rect 1907 17496 1952 17524
rect 1946 17484 1952 17496
rect 2004 17484 2010 17536
rect 2409 17527 2467 17533
rect 2409 17493 2421 17527
rect 2455 17524 2467 17527
rect 2682 17524 2688 17536
rect 2455 17496 2688 17524
rect 2455 17493 2467 17496
rect 2409 17487 2467 17493
rect 2682 17484 2688 17496
rect 2740 17484 2746 17536
rect 3513 17527 3571 17533
rect 3513 17493 3525 17527
rect 3559 17524 3571 17527
rect 3602 17524 3608 17536
rect 3559 17496 3608 17524
rect 3559 17493 3571 17496
rect 3513 17487 3571 17493
rect 3602 17484 3608 17496
rect 3660 17484 3666 17536
rect 5537 17527 5595 17533
rect 5537 17493 5549 17527
rect 5583 17524 5595 17527
rect 6178 17524 6184 17536
rect 5583 17496 6184 17524
rect 5583 17493 5595 17496
rect 5537 17487 5595 17493
rect 6178 17484 6184 17496
rect 6236 17484 6242 17536
rect 6454 17524 6460 17536
rect 6415 17496 6460 17524
rect 6454 17484 6460 17496
rect 6512 17484 6518 17536
rect 6656 17524 6684 17623
rect 7834 17620 7840 17672
rect 7892 17660 7898 17672
rect 9490 17660 9496 17672
rect 7892 17632 9496 17660
rect 7892 17620 7898 17632
rect 9490 17620 9496 17632
rect 9548 17620 9554 17672
rect 11146 17660 11152 17672
rect 11107 17632 11152 17660
rect 11146 17620 11152 17632
rect 11204 17620 11210 17672
rect 10318 17592 10324 17604
rect 10279 17564 10324 17592
rect 10318 17552 10324 17564
rect 10376 17552 10382 17604
rect 6822 17524 6828 17536
rect 6656 17496 6828 17524
rect 6822 17484 6828 17496
rect 6880 17484 6886 17536
rect 7374 17484 7380 17536
rect 7432 17524 7438 17536
rect 8021 17527 8079 17533
rect 8021 17524 8033 17527
rect 7432 17496 8033 17524
rect 7432 17484 7438 17496
rect 8021 17493 8033 17496
rect 8067 17493 8079 17527
rect 12526 17524 12532 17536
rect 12487 17496 12532 17524
rect 8021 17487 8079 17493
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 13170 17484 13176 17536
rect 13228 17524 13234 17536
rect 13265 17527 13323 17533
rect 13265 17524 13277 17527
rect 13228 17496 13277 17524
rect 13228 17484 13234 17496
rect 13265 17493 13277 17496
rect 13311 17493 13323 17527
rect 13265 17487 13323 17493
rect 14093 17527 14151 17533
rect 14093 17493 14105 17527
rect 14139 17524 14151 17527
rect 14182 17524 14188 17536
rect 14139 17496 14188 17524
rect 14139 17493 14151 17496
rect 14093 17487 14151 17493
rect 14182 17484 14188 17496
rect 14240 17484 14246 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 2133 17323 2191 17329
rect 2133 17289 2145 17323
rect 2179 17320 2191 17323
rect 2222 17320 2228 17332
rect 2179 17292 2228 17320
rect 2179 17289 2191 17292
rect 2133 17283 2191 17289
rect 2222 17280 2228 17292
rect 2280 17280 2286 17332
rect 4614 17280 4620 17332
rect 4672 17320 4678 17332
rect 4893 17323 4951 17329
rect 4893 17320 4905 17323
rect 4672 17292 4905 17320
rect 4672 17280 4678 17292
rect 4893 17289 4905 17292
rect 4939 17289 4951 17323
rect 4893 17283 4951 17289
rect 5166 17280 5172 17332
rect 5224 17320 5230 17332
rect 5261 17323 5319 17329
rect 5261 17320 5273 17323
rect 5224 17292 5273 17320
rect 5224 17280 5230 17292
rect 5261 17289 5273 17292
rect 5307 17289 5319 17323
rect 5261 17283 5319 17289
rect 6273 17323 6331 17329
rect 6273 17289 6285 17323
rect 6319 17320 6331 17323
rect 6454 17320 6460 17332
rect 6319 17292 6460 17320
rect 6319 17289 6331 17292
rect 6273 17283 6331 17289
rect 6454 17280 6460 17292
rect 6512 17280 6518 17332
rect 6641 17323 6699 17329
rect 6641 17289 6653 17323
rect 6687 17320 6699 17323
rect 6822 17320 6828 17332
rect 6687 17292 6828 17320
rect 6687 17289 6699 17292
rect 6641 17283 6699 17289
rect 6822 17280 6828 17292
rect 6880 17280 6886 17332
rect 8570 17320 8576 17332
rect 8531 17292 8576 17320
rect 8570 17280 8576 17292
rect 8628 17280 8634 17332
rect 10505 17323 10563 17329
rect 10505 17289 10517 17323
rect 10551 17320 10563 17323
rect 10778 17320 10784 17332
rect 10551 17292 10784 17320
rect 10551 17289 10563 17292
rect 10505 17283 10563 17289
rect 10778 17280 10784 17292
rect 10836 17280 10842 17332
rect 12802 17320 12808 17332
rect 12763 17292 12808 17320
rect 12802 17280 12808 17292
rect 12860 17280 12866 17332
rect 13906 17280 13912 17332
rect 13964 17320 13970 17332
rect 14645 17323 14703 17329
rect 14645 17320 14657 17323
rect 13964 17292 14657 17320
rect 13964 17280 13970 17292
rect 14645 17289 14657 17292
rect 14691 17289 14703 17323
rect 14645 17283 14703 17289
rect 5626 17252 5632 17264
rect 5587 17224 5632 17252
rect 5626 17212 5632 17224
rect 5684 17212 5690 17264
rect 8297 17255 8355 17261
rect 8297 17252 8309 17255
rect 7300 17224 8309 17252
rect 7300 17193 7328 17224
rect 8297 17221 8309 17224
rect 8343 17252 8355 17255
rect 9401 17255 9459 17261
rect 9401 17252 9413 17255
rect 8343 17224 9413 17252
rect 8343 17221 8355 17224
rect 8297 17215 8355 17221
rect 9401 17221 9413 17224
rect 9447 17221 9459 17255
rect 9401 17215 9459 17221
rect 11146 17212 11152 17264
rect 11204 17252 11210 17264
rect 11241 17255 11299 17261
rect 11241 17252 11253 17255
rect 11204 17224 11253 17252
rect 11204 17212 11210 17224
rect 11241 17221 11253 17224
rect 11287 17252 11299 17255
rect 11790 17252 11796 17264
rect 11287 17224 11796 17252
rect 11287 17221 11299 17224
rect 11241 17215 11299 17221
rect 11790 17212 11796 17224
rect 11848 17252 11854 17264
rect 12710 17252 12716 17264
rect 11848 17224 12716 17252
rect 11848 17212 11854 17224
rect 12710 17212 12716 17224
rect 12768 17252 12774 17264
rect 13081 17255 13139 17261
rect 13081 17252 13093 17255
rect 12768 17224 13093 17252
rect 12768 17212 12774 17224
rect 13081 17221 13093 17224
rect 13127 17252 13139 17255
rect 13127 17224 13308 17252
rect 13127 17221 13139 17224
rect 13081 17215 13139 17221
rect 7285 17187 7343 17193
rect 7285 17153 7297 17187
rect 7331 17153 7343 17187
rect 7285 17147 7343 17153
rect 7374 17144 7380 17196
rect 7432 17184 7438 17196
rect 7929 17187 7987 17193
rect 7432 17156 7525 17184
rect 7432 17144 7438 17156
rect 7929 17153 7941 17187
rect 7975 17184 7987 17187
rect 8202 17184 8208 17196
rect 7975 17156 8208 17184
rect 7975 17153 7987 17156
rect 7929 17147 7987 17153
rect 8202 17144 8208 17156
rect 8260 17184 8266 17196
rect 9490 17184 9496 17196
rect 8260 17156 9496 17184
rect 8260 17144 8266 17156
rect 9490 17144 9496 17156
rect 9548 17184 9554 17196
rect 9953 17187 10011 17193
rect 9953 17184 9965 17187
rect 9548 17156 9965 17184
rect 9548 17144 9554 17156
rect 9953 17153 9965 17156
rect 9999 17184 10011 17187
rect 10870 17184 10876 17196
rect 9999 17156 10876 17184
rect 9999 17153 10011 17156
rect 9953 17147 10011 17153
rect 10870 17144 10876 17156
rect 10928 17144 10934 17196
rect 11333 17187 11391 17193
rect 11333 17153 11345 17187
rect 11379 17184 11391 17187
rect 12342 17184 12348 17196
rect 11379 17156 12348 17184
rect 11379 17153 11391 17156
rect 11333 17147 11391 17153
rect 12342 17144 12348 17156
rect 12400 17144 12406 17196
rect 13280 17193 13308 17224
rect 13265 17187 13323 17193
rect 13265 17153 13277 17187
rect 13311 17153 13323 17187
rect 13265 17147 13323 17153
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17116 1455 17119
rect 1946 17116 1952 17128
rect 1443 17088 1952 17116
rect 1443 17085 1455 17088
rect 1397 17079 1455 17085
rect 1946 17076 1952 17088
rect 2004 17076 2010 17128
rect 2866 17116 2872 17128
rect 2779 17088 2872 17116
rect 2866 17076 2872 17088
rect 2924 17116 2930 17128
rect 2961 17119 3019 17125
rect 2961 17116 2973 17119
rect 2924 17088 2973 17116
rect 2924 17076 2930 17088
rect 2961 17085 2973 17088
rect 3007 17116 3019 17119
rect 4062 17116 4068 17128
rect 3007 17088 4068 17116
rect 3007 17085 3019 17088
rect 2961 17079 3019 17085
rect 4062 17076 4068 17088
rect 4120 17076 4126 17128
rect 5445 17119 5503 17125
rect 5445 17085 5457 17119
rect 5491 17116 5503 17119
rect 5534 17116 5540 17128
rect 5491 17088 5540 17116
rect 5491 17085 5503 17088
rect 5445 17079 5503 17085
rect 5534 17076 5540 17088
rect 5592 17076 5598 17128
rect 6454 17076 6460 17128
rect 6512 17116 6518 17128
rect 7392 17116 7420 17144
rect 6512 17088 7420 17116
rect 8389 17119 8447 17125
rect 6512 17076 6518 17088
rect 8389 17085 8401 17119
rect 8435 17116 8447 17119
rect 8662 17116 8668 17128
rect 8435 17088 8668 17116
rect 8435 17085 8447 17088
rect 8389 17079 8447 17085
rect 8662 17076 8668 17088
rect 8720 17116 8726 17128
rect 9214 17116 9220 17128
rect 8720 17088 9220 17116
rect 8720 17076 8726 17088
rect 9214 17076 9220 17088
rect 9272 17076 9278 17128
rect 9309 17119 9367 17125
rect 9309 17085 9321 17119
rect 9355 17116 9367 17119
rect 9769 17119 9827 17125
rect 9769 17116 9781 17119
rect 9355 17088 9781 17116
rect 9355 17085 9367 17088
rect 9309 17079 9367 17085
rect 9769 17085 9781 17088
rect 9815 17116 9827 17119
rect 10042 17116 10048 17128
rect 9815 17088 10048 17116
rect 9815 17085 9827 17088
rect 9769 17079 9827 17085
rect 10042 17076 10048 17088
rect 10100 17076 10106 17128
rect 3234 17057 3240 17060
rect 2501 17051 2559 17057
rect 2501 17017 2513 17051
rect 2547 17048 2559 17051
rect 3228 17048 3240 17057
rect 2547 17020 3240 17048
rect 2547 17017 2559 17020
rect 2501 17011 2559 17017
rect 3228 17011 3240 17020
rect 3234 17008 3240 17011
rect 3292 17008 3298 17060
rect 7193 17051 7251 17057
rect 7193 17017 7205 17051
rect 7239 17048 7251 17051
rect 7650 17048 7656 17060
rect 7239 17020 7656 17048
rect 7239 17017 7251 17020
rect 7193 17011 7251 17017
rect 7650 17008 7656 17020
rect 7708 17048 7714 17060
rect 8202 17048 8208 17060
rect 7708 17020 8208 17048
rect 7708 17008 7714 17020
rect 8202 17008 8208 17020
rect 8260 17008 8266 17060
rect 8941 17051 8999 17057
rect 8941 17017 8953 17051
rect 8987 17048 8999 17051
rect 9861 17051 9919 17057
rect 9861 17048 9873 17051
rect 8987 17020 9873 17048
rect 8987 17017 8999 17020
rect 8941 17011 8999 17017
rect 9861 17017 9873 17020
rect 9907 17048 9919 17051
rect 9950 17048 9956 17060
rect 9907 17020 9956 17048
rect 9907 17017 9919 17020
rect 9861 17011 9919 17017
rect 9950 17008 9956 17020
rect 10008 17008 10014 17060
rect 13170 17008 13176 17060
rect 13228 17048 13234 17060
rect 13510 17051 13568 17057
rect 13510 17048 13522 17051
rect 13228 17020 13522 17048
rect 13228 17008 13234 17020
rect 13510 17017 13522 17020
rect 13556 17017 13568 17051
rect 13510 17011 13568 17017
rect 1486 16940 1492 16992
rect 1544 16980 1550 16992
rect 1581 16983 1639 16989
rect 1581 16980 1593 16983
rect 1544 16952 1593 16980
rect 1544 16940 1550 16952
rect 1581 16949 1593 16952
rect 1627 16949 1639 16983
rect 1581 16943 1639 16949
rect 3050 16940 3056 16992
rect 3108 16980 3114 16992
rect 4341 16983 4399 16989
rect 4341 16980 4353 16983
rect 3108 16952 4353 16980
rect 3108 16940 3114 16952
rect 4341 16949 4353 16952
rect 4387 16980 4399 16983
rect 4706 16980 4712 16992
rect 4387 16952 4712 16980
rect 4387 16949 4399 16952
rect 4341 16943 4399 16949
rect 4706 16940 4712 16952
rect 4764 16940 4770 16992
rect 6822 16980 6828 16992
rect 6783 16952 6828 16980
rect 6822 16940 6828 16952
rect 6880 16940 6886 16992
rect 11422 16940 11428 16992
rect 11480 16980 11486 16992
rect 11793 16983 11851 16989
rect 11793 16980 11805 16983
rect 11480 16952 11805 16980
rect 11480 16940 11486 16952
rect 11793 16949 11805 16952
rect 11839 16949 11851 16983
rect 11793 16943 11851 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1581 16779 1639 16785
rect 1581 16745 1593 16779
rect 1627 16776 1639 16779
rect 1670 16776 1676 16788
rect 1627 16748 1676 16776
rect 1627 16745 1639 16748
rect 1581 16739 1639 16745
rect 1670 16736 1676 16748
rect 1728 16736 1734 16788
rect 2409 16779 2467 16785
rect 2409 16745 2421 16779
rect 2455 16776 2467 16779
rect 2590 16776 2596 16788
rect 2455 16748 2596 16776
rect 2455 16745 2467 16748
rect 2409 16739 2467 16745
rect 2590 16736 2596 16748
rect 2648 16736 2654 16788
rect 3418 16776 3424 16788
rect 3379 16748 3424 16776
rect 3418 16736 3424 16748
rect 3476 16736 3482 16788
rect 3970 16736 3976 16788
rect 4028 16776 4034 16788
rect 4433 16779 4491 16785
rect 4433 16776 4445 16779
rect 4028 16748 4445 16776
rect 4028 16736 4034 16748
rect 4433 16745 4445 16748
rect 4479 16776 4491 16779
rect 5629 16779 5687 16785
rect 5629 16776 5641 16779
rect 4479 16748 5641 16776
rect 4479 16745 4491 16748
rect 4433 16739 4491 16745
rect 5629 16745 5641 16748
rect 5675 16745 5687 16779
rect 6730 16776 6736 16788
rect 6691 16748 6736 16776
rect 5629 16739 5687 16745
rect 6730 16736 6736 16748
rect 6788 16736 6794 16788
rect 7193 16779 7251 16785
rect 7193 16745 7205 16779
rect 7239 16745 7251 16779
rect 8202 16776 8208 16788
rect 8163 16748 8208 16776
rect 7193 16739 7251 16745
rect 4525 16711 4583 16717
rect 4525 16677 4537 16711
rect 4571 16708 4583 16711
rect 5166 16708 5172 16720
rect 4571 16680 5172 16708
rect 4571 16677 4583 16680
rect 4525 16671 4583 16677
rect 5166 16668 5172 16680
rect 5224 16708 5230 16720
rect 7208 16708 7236 16739
rect 8202 16736 8208 16748
rect 8260 16736 8266 16788
rect 8662 16776 8668 16788
rect 8623 16748 8668 16776
rect 8662 16736 8668 16748
rect 8720 16736 8726 16788
rect 9490 16776 9496 16788
rect 9451 16748 9496 16776
rect 9490 16736 9496 16748
rect 9548 16736 9554 16788
rect 9950 16776 9956 16788
rect 9911 16748 9956 16776
rect 9950 16736 9956 16748
rect 10008 16736 10014 16788
rect 10042 16736 10048 16788
rect 10100 16776 10106 16788
rect 10321 16779 10379 16785
rect 10321 16776 10333 16779
rect 10100 16748 10333 16776
rect 10100 16736 10106 16748
rect 10321 16745 10333 16748
rect 10367 16776 10379 16779
rect 10686 16776 10692 16788
rect 10367 16748 10692 16776
rect 10367 16745 10379 16748
rect 10321 16739 10379 16745
rect 10686 16736 10692 16748
rect 10744 16736 10750 16788
rect 11698 16776 11704 16788
rect 10888 16748 11704 16776
rect 5224 16680 7236 16708
rect 5224 16668 5230 16680
rect 7466 16668 7472 16720
rect 7524 16708 7530 16720
rect 7653 16711 7711 16717
rect 7653 16708 7665 16711
rect 7524 16680 7665 16708
rect 7524 16668 7530 16680
rect 7653 16677 7665 16680
rect 7699 16708 7711 16711
rect 7742 16708 7748 16720
rect 7699 16680 7748 16708
rect 7699 16677 7711 16680
rect 7653 16671 7711 16677
rect 7742 16668 7748 16680
rect 7800 16668 7806 16720
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16640 1455 16643
rect 2222 16640 2228 16652
rect 1443 16612 2228 16640
rect 1443 16609 1455 16612
rect 1397 16603 1455 16609
rect 2222 16600 2228 16612
rect 2280 16600 2286 16652
rect 2501 16643 2559 16649
rect 2501 16609 2513 16643
rect 2547 16640 2559 16643
rect 3053 16643 3111 16649
rect 3053 16640 3065 16643
rect 2547 16612 3065 16640
rect 2547 16609 2559 16612
rect 2501 16603 2559 16609
rect 3053 16609 3065 16612
rect 3099 16609 3111 16643
rect 3053 16603 3111 16609
rect 2038 16532 2044 16584
rect 2096 16572 2102 16584
rect 2516 16572 2544 16603
rect 3234 16600 3240 16652
rect 3292 16640 3298 16652
rect 3881 16643 3939 16649
rect 3881 16640 3893 16643
rect 3292 16612 3893 16640
rect 3292 16600 3298 16612
rect 3881 16609 3893 16612
rect 3927 16640 3939 16643
rect 4890 16640 4896 16652
rect 3927 16612 4896 16640
rect 3927 16609 3939 16612
rect 3881 16603 3939 16609
rect 4706 16572 4712 16584
rect 2096 16544 2544 16572
rect 4667 16544 4712 16572
rect 2096 16532 2102 16544
rect 4706 16532 4712 16544
rect 4764 16532 4770 16584
rect 2406 16464 2412 16516
rect 2464 16504 2470 16516
rect 2590 16504 2596 16516
rect 2464 16476 2596 16504
rect 2464 16464 2470 16476
rect 2590 16464 2596 16476
rect 2648 16464 2654 16516
rect 4816 16504 4844 16612
rect 4890 16600 4896 16612
rect 4948 16600 4954 16652
rect 4982 16600 4988 16652
rect 5040 16640 5046 16652
rect 5077 16643 5135 16649
rect 5077 16640 5089 16643
rect 5040 16612 5089 16640
rect 5040 16600 5046 16612
rect 5077 16609 5089 16612
rect 5123 16609 5135 16643
rect 5534 16640 5540 16652
rect 5495 16612 5540 16640
rect 5077 16603 5135 16609
rect 5534 16600 5540 16612
rect 5592 16600 5598 16652
rect 5994 16640 6000 16652
rect 5955 16612 6000 16640
rect 5994 16600 6000 16612
rect 6052 16600 6058 16652
rect 7561 16643 7619 16649
rect 7561 16609 7573 16643
rect 7607 16640 7619 16643
rect 7834 16640 7840 16652
rect 7607 16612 7840 16640
rect 7607 16609 7619 16612
rect 7561 16603 7619 16609
rect 7834 16600 7840 16612
rect 7892 16600 7898 16652
rect 10888 16640 10916 16748
rect 11698 16736 11704 16748
rect 11756 16736 11762 16788
rect 13078 16776 13084 16788
rect 13039 16748 13084 16776
rect 13078 16736 13084 16748
rect 13136 16736 13142 16788
rect 15746 16736 15752 16788
rect 15804 16776 15810 16788
rect 15804 16748 15849 16776
rect 15804 16736 15810 16748
rect 12526 16708 12532 16720
rect 10428 16612 10916 16640
rect 10980 16680 12532 16708
rect 6086 16572 6092 16584
rect 6047 16544 6092 16572
rect 6086 16532 6092 16544
rect 6144 16532 6150 16584
rect 6273 16575 6331 16581
rect 6273 16541 6285 16575
rect 6319 16541 6331 16575
rect 7742 16572 7748 16584
rect 7703 16544 7748 16572
rect 6273 16535 6331 16541
rect 5350 16504 5356 16516
rect 4816 16476 5356 16504
rect 5350 16464 5356 16476
rect 5408 16504 5414 16516
rect 6288 16504 6316 16535
rect 7742 16532 7748 16544
rect 7800 16532 7806 16584
rect 10226 16532 10232 16584
rect 10284 16572 10290 16584
rect 10428 16581 10456 16612
rect 10413 16575 10471 16581
rect 10413 16572 10425 16575
rect 10284 16544 10425 16572
rect 10284 16532 10290 16544
rect 10413 16541 10425 16544
rect 10459 16541 10471 16575
rect 10413 16535 10471 16541
rect 10505 16575 10563 16581
rect 10505 16541 10517 16575
rect 10551 16572 10563 16575
rect 10980 16572 11008 16680
rect 12526 16668 12532 16680
rect 12584 16668 12590 16720
rect 11701 16643 11759 16649
rect 11701 16609 11713 16643
rect 11747 16640 11759 16643
rect 11790 16640 11796 16652
rect 11747 16612 11796 16640
rect 11747 16609 11759 16612
rect 11701 16603 11759 16609
rect 11790 16600 11796 16612
rect 11848 16600 11854 16652
rect 11974 16649 11980 16652
rect 11968 16640 11980 16649
rect 11935 16612 11980 16640
rect 11968 16603 11980 16612
rect 11974 16600 11980 16603
rect 12032 16600 12038 16652
rect 15654 16640 15660 16652
rect 15615 16612 15660 16640
rect 15654 16600 15660 16612
rect 15712 16600 15718 16652
rect 15930 16572 15936 16584
rect 10551 16544 11008 16572
rect 15891 16544 15936 16572
rect 10551 16541 10563 16544
rect 10505 16535 10563 16541
rect 7760 16504 7788 16532
rect 5408 16476 7788 16504
rect 5408 16464 5414 16476
rect 9398 16464 9404 16516
rect 9456 16504 9462 16516
rect 10520 16504 10548 16535
rect 15930 16532 15936 16544
rect 15988 16532 15994 16584
rect 9456 16476 10548 16504
rect 9456 16464 9462 16476
rect 1762 16396 1768 16448
rect 1820 16436 1826 16448
rect 1949 16439 2007 16445
rect 1949 16436 1961 16439
rect 1820 16408 1961 16436
rect 1820 16396 1826 16408
rect 1949 16405 1961 16408
rect 1995 16405 2007 16439
rect 1949 16399 2007 16405
rect 2685 16439 2743 16445
rect 2685 16405 2697 16439
rect 2731 16436 2743 16439
rect 2774 16436 2780 16448
rect 2731 16408 2780 16436
rect 2731 16405 2743 16408
rect 2685 16399 2743 16405
rect 2774 16396 2780 16408
rect 2832 16396 2838 16448
rect 4062 16436 4068 16448
rect 4023 16408 4068 16436
rect 4062 16396 4068 16408
rect 4120 16396 4126 16448
rect 6914 16396 6920 16448
rect 6972 16436 6978 16448
rect 7009 16439 7067 16445
rect 7009 16436 7021 16439
rect 6972 16408 7021 16436
rect 6972 16396 6978 16408
rect 7009 16405 7021 16408
rect 7055 16405 7067 16439
rect 7009 16399 7067 16405
rect 10134 16396 10140 16448
rect 10192 16436 10198 16448
rect 10686 16436 10692 16448
rect 10192 16408 10692 16436
rect 10192 16396 10198 16408
rect 10686 16396 10692 16408
rect 10744 16396 10750 16448
rect 15286 16436 15292 16448
rect 15247 16408 15292 16436
rect 15286 16396 15292 16408
rect 15344 16396 15350 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 1854 16192 1860 16244
rect 1912 16232 1918 16244
rect 4706 16232 4712 16244
rect 1912 16204 4568 16232
rect 4667 16204 4712 16232
rect 1912 16192 1918 16204
rect 4540 16164 4568 16204
rect 4706 16192 4712 16204
rect 4764 16192 4770 16244
rect 5261 16235 5319 16241
rect 5261 16201 5273 16235
rect 5307 16232 5319 16235
rect 5350 16232 5356 16244
rect 5307 16204 5356 16232
rect 5307 16201 5319 16204
rect 5261 16195 5319 16201
rect 5350 16192 5356 16204
rect 5408 16192 5414 16244
rect 6086 16192 6092 16244
rect 6144 16232 6150 16244
rect 6181 16235 6239 16241
rect 6181 16232 6193 16235
rect 6144 16204 6193 16232
rect 6144 16192 6150 16204
rect 6181 16201 6193 16204
rect 6227 16201 6239 16235
rect 6638 16232 6644 16244
rect 6599 16204 6644 16232
rect 6181 16195 6239 16201
rect 6638 16192 6644 16204
rect 6696 16192 6702 16244
rect 8573 16235 8631 16241
rect 8573 16201 8585 16235
rect 8619 16232 8631 16235
rect 9306 16232 9312 16244
rect 8619 16204 9312 16232
rect 8619 16201 8631 16204
rect 8573 16195 8631 16201
rect 9306 16192 9312 16204
rect 9364 16192 9370 16244
rect 9769 16235 9827 16241
rect 9769 16201 9781 16235
rect 9815 16232 9827 16235
rect 10042 16232 10048 16244
rect 9815 16204 10048 16232
rect 9815 16201 9827 16204
rect 9769 16195 9827 16201
rect 10042 16192 10048 16204
rect 10100 16192 10106 16244
rect 11790 16232 11796 16244
rect 11751 16204 11796 16232
rect 11790 16192 11796 16204
rect 11848 16192 11854 16244
rect 15930 16192 15936 16244
rect 15988 16232 15994 16244
rect 16393 16235 16451 16241
rect 16393 16232 16405 16235
rect 15988 16204 16405 16232
rect 15988 16192 15994 16204
rect 16393 16201 16405 16204
rect 16439 16201 16451 16235
rect 16393 16195 16451 16201
rect 6730 16164 6736 16176
rect 4540 16136 6736 16164
rect 6730 16124 6736 16136
rect 6788 16124 6794 16176
rect 15746 16124 15752 16176
rect 15804 16164 15810 16176
rect 16025 16167 16083 16173
rect 16025 16164 16037 16167
rect 15804 16136 16037 16164
rect 15804 16124 15810 16136
rect 16025 16133 16037 16136
rect 16071 16164 16083 16167
rect 16114 16164 16120 16176
rect 16071 16136 16120 16164
rect 16071 16133 16083 16136
rect 16025 16127 16083 16133
rect 16114 16124 16120 16136
rect 16172 16124 16178 16176
rect 2314 16096 2320 16108
rect 2275 16068 2320 16096
rect 2314 16056 2320 16068
rect 2372 16096 2378 16108
rect 2372 16068 2912 16096
rect 2372 16056 2378 16068
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 1762 16028 1768 16040
rect 1443 16000 1768 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 1762 15988 1768 16000
rect 1820 15988 1826 16040
rect 2777 16031 2835 16037
rect 2777 15997 2789 16031
rect 2823 15997 2835 16031
rect 2884 16028 2912 16068
rect 9030 16056 9036 16108
rect 9088 16096 9094 16108
rect 9309 16099 9367 16105
rect 9309 16096 9321 16099
rect 9088 16068 9321 16096
rect 9088 16056 9094 16068
rect 9309 16065 9321 16068
rect 9355 16096 9367 16099
rect 9861 16099 9919 16105
rect 9861 16096 9873 16099
rect 9355 16068 9873 16096
rect 9355 16065 9367 16068
rect 9309 16059 9367 16065
rect 9861 16065 9873 16068
rect 9907 16065 9919 16099
rect 9861 16059 9919 16065
rect 3033 16031 3091 16037
rect 3033 16028 3045 16031
rect 2884 16000 3045 16028
rect 2777 15991 2835 15997
rect 3033 15997 3045 16000
rect 3079 15997 3091 16031
rect 3033 15991 3091 15997
rect 2792 15960 2820 15991
rect 6638 15988 6644 16040
rect 6696 16028 6702 16040
rect 7193 16031 7251 16037
rect 7193 16028 7205 16031
rect 6696 16000 7205 16028
rect 6696 15988 6702 16000
rect 7193 15997 7205 16000
rect 7239 16028 7251 16031
rect 7926 16028 7932 16040
rect 7239 16000 7932 16028
rect 7239 15997 7251 16000
rect 7193 15991 7251 15997
rect 7926 15988 7932 16000
rect 7984 16028 7990 16040
rect 8570 16028 8576 16040
rect 7984 16000 8576 16028
rect 7984 15988 7990 16000
rect 8570 15988 8576 16000
rect 8628 16028 8634 16040
rect 9048 16028 9076 16056
rect 8628 16000 9076 16028
rect 9876 16028 9904 16059
rect 13541 16031 13599 16037
rect 13541 16028 13553 16031
rect 9876 16000 13553 16028
rect 8628 15988 8634 16000
rect 13541 15997 13553 16000
rect 13587 16028 13599 16031
rect 13725 16031 13783 16037
rect 13725 16028 13737 16031
rect 13587 16000 13737 16028
rect 13587 15997 13599 16000
rect 13541 15991 13599 15997
rect 13725 15997 13737 16000
rect 13771 15997 13783 16031
rect 15654 16028 15660 16040
rect 13725 15991 13783 15997
rect 13832 16000 15660 16028
rect 2866 15960 2872 15972
rect 2792 15932 2872 15960
rect 1578 15892 1584 15904
rect 1539 15864 1584 15892
rect 1578 15852 1584 15864
rect 1636 15852 1642 15904
rect 2685 15895 2743 15901
rect 2685 15861 2697 15895
rect 2731 15892 2743 15895
rect 2792 15892 2820 15932
rect 2866 15920 2872 15932
rect 2924 15920 2930 15972
rect 5629 15963 5687 15969
rect 5629 15929 5641 15963
rect 5675 15960 5687 15963
rect 6086 15960 6092 15972
rect 5675 15932 6092 15960
rect 5675 15929 5687 15932
rect 5629 15923 5687 15929
rect 6086 15920 6092 15932
rect 6144 15920 6150 15972
rect 6914 15920 6920 15972
rect 6972 15960 6978 15972
rect 10134 15969 10140 15972
rect 7438 15963 7496 15969
rect 7438 15960 7450 15963
rect 6972 15932 7450 15960
rect 6972 15920 6978 15932
rect 7438 15929 7450 15932
rect 7484 15929 7496 15963
rect 7438 15923 7496 15929
rect 10128 15923 10140 15969
rect 10192 15960 10198 15972
rect 10192 15932 10228 15960
rect 10134 15920 10140 15923
rect 10192 15920 10198 15932
rect 11790 15920 11796 15972
rect 11848 15960 11854 15972
rect 13832 15960 13860 16000
rect 15654 15988 15660 16000
rect 15712 15988 15718 16040
rect 11848 15932 13860 15960
rect 11848 15920 11854 15932
rect 13906 15920 13912 15972
rect 13964 15969 13970 15972
rect 13964 15963 14028 15969
rect 13964 15929 13982 15963
rect 14016 15929 14028 15963
rect 13964 15923 14028 15929
rect 13964 15920 13970 15923
rect 2731 15864 2820 15892
rect 4157 15895 4215 15901
rect 2731 15861 2743 15864
rect 2685 15855 2743 15861
rect 4157 15861 4169 15895
rect 4203 15892 4215 15895
rect 4522 15892 4528 15904
rect 4203 15864 4528 15892
rect 4203 15861 4215 15864
rect 4157 15855 4215 15861
rect 4522 15852 4528 15864
rect 4580 15852 4586 15904
rect 5718 15892 5724 15904
rect 5679 15864 5724 15892
rect 5718 15852 5724 15864
rect 5776 15852 5782 15904
rect 7101 15895 7159 15901
rect 7101 15861 7113 15895
rect 7147 15892 7159 15895
rect 7834 15892 7840 15904
rect 7147 15864 7840 15892
rect 7147 15861 7159 15864
rect 7101 15855 7159 15861
rect 7834 15852 7840 15864
rect 7892 15852 7898 15904
rect 11241 15895 11299 15901
rect 11241 15861 11253 15895
rect 11287 15892 11299 15895
rect 11330 15892 11336 15904
rect 11287 15864 11336 15892
rect 11287 15861 11299 15864
rect 11241 15855 11299 15861
rect 11330 15852 11336 15864
rect 11388 15892 11394 15904
rect 11974 15892 11980 15904
rect 11388 15864 11980 15892
rect 11388 15852 11394 15864
rect 11974 15852 11980 15864
rect 12032 15892 12038 15904
rect 12161 15895 12219 15901
rect 12161 15892 12173 15895
rect 12032 15864 12173 15892
rect 12032 15852 12038 15864
rect 12161 15861 12173 15864
rect 12207 15861 12219 15895
rect 15102 15892 15108 15904
rect 15063 15864 15108 15892
rect 12161 15855 12219 15861
rect 15102 15852 15108 15864
rect 15160 15852 15166 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1581 15691 1639 15697
rect 1581 15657 1593 15691
rect 1627 15688 1639 15691
rect 2038 15688 2044 15700
rect 1627 15660 2044 15688
rect 1627 15657 1639 15660
rect 1581 15651 1639 15657
rect 2038 15648 2044 15660
rect 2096 15648 2102 15700
rect 2222 15688 2228 15700
rect 2183 15660 2228 15688
rect 2222 15648 2228 15660
rect 2280 15648 2286 15700
rect 2406 15688 2412 15700
rect 2367 15660 2412 15688
rect 2406 15648 2412 15660
rect 2464 15648 2470 15700
rect 2869 15691 2927 15697
rect 2869 15657 2881 15691
rect 2915 15688 2927 15691
rect 3513 15691 3571 15697
rect 3513 15688 3525 15691
rect 2915 15660 3525 15688
rect 2915 15657 2927 15660
rect 2869 15651 2927 15657
rect 3513 15657 3525 15660
rect 3559 15688 3571 15691
rect 4062 15688 4068 15700
rect 3559 15660 4068 15688
rect 3559 15657 3571 15660
rect 3513 15651 3571 15657
rect 4062 15648 4068 15660
rect 4120 15648 4126 15700
rect 4246 15688 4252 15700
rect 4207 15660 4252 15688
rect 4246 15648 4252 15660
rect 4304 15648 4310 15700
rect 4617 15691 4675 15697
rect 4617 15657 4629 15691
rect 4663 15688 4675 15691
rect 5166 15688 5172 15700
rect 4663 15660 5172 15688
rect 4663 15657 4675 15660
rect 4617 15651 4675 15657
rect 5166 15648 5172 15660
rect 5224 15648 5230 15700
rect 5261 15691 5319 15697
rect 5261 15657 5273 15691
rect 5307 15688 5319 15691
rect 5534 15688 5540 15700
rect 5307 15660 5540 15688
rect 5307 15657 5319 15660
rect 5261 15651 5319 15657
rect 5534 15648 5540 15660
rect 5592 15688 5598 15700
rect 5718 15688 5724 15700
rect 5592 15660 5724 15688
rect 5592 15648 5598 15660
rect 5718 15648 5724 15660
rect 5776 15648 5782 15700
rect 7742 15648 7748 15700
rect 7800 15688 7806 15700
rect 8113 15691 8171 15697
rect 8113 15688 8125 15691
rect 7800 15660 8125 15688
rect 7800 15648 7806 15660
rect 8113 15657 8125 15660
rect 8159 15657 8171 15691
rect 9398 15688 9404 15700
rect 9359 15660 9404 15688
rect 8113 15651 8171 15657
rect 9398 15648 9404 15660
rect 9456 15648 9462 15700
rect 10134 15648 10140 15700
rect 10192 15688 10198 15700
rect 10321 15691 10379 15697
rect 10321 15688 10333 15691
rect 10192 15660 10333 15688
rect 10192 15648 10198 15660
rect 10321 15657 10333 15660
rect 10367 15657 10379 15691
rect 10778 15688 10784 15700
rect 10739 15660 10784 15688
rect 10321 15651 10379 15657
rect 10778 15648 10784 15660
rect 10836 15648 10842 15700
rect 11238 15688 11244 15700
rect 11151 15660 11244 15688
rect 11238 15648 11244 15660
rect 11296 15688 11302 15700
rect 12345 15691 12403 15697
rect 12345 15688 12357 15691
rect 11296 15660 12357 15688
rect 11296 15648 11302 15660
rect 12345 15657 12357 15660
rect 12391 15657 12403 15691
rect 12345 15651 12403 15657
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 12802 15688 12808 15700
rect 12492 15660 12808 15688
rect 12492 15648 12498 15660
rect 12802 15648 12808 15660
rect 12860 15648 12866 15700
rect 13817 15691 13875 15697
rect 13817 15657 13829 15691
rect 13863 15688 13875 15691
rect 13906 15688 13912 15700
rect 13863 15660 13912 15688
rect 13863 15657 13875 15660
rect 13817 15651 13875 15657
rect 3881 15623 3939 15629
rect 3881 15589 3893 15623
rect 3927 15620 3939 15623
rect 3970 15620 3976 15632
rect 3927 15592 3976 15620
rect 3927 15589 3939 15592
rect 3881 15583 3939 15589
rect 3970 15580 3976 15592
rect 4028 15580 4034 15632
rect 5994 15580 6000 15632
rect 6052 15629 6058 15632
rect 6052 15623 6116 15629
rect 6052 15589 6070 15623
rect 6104 15589 6116 15623
rect 6052 15583 6116 15589
rect 7837 15623 7895 15629
rect 7837 15589 7849 15623
rect 7883 15620 7895 15623
rect 7926 15620 7932 15632
rect 7883 15592 7932 15620
rect 7883 15589 7895 15592
rect 7837 15583 7895 15589
rect 6052 15580 6058 15583
rect 7926 15580 7932 15592
rect 7984 15580 7990 15632
rect 11149 15623 11207 15629
rect 11149 15589 11161 15623
rect 11195 15620 11207 15623
rect 11514 15620 11520 15632
rect 11195 15592 11520 15620
rect 11195 15589 11207 15592
rect 11149 15583 11207 15589
rect 11514 15580 11520 15592
rect 11572 15580 11578 15632
rect 13832 15620 13860 15651
rect 13906 15648 13912 15660
rect 13964 15648 13970 15700
rect 14369 15691 14427 15697
rect 14369 15657 14381 15691
rect 14415 15688 14427 15691
rect 14550 15688 14556 15700
rect 14415 15660 14556 15688
rect 14415 15657 14427 15660
rect 14369 15651 14427 15657
rect 14550 15648 14556 15660
rect 14608 15648 14614 15700
rect 15746 15620 15752 15632
rect 13372 15592 13860 15620
rect 15707 15592 15752 15620
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15552 1455 15555
rect 1949 15555 2007 15561
rect 1949 15552 1961 15555
rect 1443 15524 1961 15552
rect 1443 15521 1455 15524
rect 1397 15515 1455 15521
rect 1949 15521 1961 15524
rect 1995 15552 2007 15555
rect 2038 15552 2044 15564
rect 1995 15524 2044 15552
rect 1995 15521 2007 15524
rect 1949 15515 2007 15521
rect 2038 15512 2044 15524
rect 2096 15512 2102 15564
rect 2682 15512 2688 15564
rect 2740 15552 2746 15564
rect 2777 15555 2835 15561
rect 2777 15552 2789 15555
rect 2740 15524 2789 15552
rect 2740 15512 2746 15524
rect 2777 15521 2789 15524
rect 2823 15552 2835 15555
rect 3786 15552 3792 15564
rect 2823 15524 3792 15552
rect 2823 15521 2835 15524
rect 2777 15515 2835 15521
rect 3786 15512 3792 15524
rect 3844 15512 3850 15564
rect 4062 15552 4068 15564
rect 4023 15524 4068 15552
rect 4062 15512 4068 15524
rect 4120 15512 4126 15564
rect 5813 15555 5871 15561
rect 5813 15521 5825 15555
rect 5859 15552 5871 15555
rect 6638 15552 6644 15564
rect 5859 15524 6644 15552
rect 5859 15521 5871 15524
rect 5813 15515 5871 15521
rect 6638 15512 6644 15524
rect 6696 15512 6702 15564
rect 12710 15552 12716 15564
rect 12671 15524 12716 15552
rect 12710 15512 12716 15524
rect 12768 15512 12774 15564
rect 2590 15444 2596 15496
rect 2648 15484 2654 15496
rect 3053 15487 3111 15493
rect 3053 15484 3065 15487
rect 2648 15456 3065 15484
rect 2648 15444 2654 15456
rect 3053 15453 3065 15456
rect 3099 15484 3111 15487
rect 4522 15484 4528 15496
rect 3099 15456 4528 15484
rect 3099 15453 3111 15456
rect 3053 15447 3111 15453
rect 4522 15444 4528 15456
rect 4580 15444 4586 15496
rect 8573 15487 8631 15493
rect 8573 15453 8585 15487
rect 8619 15484 8631 15487
rect 9858 15484 9864 15496
rect 8619 15456 9864 15484
rect 8619 15453 8631 15456
rect 8573 15447 8631 15453
rect 9858 15444 9864 15456
rect 9916 15444 9922 15496
rect 10962 15444 10968 15496
rect 11020 15484 11026 15496
rect 11422 15484 11428 15496
rect 11020 15456 11428 15484
rect 11020 15444 11026 15456
rect 11422 15444 11428 15456
rect 11480 15444 11486 15496
rect 12989 15487 13047 15493
rect 12989 15453 13001 15487
rect 13035 15484 13047 15487
rect 13078 15484 13084 15496
rect 13035 15456 13084 15484
rect 13035 15453 13047 15456
rect 12989 15447 13047 15453
rect 13078 15444 13084 15456
rect 13136 15484 13142 15496
rect 13372 15484 13400 15592
rect 15746 15580 15752 15592
rect 15804 15580 15810 15632
rect 13814 15512 13820 15564
rect 13872 15552 13878 15564
rect 14185 15555 14243 15561
rect 14185 15552 14197 15555
rect 13872 15524 14197 15552
rect 13872 15512 13878 15524
rect 14185 15521 14197 15524
rect 14231 15552 14243 15555
rect 14645 15555 14703 15561
rect 14645 15552 14657 15555
rect 14231 15524 14657 15552
rect 14231 15521 14243 15524
rect 14185 15515 14243 15521
rect 14645 15521 14657 15524
rect 14691 15521 14703 15555
rect 14645 15515 14703 15521
rect 15657 15555 15715 15561
rect 15657 15521 15669 15555
rect 15703 15552 15715 15555
rect 15930 15552 15936 15564
rect 15703 15524 15936 15552
rect 15703 15521 15715 15524
rect 15657 15515 15715 15521
rect 15930 15512 15936 15524
rect 15988 15512 15994 15564
rect 15838 15484 15844 15496
rect 13136 15456 13400 15484
rect 15799 15456 15844 15484
rect 13136 15444 13142 15456
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 3234 15376 3240 15428
rect 3292 15416 3298 15428
rect 9033 15419 9091 15425
rect 9033 15416 9045 15419
rect 3292 15388 5663 15416
rect 3292 15376 3298 15388
rect 5442 15308 5448 15360
rect 5500 15348 5506 15360
rect 5537 15351 5595 15357
rect 5537 15348 5549 15351
rect 5500 15320 5549 15348
rect 5500 15308 5506 15320
rect 5537 15317 5549 15320
rect 5583 15317 5595 15351
rect 5635 15348 5663 15388
rect 6748 15388 9045 15416
rect 6748 15348 6776 15388
rect 9033 15385 9045 15388
rect 9079 15385 9091 15419
rect 10042 15416 10048 15428
rect 10003 15388 10048 15416
rect 9033 15379 9091 15385
rect 10042 15376 10048 15388
rect 10100 15376 10106 15428
rect 5635 15320 6776 15348
rect 5537 15311 5595 15317
rect 6914 15308 6920 15360
rect 6972 15348 6978 15360
rect 7193 15351 7251 15357
rect 7193 15348 7205 15351
rect 6972 15320 7205 15348
rect 6972 15308 6978 15320
rect 7193 15317 7205 15320
rect 7239 15317 7251 15351
rect 7193 15311 7251 15317
rect 14458 15308 14464 15360
rect 14516 15348 14522 15360
rect 15289 15351 15347 15357
rect 15289 15348 15301 15351
rect 14516 15320 15301 15348
rect 14516 15308 14522 15320
rect 15289 15317 15301 15320
rect 15335 15317 15347 15351
rect 15289 15311 15347 15317
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1949 15147 2007 15153
rect 1949 15113 1961 15147
rect 1995 15144 2007 15147
rect 2590 15144 2596 15156
rect 1995 15116 2596 15144
rect 1995 15113 2007 15116
rect 1949 15107 2007 15113
rect 2590 15104 2596 15116
rect 2648 15104 2654 15156
rect 3881 15147 3939 15153
rect 3881 15113 3893 15147
rect 3927 15144 3939 15147
rect 4062 15144 4068 15156
rect 3927 15116 4068 15144
rect 3927 15113 3939 15116
rect 3881 15107 3939 15113
rect 4062 15104 4068 15116
rect 4120 15104 4126 15156
rect 6086 15104 6092 15156
rect 6144 15144 6150 15156
rect 6914 15144 6920 15156
rect 6144 15116 6920 15144
rect 6144 15104 6150 15116
rect 6914 15104 6920 15116
rect 6972 15104 6978 15156
rect 8570 15144 8576 15156
rect 8531 15116 8576 15144
rect 8570 15104 8576 15116
rect 8628 15104 8634 15156
rect 10134 15144 10140 15156
rect 10095 15116 10140 15144
rect 10134 15104 10140 15116
rect 10192 15104 10198 15156
rect 10873 15147 10931 15153
rect 10873 15113 10885 15147
rect 10919 15144 10931 15147
rect 10962 15144 10968 15156
rect 10919 15116 10968 15144
rect 10919 15113 10931 15116
rect 10873 15107 10931 15113
rect 10962 15104 10968 15116
rect 11020 15104 11026 15156
rect 11238 15144 11244 15156
rect 11199 15116 11244 15144
rect 11238 15104 11244 15116
rect 11296 15104 11302 15156
rect 11514 15144 11520 15156
rect 11475 15116 11520 15144
rect 11514 15104 11520 15116
rect 11572 15104 11578 15156
rect 12253 15147 12311 15153
rect 12253 15113 12265 15147
rect 12299 15144 12311 15147
rect 12342 15144 12348 15156
rect 12299 15116 12348 15144
rect 12299 15113 12311 15116
rect 12253 15107 12311 15113
rect 12342 15104 12348 15116
rect 12400 15104 12406 15156
rect 13078 15144 13084 15156
rect 13039 15116 13084 15144
rect 13078 15104 13084 15116
rect 13136 15104 13142 15156
rect 1581 15079 1639 15085
rect 1581 15045 1593 15079
rect 1627 15076 1639 15079
rect 3970 15076 3976 15088
rect 1627 15048 3976 15076
rect 1627 15045 1639 15048
rect 1581 15039 1639 15045
rect 3970 15036 3976 15048
rect 4028 15036 4034 15088
rect 6273 15079 6331 15085
rect 6273 15045 6285 15079
rect 6319 15076 6331 15079
rect 6638 15076 6644 15088
rect 6319 15048 6644 15076
rect 6319 15045 6331 15048
rect 6273 15039 6331 15045
rect 6638 15036 6644 15048
rect 6696 15036 6702 15088
rect 2866 15008 2872 15020
rect 2827 14980 2872 15008
rect 2866 14968 2872 14980
rect 2924 14968 2930 15020
rect 3053 15011 3111 15017
rect 3053 14977 3065 15011
rect 3099 15008 3111 15011
rect 3510 15008 3516 15020
rect 3099 14980 3516 15008
rect 3099 14977 3111 14980
rect 3053 14971 3111 14977
rect 3510 14968 3516 14980
rect 3568 14968 3574 15020
rect 4709 15011 4767 15017
rect 4709 14977 4721 15011
rect 4755 15008 4767 15011
rect 5721 15011 5779 15017
rect 5721 15008 5733 15011
rect 4755 14980 5733 15008
rect 4755 14977 4767 14980
rect 4709 14971 4767 14977
rect 5721 14977 5733 14980
rect 5767 15008 5779 15011
rect 5994 15008 6000 15020
rect 5767 14980 6000 15008
rect 5767 14977 5779 14980
rect 5721 14971 5779 14977
rect 5994 14968 6000 14980
rect 6052 15008 6058 15020
rect 7377 15011 7435 15017
rect 7377 15008 7389 15011
rect 6052 14980 7389 15008
rect 6052 14968 6058 14980
rect 7377 14977 7389 14980
rect 7423 15008 7435 15011
rect 7837 15011 7895 15017
rect 7837 15008 7849 15011
rect 7423 14980 7849 15008
rect 7423 14977 7435 14980
rect 7377 14971 7435 14977
rect 7837 14977 7849 14980
rect 7883 15008 7895 15011
rect 7926 15008 7932 15020
rect 7883 14980 7932 15008
rect 7883 14977 7895 14980
rect 7837 14971 7895 14977
rect 7926 14968 7932 14980
rect 7984 14968 7990 15020
rect 8297 15011 8355 15017
rect 8297 14977 8309 15011
rect 8343 15008 8355 15011
rect 8343 14980 8892 15008
rect 8343 14977 8355 14980
rect 8297 14971 8355 14977
rect 1394 14940 1400 14952
rect 1355 14912 1400 14940
rect 1394 14900 1400 14912
rect 1452 14900 1458 14952
rect 3970 14940 3976 14952
rect 3931 14912 3976 14940
rect 3970 14900 3976 14912
rect 4028 14900 4034 14952
rect 5534 14940 5540 14952
rect 5495 14912 5540 14940
rect 5534 14900 5540 14912
rect 5592 14900 5598 14952
rect 5629 14943 5687 14949
rect 5629 14909 5641 14943
rect 5675 14940 5687 14943
rect 6454 14940 6460 14952
rect 5675 14912 6460 14940
rect 5675 14909 5687 14912
rect 5629 14903 5687 14909
rect 2317 14875 2375 14881
rect 2317 14841 2329 14875
rect 2363 14872 2375 14875
rect 2774 14872 2780 14884
rect 2363 14844 2780 14872
rect 2363 14841 2375 14844
rect 2317 14835 2375 14841
rect 2774 14832 2780 14844
rect 2832 14832 2838 14884
rect 5077 14875 5135 14881
rect 5077 14841 5089 14875
rect 5123 14872 5135 14875
rect 5644 14872 5672 14903
rect 6454 14900 6460 14912
rect 6512 14900 6518 14952
rect 6641 14943 6699 14949
rect 6641 14909 6653 14943
rect 6687 14940 6699 14943
rect 7190 14940 7196 14952
rect 6687 14912 7196 14940
rect 6687 14909 6699 14912
rect 6641 14903 6699 14909
rect 7190 14900 7196 14912
rect 7248 14900 7254 14952
rect 8570 14900 8576 14952
rect 8628 14940 8634 14952
rect 8757 14943 8815 14949
rect 8757 14940 8769 14943
rect 8628 14912 8769 14940
rect 8628 14900 8634 14912
rect 8757 14909 8769 14912
rect 8803 14909 8815 14943
rect 8864 14940 8892 14980
rect 9024 14943 9082 14949
rect 9024 14940 9036 14943
rect 8864 14912 9036 14940
rect 8757 14903 8815 14909
rect 9024 14909 9036 14912
rect 9070 14940 9082 14943
rect 9306 14940 9312 14952
rect 9070 14912 9312 14940
rect 9070 14909 9082 14912
rect 9024 14903 9082 14909
rect 9306 14900 9312 14912
rect 9364 14900 9370 14952
rect 12802 14900 12808 14952
rect 12860 14940 12866 14952
rect 13817 14943 13875 14949
rect 13817 14940 13829 14943
rect 12860 14912 13829 14940
rect 12860 14900 12866 14912
rect 13817 14909 13829 14912
rect 13863 14940 13875 14943
rect 13909 14943 13967 14949
rect 13909 14940 13921 14943
rect 13863 14912 13921 14940
rect 13863 14909 13875 14912
rect 13817 14903 13875 14909
rect 13909 14909 13921 14912
rect 13955 14909 13967 14943
rect 13909 14903 13967 14909
rect 12710 14872 12716 14884
rect 5123 14844 5672 14872
rect 12623 14844 12716 14872
rect 5123 14841 5135 14844
rect 5077 14835 5135 14841
rect 12710 14832 12716 14844
rect 12768 14872 12774 14884
rect 13262 14872 13268 14884
rect 12768 14844 13268 14872
rect 12768 14832 12774 14844
rect 13262 14832 13268 14844
rect 13320 14832 13326 14884
rect 13446 14872 13452 14884
rect 13359 14844 13452 14872
rect 13446 14832 13452 14844
rect 13504 14872 13510 14884
rect 14090 14872 14096 14884
rect 13504 14844 14096 14872
rect 13504 14832 13510 14844
rect 14090 14832 14096 14844
rect 14148 14881 14154 14884
rect 14148 14875 14212 14881
rect 14148 14841 14166 14875
rect 14200 14841 14212 14875
rect 14148 14835 14212 14841
rect 14148 14832 14154 14835
rect 2409 14807 2467 14813
rect 2409 14773 2421 14807
rect 2455 14804 2467 14807
rect 3142 14804 3148 14816
rect 2455 14776 3148 14804
rect 2455 14773 2467 14776
rect 2409 14767 2467 14773
rect 3142 14764 3148 14776
rect 3200 14764 3206 14816
rect 3510 14804 3516 14816
rect 3471 14776 3516 14804
rect 3510 14764 3516 14776
rect 3568 14764 3574 14816
rect 4154 14804 4160 14816
rect 4115 14776 4160 14804
rect 4154 14764 4160 14776
rect 4212 14764 4218 14816
rect 5169 14807 5227 14813
rect 5169 14773 5181 14807
rect 5215 14804 5227 14807
rect 5442 14804 5448 14816
rect 5215 14776 5448 14804
rect 5215 14773 5227 14776
rect 5169 14767 5227 14773
rect 5442 14764 5448 14776
rect 5500 14764 5506 14816
rect 6822 14804 6828 14816
rect 6783 14776 6828 14804
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 7282 14764 7288 14816
rect 7340 14804 7346 14816
rect 7340 14776 7385 14804
rect 7340 14764 7346 14776
rect 14918 14764 14924 14816
rect 14976 14804 14982 14816
rect 15289 14807 15347 14813
rect 15289 14804 15301 14807
rect 14976 14776 15301 14804
rect 14976 14764 14982 14776
rect 15289 14773 15301 14776
rect 15335 14804 15347 14807
rect 15378 14804 15384 14816
rect 15335 14776 15384 14804
rect 15335 14773 15347 14776
rect 15289 14767 15347 14773
rect 15378 14764 15384 14776
rect 15436 14764 15442 14816
rect 15746 14764 15752 14816
rect 15804 14804 15810 14816
rect 15841 14807 15899 14813
rect 15841 14804 15853 14807
rect 15804 14776 15853 14804
rect 15804 14764 15810 14776
rect 15841 14773 15853 14776
rect 15887 14773 15899 14807
rect 15841 14767 15899 14773
rect 15930 14764 15936 14816
rect 15988 14804 15994 14816
rect 16209 14807 16267 14813
rect 16209 14804 16221 14807
rect 15988 14776 16221 14804
rect 15988 14764 15994 14776
rect 16209 14773 16221 14776
rect 16255 14773 16267 14807
rect 16666 14804 16672 14816
rect 16627 14776 16672 14804
rect 16209 14767 16267 14773
rect 16666 14764 16672 14776
rect 16724 14764 16730 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1581 14603 1639 14609
rect 1581 14569 1593 14603
rect 1627 14600 1639 14603
rect 2222 14600 2228 14612
rect 1627 14572 2228 14600
rect 1627 14569 1639 14572
rect 1581 14563 1639 14569
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 3786 14600 3792 14612
rect 3747 14572 3792 14600
rect 3786 14560 3792 14572
rect 3844 14560 3850 14612
rect 5994 14600 6000 14612
rect 5955 14572 6000 14600
rect 5994 14560 6000 14572
rect 6052 14560 6058 14612
rect 7926 14600 7932 14612
rect 7887 14572 7932 14600
rect 7926 14560 7932 14572
rect 7984 14560 7990 14612
rect 9674 14600 9680 14612
rect 9635 14572 9680 14600
rect 9674 14560 9680 14572
rect 9732 14560 9738 14612
rect 14090 14600 14096 14612
rect 14051 14572 14096 14600
rect 14090 14560 14096 14572
rect 14148 14560 14154 14612
rect 14918 14600 14924 14612
rect 14879 14572 14924 14600
rect 14918 14560 14924 14572
rect 14976 14560 14982 14612
rect 2866 14532 2872 14544
rect 2827 14504 2872 14532
rect 2866 14492 2872 14504
rect 2924 14492 2930 14544
rect 4332 14535 4390 14541
rect 4332 14501 4344 14535
rect 4378 14532 4390 14535
rect 4522 14532 4528 14544
rect 4378 14504 4528 14532
rect 4378 14501 4390 14504
rect 4332 14495 4390 14501
rect 4522 14492 4528 14504
rect 4580 14492 4586 14544
rect 15562 14492 15568 14544
rect 15620 14532 15626 14544
rect 15749 14535 15807 14541
rect 15749 14532 15761 14535
rect 15620 14504 15761 14532
rect 15620 14492 15626 14504
rect 15749 14501 15761 14504
rect 15795 14501 15807 14535
rect 15749 14495 15807 14501
rect 15838 14492 15844 14544
rect 15896 14492 15902 14544
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14464 1455 14467
rect 2406 14464 2412 14476
rect 1443 14436 2412 14464
rect 1443 14433 1455 14436
rect 1397 14427 1455 14433
rect 2406 14424 2412 14436
rect 2464 14424 2470 14476
rect 2777 14467 2835 14473
rect 2777 14433 2789 14467
rect 2823 14464 2835 14467
rect 3234 14464 3240 14476
rect 2823 14436 3240 14464
rect 2823 14433 2835 14436
rect 2777 14427 2835 14433
rect 2498 14356 2504 14408
rect 2556 14396 2562 14408
rect 2792 14396 2820 14427
rect 3234 14424 3240 14436
rect 3292 14424 3298 14476
rect 4062 14464 4068 14476
rect 3975 14436 4068 14464
rect 4062 14424 4068 14436
rect 4120 14464 4126 14476
rect 4120 14436 5120 14464
rect 4120 14424 4126 14436
rect 2556 14368 2820 14396
rect 3053 14399 3111 14405
rect 2556 14356 2562 14368
rect 3053 14365 3065 14399
rect 3099 14396 3111 14399
rect 3510 14396 3516 14408
rect 3099 14368 3516 14396
rect 3099 14365 3111 14368
rect 3053 14359 3111 14365
rect 3510 14356 3516 14368
rect 3568 14396 3574 14408
rect 3786 14396 3792 14408
rect 3568 14368 3792 14396
rect 3568 14356 3574 14368
rect 3786 14356 3792 14368
rect 3844 14356 3850 14408
rect 5092 14396 5120 14436
rect 6178 14424 6184 14476
rect 6236 14464 6242 14476
rect 6805 14467 6863 14473
rect 6805 14464 6817 14467
rect 6236 14436 6817 14464
rect 6236 14424 6242 14436
rect 6805 14433 6817 14436
rect 6851 14433 6863 14467
rect 6805 14427 6863 14433
rect 10045 14467 10103 14473
rect 10045 14433 10057 14467
rect 10091 14464 10103 14467
rect 10318 14464 10324 14476
rect 10091 14436 10324 14464
rect 10091 14433 10103 14436
rect 10045 14427 10103 14433
rect 10318 14424 10324 14436
rect 10376 14464 10382 14476
rect 10689 14467 10747 14473
rect 10689 14464 10701 14467
rect 10376 14436 10701 14464
rect 10376 14424 10382 14436
rect 10689 14433 10701 14436
rect 10735 14433 10747 14467
rect 10689 14427 10747 14433
rect 12250 14424 12256 14476
rect 12308 14464 12314 14476
rect 12969 14467 13027 14473
rect 12969 14464 12981 14467
rect 12308 14436 12981 14464
rect 12308 14424 12314 14436
rect 12969 14433 12981 14436
rect 13015 14464 13027 14467
rect 13538 14464 13544 14476
rect 13015 14436 13544 14464
rect 13015 14433 13027 14436
rect 12969 14427 13027 14433
rect 13538 14424 13544 14436
rect 13596 14424 13602 14476
rect 15654 14464 15660 14476
rect 15615 14436 15660 14464
rect 15654 14424 15660 14436
rect 15712 14424 15718 14476
rect 6454 14396 6460 14408
rect 5092 14368 6460 14396
rect 6454 14356 6460 14368
rect 6512 14396 6518 14408
rect 6549 14399 6607 14405
rect 6549 14396 6561 14399
rect 6512 14368 6561 14396
rect 6512 14356 6518 14368
rect 6549 14365 6561 14368
rect 6595 14365 6607 14399
rect 6549 14359 6607 14365
rect 9493 14399 9551 14405
rect 9493 14365 9505 14399
rect 9539 14396 9551 14399
rect 9674 14396 9680 14408
rect 9539 14368 9680 14396
rect 9539 14365 9551 14368
rect 9493 14359 9551 14365
rect 9674 14356 9680 14368
rect 9732 14396 9738 14408
rect 10137 14399 10195 14405
rect 10137 14396 10149 14399
rect 9732 14368 10149 14396
rect 9732 14356 9738 14368
rect 10137 14365 10149 14368
rect 10183 14365 10195 14399
rect 10137 14359 10195 14365
rect 10229 14399 10287 14405
rect 10229 14365 10241 14399
rect 10275 14396 10287 14399
rect 11330 14396 11336 14408
rect 10275 14368 11336 14396
rect 10275 14365 10287 14368
rect 10229 14359 10287 14365
rect 11330 14356 11336 14368
rect 11388 14356 11394 14408
rect 12710 14396 12716 14408
rect 12671 14368 12716 14396
rect 12710 14356 12716 14368
rect 12768 14356 12774 14408
rect 13906 14356 13912 14408
rect 13964 14396 13970 14408
rect 15856 14396 15884 14492
rect 15933 14399 15991 14405
rect 15933 14396 15945 14399
rect 13964 14368 15945 14396
rect 13964 14356 13970 14368
rect 15933 14365 15945 14368
rect 15979 14396 15991 14399
rect 16666 14396 16672 14408
rect 15979 14368 16672 14396
rect 15979 14365 15991 14368
rect 15933 14359 15991 14365
rect 16666 14356 16672 14368
rect 16724 14356 16730 14408
rect 12253 14331 12311 14337
rect 12253 14297 12265 14331
rect 12299 14328 12311 14331
rect 12434 14328 12440 14340
rect 12299 14300 12440 14328
rect 12299 14297 12311 14300
rect 12253 14291 12311 14297
rect 12434 14288 12440 14300
rect 12492 14288 12498 14340
rect 1946 14260 1952 14272
rect 1907 14232 1952 14260
rect 1946 14220 1952 14232
rect 2004 14220 2010 14272
rect 2222 14260 2228 14272
rect 2183 14232 2228 14260
rect 2222 14220 2228 14232
rect 2280 14220 2286 14272
rect 2409 14263 2467 14269
rect 2409 14229 2421 14263
rect 2455 14260 2467 14263
rect 2958 14260 2964 14272
rect 2455 14232 2964 14260
rect 2455 14229 2467 14232
rect 2409 14223 2467 14229
rect 2958 14220 2964 14232
rect 3016 14220 3022 14272
rect 5445 14263 5503 14269
rect 5445 14229 5457 14263
rect 5491 14260 5503 14263
rect 5534 14260 5540 14272
rect 5491 14232 5540 14260
rect 5491 14229 5503 14232
rect 5445 14223 5503 14229
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 6457 14263 6515 14269
rect 6457 14229 6469 14263
rect 6503 14260 6515 14263
rect 7282 14260 7288 14272
rect 6503 14232 7288 14260
rect 6503 14229 6515 14232
rect 6457 14223 6515 14229
rect 7282 14220 7288 14232
rect 7340 14220 7346 14272
rect 8846 14260 8852 14272
rect 8807 14232 8852 14260
rect 8846 14220 8852 14232
rect 8904 14220 8910 14272
rect 11885 14263 11943 14269
rect 11885 14229 11897 14263
rect 11931 14260 11943 14263
rect 12158 14260 12164 14272
rect 11931 14232 12164 14260
rect 11931 14229 11943 14232
rect 11885 14223 11943 14229
rect 12158 14220 12164 14232
rect 12216 14220 12222 14272
rect 12526 14260 12532 14272
rect 12487 14232 12532 14260
rect 12526 14220 12532 14232
rect 12584 14220 12590 14272
rect 15289 14263 15347 14269
rect 15289 14229 15301 14263
rect 15335 14260 15347 14263
rect 15470 14260 15476 14272
rect 15335 14232 15476 14260
rect 15335 14229 15347 14232
rect 15289 14223 15347 14229
rect 15470 14220 15476 14232
rect 15528 14220 15534 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 3326 14056 3332 14068
rect 1627 14028 3332 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 3326 14016 3332 14028
rect 3384 14016 3390 14068
rect 4062 14016 4068 14068
rect 4120 14056 4126 14068
rect 4157 14059 4215 14065
rect 4157 14056 4169 14059
rect 4120 14028 4169 14056
rect 4120 14016 4126 14028
rect 4157 14025 4169 14028
rect 4203 14025 4215 14059
rect 4522 14056 4528 14068
rect 4483 14028 4528 14056
rect 4157 14019 4215 14025
rect 4522 14016 4528 14028
rect 4580 14016 4586 14068
rect 5166 14056 5172 14068
rect 5127 14028 5172 14056
rect 5166 14016 5172 14028
rect 5224 14016 5230 14068
rect 5534 14016 5540 14068
rect 5592 14056 5598 14068
rect 6178 14056 6184 14068
rect 5592 14028 6184 14056
rect 5592 14016 5598 14028
rect 6178 14016 6184 14028
rect 6236 14016 6242 14068
rect 6454 14016 6460 14068
rect 6512 14056 6518 14068
rect 6638 14056 6644 14068
rect 6512 14028 6644 14056
rect 6512 14016 6518 14028
rect 6638 14016 6644 14028
rect 6696 14016 6702 14068
rect 7193 14059 7251 14065
rect 7193 14025 7205 14059
rect 7239 14056 7251 14059
rect 7282 14056 7288 14068
rect 7239 14028 7288 14056
rect 7239 14025 7251 14028
rect 7193 14019 7251 14025
rect 7282 14016 7288 14028
rect 7340 14016 7346 14068
rect 8478 14016 8484 14068
rect 8536 14056 8542 14068
rect 8573 14059 8631 14065
rect 8573 14056 8585 14059
rect 8536 14028 8585 14056
rect 8536 14016 8542 14028
rect 8573 14025 8585 14028
rect 8619 14025 8631 14059
rect 9858 14056 9864 14068
rect 9819 14028 9864 14056
rect 8573 14019 8631 14025
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 10042 14016 10048 14068
rect 10100 14056 10106 14068
rect 10137 14059 10195 14065
rect 10137 14056 10149 14059
rect 10100 14028 10149 14056
rect 10100 14016 10106 14028
rect 10137 14025 10149 14028
rect 10183 14025 10195 14059
rect 10318 14056 10324 14068
rect 10279 14028 10324 14056
rect 10137 14019 10195 14025
rect 10318 14016 10324 14028
rect 10376 14016 10382 14068
rect 11330 14056 11336 14068
rect 11291 14028 11336 14056
rect 11330 14016 11336 14028
rect 11388 14016 11394 14068
rect 12250 14056 12256 14068
rect 12211 14028 12256 14056
rect 12250 14016 12256 14028
rect 12308 14016 12314 14068
rect 12710 14056 12716 14068
rect 12671 14028 12716 14056
rect 12710 14016 12716 14028
rect 12768 14016 12774 14068
rect 13265 14059 13323 14065
rect 13265 14025 13277 14059
rect 13311 14056 13323 14059
rect 13814 14056 13820 14068
rect 13311 14028 13820 14056
rect 13311 14025 13323 14028
rect 13265 14019 13323 14025
rect 13814 14016 13820 14028
rect 13872 14016 13878 14068
rect 13906 14016 13912 14068
rect 13964 14056 13970 14068
rect 14277 14059 14335 14065
rect 14277 14056 14289 14059
rect 13964 14028 14289 14056
rect 13964 14016 13970 14028
rect 14277 14025 14289 14028
rect 14323 14025 14335 14059
rect 14277 14019 14335 14025
rect 3145 13991 3203 13997
rect 3145 13957 3157 13991
rect 3191 13988 3203 13991
rect 3191 13960 4108 13988
rect 3191 13957 3203 13960
rect 3145 13951 3203 13957
rect 2222 13920 2228 13932
rect 2183 13892 2228 13920
rect 2222 13880 2228 13892
rect 2280 13880 2286 13932
rect 3694 13920 3700 13932
rect 3655 13892 3700 13920
rect 3694 13880 3700 13892
rect 3752 13880 3758 13932
rect 2038 13852 2044 13864
rect 1999 13824 2044 13852
rect 2038 13812 2044 13824
rect 2096 13812 2102 13864
rect 2685 13855 2743 13861
rect 2685 13821 2697 13855
rect 2731 13852 2743 13855
rect 3050 13852 3056 13864
rect 2731 13824 2912 13852
rect 2963 13824 3056 13852
rect 2731 13821 2743 13824
rect 2685 13815 2743 13821
rect 2884 13784 2912 13824
rect 3050 13812 3056 13824
rect 3108 13852 3114 13864
rect 3602 13852 3608 13864
rect 3108 13824 3608 13852
rect 3108 13812 3114 13824
rect 3602 13812 3608 13824
rect 3660 13812 3666 13864
rect 3510 13784 3516 13796
rect 2884 13756 3516 13784
rect 3510 13744 3516 13756
rect 3568 13744 3574 13796
rect 4080 13784 4108 13960
rect 5077 13923 5135 13929
rect 5077 13889 5089 13923
rect 5123 13920 5135 13923
rect 5721 13923 5779 13929
rect 5721 13920 5733 13923
rect 5123 13892 5733 13920
rect 5123 13889 5135 13892
rect 5077 13883 5135 13889
rect 5721 13889 5733 13892
rect 5767 13920 5779 13923
rect 6086 13920 6092 13932
rect 5767 13892 6092 13920
rect 5767 13889 5779 13892
rect 5721 13883 5779 13889
rect 6086 13880 6092 13892
rect 6144 13880 6150 13932
rect 6196 13920 6224 14016
rect 8754 13948 8760 14000
rect 8812 13988 8818 14000
rect 9306 13988 9312 14000
rect 8812 13960 9312 13988
rect 8812 13948 8818 13960
rect 9306 13948 9312 13960
rect 9364 13948 9370 14000
rect 12728 13988 12756 14016
rect 14553 13991 14611 13997
rect 14553 13988 14565 13991
rect 12728 13960 14565 13988
rect 14553 13957 14565 13960
rect 14599 13988 14611 13991
rect 14645 13991 14703 13997
rect 14645 13988 14657 13991
rect 14599 13960 14657 13988
rect 14599 13957 14611 13960
rect 14553 13951 14611 13957
rect 14645 13957 14657 13960
rect 14691 13957 14703 13991
rect 14645 13951 14703 13957
rect 7558 13920 7564 13932
rect 6196 13892 7564 13920
rect 7558 13880 7564 13892
rect 7616 13920 7622 13932
rect 7745 13923 7803 13929
rect 7745 13920 7757 13923
rect 7616 13892 7757 13920
rect 7616 13880 7622 13892
rect 7745 13889 7757 13892
rect 7791 13889 7803 13923
rect 9398 13920 9404 13932
rect 9359 13892 9404 13920
rect 7745 13883 7803 13889
rect 9398 13880 9404 13892
rect 9456 13880 9462 13932
rect 10134 13880 10140 13932
rect 10192 13920 10198 13932
rect 10686 13920 10692 13932
rect 10192 13892 10692 13920
rect 10192 13880 10198 13892
rect 10686 13880 10692 13892
rect 10744 13920 10750 13932
rect 10873 13923 10931 13929
rect 10873 13920 10885 13923
rect 10744 13892 10885 13920
rect 10744 13880 10750 13892
rect 10873 13889 10885 13892
rect 10919 13889 10931 13923
rect 10873 13883 10931 13889
rect 13173 13923 13231 13929
rect 13173 13889 13185 13923
rect 13219 13920 13231 13923
rect 13909 13923 13967 13929
rect 13909 13920 13921 13923
rect 13219 13892 13921 13920
rect 13219 13889 13231 13892
rect 13173 13883 13231 13889
rect 13909 13889 13921 13892
rect 13955 13920 13967 13923
rect 13955 13892 14964 13920
rect 13955 13889 13967 13892
rect 13909 13883 13967 13889
rect 5629 13855 5687 13861
rect 5629 13821 5641 13855
rect 5675 13852 5687 13855
rect 5902 13852 5908 13864
rect 5675 13824 5908 13852
rect 5675 13821 5687 13824
rect 5629 13815 5687 13821
rect 5902 13812 5908 13824
rect 5960 13852 5966 13864
rect 6822 13852 6828 13864
rect 5960 13824 6828 13852
rect 5960 13812 5966 13824
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 7653 13855 7711 13861
rect 7653 13821 7665 13855
rect 7699 13852 7711 13855
rect 7926 13852 7932 13864
rect 7699 13824 7932 13852
rect 7699 13821 7711 13824
rect 7653 13815 7711 13821
rect 7926 13812 7932 13824
rect 7984 13812 7990 13864
rect 8846 13812 8852 13864
rect 8904 13852 8910 13864
rect 9125 13855 9183 13861
rect 9125 13852 9137 13855
rect 8904 13824 9137 13852
rect 8904 13812 8910 13824
rect 9125 13821 9137 13824
rect 9171 13821 9183 13855
rect 9125 13815 9183 13821
rect 10042 13812 10048 13864
rect 10100 13852 10106 13864
rect 10781 13855 10839 13861
rect 10781 13852 10793 13855
rect 10100 13824 10793 13852
rect 10100 13812 10106 13824
rect 10781 13821 10793 13824
rect 10827 13821 10839 13855
rect 10781 13815 10839 13821
rect 14553 13855 14611 13861
rect 14553 13821 14565 13855
rect 14599 13852 14611 13855
rect 14829 13855 14887 13861
rect 14829 13852 14841 13855
rect 14599 13824 14841 13852
rect 14599 13821 14611 13824
rect 14553 13815 14611 13821
rect 14829 13821 14841 13824
rect 14875 13821 14887 13855
rect 14936 13852 14964 13892
rect 15096 13855 15154 13861
rect 15096 13852 15108 13855
rect 14936 13824 15108 13852
rect 14829 13815 14887 13821
rect 15096 13821 15108 13824
rect 15142 13852 15154 13855
rect 15378 13852 15384 13864
rect 15142 13824 15384 13852
rect 15142 13821 15154 13824
rect 15096 13815 15154 13821
rect 15378 13812 15384 13824
rect 15436 13812 15442 13864
rect 15562 13812 15568 13864
rect 15620 13852 15626 13864
rect 16761 13855 16819 13861
rect 16761 13852 16773 13855
rect 15620 13824 16773 13852
rect 15620 13812 15626 13824
rect 16761 13821 16773 13824
rect 16807 13821 16819 13855
rect 16761 13815 16819 13821
rect 4890 13784 4896 13796
rect 4080 13756 4896 13784
rect 4890 13744 4896 13756
rect 4948 13744 4954 13796
rect 5534 13784 5540 13796
rect 5495 13756 5540 13784
rect 5534 13744 5540 13756
rect 5592 13744 5598 13796
rect 8478 13744 8484 13796
rect 8536 13784 8542 13796
rect 9214 13784 9220 13796
rect 8536 13756 9220 13784
rect 8536 13744 8542 13756
rect 9214 13744 9220 13756
rect 9272 13744 9278 13796
rect 9858 13744 9864 13796
rect 9916 13784 9922 13796
rect 10689 13787 10747 13793
rect 10689 13784 10701 13787
rect 9916 13756 10701 13784
rect 9916 13744 9922 13756
rect 10689 13753 10701 13756
rect 10735 13753 10747 13787
rect 10689 13747 10747 13753
rect 11146 13744 11152 13796
rect 11204 13784 11210 13796
rect 11793 13787 11851 13793
rect 11793 13784 11805 13787
rect 11204 13756 11805 13784
rect 11204 13744 11210 13756
rect 11793 13753 11805 13756
rect 11839 13753 11851 13787
rect 11793 13747 11851 13753
rect 12526 13744 12532 13796
rect 12584 13784 12590 13796
rect 13633 13787 13691 13793
rect 13633 13784 13645 13787
rect 12584 13756 13645 13784
rect 12584 13744 12590 13756
rect 13633 13753 13645 13756
rect 13679 13753 13691 13787
rect 13633 13747 13691 13753
rect 1949 13719 2007 13725
rect 1949 13685 1961 13719
rect 1995 13716 2007 13719
rect 2038 13716 2044 13728
rect 1995 13688 2044 13716
rect 1995 13685 2007 13688
rect 1949 13679 2007 13685
rect 2038 13676 2044 13688
rect 2096 13676 2102 13728
rect 7101 13719 7159 13725
rect 7101 13685 7113 13719
rect 7147 13716 7159 13719
rect 7374 13716 7380 13728
rect 7147 13688 7380 13716
rect 7147 13685 7159 13688
rect 7101 13679 7159 13685
rect 7374 13676 7380 13688
rect 7432 13716 7438 13728
rect 7561 13719 7619 13725
rect 7561 13716 7573 13719
rect 7432 13688 7573 13716
rect 7432 13676 7438 13688
rect 7561 13685 7573 13688
rect 7607 13685 7619 13719
rect 8294 13716 8300 13728
rect 8255 13688 8300 13716
rect 7561 13679 7619 13685
rect 8294 13676 8300 13688
rect 8352 13676 8358 13728
rect 8754 13716 8760 13728
rect 8715 13688 8760 13716
rect 8754 13676 8760 13688
rect 8812 13676 8818 13728
rect 13722 13676 13728 13728
rect 13780 13716 13786 13728
rect 16206 13716 16212 13728
rect 13780 13688 13825 13716
rect 16167 13688 16212 13716
rect 13780 13676 13786 13688
rect 16206 13676 16212 13688
rect 16264 13676 16270 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 2869 13515 2927 13521
rect 2869 13481 2881 13515
rect 2915 13512 2927 13515
rect 3050 13512 3056 13524
rect 2915 13484 3056 13512
rect 2915 13481 2927 13484
rect 2869 13475 2927 13481
rect 3050 13472 3056 13484
rect 3108 13472 3114 13524
rect 3510 13512 3516 13524
rect 3423 13484 3516 13512
rect 3510 13472 3516 13484
rect 3568 13512 3574 13524
rect 3694 13512 3700 13524
rect 3568 13484 3700 13512
rect 3568 13472 3574 13484
rect 3694 13472 3700 13484
rect 3752 13472 3758 13524
rect 3970 13472 3976 13524
rect 4028 13512 4034 13524
rect 4249 13515 4307 13521
rect 4249 13512 4261 13515
rect 4028 13484 4261 13512
rect 4028 13472 4034 13484
rect 4249 13481 4261 13484
rect 4295 13481 4307 13515
rect 4249 13475 4307 13481
rect 4338 13472 4344 13524
rect 4396 13512 4402 13524
rect 4614 13512 4620 13524
rect 4396 13484 4620 13512
rect 4396 13472 4402 13484
rect 4614 13472 4620 13484
rect 4672 13512 4678 13524
rect 4801 13515 4859 13521
rect 4801 13512 4813 13515
rect 4672 13484 4813 13512
rect 4672 13472 4678 13484
rect 4801 13481 4813 13484
rect 4847 13481 4859 13515
rect 5534 13512 5540 13524
rect 5495 13484 5540 13512
rect 4801 13475 4859 13481
rect 5534 13472 5540 13484
rect 5592 13472 5598 13524
rect 5902 13512 5908 13524
rect 5863 13484 5908 13512
rect 5902 13472 5908 13484
rect 5960 13472 5966 13524
rect 5997 13515 6055 13521
rect 5997 13481 6009 13515
rect 6043 13512 6055 13515
rect 6546 13512 6552 13524
rect 6043 13484 6552 13512
rect 6043 13481 6055 13484
rect 5997 13475 6055 13481
rect 6546 13472 6552 13484
rect 6604 13472 6610 13524
rect 7558 13512 7564 13524
rect 7519 13484 7564 13512
rect 7558 13472 7564 13484
rect 7616 13472 7622 13524
rect 8386 13472 8392 13524
rect 8444 13512 8450 13524
rect 8938 13512 8944 13524
rect 8444 13484 8944 13512
rect 8444 13472 8450 13484
rect 8938 13472 8944 13484
rect 8996 13472 9002 13524
rect 9674 13512 9680 13524
rect 9635 13484 9680 13512
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 9950 13472 9956 13524
rect 10008 13512 10014 13524
rect 10137 13515 10195 13521
rect 10137 13512 10149 13515
rect 10008 13484 10149 13512
rect 10008 13472 10014 13484
rect 10137 13481 10149 13484
rect 10183 13481 10195 13515
rect 10686 13512 10692 13524
rect 10647 13484 10692 13512
rect 10137 13475 10195 13481
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 11793 13515 11851 13521
rect 11793 13481 11805 13515
rect 11839 13512 11851 13515
rect 13265 13515 13323 13521
rect 13265 13512 13277 13515
rect 11839 13484 13277 13512
rect 11839 13481 11851 13484
rect 11793 13475 11851 13481
rect 13265 13481 13277 13484
rect 13311 13512 13323 13515
rect 13722 13512 13728 13524
rect 13311 13484 13728 13512
rect 13311 13481 13323 13484
rect 13265 13475 13323 13481
rect 13722 13472 13728 13484
rect 13780 13472 13786 13524
rect 13817 13515 13875 13521
rect 13817 13481 13829 13515
rect 13863 13512 13875 13515
rect 13998 13512 14004 13524
rect 13863 13484 14004 13512
rect 13863 13481 13875 13484
rect 13817 13475 13875 13481
rect 13998 13472 14004 13484
rect 14056 13512 14062 13524
rect 15470 13512 15476 13524
rect 14056 13484 15476 13512
rect 14056 13472 14062 13484
rect 15470 13472 15476 13484
rect 15528 13472 15534 13524
rect 15654 13472 15660 13524
rect 15712 13472 15718 13524
rect 16666 13512 16672 13524
rect 16627 13484 16672 13512
rect 16666 13472 16672 13484
rect 16724 13472 16730 13524
rect 17310 13512 17316 13524
rect 17271 13484 17316 13512
rect 17310 13472 17316 13484
rect 17368 13472 17374 13524
rect 7285 13447 7343 13453
rect 4908 13416 7236 13444
rect 1394 13376 1400 13388
rect 1355 13348 1400 13376
rect 1394 13336 1400 13348
rect 1452 13336 1458 13388
rect 2317 13379 2375 13385
rect 2317 13345 2329 13379
rect 2363 13376 2375 13379
rect 2682 13376 2688 13388
rect 2363 13348 2688 13376
rect 2363 13345 2375 13348
rect 2317 13339 2375 13345
rect 2682 13336 2688 13348
rect 2740 13376 2746 13388
rect 2777 13379 2835 13385
rect 2777 13376 2789 13379
rect 2740 13348 2789 13376
rect 2740 13336 2746 13348
rect 2777 13345 2789 13348
rect 2823 13345 2835 13379
rect 2777 13339 2835 13345
rect 3694 13336 3700 13388
rect 3752 13376 3758 13388
rect 4908 13385 4936 13416
rect 4893 13379 4951 13385
rect 4893 13376 4905 13379
rect 3752 13348 4905 13376
rect 3752 13336 3758 13348
rect 4893 13345 4905 13348
rect 4939 13345 4951 13379
rect 4893 13339 4951 13345
rect 5350 13336 5356 13388
rect 5408 13376 5414 13388
rect 6362 13376 6368 13388
rect 5408 13348 6368 13376
rect 5408 13336 5414 13348
rect 6362 13336 6368 13348
rect 6420 13336 6426 13388
rect 7208 13376 7236 13416
rect 7285 13413 7297 13447
rect 7331 13444 7343 13447
rect 7926 13444 7932 13456
rect 7331 13416 7932 13444
rect 7331 13413 7343 13416
rect 7285 13407 7343 13413
rect 7926 13404 7932 13416
rect 7984 13404 7990 13456
rect 11054 13444 11060 13456
rect 11015 13416 11060 13444
rect 11054 13404 11060 13416
rect 11112 13404 11118 13456
rect 12158 13444 12164 13456
rect 12119 13416 12164 13444
rect 12158 13404 12164 13416
rect 12216 13404 12222 13456
rect 12802 13404 12808 13456
rect 12860 13444 12866 13456
rect 15105 13447 15163 13453
rect 15105 13444 15117 13447
rect 12860 13416 15117 13444
rect 12860 13404 12866 13416
rect 15105 13413 15117 13416
rect 15151 13444 15163 13447
rect 15672 13444 15700 13472
rect 15151 13416 15700 13444
rect 17221 13447 17279 13453
rect 15151 13413 15163 13416
rect 15105 13407 15163 13413
rect 17221 13413 17233 13447
rect 17267 13444 17279 13447
rect 17402 13444 17408 13456
rect 17267 13416 17408 13444
rect 17267 13413 17279 13416
rect 17221 13407 17279 13413
rect 17402 13404 17408 13416
rect 17460 13404 17466 13456
rect 8386 13376 8392 13388
rect 7208 13348 8392 13376
rect 8386 13336 8392 13348
rect 8444 13336 8450 13388
rect 9030 13336 9036 13388
rect 9088 13376 9094 13388
rect 10045 13379 10103 13385
rect 10045 13376 10057 13379
rect 9088 13348 10057 13376
rect 9088 13336 9094 13348
rect 10045 13345 10057 13348
rect 10091 13376 10103 13379
rect 11514 13376 11520 13388
rect 10091 13348 11520 13376
rect 10091 13345 10103 13348
rect 10045 13339 10103 13345
rect 11514 13336 11520 13348
rect 11572 13336 11578 13388
rect 13722 13376 13728 13388
rect 13683 13348 13728 13376
rect 13722 13336 13728 13348
rect 13780 13376 13786 13388
rect 14369 13379 14427 13385
rect 14369 13376 14381 13379
rect 13780 13348 14381 13376
rect 13780 13336 13786 13348
rect 14369 13345 14381 13348
rect 14415 13345 14427 13379
rect 14369 13339 14427 13345
rect 14550 13336 14556 13388
rect 14608 13376 14614 13388
rect 15562 13376 15568 13388
rect 14608 13348 15568 13376
rect 14608 13336 14614 13348
rect 15562 13336 15568 13348
rect 15620 13376 15626 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 15620 13348 15669 13376
rect 15620 13336 15626 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 15746 13336 15752 13388
rect 15804 13376 15810 13388
rect 15804 13348 15897 13376
rect 15804 13336 15810 13348
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13308 3111 13311
rect 5077 13311 5135 13317
rect 3099 13280 3924 13308
rect 3099 13277 3111 13280
rect 3053 13271 3111 13277
rect 1581 13243 1639 13249
rect 1581 13209 1593 13243
rect 1627 13240 1639 13243
rect 1762 13240 1768 13252
rect 1627 13212 1768 13240
rect 1627 13209 1639 13212
rect 1581 13203 1639 13209
rect 1762 13200 1768 13212
rect 1820 13200 1826 13252
rect 1949 13243 2007 13249
rect 1949 13209 1961 13243
rect 1995 13240 2007 13243
rect 2038 13240 2044 13252
rect 1995 13212 2044 13240
rect 1995 13209 2007 13212
rect 1949 13203 2007 13209
rect 2038 13200 2044 13212
rect 2096 13240 2102 13252
rect 3234 13240 3240 13252
rect 2096 13212 3240 13240
rect 2096 13200 2102 13212
rect 3234 13200 3240 13212
rect 3292 13200 3298 13252
rect 3896 13249 3924 13280
rect 5077 13277 5089 13311
rect 5123 13308 5135 13311
rect 5534 13308 5540 13320
rect 5123 13280 5540 13308
rect 5123 13277 5135 13280
rect 5077 13271 5135 13277
rect 3881 13243 3939 13249
rect 3881 13209 3893 13243
rect 3927 13240 3939 13243
rect 5092 13240 5120 13271
rect 5534 13268 5540 13280
rect 5592 13268 5598 13320
rect 6454 13308 6460 13320
rect 6415 13280 6460 13308
rect 6454 13268 6460 13280
rect 6512 13268 6518 13320
rect 6546 13268 6552 13320
rect 6604 13308 6610 13320
rect 6604 13280 6649 13308
rect 6604 13268 6610 13280
rect 6730 13268 6736 13320
rect 6788 13308 6794 13320
rect 7926 13308 7932 13320
rect 6788 13280 7932 13308
rect 6788 13268 6794 13280
rect 7926 13268 7932 13280
rect 7984 13308 7990 13320
rect 8478 13308 8484 13320
rect 7984 13280 8484 13308
rect 7984 13268 7990 13280
rect 8478 13268 8484 13280
rect 8536 13268 8542 13320
rect 8665 13311 8723 13317
rect 8665 13277 8677 13311
rect 8711 13308 8723 13311
rect 10321 13311 10379 13317
rect 8711 13280 9260 13308
rect 8711 13277 8723 13280
rect 8665 13271 8723 13277
rect 3927 13212 5120 13240
rect 3927 13209 3939 13212
rect 3881 13203 3939 13209
rect 8202 13200 8208 13252
rect 8260 13240 8266 13252
rect 8680 13240 8708 13271
rect 8260 13212 8708 13240
rect 8260 13200 8266 13212
rect 2406 13172 2412 13184
rect 2367 13144 2412 13172
rect 2406 13132 2412 13144
rect 2464 13132 2470 13184
rect 4430 13172 4436 13184
rect 4391 13144 4436 13172
rect 4430 13132 4436 13144
rect 4488 13132 4494 13184
rect 8018 13172 8024 13184
rect 7979 13144 8024 13172
rect 8018 13132 8024 13144
rect 8076 13132 8082 13184
rect 9232 13181 9260 13280
rect 10321 13277 10333 13311
rect 10367 13308 10379 13311
rect 10686 13308 10692 13320
rect 10367 13280 10692 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 10686 13268 10692 13280
rect 10744 13268 10750 13320
rect 11146 13268 11152 13320
rect 11204 13308 11210 13320
rect 12253 13311 12311 13317
rect 12253 13308 12265 13311
rect 11204 13280 12265 13308
rect 11204 13268 11210 13280
rect 12253 13277 12265 13280
rect 12299 13277 12311 13311
rect 12253 13271 12311 13277
rect 12437 13311 12495 13317
rect 12437 13277 12449 13311
rect 12483 13308 12495 13311
rect 13446 13308 13452 13320
rect 12483 13280 13452 13308
rect 12483 13277 12495 13280
rect 12437 13271 12495 13277
rect 13446 13268 13452 13280
rect 13504 13268 13510 13320
rect 13538 13268 13544 13320
rect 13596 13308 13602 13320
rect 13909 13311 13967 13317
rect 13909 13308 13921 13311
rect 13596 13280 13921 13308
rect 13596 13268 13602 13280
rect 13909 13277 13921 13280
rect 13955 13277 13967 13311
rect 13909 13271 13967 13277
rect 14734 13268 14740 13320
rect 14792 13308 14798 13320
rect 15764 13308 15792 13336
rect 14792 13280 15792 13308
rect 15933 13311 15991 13317
rect 14792 13268 14798 13280
rect 15933 13277 15945 13311
rect 15979 13308 15991 13311
rect 16206 13308 16212 13320
rect 15979 13280 16212 13308
rect 15979 13277 15991 13280
rect 15933 13271 15991 13277
rect 16206 13268 16212 13280
rect 16264 13308 16270 13320
rect 16301 13311 16359 13317
rect 16301 13308 16313 13311
rect 16264 13280 16313 13308
rect 16264 13268 16270 13280
rect 16301 13277 16313 13280
rect 16347 13277 16359 13311
rect 16301 13271 16359 13277
rect 16666 13268 16672 13320
rect 16724 13308 16730 13320
rect 17405 13311 17463 13317
rect 17405 13308 17417 13311
rect 16724 13280 17417 13308
rect 16724 13268 16730 13280
rect 17405 13277 17417 13280
rect 17451 13308 17463 13311
rect 17678 13308 17684 13320
rect 17451 13280 17684 13308
rect 17451 13277 17463 13280
rect 17405 13271 17463 13277
rect 17678 13268 17684 13280
rect 17736 13268 17742 13320
rect 12158 13200 12164 13252
rect 12216 13240 12222 13252
rect 13357 13243 13415 13249
rect 13357 13240 13369 13243
rect 12216 13212 13369 13240
rect 12216 13200 12222 13212
rect 13357 13209 13369 13212
rect 13403 13209 13415 13243
rect 13357 13203 13415 13209
rect 15562 13200 15568 13252
rect 15620 13240 15626 13252
rect 16022 13240 16028 13252
rect 15620 13212 16028 13240
rect 15620 13200 15626 13212
rect 16022 13200 16028 13212
rect 16080 13200 16086 13252
rect 9217 13175 9275 13181
rect 9217 13141 9229 13175
rect 9263 13172 9275 13175
rect 9398 13172 9404 13184
rect 9263 13144 9404 13172
rect 9263 13141 9275 13144
rect 9217 13135 9275 13141
rect 9398 13132 9404 13144
rect 9456 13132 9462 13184
rect 11422 13172 11428 13184
rect 11383 13144 11428 13172
rect 11422 13132 11428 13144
rect 11480 13132 11486 13184
rect 12894 13172 12900 13184
rect 12855 13144 12900 13172
rect 12894 13132 12900 13144
rect 12952 13132 12958 13184
rect 15289 13175 15347 13181
rect 15289 13141 15301 13175
rect 15335 13172 15347 13175
rect 15838 13172 15844 13184
rect 15335 13144 15844 13172
rect 15335 13141 15347 13144
rect 15289 13135 15347 13141
rect 15838 13132 15844 13144
rect 15896 13132 15902 13184
rect 16758 13132 16764 13184
rect 16816 13172 16822 13184
rect 16853 13175 16911 13181
rect 16853 13172 16865 13175
rect 16816 13144 16865 13172
rect 16816 13132 16822 13144
rect 16853 13141 16865 13144
rect 16899 13141 16911 13175
rect 16853 13135 16911 13141
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 2038 12928 2044 12980
rect 2096 12968 2102 12980
rect 2314 12968 2320 12980
rect 2096 12940 2320 12968
rect 2096 12928 2102 12940
rect 2314 12928 2320 12940
rect 2372 12928 2378 12980
rect 3694 12928 3700 12980
rect 3752 12968 3758 12980
rect 4341 12971 4399 12977
rect 4341 12968 4353 12971
rect 3752 12940 4353 12968
rect 3752 12928 3758 12940
rect 4341 12937 4353 12940
rect 4387 12937 4399 12971
rect 4341 12931 4399 12937
rect 6089 12971 6147 12977
rect 6089 12937 6101 12971
rect 6135 12968 6147 12971
rect 6546 12968 6552 12980
rect 6135 12940 6552 12968
rect 6135 12937 6147 12940
rect 6089 12931 6147 12937
rect 6546 12928 6552 12940
rect 6604 12928 6610 12980
rect 7926 12928 7932 12980
rect 7984 12968 7990 12980
rect 8021 12971 8079 12977
rect 8021 12968 8033 12971
rect 7984 12940 8033 12968
rect 7984 12928 7990 12940
rect 8021 12937 8033 12940
rect 8067 12937 8079 12971
rect 8386 12968 8392 12980
rect 8347 12940 8392 12968
rect 8021 12931 8079 12937
rect 8386 12928 8392 12940
rect 8444 12928 8450 12980
rect 9030 12968 9036 12980
rect 8991 12940 9036 12968
rect 9030 12928 9036 12940
rect 9088 12928 9094 12980
rect 10686 12928 10692 12980
rect 10744 12968 10750 12980
rect 11057 12971 11115 12977
rect 11057 12968 11069 12971
rect 10744 12940 11069 12968
rect 10744 12928 10750 12940
rect 11057 12937 11069 12940
rect 11103 12937 11115 12971
rect 12526 12968 12532 12980
rect 12487 12940 12532 12968
rect 11057 12931 11115 12937
rect 12526 12928 12532 12940
rect 12584 12928 12590 12980
rect 13538 12968 13544 12980
rect 13499 12940 13544 12968
rect 13538 12928 13544 12940
rect 13596 12928 13602 12980
rect 13998 12968 14004 12980
rect 13959 12940 14004 12968
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 14550 12968 14556 12980
rect 14511 12940 14556 12968
rect 14550 12928 14556 12940
rect 14608 12928 14614 12980
rect 14734 12928 14740 12980
rect 14792 12968 14798 12980
rect 14921 12971 14979 12977
rect 14921 12968 14933 12971
rect 14792 12940 14933 12968
rect 14792 12928 14798 12940
rect 14921 12937 14933 12940
rect 14967 12937 14979 12971
rect 17402 12968 17408 12980
rect 17363 12940 17408 12968
rect 14921 12931 14979 12937
rect 17402 12928 17408 12940
rect 17460 12928 17466 12980
rect 4062 12900 4068 12912
rect 4023 12872 4068 12900
rect 4062 12860 4068 12872
rect 4120 12860 4126 12912
rect 6454 12860 6460 12912
rect 6512 12900 6518 12912
rect 6825 12903 6883 12909
rect 6825 12900 6837 12903
rect 6512 12872 6837 12900
rect 6512 12860 6518 12872
rect 6825 12869 6837 12872
rect 6871 12869 6883 12903
rect 6825 12863 6883 12869
rect 12176 12872 13216 12900
rect 4982 12832 4988 12844
rect 4943 12804 4988 12832
rect 4982 12792 4988 12804
rect 5040 12792 5046 12844
rect 5166 12832 5172 12844
rect 5127 12804 5172 12832
rect 5166 12792 5172 12804
rect 5224 12792 5230 12844
rect 6641 12835 6699 12841
rect 6641 12801 6653 12835
rect 6687 12832 6699 12835
rect 6730 12832 6736 12844
rect 6687 12804 6736 12832
rect 6687 12801 6699 12804
rect 6641 12795 6699 12801
rect 6730 12792 6736 12804
rect 6788 12832 6794 12844
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 6788 12804 7389 12832
rect 6788 12792 6794 12804
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 8662 12792 8668 12844
rect 8720 12832 8726 12844
rect 9122 12832 9128 12844
rect 8720 12804 9128 12832
rect 8720 12792 8726 12804
rect 9122 12792 9128 12804
rect 9180 12792 9186 12844
rect 2041 12767 2099 12773
rect 2041 12764 2053 12767
rect 1872 12736 2053 12764
rect 1872 12640 1900 12736
rect 2041 12733 2053 12736
rect 2087 12733 2099 12767
rect 4890 12764 4896 12776
rect 4851 12736 4896 12764
rect 2041 12727 2099 12733
rect 4890 12724 4896 12736
rect 4948 12724 4954 12776
rect 9398 12773 9404 12776
rect 9392 12764 9404 12773
rect 9359 12736 9404 12764
rect 9392 12727 9404 12736
rect 9398 12724 9404 12727
rect 9456 12724 9462 12776
rect 9950 12724 9956 12776
rect 10008 12764 10014 12776
rect 11425 12767 11483 12773
rect 11425 12764 11437 12767
rect 10008 12736 11437 12764
rect 10008 12724 10014 12736
rect 11425 12733 11437 12736
rect 11471 12733 11483 12767
rect 11425 12727 11483 12733
rect 2308 12699 2366 12705
rect 2308 12665 2320 12699
rect 2354 12696 2366 12699
rect 2682 12696 2688 12708
rect 2354 12668 2688 12696
rect 2354 12665 2366 12668
rect 2308 12659 2366 12665
rect 2682 12656 2688 12668
rect 2740 12656 2746 12708
rect 12176 12705 12204 12872
rect 12434 12792 12440 12844
rect 12492 12832 12498 12844
rect 13188 12841 13216 12872
rect 12989 12835 13047 12841
rect 12989 12832 13001 12835
rect 12492 12804 13001 12832
rect 12492 12792 12498 12804
rect 12989 12801 13001 12804
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 13173 12835 13231 12841
rect 13173 12801 13185 12835
rect 13219 12832 13231 12835
rect 13446 12832 13452 12844
rect 13219 12804 13452 12832
rect 13219 12801 13231 12804
rect 13173 12795 13231 12801
rect 13446 12792 13452 12804
rect 13504 12792 13510 12844
rect 15194 12792 15200 12844
rect 15252 12832 15258 12844
rect 17865 12835 17923 12841
rect 15252 12804 15608 12832
rect 15252 12792 15258 12804
rect 12894 12764 12900 12776
rect 12855 12736 12900 12764
rect 12894 12724 12900 12736
rect 12952 12724 12958 12776
rect 15473 12767 15531 12773
rect 15473 12733 15485 12767
rect 15519 12733 15531 12767
rect 15580 12764 15608 12804
rect 17865 12801 17877 12835
rect 17911 12832 17923 12835
rect 17911 12804 18184 12832
rect 17911 12801 17923 12804
rect 17865 12795 17923 12801
rect 15729 12767 15787 12773
rect 15729 12764 15741 12767
rect 15580 12736 15741 12764
rect 15473 12727 15531 12733
rect 15729 12733 15741 12736
rect 15775 12764 15787 12767
rect 16206 12764 16212 12776
rect 15775 12736 16212 12764
rect 15775 12733 15787 12736
rect 15729 12727 15787 12733
rect 11885 12699 11943 12705
rect 11885 12665 11897 12699
rect 11931 12696 11943 12699
rect 12161 12699 12219 12705
rect 12161 12696 12173 12699
rect 11931 12668 12173 12696
rect 11931 12665 11943 12668
rect 11885 12659 11943 12665
rect 12161 12665 12173 12668
rect 12207 12665 12219 12699
rect 12161 12659 12219 12665
rect 15381 12699 15439 12705
rect 15381 12665 15393 12699
rect 15427 12696 15439 12699
rect 15488 12696 15516 12727
rect 16206 12724 16212 12736
rect 16264 12724 16270 12776
rect 18046 12764 18052 12776
rect 18007 12736 18052 12764
rect 18046 12724 18052 12736
rect 18104 12724 18110 12776
rect 18156 12764 18184 12804
rect 18322 12773 18328 12776
rect 18316 12764 18328 12773
rect 18156 12736 18328 12764
rect 18316 12727 18328 12736
rect 18322 12724 18328 12727
rect 18380 12724 18386 12776
rect 16482 12696 16488 12708
rect 15427 12668 16488 12696
rect 15427 12665 15439 12668
rect 15381 12659 15439 12665
rect 16482 12656 16488 12668
rect 16540 12696 16546 12708
rect 18064 12696 18092 12724
rect 16540 12668 18092 12696
rect 16540 12656 16546 12668
rect 1854 12628 1860 12640
rect 1815 12600 1860 12628
rect 1854 12588 1860 12600
rect 1912 12588 1918 12640
rect 3418 12628 3424 12640
rect 3379 12600 3424 12628
rect 3418 12588 3424 12600
rect 3476 12588 3482 12640
rect 4522 12628 4528 12640
rect 4483 12600 4528 12628
rect 4522 12588 4528 12600
rect 4580 12588 4586 12640
rect 5626 12628 5632 12640
rect 5587 12600 5632 12628
rect 5626 12588 5632 12600
rect 5684 12588 5690 12640
rect 7190 12628 7196 12640
rect 7151 12600 7196 12628
rect 7190 12588 7196 12600
rect 7248 12588 7254 12640
rect 7282 12588 7288 12640
rect 7340 12628 7346 12640
rect 10505 12631 10563 12637
rect 7340 12600 7385 12628
rect 7340 12588 7346 12600
rect 10505 12597 10517 12631
rect 10551 12628 10563 12631
rect 10778 12628 10784 12640
rect 10551 12600 10784 12628
rect 10551 12597 10563 12600
rect 10505 12591 10563 12597
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 14090 12628 14096 12640
rect 14051 12600 14096 12628
rect 14090 12588 14096 12600
rect 14148 12588 14154 12640
rect 16850 12628 16856 12640
rect 16811 12600 16856 12628
rect 16850 12588 16856 12600
rect 16908 12588 16914 12640
rect 19426 12628 19432 12640
rect 19387 12600 19432 12628
rect 19426 12588 19432 12600
rect 19484 12588 19490 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1670 12384 1676 12436
rect 1728 12424 1734 12436
rect 1946 12424 1952 12436
rect 1728 12396 1952 12424
rect 1728 12384 1734 12396
rect 1946 12384 1952 12396
rect 2004 12384 2010 12436
rect 2314 12384 2320 12436
rect 2372 12424 2378 12436
rect 2590 12424 2596 12436
rect 2372 12396 2596 12424
rect 2372 12384 2378 12396
rect 2590 12384 2596 12396
rect 2648 12384 2654 12436
rect 2682 12384 2688 12436
rect 2740 12424 2746 12436
rect 2777 12427 2835 12433
rect 2777 12424 2789 12427
rect 2740 12396 2789 12424
rect 2740 12384 2746 12396
rect 2777 12393 2789 12396
rect 2823 12424 2835 12427
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 2823 12396 3801 12424
rect 2823 12393 2835 12396
rect 2777 12387 2835 12393
rect 3789 12393 3801 12396
rect 3835 12424 3847 12427
rect 5077 12427 5135 12433
rect 5077 12424 5089 12427
rect 3835 12396 5089 12424
rect 3835 12393 3847 12396
rect 3789 12387 3847 12393
rect 5077 12393 5089 12396
rect 5123 12424 5135 12427
rect 5166 12424 5172 12436
rect 5123 12396 5172 12424
rect 5123 12393 5135 12396
rect 5077 12387 5135 12393
rect 5166 12384 5172 12396
rect 5224 12384 5230 12436
rect 6730 12424 6736 12436
rect 6691 12396 6736 12424
rect 6730 12384 6736 12396
rect 6788 12384 6794 12436
rect 7282 12424 7288 12436
rect 7243 12396 7288 12424
rect 7282 12384 7288 12396
rect 7340 12424 7346 12436
rect 7837 12427 7895 12433
rect 7837 12424 7849 12427
rect 7340 12396 7849 12424
rect 7340 12384 7346 12396
rect 7837 12393 7849 12396
rect 7883 12393 7895 12427
rect 7837 12387 7895 12393
rect 8202 12384 8208 12436
rect 8260 12384 8266 12436
rect 9122 12424 9128 12436
rect 9083 12396 9128 12424
rect 9122 12384 9128 12396
rect 9180 12384 9186 12436
rect 9674 12424 9680 12436
rect 9635 12396 9680 12424
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 10134 12424 10140 12436
rect 10047 12396 10140 12424
rect 10134 12384 10140 12396
rect 10192 12424 10198 12436
rect 11241 12427 11299 12433
rect 11241 12424 11253 12427
rect 10192 12396 11253 12424
rect 10192 12384 10198 12396
rect 11241 12393 11253 12396
rect 11287 12393 11299 12427
rect 11241 12387 11299 12393
rect 12805 12427 12863 12433
rect 12805 12393 12817 12427
rect 12851 12424 12863 12427
rect 12894 12424 12900 12436
rect 12851 12396 12900 12424
rect 12851 12393 12863 12396
rect 12805 12387 12863 12393
rect 12894 12384 12900 12396
rect 12952 12384 12958 12436
rect 13633 12427 13691 12433
rect 13633 12393 13645 12427
rect 13679 12424 13691 12427
rect 14277 12427 14335 12433
rect 14277 12424 14289 12427
rect 13679 12396 14289 12424
rect 13679 12393 13691 12396
rect 13633 12387 13691 12393
rect 14277 12393 14289 12396
rect 14323 12424 14335 12427
rect 14458 12424 14464 12436
rect 14323 12396 14464 12424
rect 14323 12393 14335 12396
rect 14277 12387 14335 12393
rect 14458 12384 14464 12396
rect 14516 12384 14522 12436
rect 14737 12427 14795 12433
rect 14737 12393 14749 12427
rect 14783 12424 14795 12427
rect 15102 12424 15108 12436
rect 14783 12396 15108 12424
rect 14783 12393 14795 12396
rect 14737 12387 14795 12393
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 15838 12424 15844 12436
rect 15799 12396 15844 12424
rect 15838 12384 15844 12396
rect 15896 12384 15902 12436
rect 17402 12384 17408 12436
rect 17460 12424 17466 12436
rect 17586 12424 17592 12436
rect 17460 12396 17592 12424
rect 17460 12384 17466 12396
rect 17586 12384 17592 12396
rect 17644 12384 17650 12436
rect 18046 12424 18052 12436
rect 18007 12396 18052 12424
rect 18046 12384 18052 12396
rect 18104 12384 18110 12436
rect 7745 12359 7803 12365
rect 7745 12325 7757 12359
rect 7791 12356 7803 12359
rect 8220 12356 8248 12384
rect 7791 12328 8248 12356
rect 7791 12325 7803 12328
rect 7745 12319 7803 12325
rect 9490 12316 9496 12368
rect 9548 12356 9554 12368
rect 12621 12359 12679 12365
rect 12621 12356 12633 12359
rect 9548 12328 12633 12356
rect 9548 12316 9554 12328
rect 12621 12325 12633 12328
rect 12667 12356 12679 12359
rect 13078 12356 13084 12368
rect 12667 12328 13084 12356
rect 12667 12325 12679 12328
rect 12621 12319 12679 12325
rect 13078 12316 13084 12328
rect 13136 12356 13142 12368
rect 13722 12356 13728 12368
rect 13136 12328 13728 12356
rect 13136 12316 13142 12328
rect 13722 12316 13728 12328
rect 13780 12316 13786 12368
rect 17313 12359 17371 12365
rect 17313 12325 17325 12359
rect 17359 12325 17371 12359
rect 17313 12319 17371 12325
rect 1664 12291 1722 12297
rect 1664 12257 1676 12291
rect 1710 12288 1722 12291
rect 1946 12288 1952 12300
rect 1710 12260 1952 12288
rect 1710 12257 1722 12260
rect 1664 12251 1722 12257
rect 1946 12248 1952 12260
rect 2004 12288 2010 12300
rect 4062 12288 4068 12300
rect 2004 12260 3464 12288
rect 4023 12260 4068 12288
rect 2004 12248 2010 12260
rect 1394 12220 1400 12232
rect 1355 12192 1400 12220
rect 1394 12180 1400 12192
rect 1452 12180 1458 12232
rect 3436 12229 3464 12260
rect 4062 12248 4068 12260
rect 4120 12248 4126 12300
rect 4430 12248 4436 12300
rect 4488 12288 4494 12300
rect 5074 12288 5080 12300
rect 4488 12260 5080 12288
rect 4488 12248 4494 12260
rect 5074 12248 5080 12260
rect 5132 12248 5138 12300
rect 5620 12291 5678 12297
rect 5620 12257 5632 12291
rect 5666 12288 5678 12291
rect 5994 12288 6000 12300
rect 5666 12260 6000 12288
rect 5666 12257 5678 12260
rect 5620 12251 5678 12257
rect 5994 12248 6000 12260
rect 6052 12248 6058 12300
rect 7466 12248 7472 12300
rect 7524 12288 7530 12300
rect 8018 12288 8024 12300
rect 7524 12260 8024 12288
rect 7524 12248 7530 12260
rect 8018 12248 8024 12260
rect 8076 12288 8082 12300
rect 8205 12291 8263 12297
rect 8205 12288 8217 12291
rect 8076 12260 8217 12288
rect 8076 12248 8082 12260
rect 8205 12257 8217 12260
rect 8251 12257 8263 12291
rect 10042 12288 10048 12300
rect 9955 12260 10048 12288
rect 8205 12251 8263 12257
rect 10042 12248 10048 12260
rect 10100 12288 10106 12300
rect 10870 12288 10876 12300
rect 10100 12260 10876 12288
rect 10100 12248 10106 12260
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 11606 12288 11612 12300
rect 11567 12260 11612 12288
rect 11606 12248 11612 12260
rect 11664 12248 11670 12300
rect 11698 12248 11704 12300
rect 11756 12288 11762 12300
rect 13173 12291 13231 12297
rect 11756 12260 11801 12288
rect 11756 12248 11762 12260
rect 13173 12257 13185 12291
rect 13219 12288 13231 12291
rect 14090 12288 14096 12300
rect 13219 12260 14096 12288
rect 13219 12257 13231 12260
rect 13173 12251 13231 12257
rect 14090 12248 14096 12260
rect 14148 12248 14154 12300
rect 15746 12288 15752 12300
rect 15707 12260 15752 12288
rect 15746 12248 15752 12260
rect 15804 12288 15810 12300
rect 16761 12291 16819 12297
rect 16761 12288 16773 12291
rect 15804 12260 16773 12288
rect 15804 12248 15810 12260
rect 16761 12257 16773 12260
rect 16807 12288 16819 12291
rect 17034 12288 17040 12300
rect 16807 12260 17040 12288
rect 16807 12257 16819 12260
rect 16761 12251 16819 12257
rect 17034 12248 17040 12260
rect 17092 12248 17098 12300
rect 17328 12232 17356 12319
rect 3421 12223 3479 12229
rect 3421 12189 3433 12223
rect 3467 12220 3479 12223
rect 3510 12220 3516 12232
rect 3467 12192 3516 12220
rect 3467 12189 3479 12192
rect 3421 12183 3479 12189
rect 3510 12180 3516 12192
rect 3568 12180 3574 12232
rect 5353 12223 5411 12229
rect 5353 12189 5365 12223
rect 5399 12189 5411 12223
rect 8294 12220 8300 12232
rect 8255 12192 8300 12220
rect 5353 12183 5411 12189
rect 3142 12044 3148 12096
rect 3200 12084 3206 12096
rect 3602 12084 3608 12096
rect 3200 12056 3608 12084
rect 3200 12044 3206 12056
rect 3602 12044 3608 12056
rect 3660 12044 3666 12096
rect 4246 12084 4252 12096
rect 4207 12056 4252 12084
rect 4246 12044 4252 12056
rect 4304 12044 4310 12096
rect 4614 12044 4620 12096
rect 4672 12084 4678 12096
rect 4709 12087 4767 12093
rect 4709 12084 4721 12087
rect 4672 12056 4721 12084
rect 4672 12044 4678 12056
rect 4709 12053 4721 12056
rect 4755 12084 4767 12087
rect 4890 12084 4896 12096
rect 4755 12056 4896 12084
rect 4755 12053 4767 12056
rect 4709 12047 4767 12053
rect 4890 12044 4896 12056
rect 4948 12044 4954 12096
rect 5368 12084 5396 12183
rect 8294 12180 8300 12192
rect 8352 12180 8358 12232
rect 8478 12220 8484 12232
rect 8439 12192 8484 12220
rect 8478 12180 8484 12192
rect 8536 12180 8542 12232
rect 10318 12220 10324 12232
rect 10231 12192 10324 12220
rect 10318 12180 10324 12192
rect 10376 12220 10382 12232
rect 10778 12220 10784 12232
rect 10376 12192 10784 12220
rect 10376 12180 10382 12192
rect 10778 12180 10784 12192
rect 10836 12180 10842 12232
rect 11882 12220 11888 12232
rect 11843 12192 11888 12220
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 13265 12223 13323 12229
rect 13265 12189 13277 12223
rect 13311 12189 13323 12223
rect 13446 12220 13452 12232
rect 13359 12192 13452 12220
rect 13265 12183 13323 12189
rect 11149 12155 11207 12161
rect 11149 12121 11161 12155
rect 11195 12152 11207 12155
rect 11900 12152 11928 12180
rect 11195 12124 11928 12152
rect 13280 12152 13308 12183
rect 13446 12180 13452 12192
rect 13504 12220 13510 12232
rect 16022 12220 16028 12232
rect 13504 12192 13860 12220
rect 15983 12192 16028 12220
rect 13504 12180 13510 12192
rect 13722 12152 13728 12164
rect 13280 12124 13728 12152
rect 11195 12121 11207 12124
rect 11149 12115 11207 12121
rect 13722 12112 13728 12124
rect 13780 12112 13786 12164
rect 13832 12096 13860 12192
rect 16022 12180 16028 12192
rect 16080 12220 16086 12232
rect 16850 12220 16856 12232
rect 16080 12192 16856 12220
rect 16080 12180 16086 12192
rect 16850 12180 16856 12192
rect 16908 12180 16914 12232
rect 17310 12180 17316 12232
rect 17368 12180 17374 12232
rect 17405 12223 17463 12229
rect 17405 12189 17417 12223
rect 17451 12189 17463 12223
rect 17586 12220 17592 12232
rect 17547 12192 17592 12220
rect 17405 12183 17463 12189
rect 17034 12112 17040 12164
rect 17092 12152 17098 12164
rect 17420 12152 17448 12183
rect 17586 12180 17592 12192
rect 17644 12180 17650 12232
rect 17092 12124 17448 12152
rect 17092 12112 17098 12124
rect 5534 12084 5540 12096
rect 5368 12056 5540 12084
rect 5534 12044 5540 12056
rect 5592 12044 5598 12096
rect 10778 12084 10784 12096
rect 10739 12056 10784 12084
rect 10778 12044 10784 12056
rect 10836 12044 10842 12096
rect 11238 12044 11244 12096
rect 11296 12084 11302 12096
rect 13633 12087 13691 12093
rect 13633 12084 13645 12087
rect 11296 12056 13645 12084
rect 11296 12044 11302 12056
rect 13633 12053 13645 12056
rect 13679 12053 13691 12087
rect 13814 12084 13820 12096
rect 13775 12056 13820 12084
rect 13633 12047 13691 12053
rect 13814 12044 13820 12056
rect 13872 12044 13878 12096
rect 14734 12044 14740 12096
rect 14792 12084 14798 12096
rect 15013 12087 15071 12093
rect 15013 12084 15025 12087
rect 14792 12056 15025 12084
rect 14792 12044 14798 12056
rect 15013 12053 15025 12056
rect 15059 12053 15071 12087
rect 15013 12047 15071 12053
rect 15286 12044 15292 12096
rect 15344 12084 15350 12096
rect 15381 12087 15439 12093
rect 15381 12084 15393 12087
rect 15344 12056 15393 12084
rect 15344 12044 15350 12056
rect 15381 12053 15393 12056
rect 15427 12053 15439 12087
rect 16390 12084 16396 12096
rect 16351 12056 16396 12084
rect 15381 12047 15439 12053
rect 16390 12044 16396 12056
rect 16448 12044 16454 12096
rect 16942 12084 16948 12096
rect 16903 12056 16948 12084
rect 16942 12044 16948 12056
rect 17000 12044 17006 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1578 11880 1584 11892
rect 1539 11852 1584 11880
rect 1578 11840 1584 11852
rect 1636 11840 1642 11892
rect 4062 11840 4068 11892
rect 4120 11880 4126 11892
rect 4801 11883 4859 11889
rect 4801 11880 4813 11883
rect 4120 11852 4813 11880
rect 4120 11840 4126 11852
rect 4801 11849 4813 11852
rect 4847 11849 4859 11883
rect 4801 11843 4859 11849
rect 6273 11883 6331 11889
rect 6273 11849 6285 11883
rect 6319 11880 6331 11883
rect 6546 11880 6552 11892
rect 6319 11852 6552 11880
rect 6319 11849 6331 11852
rect 6273 11843 6331 11849
rect 6546 11840 6552 11852
rect 6604 11840 6610 11892
rect 8294 11840 8300 11892
rect 8352 11880 8358 11892
rect 8754 11880 8760 11892
rect 8352 11852 8760 11880
rect 8352 11840 8358 11852
rect 8754 11840 8760 11852
rect 8812 11880 8818 11892
rect 9125 11883 9183 11889
rect 9125 11880 9137 11883
rect 8812 11852 9137 11880
rect 8812 11840 8818 11852
rect 9125 11849 9137 11852
rect 9171 11849 9183 11883
rect 9125 11843 9183 11849
rect 9769 11883 9827 11889
rect 9769 11849 9781 11883
rect 9815 11880 9827 11883
rect 10042 11880 10048 11892
rect 9815 11852 10048 11880
rect 9815 11849 9827 11852
rect 9769 11843 9827 11849
rect 10042 11840 10048 11852
rect 10100 11840 10106 11892
rect 10137 11883 10195 11889
rect 10137 11849 10149 11883
rect 10183 11880 10195 11883
rect 10318 11880 10324 11892
rect 10183 11852 10324 11880
rect 10183 11849 10195 11852
rect 10137 11843 10195 11849
rect 1394 11772 1400 11824
rect 1452 11812 1458 11824
rect 1854 11812 1860 11824
rect 1452 11784 1860 11812
rect 1452 11772 1458 11784
rect 1854 11772 1860 11784
rect 1912 11812 1918 11824
rect 1949 11815 2007 11821
rect 1949 11812 1961 11815
rect 1912 11784 1961 11812
rect 1912 11772 1918 11784
rect 1949 11781 1961 11784
rect 1995 11781 2007 11815
rect 1949 11775 2007 11781
rect 1394 11676 1400 11688
rect 1355 11648 1400 11676
rect 1394 11636 1400 11648
rect 1452 11636 1458 11688
rect 1964 11676 1992 11775
rect 6564 11744 6592 11840
rect 8478 11772 8484 11824
rect 8536 11812 8542 11824
rect 8849 11815 8907 11821
rect 8849 11812 8861 11815
rect 8536 11784 8861 11812
rect 8536 11772 8542 11784
rect 8849 11781 8861 11784
rect 8895 11812 8907 11815
rect 10152 11812 10180 11843
rect 10318 11840 10324 11852
rect 10376 11840 10382 11892
rect 10781 11883 10839 11889
rect 10781 11849 10793 11883
rect 10827 11880 10839 11883
rect 10962 11880 10968 11892
rect 10827 11852 10968 11880
rect 10827 11849 10839 11852
rect 10781 11843 10839 11849
rect 10962 11840 10968 11852
rect 11020 11840 11026 11892
rect 11606 11840 11612 11892
rect 11664 11880 11670 11892
rect 11793 11883 11851 11889
rect 11793 11880 11805 11883
rect 11664 11852 11805 11880
rect 11664 11840 11670 11852
rect 11793 11849 11805 11852
rect 11839 11849 11851 11883
rect 11793 11843 11851 11849
rect 12526 11840 12532 11892
rect 12584 11880 12590 11892
rect 12802 11880 12808 11892
rect 12584 11852 12808 11880
rect 12584 11840 12590 11852
rect 12802 11840 12808 11852
rect 12860 11840 12866 11892
rect 14090 11840 14096 11892
rect 14148 11880 14154 11892
rect 14461 11883 14519 11889
rect 14461 11880 14473 11883
rect 14148 11852 14473 11880
rect 14148 11840 14154 11852
rect 14461 11849 14473 11852
rect 14507 11849 14519 11883
rect 14461 11843 14519 11849
rect 14642 11840 14648 11892
rect 14700 11880 14706 11892
rect 15013 11883 15071 11889
rect 15013 11880 15025 11883
rect 14700 11852 15025 11880
rect 14700 11840 14706 11852
rect 15013 11849 15025 11852
rect 15059 11849 15071 11883
rect 15013 11843 15071 11849
rect 15838 11840 15844 11892
rect 15896 11880 15902 11892
rect 16393 11883 16451 11889
rect 16393 11880 16405 11883
rect 15896 11852 16405 11880
rect 15896 11840 15902 11852
rect 16393 11849 16405 11852
rect 16439 11849 16451 11883
rect 16393 11843 16451 11849
rect 8895 11784 10180 11812
rect 10689 11815 10747 11821
rect 8895 11781 8907 11784
rect 8849 11775 8907 11781
rect 10689 11781 10701 11815
rect 10735 11812 10747 11815
rect 11698 11812 11704 11824
rect 10735 11784 11704 11812
rect 10735 11781 10747 11784
rect 10689 11775 10747 11781
rect 11698 11772 11704 11784
rect 11756 11772 11762 11824
rect 15746 11772 15752 11824
rect 15804 11812 15810 11824
rect 16025 11815 16083 11821
rect 16025 11812 16037 11815
rect 15804 11784 16037 11812
rect 15804 11772 15810 11784
rect 16025 11781 16037 11784
rect 16071 11781 16083 11815
rect 16025 11775 16083 11781
rect 6564 11716 6960 11744
rect 6932 11688 6960 11716
rect 10778 11704 10784 11756
rect 10836 11744 10842 11756
rect 11333 11747 11391 11753
rect 11333 11744 11345 11747
rect 10836 11716 11345 11744
rect 10836 11704 10842 11716
rect 11333 11713 11345 11716
rect 11379 11744 11391 11747
rect 12437 11747 12495 11753
rect 12437 11744 12449 11747
rect 11379 11716 12449 11744
rect 11379 11713 11391 11716
rect 11333 11707 11391 11713
rect 12437 11713 12449 11716
rect 12483 11713 12495 11747
rect 12437 11707 12495 11713
rect 14734 11704 14740 11756
rect 14792 11744 14798 11756
rect 15378 11744 15384 11756
rect 14792 11716 15384 11744
rect 14792 11704 14798 11716
rect 15378 11704 15384 11716
rect 15436 11744 15442 11756
rect 15565 11747 15623 11753
rect 15565 11744 15577 11747
rect 15436 11716 15577 11744
rect 15436 11704 15442 11716
rect 15565 11713 15577 11716
rect 15611 11713 15623 11747
rect 15565 11707 15623 11713
rect 2774 11676 2780 11688
rect 1964 11648 2780 11676
rect 2774 11636 2780 11648
rect 2832 11676 2838 11688
rect 2869 11679 2927 11685
rect 2869 11676 2881 11679
rect 2832 11648 2881 11676
rect 2832 11636 2838 11648
rect 2869 11645 2881 11648
rect 2915 11645 2927 11679
rect 3136 11679 3194 11685
rect 3136 11676 3148 11679
rect 2869 11639 2927 11645
rect 2976 11648 3148 11676
rect 2976 11620 3004 11648
rect 3136 11645 3148 11648
rect 3182 11676 3194 11679
rect 3418 11676 3424 11688
rect 3182 11648 3424 11676
rect 3182 11645 3194 11648
rect 3136 11639 3194 11645
rect 3418 11636 3424 11648
rect 3476 11636 3482 11688
rect 6638 11636 6644 11688
rect 6696 11676 6702 11688
rect 6825 11679 6883 11685
rect 6825 11676 6837 11679
rect 6696 11648 6837 11676
rect 6696 11636 6702 11648
rect 6825 11645 6837 11648
rect 6871 11645 6883 11679
rect 6825 11639 6883 11645
rect 6914 11636 6920 11688
rect 6972 11676 6978 11688
rect 7081 11679 7139 11685
rect 7081 11676 7093 11679
rect 6972 11648 7093 11676
rect 6972 11636 6978 11648
rect 7081 11645 7093 11648
rect 7127 11645 7139 11679
rect 11238 11676 11244 11688
rect 11199 11648 11244 11676
rect 7081 11639 7139 11645
rect 11238 11636 11244 11648
rect 11296 11636 11302 11688
rect 11422 11636 11428 11688
rect 11480 11676 11486 11688
rect 12253 11679 12311 11685
rect 12253 11676 12265 11679
rect 11480 11648 12265 11676
rect 11480 11636 11486 11648
rect 12253 11645 12265 11648
rect 12299 11676 12311 11679
rect 12529 11679 12587 11685
rect 12529 11676 12541 11679
rect 12299 11648 12541 11676
rect 12299 11645 12311 11648
rect 12253 11639 12311 11645
rect 12529 11645 12541 11648
rect 12575 11676 12587 11679
rect 12618 11676 12624 11688
rect 12575 11648 12624 11676
rect 12575 11645 12587 11648
rect 12529 11639 12587 11645
rect 12618 11636 12624 11648
rect 12676 11636 12682 11688
rect 12796 11679 12854 11685
rect 12796 11676 12808 11679
rect 12728 11648 12808 11676
rect 12728 11620 12756 11648
rect 12796 11645 12808 11648
rect 12842 11676 12854 11679
rect 13078 11676 13084 11688
rect 12842 11648 13084 11676
rect 12842 11645 12854 11648
rect 12796 11639 12854 11645
rect 13078 11636 13084 11648
rect 13136 11636 13142 11688
rect 17037 11679 17095 11685
rect 17037 11645 17049 11679
rect 17083 11676 17095 11679
rect 17310 11676 17316 11688
rect 17083 11648 17316 11676
rect 17083 11645 17095 11648
rect 17037 11639 17095 11645
rect 17310 11636 17316 11648
rect 17368 11636 17374 11688
rect 2409 11611 2467 11617
rect 2409 11577 2421 11611
rect 2455 11608 2467 11611
rect 2958 11608 2964 11620
rect 2455 11580 2964 11608
rect 2455 11577 2467 11580
rect 2409 11571 2467 11577
rect 2958 11568 2964 11580
rect 3016 11568 3022 11620
rect 3068 11580 5488 11608
rect 2774 11500 2780 11552
rect 2832 11540 2838 11552
rect 3068 11540 3096 11580
rect 2832 11512 3096 11540
rect 2832 11500 2838 11512
rect 3418 11500 3424 11552
rect 3476 11540 3482 11552
rect 5460 11549 5488 11580
rect 5534 11568 5540 11620
rect 5592 11608 5598 11620
rect 5813 11611 5871 11617
rect 5813 11608 5825 11611
rect 5592 11580 5825 11608
rect 5592 11568 5598 11580
rect 5813 11577 5825 11580
rect 5859 11608 5871 11611
rect 5994 11608 6000 11620
rect 5859 11580 6000 11608
rect 5859 11577 5871 11580
rect 5813 11571 5871 11577
rect 5994 11568 6000 11580
rect 6052 11608 6058 11620
rect 8478 11608 8484 11620
rect 6052 11580 8484 11608
rect 6052 11568 6058 11580
rect 8478 11568 8484 11580
rect 8536 11568 8542 11620
rect 11146 11608 11152 11620
rect 11107 11580 11152 11608
rect 11146 11568 11152 11580
rect 11204 11568 11210 11620
rect 12710 11568 12716 11620
rect 12768 11568 12774 11620
rect 15381 11611 15439 11617
rect 15381 11608 15393 11611
rect 14844 11580 15393 11608
rect 14844 11552 14872 11580
rect 15381 11577 15393 11580
rect 15427 11577 15439 11611
rect 15381 11571 15439 11577
rect 4249 11543 4307 11549
rect 4249 11540 4261 11543
rect 3476 11512 4261 11540
rect 3476 11500 3482 11512
rect 4249 11509 4261 11512
rect 4295 11509 4307 11543
rect 4249 11503 4307 11509
rect 5445 11543 5503 11549
rect 5445 11509 5457 11543
rect 5491 11540 5503 11543
rect 5626 11540 5632 11552
rect 5491 11512 5632 11540
rect 5491 11509 5503 11512
rect 5445 11503 5503 11509
rect 5626 11500 5632 11512
rect 5684 11540 5690 11552
rect 6638 11540 6644 11552
rect 5684 11512 6644 11540
rect 5684 11500 5690 11512
rect 6638 11500 6644 11512
rect 6696 11500 6702 11552
rect 8202 11540 8208 11552
rect 8163 11512 8208 11540
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 12437 11543 12495 11549
rect 12437 11509 12449 11543
rect 12483 11540 12495 11543
rect 13446 11540 13452 11552
rect 12483 11512 13452 11540
rect 12483 11509 12495 11512
rect 12437 11503 12495 11509
rect 13446 11500 13452 11512
rect 13504 11540 13510 11552
rect 13814 11540 13820 11552
rect 13504 11512 13820 11540
rect 13504 11500 13510 11512
rect 13814 11500 13820 11512
rect 13872 11540 13878 11552
rect 13909 11543 13967 11549
rect 13909 11540 13921 11543
rect 13872 11512 13921 11540
rect 13872 11500 13878 11512
rect 13909 11509 13921 11512
rect 13955 11509 13967 11543
rect 14826 11540 14832 11552
rect 14787 11512 14832 11540
rect 13909 11503 13967 11509
rect 14826 11500 14832 11512
rect 14884 11500 14890 11552
rect 15470 11540 15476 11552
rect 15431 11512 15476 11540
rect 15470 11500 15476 11512
rect 15528 11500 15534 11552
rect 17034 11500 17040 11552
rect 17092 11540 17098 11552
rect 17313 11543 17371 11549
rect 17313 11540 17325 11543
rect 17092 11512 17325 11540
rect 17092 11500 17098 11512
rect 17313 11509 17325 11512
rect 17359 11509 17371 11543
rect 17313 11503 17371 11509
rect 17586 11500 17592 11552
rect 17644 11540 17650 11552
rect 17773 11543 17831 11549
rect 17773 11540 17785 11543
rect 17644 11512 17785 11540
rect 17644 11500 17650 11512
rect 17773 11509 17785 11512
rect 17819 11540 17831 11543
rect 18598 11540 18604 11552
rect 17819 11512 18604 11540
rect 17819 11509 17831 11512
rect 17773 11503 17831 11509
rect 18598 11500 18604 11512
rect 18656 11500 18662 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1394 11296 1400 11348
rect 1452 11336 1458 11348
rect 1581 11339 1639 11345
rect 1581 11336 1593 11339
rect 1452 11308 1593 11336
rect 1452 11296 1458 11308
rect 1581 11305 1593 11308
rect 1627 11305 1639 11339
rect 1946 11336 1952 11348
rect 1907 11308 1952 11336
rect 1581 11299 1639 11305
rect 1596 11268 1624 11299
rect 1946 11296 1952 11308
rect 2004 11296 2010 11348
rect 2038 11296 2044 11348
rect 2096 11336 2102 11348
rect 2409 11339 2467 11345
rect 2409 11336 2421 11339
rect 2096 11308 2421 11336
rect 2096 11296 2102 11308
rect 2409 11305 2421 11308
rect 2455 11305 2467 11339
rect 3789 11339 3847 11345
rect 3789 11336 3801 11339
rect 2409 11299 2467 11305
rect 2516 11308 3801 11336
rect 2516 11268 2544 11308
rect 3789 11305 3801 11308
rect 3835 11305 3847 11339
rect 3789 11299 3847 11305
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 4341 11339 4399 11345
rect 4341 11336 4353 11339
rect 4120 11308 4353 11336
rect 4120 11296 4126 11308
rect 4341 11305 4353 11308
rect 4387 11305 4399 11339
rect 4341 11299 4399 11305
rect 5261 11339 5319 11345
rect 5261 11305 5273 11339
rect 5307 11336 5319 11339
rect 5442 11336 5448 11348
rect 5307 11308 5448 11336
rect 5307 11305 5319 11308
rect 5261 11299 5319 11305
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 5626 11296 5632 11348
rect 5684 11296 5690 11348
rect 6825 11339 6883 11345
rect 6825 11305 6837 11339
rect 6871 11336 6883 11339
rect 6914 11336 6920 11348
rect 6871 11308 6920 11336
rect 6871 11305 6883 11308
rect 6825 11299 6883 11305
rect 6914 11296 6920 11308
rect 6972 11296 6978 11348
rect 7466 11336 7472 11348
rect 7427 11308 7472 11336
rect 7466 11296 7472 11308
rect 7524 11296 7530 11348
rect 7837 11339 7895 11345
rect 7837 11305 7849 11339
rect 7883 11336 7895 11339
rect 8202 11336 8208 11348
rect 7883 11308 8208 11336
rect 7883 11305 7895 11308
rect 7837 11299 7895 11305
rect 8202 11296 8208 11308
rect 8260 11296 8266 11348
rect 8294 11296 8300 11348
rect 8352 11336 8358 11348
rect 8938 11336 8944 11348
rect 8352 11308 8800 11336
rect 8899 11308 8944 11336
rect 8352 11296 8358 11308
rect 1596 11240 2544 11268
rect 2869 11271 2927 11277
rect 2869 11237 2881 11271
rect 2915 11268 2927 11271
rect 3142 11268 3148 11280
rect 2915 11240 3148 11268
rect 2915 11237 2927 11240
rect 2869 11231 2927 11237
rect 3142 11228 3148 11240
rect 3200 11228 3206 11280
rect 3418 11268 3424 11280
rect 3379 11240 3424 11268
rect 3418 11228 3424 11240
rect 3476 11228 3482 11280
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 2130 11200 2136 11212
rect 1443 11172 2136 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 2130 11160 2136 11172
rect 2188 11160 2194 11212
rect 2774 11160 2780 11212
rect 2832 11200 2838 11212
rect 4157 11203 4215 11209
rect 2832 11172 2877 11200
rect 2832 11160 2838 11172
rect 4157 11169 4169 11203
rect 4203 11200 4215 11203
rect 4338 11200 4344 11212
rect 4203 11172 4344 11200
rect 4203 11169 4215 11172
rect 4157 11163 4215 11169
rect 4338 11160 4344 11172
rect 4396 11200 4402 11212
rect 4798 11200 4804 11212
rect 4396 11172 4804 11200
rect 4396 11160 4402 11172
rect 4798 11160 4804 11172
rect 4856 11160 4862 11212
rect 5445 11203 5503 11209
rect 5445 11169 5457 11203
rect 5491 11200 5503 11203
rect 5644 11200 5672 11296
rect 5712 11271 5770 11277
rect 5712 11237 5724 11271
rect 5758 11268 5770 11271
rect 5994 11268 6000 11280
rect 5758 11240 6000 11268
rect 5758 11237 5770 11240
rect 5712 11231 5770 11237
rect 5994 11228 6000 11240
rect 6052 11268 6058 11280
rect 6730 11268 6736 11280
rect 6052 11240 6736 11268
rect 6052 11228 6058 11240
rect 6730 11228 6736 11240
rect 6788 11228 6794 11280
rect 8220 11268 8248 11296
rect 8772 11268 8800 11308
rect 8938 11296 8944 11308
rect 8996 11296 9002 11348
rect 9493 11339 9551 11345
rect 9493 11305 9505 11339
rect 9539 11336 9551 11339
rect 10134 11336 10140 11348
rect 9539 11308 10140 11336
rect 9539 11305 9551 11308
rect 9493 11299 9551 11305
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 12897 11339 12955 11345
rect 12897 11336 12909 11339
rect 12492 11308 12909 11336
rect 12492 11296 12498 11308
rect 12897 11305 12909 11308
rect 12943 11305 12955 11339
rect 13262 11336 13268 11348
rect 13223 11308 13268 11336
rect 12897 11299 12955 11305
rect 13262 11296 13268 11308
rect 13320 11296 13326 11348
rect 13722 11296 13728 11348
rect 13780 11336 13786 11348
rect 14274 11336 14280 11348
rect 13780 11308 14044 11336
rect 14235 11308 14280 11336
rect 13780 11296 13786 11308
rect 9582 11268 9588 11280
rect 8220 11240 8432 11268
rect 8772 11240 9588 11268
rect 5491 11172 5672 11200
rect 5491 11169 5503 11172
rect 5445 11163 5503 11169
rect 7742 11160 7748 11212
rect 7800 11200 7806 11212
rect 8294 11200 8300 11212
rect 7800 11172 8300 11200
rect 7800 11160 7806 11172
rect 8294 11160 8300 11172
rect 8352 11160 8358 11212
rect 8404 11200 8432 11240
rect 9582 11228 9588 11240
rect 9640 11228 9646 11280
rect 10042 11228 10048 11280
rect 10100 11268 10106 11280
rect 11330 11268 11336 11280
rect 10100 11240 11336 11268
rect 10100 11228 10106 11240
rect 11330 11228 11336 11240
rect 11388 11268 11394 11280
rect 13906 11268 13912 11280
rect 11388 11240 13768 11268
rect 13867 11240 13912 11268
rect 11388 11228 11394 11240
rect 10680 11203 10738 11209
rect 8404 11172 8524 11200
rect 2958 11092 2964 11144
rect 3016 11132 3022 11144
rect 4614 11132 4620 11144
rect 3016 11104 3061 11132
rect 4575 11104 4620 11132
rect 3016 11092 3022 11104
rect 4614 11092 4620 11104
rect 4672 11092 4678 11144
rect 8386 11132 8392 11144
rect 8347 11104 8392 11132
rect 8386 11092 8392 11104
rect 8444 11092 8450 11144
rect 8496 11141 8524 11172
rect 10680 11169 10692 11203
rect 10726 11200 10738 11203
rect 10962 11200 10968 11212
rect 10726 11172 10968 11200
rect 10726 11169 10738 11172
rect 10680 11163 10738 11169
rect 10962 11160 10968 11172
rect 11020 11160 11026 11212
rect 13740 11200 13768 11240
rect 13906 11228 13912 11240
rect 13964 11228 13970 11280
rect 14016 11268 14044 11308
rect 14274 11296 14280 11308
rect 14332 11296 14338 11348
rect 14737 11339 14795 11345
rect 14737 11305 14749 11339
rect 14783 11336 14795 11339
rect 14918 11336 14924 11348
rect 14783 11308 14924 11336
rect 14783 11305 14795 11308
rect 14737 11299 14795 11305
rect 14752 11268 14780 11299
rect 14918 11296 14924 11308
rect 14976 11296 14982 11348
rect 16025 11339 16083 11345
rect 16025 11305 16037 11339
rect 16071 11336 16083 11339
rect 16390 11336 16396 11348
rect 16071 11308 16396 11336
rect 16071 11305 16083 11308
rect 16025 11299 16083 11305
rect 16390 11296 16396 11308
rect 16448 11336 16454 11348
rect 17221 11339 17279 11345
rect 17221 11336 17233 11339
rect 16448 11308 17233 11336
rect 16448 11296 16454 11308
rect 17221 11305 17233 11308
rect 17267 11305 17279 11339
rect 17221 11299 17279 11305
rect 17126 11268 17132 11280
rect 14016 11240 14780 11268
rect 17087 11240 17132 11268
rect 17126 11228 17132 11240
rect 17184 11268 17190 11280
rect 17681 11271 17739 11277
rect 17681 11268 17693 11271
rect 17184 11240 17693 11268
rect 17184 11228 17190 11240
rect 17681 11237 17693 11240
rect 17727 11237 17739 11271
rect 17681 11231 17739 11237
rect 15013 11203 15071 11209
rect 15013 11200 15025 11203
rect 13740 11172 15025 11200
rect 15013 11169 15025 11172
rect 15059 11200 15071 11203
rect 15470 11200 15476 11212
rect 15059 11172 15476 11200
rect 15059 11169 15071 11172
rect 15013 11163 15071 11169
rect 15470 11160 15476 11172
rect 15528 11160 15534 11212
rect 15565 11203 15623 11209
rect 15565 11169 15577 11203
rect 15611 11200 15623 11203
rect 15746 11200 15752 11212
rect 15611 11172 15752 11200
rect 15611 11169 15623 11172
rect 15565 11163 15623 11169
rect 15746 11160 15752 11172
rect 15804 11200 15810 11212
rect 16022 11200 16028 11212
rect 15804 11172 16028 11200
rect 15804 11160 15810 11172
rect 16022 11160 16028 11172
rect 16080 11200 16086 11212
rect 16080 11172 16804 11200
rect 16080 11160 16086 11172
rect 8481 11135 8539 11141
rect 8481 11101 8493 11135
rect 8527 11101 8539 11135
rect 8481 11095 8539 11101
rect 10413 11135 10471 11141
rect 10413 11101 10425 11135
rect 10459 11101 10471 11135
rect 10413 11095 10471 11101
rect 13357 11135 13415 11141
rect 13357 11101 13369 11135
rect 13403 11101 13415 11135
rect 13357 11095 13415 11101
rect 2317 11067 2375 11073
rect 2317 11033 2329 11067
rect 2363 11064 2375 11067
rect 2976 11064 3004 11092
rect 2363 11036 3004 11064
rect 2363 11033 2375 11036
rect 2317 11027 2375 11033
rect 4062 11024 4068 11076
rect 4120 11064 4126 11076
rect 4890 11064 4896 11076
rect 4120 11036 4896 11064
rect 4120 11024 4126 11036
rect 4890 11024 4896 11036
rect 4948 11024 4954 11076
rect 6914 11024 6920 11076
rect 6972 11064 6978 11076
rect 7929 11067 7987 11073
rect 7929 11064 7941 11067
rect 6972 11036 7941 11064
rect 6972 11024 6978 11036
rect 7929 11033 7941 11036
rect 7975 11064 7987 11067
rect 7975 11036 8340 11064
rect 7975 11033 7987 11036
rect 7929 11027 7987 11033
rect 8312 10996 8340 11036
rect 10226 11024 10232 11076
rect 10284 11064 10290 11076
rect 10428 11064 10456 11095
rect 10284 11036 10456 11064
rect 10284 11024 10290 11036
rect 8570 10996 8576 11008
rect 8312 10968 8576 10996
rect 8570 10956 8576 10968
rect 8628 10956 8634 11008
rect 9950 10996 9956 11008
rect 9911 10968 9956 10996
rect 9950 10956 9956 10968
rect 10008 10956 10014 11008
rect 10318 10996 10324 11008
rect 10279 10968 10324 10996
rect 10318 10956 10324 10968
rect 10376 10956 10382 11008
rect 10428 10996 10456 11036
rect 11793 11067 11851 11073
rect 11793 11033 11805 11067
rect 11839 11064 11851 11067
rect 12710 11064 12716 11076
rect 11839 11036 12716 11064
rect 11839 11033 11851 11036
rect 11793 11027 11851 11033
rect 12710 11024 12716 11036
rect 12768 11024 12774 11076
rect 13372 11064 13400 11095
rect 13446 11092 13452 11144
rect 13504 11132 13510 11144
rect 13504 11104 13549 11132
rect 13504 11092 13510 11104
rect 15286 11092 15292 11144
rect 15344 11132 15350 11144
rect 16117 11135 16175 11141
rect 16117 11132 16129 11135
rect 15344 11104 16129 11132
rect 15344 11092 15350 11104
rect 16117 11101 16129 11104
rect 16163 11101 16175 11135
rect 16298 11132 16304 11144
rect 16259 11104 16304 11132
rect 16117 11095 16175 11101
rect 16298 11092 16304 11104
rect 16356 11092 16362 11144
rect 16776 11141 16804 11172
rect 17402 11160 17408 11212
rect 17460 11200 17466 11212
rect 17589 11203 17647 11209
rect 17589 11200 17601 11203
rect 17460 11172 17601 11200
rect 17460 11160 17466 11172
rect 17589 11169 17601 11172
rect 17635 11169 17647 11203
rect 17589 11163 17647 11169
rect 16761 11135 16819 11141
rect 16761 11101 16773 11135
rect 16807 11132 16819 11135
rect 17862 11132 17868 11144
rect 16807 11104 17868 11132
rect 16807 11101 16819 11104
rect 16761 11095 16819 11101
rect 17862 11092 17868 11104
rect 17920 11092 17926 11144
rect 15654 11064 15660 11076
rect 13372 11036 13768 11064
rect 15615 11036 15660 11064
rect 11422 10996 11428 11008
rect 10428 10968 11428 10996
rect 11422 10956 11428 10968
rect 11480 10956 11486 11008
rect 12529 10999 12587 11005
rect 12529 10965 12541 10999
rect 12575 10996 12587 10999
rect 13078 10996 13084 11008
rect 12575 10968 13084 10996
rect 12575 10965 12587 10968
rect 12529 10959 12587 10965
rect 13078 10956 13084 10968
rect 13136 10956 13142 11008
rect 13740 10996 13768 11036
rect 15654 11024 15660 11036
rect 15712 11024 15718 11076
rect 14642 10996 14648 11008
rect 13740 10968 14648 10996
rect 14642 10956 14648 10968
rect 14700 10956 14706 11008
rect 18325 10999 18383 11005
rect 18325 10965 18337 10999
rect 18371 10996 18383 10999
rect 18598 10996 18604 11008
rect 18371 10968 18604 10996
rect 18371 10965 18383 10968
rect 18325 10959 18383 10965
rect 18598 10956 18604 10968
rect 18656 10956 18662 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1397 10795 1455 10801
rect 1397 10761 1409 10795
rect 1443 10792 1455 10795
rect 2682 10792 2688 10804
rect 1443 10764 2688 10792
rect 1443 10761 1455 10764
rect 1397 10755 1455 10761
rect 2682 10752 2688 10764
rect 2740 10752 2746 10804
rect 3050 10752 3056 10804
rect 3108 10792 3114 10804
rect 3237 10795 3295 10801
rect 3237 10792 3249 10795
rect 3108 10764 3249 10792
rect 3108 10752 3114 10764
rect 3237 10761 3249 10764
rect 3283 10761 3295 10795
rect 4338 10792 4344 10804
rect 4299 10764 4344 10792
rect 3237 10755 3295 10761
rect 4338 10752 4344 10764
rect 4396 10752 4402 10804
rect 5169 10795 5227 10801
rect 5169 10761 5181 10795
rect 5215 10792 5227 10795
rect 5350 10792 5356 10804
rect 5215 10764 5356 10792
rect 5215 10761 5227 10764
rect 5169 10755 5227 10761
rect 5350 10752 5356 10764
rect 5408 10752 5414 10804
rect 6641 10795 6699 10801
rect 6641 10761 6653 10795
rect 6687 10792 6699 10795
rect 7190 10792 7196 10804
rect 6687 10764 7196 10792
rect 6687 10761 6699 10764
rect 6641 10755 6699 10761
rect 7190 10752 7196 10764
rect 7248 10752 7254 10804
rect 7285 10795 7343 10801
rect 7285 10761 7297 10795
rect 7331 10792 7343 10795
rect 8386 10792 8392 10804
rect 7331 10764 8392 10792
rect 7331 10761 7343 10764
rect 7285 10755 7343 10761
rect 8386 10752 8392 10764
rect 8444 10752 8450 10804
rect 9674 10792 9680 10804
rect 9635 10764 9680 10792
rect 9674 10752 9680 10764
rect 9732 10752 9738 10804
rect 11333 10795 11391 10801
rect 11333 10761 11345 10795
rect 11379 10792 11391 10795
rect 11422 10792 11428 10804
rect 11379 10764 11428 10792
rect 11379 10761 11391 10764
rect 11333 10755 11391 10761
rect 11422 10752 11428 10764
rect 11480 10752 11486 10804
rect 13446 10792 13452 10804
rect 13407 10764 13452 10792
rect 13446 10752 13452 10764
rect 13504 10752 13510 10804
rect 14642 10792 14648 10804
rect 14603 10764 14648 10792
rect 14642 10752 14648 10764
rect 14700 10752 14706 10804
rect 14734 10752 14740 10804
rect 14792 10792 14798 10804
rect 14921 10795 14979 10801
rect 14921 10792 14933 10795
rect 14792 10764 14933 10792
rect 14792 10752 14798 10764
rect 14921 10761 14933 10764
rect 14967 10761 14979 10795
rect 14921 10755 14979 10761
rect 15381 10795 15439 10801
rect 15381 10761 15393 10795
rect 15427 10792 15439 10795
rect 15838 10792 15844 10804
rect 15427 10764 15844 10792
rect 15427 10761 15439 10764
rect 15381 10755 15439 10761
rect 7742 10724 7748 10736
rect 4632 10696 7748 10724
rect 2038 10656 2044 10668
rect 1999 10628 2044 10656
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 2314 10616 2320 10668
rect 2372 10656 2378 10668
rect 3053 10659 3111 10665
rect 3053 10656 3065 10659
rect 2372 10628 3065 10656
rect 2372 10616 2378 10628
rect 3053 10625 3065 10628
rect 3099 10625 3111 10659
rect 3053 10619 3111 10625
rect 1394 10548 1400 10600
rect 1452 10588 1458 10600
rect 1765 10591 1823 10597
rect 1765 10588 1777 10591
rect 1452 10560 1777 10588
rect 1452 10548 1458 10560
rect 1765 10557 1777 10560
rect 1811 10557 1823 10591
rect 3068 10588 3096 10619
rect 3418 10616 3424 10668
rect 3476 10656 3482 10668
rect 3789 10659 3847 10665
rect 3789 10656 3801 10659
rect 3476 10628 3801 10656
rect 3476 10616 3482 10628
rect 3789 10625 3801 10628
rect 3835 10656 3847 10659
rect 3878 10656 3884 10668
rect 3835 10628 3884 10656
rect 3835 10625 3847 10628
rect 3789 10619 3847 10625
rect 3878 10616 3884 10628
rect 3936 10616 3942 10668
rect 3697 10591 3755 10597
rect 3697 10588 3709 10591
rect 3068 10560 3709 10588
rect 1765 10551 1823 10557
rect 3697 10557 3709 10560
rect 3743 10588 3755 10591
rect 4632 10588 4660 10696
rect 7742 10684 7748 10696
rect 7800 10684 7806 10736
rect 8754 10684 8760 10736
rect 8812 10724 8818 10736
rect 10229 10727 10287 10733
rect 10229 10724 10241 10727
rect 8812 10696 10241 10724
rect 8812 10684 8818 10696
rect 10229 10693 10241 10696
rect 10275 10724 10287 10727
rect 11054 10724 11060 10736
rect 10275 10696 11060 10724
rect 10275 10693 10287 10696
rect 10229 10687 10287 10693
rect 11054 10684 11060 10696
rect 11112 10684 11118 10736
rect 4709 10659 4767 10665
rect 4709 10625 4721 10659
rect 4755 10656 4767 10659
rect 5077 10659 5135 10665
rect 5077 10656 5089 10659
rect 4755 10628 5089 10656
rect 4755 10625 4767 10628
rect 4709 10619 4767 10625
rect 5077 10625 5089 10628
rect 5123 10656 5135 10659
rect 5813 10659 5871 10665
rect 5813 10656 5825 10659
rect 5123 10628 5825 10656
rect 5123 10625 5135 10628
rect 5077 10619 5135 10625
rect 5813 10625 5825 10628
rect 5859 10656 5871 10659
rect 5994 10656 6000 10668
rect 5859 10628 6000 10656
rect 5859 10625 5871 10628
rect 5813 10619 5871 10625
rect 5994 10616 6000 10628
rect 6052 10616 6058 10668
rect 9950 10616 9956 10668
rect 10008 10656 10014 10668
rect 10781 10659 10839 10665
rect 10781 10656 10793 10659
rect 10008 10628 10793 10656
rect 10008 10616 10014 10628
rect 10781 10625 10793 10628
rect 10827 10625 10839 10659
rect 13078 10656 13084 10668
rect 13039 10628 13084 10656
rect 10781 10619 10839 10625
rect 13078 10616 13084 10628
rect 13136 10616 13142 10668
rect 15488 10665 15516 10764
rect 15838 10752 15844 10764
rect 15896 10792 15902 10804
rect 16482 10792 16488 10804
rect 15896 10764 16488 10792
rect 15896 10752 15902 10764
rect 16482 10752 16488 10764
rect 16540 10752 16546 10804
rect 18046 10792 18052 10804
rect 18007 10764 18052 10792
rect 18046 10752 18052 10764
rect 18104 10752 18110 10804
rect 15473 10659 15531 10665
rect 15473 10625 15485 10659
rect 15519 10625 15531 10659
rect 18598 10656 18604 10668
rect 18559 10628 18604 10656
rect 15473 10619 15531 10625
rect 18598 10616 18604 10628
rect 18656 10616 18662 10668
rect 3743 10560 4660 10588
rect 3743 10557 3755 10560
rect 3697 10551 3755 10557
rect 5534 10548 5540 10600
rect 5592 10588 5598 10600
rect 5629 10591 5687 10597
rect 5629 10588 5641 10591
rect 5592 10560 5641 10588
rect 5592 10548 5598 10560
rect 5629 10557 5641 10560
rect 5675 10557 5687 10591
rect 5629 10551 5687 10557
rect 6273 10591 6331 10597
rect 6273 10557 6285 10591
rect 6319 10588 6331 10591
rect 6638 10588 6644 10600
rect 6319 10560 6644 10588
rect 6319 10557 6331 10560
rect 6273 10551 6331 10557
rect 6638 10548 6644 10560
rect 6696 10588 6702 10600
rect 7098 10588 7104 10600
rect 6696 10560 7104 10588
rect 6696 10548 6702 10560
rect 7098 10548 7104 10560
rect 7156 10588 7162 10600
rect 7653 10591 7711 10597
rect 7653 10588 7665 10591
rect 7156 10560 7665 10588
rect 7156 10548 7162 10560
rect 7653 10557 7665 10560
rect 7699 10588 7711 10591
rect 7745 10591 7803 10597
rect 7745 10588 7757 10591
rect 7699 10560 7757 10588
rect 7699 10557 7711 10560
rect 7653 10551 7711 10557
rect 7745 10557 7757 10560
rect 7791 10588 7803 10591
rect 9674 10588 9680 10600
rect 7791 10560 9680 10588
rect 7791 10557 7803 10560
rect 7745 10551 7803 10557
rect 9674 10548 9680 10560
rect 9732 10588 9738 10600
rect 10226 10588 10232 10600
rect 9732 10560 10232 10588
rect 9732 10548 9738 10560
rect 10226 10548 10232 10560
rect 10284 10548 10290 10600
rect 10318 10548 10324 10600
rect 10376 10588 10382 10600
rect 10689 10591 10747 10597
rect 10689 10588 10701 10591
rect 10376 10560 10701 10588
rect 10376 10548 10382 10560
rect 10689 10557 10701 10560
rect 10735 10557 10747 10591
rect 10689 10551 10747 10557
rect 12618 10548 12624 10600
rect 12676 10588 12682 10600
rect 12805 10591 12863 10597
rect 12805 10588 12817 10591
rect 12676 10560 12817 10588
rect 12676 10548 12682 10560
rect 12805 10557 12817 10560
rect 12851 10557 12863 10591
rect 12805 10551 12863 10557
rect 12897 10591 12955 10597
rect 12897 10557 12909 10591
rect 12943 10588 12955 10591
rect 13170 10588 13176 10600
rect 12943 10560 13176 10588
rect 12943 10557 12955 10560
rect 12897 10551 12955 10557
rect 1854 10520 1860 10532
rect 1815 10492 1860 10520
rect 1854 10480 1860 10492
rect 1912 10480 1918 10532
rect 2777 10523 2835 10529
rect 2777 10489 2789 10523
rect 2823 10520 2835 10523
rect 3605 10523 3663 10529
rect 3605 10520 3617 10523
rect 2823 10492 3617 10520
rect 2823 10489 2835 10492
rect 2777 10483 2835 10489
rect 3605 10489 3617 10492
rect 3651 10520 3663 10523
rect 4062 10520 4068 10532
rect 3651 10492 4068 10520
rect 3651 10489 3663 10492
rect 3605 10483 3663 10489
rect 4062 10480 4068 10492
rect 4120 10480 4126 10532
rect 8012 10523 8070 10529
rect 8012 10489 8024 10523
rect 8058 10520 8070 10523
rect 8202 10520 8208 10532
rect 8058 10492 8208 10520
rect 8058 10489 8070 10492
rect 8012 10483 8070 10489
rect 8202 10480 8208 10492
rect 8260 10480 8266 10532
rect 9306 10480 9312 10532
rect 9364 10520 9370 10532
rect 9490 10520 9496 10532
rect 9364 10492 9496 10520
rect 9364 10480 9370 10492
rect 9490 10480 9496 10492
rect 9548 10520 9554 10532
rect 10045 10523 10103 10529
rect 10045 10520 10057 10523
rect 9548 10492 10057 10520
rect 9548 10480 9554 10492
rect 10045 10489 10057 10492
rect 10091 10520 10103 10523
rect 10597 10523 10655 10529
rect 10597 10520 10609 10523
rect 10091 10492 10609 10520
rect 10091 10489 10103 10492
rect 10045 10483 10103 10489
rect 10597 10489 10609 10492
rect 10643 10489 10655 10523
rect 10597 10483 10655 10489
rect 12253 10523 12311 10529
rect 12253 10489 12265 10523
rect 12299 10520 12311 10523
rect 12912 10520 12940 10551
rect 13170 10548 13176 10560
rect 13228 10548 13234 10600
rect 13814 10588 13820 10600
rect 13775 10560 13820 10588
rect 13814 10548 13820 10560
rect 13872 10548 13878 10600
rect 15746 10529 15752 10532
rect 15740 10520 15752 10529
rect 12299 10492 12940 10520
rect 15707 10492 15752 10520
rect 12299 10489 12311 10492
rect 12253 10483 12311 10489
rect 15740 10483 15752 10492
rect 15746 10480 15752 10483
rect 15804 10480 15810 10532
rect 17865 10523 17923 10529
rect 17865 10489 17877 10523
rect 17911 10520 17923 10523
rect 18230 10520 18236 10532
rect 17911 10492 18236 10520
rect 17911 10489 17923 10492
rect 17865 10483 17923 10489
rect 18230 10480 18236 10492
rect 18288 10520 18294 10532
rect 18509 10523 18567 10529
rect 18509 10520 18521 10523
rect 18288 10492 18521 10520
rect 18288 10480 18294 10492
rect 18509 10489 18521 10492
rect 18555 10489 18567 10523
rect 18509 10483 18567 10489
rect 5537 10455 5595 10461
rect 5537 10421 5549 10455
rect 5583 10452 5595 10455
rect 5626 10452 5632 10464
rect 5583 10424 5632 10452
rect 5583 10421 5595 10424
rect 5537 10415 5595 10421
rect 5626 10412 5632 10424
rect 5684 10412 5690 10464
rect 9122 10452 9128 10464
rect 9035 10424 9128 10452
rect 9122 10412 9128 10424
rect 9180 10452 9186 10464
rect 9950 10452 9956 10464
rect 9180 10424 9956 10452
rect 9180 10412 9186 10424
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 11606 10452 11612 10464
rect 11567 10424 11612 10452
rect 11606 10412 11612 10424
rect 11664 10412 11670 10464
rect 12437 10455 12495 10461
rect 12437 10421 12449 10455
rect 12483 10452 12495 10455
rect 12710 10452 12716 10464
rect 12483 10424 12716 10452
rect 12483 10421 12495 10424
rect 12437 10415 12495 10421
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 13906 10412 13912 10464
rect 13964 10452 13970 10464
rect 14185 10455 14243 10461
rect 14185 10452 14197 10455
rect 13964 10424 14197 10452
rect 13964 10412 13970 10424
rect 14185 10421 14197 10424
rect 14231 10421 14243 10455
rect 14185 10415 14243 10421
rect 16758 10412 16764 10464
rect 16816 10452 16822 10464
rect 16853 10455 16911 10461
rect 16853 10452 16865 10455
rect 16816 10424 16865 10452
rect 16816 10412 16822 10424
rect 16853 10421 16865 10424
rect 16899 10421 16911 10455
rect 17402 10452 17408 10464
rect 17363 10424 17408 10452
rect 16853 10415 16911 10421
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 18046 10412 18052 10464
rect 18104 10452 18110 10464
rect 18417 10455 18475 10461
rect 18417 10452 18429 10455
rect 18104 10424 18429 10452
rect 18104 10412 18110 10424
rect 18417 10421 18429 10424
rect 18463 10421 18475 10455
rect 18417 10415 18475 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 2038 10208 2044 10260
rect 2096 10248 2102 10260
rect 2590 10248 2596 10260
rect 2096 10220 2596 10248
rect 2096 10208 2102 10220
rect 2590 10208 2596 10220
rect 2648 10248 2654 10260
rect 3421 10251 3479 10257
rect 3421 10248 3433 10251
rect 2648 10220 3433 10248
rect 2648 10208 2654 10220
rect 3421 10217 3433 10220
rect 3467 10217 3479 10251
rect 3786 10248 3792 10260
rect 3747 10220 3792 10248
rect 3421 10211 3479 10217
rect 3786 10208 3792 10220
rect 3844 10208 3850 10260
rect 4893 10251 4951 10257
rect 4893 10217 4905 10251
rect 4939 10248 4951 10251
rect 5626 10248 5632 10260
rect 4939 10220 5632 10248
rect 4939 10217 4951 10220
rect 4893 10211 4951 10217
rect 5626 10208 5632 10220
rect 5684 10248 5690 10260
rect 6273 10251 6331 10257
rect 6273 10248 6285 10251
rect 5684 10220 6285 10248
rect 5684 10208 5690 10220
rect 6273 10217 6285 10220
rect 6319 10217 6331 10251
rect 6273 10211 6331 10217
rect 6457 10251 6515 10257
rect 6457 10217 6469 10251
rect 6503 10248 6515 10251
rect 8481 10251 8539 10257
rect 8481 10248 8493 10251
rect 6503 10220 8493 10248
rect 6503 10217 6515 10220
rect 6457 10211 6515 10217
rect 8481 10217 8493 10220
rect 8527 10248 8539 10251
rect 9401 10251 9459 10257
rect 9401 10248 9413 10251
rect 8527 10220 9413 10248
rect 8527 10217 8539 10220
rect 8481 10211 8539 10217
rect 9401 10217 9413 10220
rect 9447 10217 9459 10251
rect 9401 10211 9459 10217
rect 10962 10208 10968 10260
rect 11020 10248 11026 10260
rect 11057 10251 11115 10257
rect 11057 10248 11069 10251
rect 11020 10220 11069 10248
rect 11020 10208 11026 10220
rect 11057 10217 11069 10220
rect 11103 10248 11115 10251
rect 11606 10248 11612 10260
rect 11103 10220 11612 10248
rect 11103 10217 11115 10220
rect 11057 10211 11115 10217
rect 11606 10208 11612 10220
rect 11664 10208 11670 10260
rect 12529 10251 12587 10257
rect 12529 10217 12541 10251
rect 12575 10248 12587 10251
rect 12618 10248 12624 10260
rect 12575 10220 12624 10248
rect 12575 10217 12587 10220
rect 12529 10211 12587 10217
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 13814 10248 13820 10260
rect 13775 10220 13820 10248
rect 13814 10208 13820 10220
rect 13872 10208 13878 10260
rect 15102 10248 15108 10260
rect 15063 10220 15108 10248
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 15565 10251 15623 10257
rect 15565 10217 15577 10251
rect 15611 10248 15623 10251
rect 15746 10248 15752 10260
rect 15611 10220 15752 10248
rect 15611 10217 15623 10220
rect 15565 10211 15623 10217
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 18046 10248 18052 10260
rect 18007 10220 18052 10248
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 18506 10248 18512 10260
rect 18467 10220 18512 10248
rect 18506 10208 18512 10220
rect 18564 10208 18570 10260
rect 18966 10248 18972 10260
rect 18927 10220 18972 10248
rect 18966 10208 18972 10220
rect 19024 10248 19030 10260
rect 19426 10248 19432 10260
rect 19024 10220 19432 10248
rect 19024 10208 19030 10220
rect 19426 10208 19432 10220
rect 19484 10208 19490 10260
rect 6914 10180 6920 10192
rect 6875 10152 6920 10180
rect 6914 10140 6920 10152
rect 6972 10140 6978 10192
rect 7929 10183 7987 10189
rect 7929 10149 7941 10183
rect 7975 10180 7987 10183
rect 8202 10180 8208 10192
rect 7975 10152 8208 10180
rect 7975 10149 7987 10152
rect 7929 10143 7987 10149
rect 8202 10140 8208 10152
rect 8260 10140 8266 10192
rect 8570 10140 8576 10192
rect 8628 10180 8634 10192
rect 9033 10183 9091 10189
rect 9033 10180 9045 10183
rect 8628 10152 9045 10180
rect 8628 10140 8634 10152
rect 9033 10149 9045 10152
rect 9079 10149 9091 10183
rect 14182 10180 14188 10192
rect 14143 10152 14188 10180
rect 9033 10143 9091 10149
rect 14182 10140 14188 10152
rect 14240 10140 14246 10192
rect 1762 10112 1768 10124
rect 1723 10084 1768 10112
rect 1762 10072 1768 10084
rect 1820 10112 1826 10124
rect 2409 10115 2467 10121
rect 2409 10112 2421 10115
rect 1820 10084 2421 10112
rect 1820 10072 1826 10084
rect 2409 10081 2421 10084
rect 2455 10081 2467 10115
rect 5258 10112 5264 10124
rect 5219 10084 5264 10112
rect 2409 10075 2467 10081
rect 5258 10072 5264 10084
rect 5316 10072 5322 10124
rect 6822 10112 6828 10124
rect 6783 10084 6828 10112
rect 6822 10072 6828 10084
rect 6880 10072 6886 10124
rect 8389 10115 8447 10121
rect 8389 10081 8401 10115
rect 8435 10112 8447 10115
rect 8754 10112 8760 10124
rect 8435 10084 8760 10112
rect 8435 10081 8447 10084
rect 8389 10075 8447 10081
rect 8754 10072 8760 10084
rect 8812 10072 8818 10124
rect 9933 10115 9991 10121
rect 9933 10112 9945 10115
rect 9600 10084 9945 10112
rect 1670 10004 1676 10056
rect 1728 10044 1734 10056
rect 1857 10047 1915 10053
rect 1857 10044 1869 10047
rect 1728 10016 1869 10044
rect 1728 10004 1734 10016
rect 1857 10013 1869 10016
rect 1903 10013 1915 10047
rect 1857 10007 1915 10013
rect 1946 10004 1952 10056
rect 2004 10044 2010 10056
rect 2004 10016 2049 10044
rect 2004 10004 2010 10016
rect 4982 10004 4988 10056
rect 5040 10044 5046 10056
rect 5353 10047 5411 10053
rect 5353 10044 5365 10047
rect 5040 10016 5365 10044
rect 5040 10004 5046 10016
rect 5353 10013 5365 10016
rect 5399 10013 5411 10047
rect 5353 10007 5411 10013
rect 5442 10004 5448 10056
rect 5500 10044 5506 10056
rect 7101 10047 7159 10053
rect 5500 10016 5545 10044
rect 5500 10004 5506 10016
rect 7101 10013 7113 10047
rect 7147 10013 7159 10047
rect 7101 10007 7159 10013
rect 1394 9976 1400 9988
rect 1355 9948 1400 9976
rect 1394 9936 1400 9948
rect 1452 9936 1458 9988
rect 6546 9936 6552 9988
rect 6604 9976 6610 9988
rect 7116 9976 7144 10007
rect 8294 10004 8300 10056
rect 8352 10044 8358 10056
rect 8573 10047 8631 10053
rect 8573 10044 8585 10047
rect 8352 10016 8585 10044
rect 8352 10004 8358 10016
rect 8573 10013 8585 10016
rect 8619 10044 8631 10047
rect 9600 10044 9628 10084
rect 9933 10081 9945 10084
rect 9979 10081 9991 10115
rect 9933 10075 9991 10081
rect 12434 10072 12440 10124
rect 12492 10112 12498 10124
rect 13173 10115 13231 10121
rect 13173 10112 13185 10115
rect 12492 10084 13185 10112
rect 12492 10072 12498 10084
rect 13173 10081 13185 10084
rect 13219 10081 13231 10115
rect 13173 10075 13231 10081
rect 15930 10072 15936 10124
rect 15988 10112 15994 10124
rect 16298 10121 16304 10124
rect 16281 10115 16304 10121
rect 16281 10112 16293 10115
rect 15988 10084 16293 10112
rect 15988 10072 15994 10084
rect 16281 10081 16293 10084
rect 16356 10112 16362 10124
rect 18874 10112 18880 10124
rect 16356 10084 16429 10112
rect 18835 10084 18880 10112
rect 16281 10075 16304 10081
rect 16298 10072 16304 10075
rect 16356 10072 16362 10084
rect 18874 10072 18880 10084
rect 18932 10072 18938 10124
rect 8619 10016 9628 10044
rect 8619 10013 8631 10016
rect 8573 10007 8631 10013
rect 9674 10004 9680 10056
rect 9732 10044 9738 10056
rect 9732 10016 9777 10044
rect 9732 10004 9738 10016
rect 12618 10004 12624 10056
rect 12676 10044 12682 10056
rect 13262 10044 13268 10056
rect 12676 10016 13268 10044
rect 12676 10004 12682 10016
rect 13262 10004 13268 10016
rect 13320 10004 13326 10056
rect 13446 10044 13452 10056
rect 13407 10016 13452 10044
rect 13446 10004 13452 10016
rect 13504 10004 13510 10056
rect 15838 10004 15844 10056
rect 15896 10044 15902 10056
rect 16022 10044 16028 10056
rect 15896 10016 16028 10044
rect 15896 10004 15902 10016
rect 16022 10004 16028 10016
rect 16080 10004 16086 10056
rect 19058 10044 19064 10056
rect 17420 10016 19064 10044
rect 9122 9976 9128 9988
rect 6604 9948 9128 9976
rect 6604 9936 6610 9948
rect 9122 9936 9128 9948
rect 9180 9936 9186 9988
rect 11790 9976 11796 9988
rect 11072 9948 11796 9976
rect 2774 9868 2780 9920
rect 2832 9908 2838 9920
rect 3053 9911 3111 9917
rect 3053 9908 3065 9911
rect 2832 9880 3065 9908
rect 2832 9868 2838 9880
rect 3053 9877 3065 9880
rect 3099 9877 3111 9911
rect 4338 9908 4344 9920
rect 4299 9880 4344 9908
rect 3053 9871 3111 9877
rect 4338 9868 4344 9880
rect 4396 9868 4402 9920
rect 4614 9908 4620 9920
rect 4575 9880 4620 9908
rect 4614 9868 4620 9880
rect 4672 9868 4678 9920
rect 5534 9868 5540 9920
rect 5592 9908 5598 9920
rect 5905 9911 5963 9917
rect 5905 9908 5917 9911
rect 5592 9880 5917 9908
rect 5592 9868 5598 9880
rect 5905 9877 5917 9880
rect 5951 9877 5963 9911
rect 7466 9908 7472 9920
rect 7427 9880 7472 9908
rect 5905 9871 5963 9877
rect 7466 9868 7472 9880
rect 7524 9868 7530 9920
rect 8018 9908 8024 9920
rect 7979 9880 8024 9908
rect 8018 9868 8024 9880
rect 8076 9868 8082 9920
rect 9858 9868 9864 9920
rect 9916 9908 9922 9920
rect 11072 9908 11100 9948
rect 11790 9936 11796 9948
rect 11848 9936 11854 9988
rect 12805 9979 12863 9985
rect 12805 9945 12817 9979
rect 12851 9976 12863 9979
rect 13630 9976 13636 9988
rect 12851 9948 13636 9976
rect 12851 9945 12863 9948
rect 12805 9939 12863 9945
rect 13630 9936 13636 9948
rect 13688 9936 13694 9988
rect 9916 9880 11100 9908
rect 9916 9868 9922 9880
rect 11146 9868 11152 9920
rect 11204 9908 11210 9920
rect 11609 9911 11667 9917
rect 11609 9908 11621 9911
rect 11204 9880 11621 9908
rect 11204 9868 11210 9880
rect 11609 9877 11621 9880
rect 11655 9877 11667 9911
rect 11974 9908 11980 9920
rect 11935 9880 11980 9908
rect 11609 9871 11667 9877
rect 11974 9868 11980 9880
rect 12032 9868 12038 9920
rect 14550 9908 14556 9920
rect 14511 9880 14556 9908
rect 14550 9868 14556 9880
rect 14608 9868 14614 9920
rect 15930 9908 15936 9920
rect 15891 9880 15936 9908
rect 15930 9868 15936 9880
rect 15988 9868 15994 9920
rect 16942 9868 16948 9920
rect 17000 9908 17006 9920
rect 17420 9917 17448 10016
rect 19058 10004 19064 10016
rect 19116 10004 19122 10056
rect 17405 9911 17463 9917
rect 17405 9908 17417 9911
rect 17000 9880 17417 9908
rect 17000 9868 17006 9880
rect 17405 9877 17417 9880
rect 17451 9877 17463 9911
rect 17405 9871 17463 9877
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 1397 9707 1455 9713
rect 1397 9673 1409 9707
rect 1443 9704 1455 9707
rect 1854 9704 1860 9716
rect 1443 9676 1860 9704
rect 1443 9673 1455 9676
rect 1397 9667 1455 9673
rect 1854 9664 1860 9676
rect 1912 9664 1918 9716
rect 5258 9664 5264 9716
rect 5316 9704 5322 9716
rect 5353 9707 5411 9713
rect 5353 9704 5365 9707
rect 5316 9676 5365 9704
rect 5316 9664 5322 9676
rect 5353 9673 5365 9676
rect 5399 9673 5411 9707
rect 5353 9667 5411 9673
rect 6273 9707 6331 9713
rect 6273 9673 6285 9707
rect 6319 9704 6331 9707
rect 6730 9704 6736 9716
rect 6319 9676 6736 9704
rect 6319 9673 6331 9676
rect 6273 9667 6331 9673
rect 1670 9596 1676 9648
rect 1728 9636 1734 9648
rect 2409 9639 2467 9645
rect 2409 9636 2421 9639
rect 1728 9608 2421 9636
rect 1728 9596 1734 9608
rect 2409 9605 2421 9608
rect 2455 9605 2467 9639
rect 2409 9599 2467 9605
rect 1946 9568 1952 9580
rect 1907 9540 1952 9568
rect 1946 9528 1952 9540
rect 2004 9568 2010 9580
rect 2958 9568 2964 9580
rect 2004 9540 2964 9568
rect 2004 9528 2010 9540
rect 2958 9528 2964 9540
rect 3016 9528 3022 9580
rect 5368 9568 5396 9667
rect 6730 9664 6736 9676
rect 6788 9664 6794 9716
rect 7098 9704 7104 9716
rect 6840 9676 7104 9704
rect 5537 9571 5595 9577
rect 5537 9568 5549 9571
rect 5368 9540 5549 9568
rect 5537 9537 5549 9540
rect 5583 9537 5595 9571
rect 5537 9531 5595 9537
rect 1486 9460 1492 9512
rect 1544 9500 1550 9512
rect 2774 9500 2780 9512
rect 1544 9472 2780 9500
rect 1544 9460 1550 9472
rect 2774 9460 2780 9472
rect 2832 9500 2838 9512
rect 3053 9503 3111 9509
rect 3053 9500 3065 9503
rect 2832 9472 3065 9500
rect 2832 9460 2838 9472
rect 3053 9469 3065 9472
rect 3099 9469 3111 9503
rect 3053 9463 3111 9469
rect 3142 9460 3148 9512
rect 3200 9500 3206 9512
rect 3320 9503 3378 9509
rect 3320 9500 3332 9503
rect 3200 9472 3332 9500
rect 3200 9460 3206 9472
rect 3320 9469 3332 9472
rect 3366 9500 3378 9503
rect 3786 9500 3792 9512
rect 3366 9472 3792 9500
rect 3366 9469 3378 9472
rect 3320 9463 3378 9469
rect 3786 9460 3792 9472
rect 3844 9460 3850 9512
rect 6840 9509 6868 9676
rect 7098 9664 7104 9676
rect 7156 9664 7162 9716
rect 9674 9664 9680 9716
rect 9732 9704 9738 9716
rect 12618 9704 12624 9716
rect 9732 9676 9777 9704
rect 12360 9676 12624 9704
rect 9732 9664 9738 9676
rect 8110 9596 8116 9648
rect 8168 9636 8174 9648
rect 8205 9639 8263 9645
rect 8205 9636 8217 9639
rect 8168 9608 8217 9636
rect 8168 9596 8174 9608
rect 8205 9605 8217 9608
rect 8251 9605 8263 9639
rect 8205 9599 8263 9605
rect 12253 9639 12311 9645
rect 12253 9605 12265 9639
rect 12299 9636 12311 9639
rect 12360 9636 12388 9676
rect 12618 9664 12624 9676
rect 12676 9664 12682 9716
rect 12710 9664 12716 9716
rect 12768 9704 12774 9716
rect 13262 9704 13268 9716
rect 12768 9676 13268 9704
rect 12768 9664 12774 9676
rect 13262 9664 13268 9676
rect 13320 9664 13326 9716
rect 19058 9704 19064 9716
rect 19019 9676 19064 9704
rect 19058 9664 19064 9676
rect 19116 9664 19122 9716
rect 19334 9664 19340 9716
rect 19392 9704 19398 9716
rect 20162 9704 20168 9716
rect 19392 9676 20168 9704
rect 19392 9664 19398 9676
rect 20162 9664 20168 9676
rect 20220 9664 20226 9716
rect 12299 9608 12388 9636
rect 15197 9639 15255 9645
rect 12299 9605 12311 9608
rect 12253 9599 12311 9605
rect 15197 9605 15209 9639
rect 15243 9636 15255 9639
rect 15378 9636 15384 9648
rect 15243 9608 15384 9636
rect 15243 9605 15255 9608
rect 15197 9599 15255 9605
rect 15378 9596 15384 9608
rect 15436 9596 15442 9648
rect 16298 9636 16304 9648
rect 16259 9608 16304 9636
rect 16298 9596 16304 9608
rect 16356 9596 16362 9648
rect 18049 9639 18107 9645
rect 18049 9636 18061 9639
rect 16684 9608 18061 9636
rect 7926 9528 7932 9580
rect 7984 9568 7990 9580
rect 9582 9568 9588 9580
rect 7984 9540 9588 9568
rect 7984 9528 7990 9540
rect 9582 9528 9588 9540
rect 9640 9528 9646 9580
rect 10321 9571 10379 9577
rect 10321 9537 10333 9571
rect 10367 9568 10379 9571
rect 11330 9568 11336 9580
rect 10367 9540 11336 9568
rect 10367 9537 10379 9540
rect 10321 9531 10379 9537
rect 11330 9528 11336 9540
rect 11388 9528 11394 9580
rect 6825 9503 6883 9509
rect 6825 9500 6837 9503
rect 6564 9472 6837 9500
rect 1857 9435 1915 9441
rect 1857 9401 1869 9435
rect 1903 9432 1915 9435
rect 2038 9432 2044 9444
rect 1903 9404 2044 9432
rect 1903 9401 1915 9404
rect 1857 9395 1915 9401
rect 2038 9392 2044 9404
rect 2096 9432 2102 9444
rect 2096 9404 2728 9432
rect 2096 9392 2102 9404
rect 1765 9367 1823 9373
rect 1765 9333 1777 9367
rect 1811 9364 1823 9367
rect 2222 9364 2228 9376
rect 1811 9336 2228 9364
rect 1811 9333 1823 9336
rect 1765 9327 1823 9333
rect 2222 9324 2228 9336
rect 2280 9324 2286 9376
rect 2700 9364 2728 9404
rect 2777 9367 2835 9373
rect 2777 9364 2789 9367
rect 2700 9336 2789 9364
rect 2777 9333 2789 9336
rect 2823 9333 2835 9367
rect 2777 9327 2835 9333
rect 4433 9367 4491 9373
rect 4433 9333 4445 9367
rect 4479 9364 4491 9367
rect 4522 9364 4528 9376
rect 4479 9336 4528 9364
rect 4479 9333 4491 9336
rect 4433 9327 4491 9333
rect 4522 9324 4528 9336
rect 4580 9324 4586 9376
rect 4982 9364 4988 9376
rect 4943 9336 4988 9364
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 6454 9324 6460 9376
rect 6512 9364 6518 9376
rect 6564 9373 6592 9472
rect 6825 9469 6837 9472
rect 6871 9469 6883 9503
rect 6825 9463 6883 9469
rect 7092 9503 7150 9509
rect 7092 9469 7104 9503
rect 7138 9500 7150 9503
rect 7466 9500 7472 9512
rect 7138 9472 7472 9500
rect 7138 9469 7150 9472
rect 7092 9463 7150 9469
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 13630 9460 13636 9512
rect 13688 9500 13694 9512
rect 13817 9503 13875 9509
rect 13817 9500 13829 9503
rect 13688 9472 13829 9500
rect 13688 9460 13694 9472
rect 13817 9469 13829 9472
rect 13863 9500 13875 9503
rect 16022 9500 16028 9512
rect 13863 9472 16028 9500
rect 13863 9469 13875 9472
rect 13817 9463 13875 9469
rect 16022 9460 16028 9472
rect 16080 9460 16086 9512
rect 16684 9509 16712 9608
rect 18049 9605 18061 9608
rect 18095 9636 18107 9639
rect 18966 9636 18972 9648
rect 18095 9608 18972 9636
rect 18095 9605 18107 9608
rect 18049 9599 18107 9605
rect 18966 9596 18972 9608
rect 19024 9596 19030 9648
rect 19426 9596 19432 9648
rect 19484 9636 19490 9648
rect 19797 9639 19855 9645
rect 19797 9636 19809 9639
rect 19484 9608 19809 9636
rect 19484 9596 19490 9608
rect 19797 9605 19809 9608
rect 19843 9605 19855 9639
rect 19797 9599 19855 9605
rect 16758 9528 16764 9580
rect 16816 9568 16822 9580
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16816 9540 16865 9568
rect 16816 9528 16822 9540
rect 16853 9537 16865 9540
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 17954 9528 17960 9580
rect 18012 9568 18018 9580
rect 18598 9568 18604 9580
rect 18012 9540 18604 9568
rect 18012 9528 18018 9540
rect 18598 9528 18604 9540
rect 18656 9528 18662 9580
rect 16669 9503 16727 9509
rect 16669 9469 16681 9503
rect 16715 9469 16727 9503
rect 17586 9500 17592 9512
rect 16669 9463 16727 9469
rect 16776 9472 17592 9500
rect 11241 9435 11299 9441
rect 11241 9432 11253 9435
rect 10612 9404 11253 9432
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 6512 9336 6561 9364
rect 6512 9324 6518 9336
rect 6549 9333 6561 9336
rect 6595 9333 6607 9367
rect 6549 9327 6607 9333
rect 8294 9324 8300 9376
rect 8352 9364 8358 9376
rect 8757 9367 8815 9373
rect 8757 9364 8769 9367
rect 8352 9336 8769 9364
rect 8352 9324 8358 9336
rect 8757 9333 8769 9336
rect 8803 9364 8815 9367
rect 9309 9367 9367 9373
rect 9309 9364 9321 9367
rect 8803 9336 9321 9364
rect 8803 9333 8815 9336
rect 8757 9327 8815 9333
rect 9309 9333 9321 9336
rect 9355 9333 9367 9367
rect 9309 9327 9367 9333
rect 10042 9324 10048 9376
rect 10100 9364 10106 9376
rect 10612 9373 10640 9404
rect 11241 9401 11253 9404
rect 11287 9432 11299 9435
rect 11606 9432 11612 9444
rect 11287 9404 11612 9432
rect 11287 9401 11299 9404
rect 11241 9395 11299 9401
rect 11606 9392 11612 9404
rect 11664 9392 11670 9444
rect 12897 9435 12955 9441
rect 12897 9401 12909 9435
rect 12943 9432 12955 9435
rect 13446 9432 13452 9444
rect 12943 9404 13452 9432
rect 12943 9401 12955 9404
rect 12897 9395 12955 9401
rect 13446 9392 13452 9404
rect 13504 9432 13510 9444
rect 13906 9432 13912 9444
rect 13504 9404 13912 9432
rect 13504 9392 13510 9404
rect 13906 9392 13912 9404
rect 13964 9432 13970 9444
rect 16776 9441 16804 9472
rect 17586 9460 17592 9472
rect 17644 9500 17650 9512
rect 19429 9503 19487 9509
rect 19429 9500 19441 9503
rect 17644 9472 19441 9500
rect 17644 9460 17650 9472
rect 19429 9469 19441 9472
rect 19475 9469 19487 9503
rect 19429 9463 19487 9469
rect 14062 9435 14120 9441
rect 14062 9432 14074 9435
rect 13964 9404 14074 9432
rect 13964 9392 13970 9404
rect 14062 9401 14074 9404
rect 14108 9401 14120 9435
rect 14062 9395 14120 9401
rect 16761 9435 16819 9441
rect 16761 9401 16773 9435
rect 16807 9401 16819 9435
rect 18417 9435 18475 9441
rect 18417 9432 18429 9435
rect 16761 9395 16819 9401
rect 17420 9404 18429 9432
rect 17420 9376 17448 9404
rect 18417 9401 18429 9404
rect 18463 9401 18475 9435
rect 18417 9395 18475 9401
rect 10597 9367 10655 9373
rect 10597 9364 10609 9367
rect 10100 9336 10609 9364
rect 10100 9324 10106 9336
rect 10597 9333 10609 9336
rect 10643 9333 10655 9367
rect 10778 9364 10784 9376
rect 10739 9336 10784 9364
rect 10597 9327 10655 9333
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 10870 9324 10876 9376
rect 10928 9364 10934 9376
rect 11149 9367 11207 9373
rect 11149 9364 11161 9367
rect 10928 9336 11161 9364
rect 10928 9324 10934 9336
rect 11149 9333 11161 9336
rect 11195 9333 11207 9367
rect 11149 9327 11207 9333
rect 11698 9324 11704 9376
rect 11756 9364 11762 9376
rect 11793 9367 11851 9373
rect 11793 9364 11805 9367
rect 11756 9336 11805 9364
rect 11756 9324 11762 9336
rect 11793 9333 11805 9336
rect 11839 9364 11851 9367
rect 12342 9364 12348 9376
rect 11839 9336 12348 9364
rect 11839 9333 11851 9336
rect 11793 9327 11851 9333
rect 12342 9324 12348 9336
rect 12400 9324 12406 9376
rect 13630 9364 13636 9376
rect 13591 9336 13636 9364
rect 13630 9324 13636 9336
rect 13688 9324 13694 9376
rect 17402 9364 17408 9376
rect 17363 9336 17408 9364
rect 17402 9324 17408 9336
rect 17460 9324 17466 9376
rect 17770 9364 17776 9376
rect 17731 9336 17776 9364
rect 17770 9324 17776 9336
rect 17828 9364 17834 9376
rect 18509 9367 18567 9373
rect 18509 9364 18521 9367
rect 17828 9336 18521 9364
rect 17828 9324 17834 9336
rect 18509 9333 18521 9336
rect 18555 9333 18567 9367
rect 18509 9327 18567 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 2958 9120 2964 9172
rect 3016 9160 3022 9172
rect 3421 9163 3479 9169
rect 3421 9160 3433 9163
rect 3016 9132 3433 9160
rect 3016 9120 3022 9132
rect 3421 9129 3433 9132
rect 3467 9129 3479 9163
rect 3421 9123 3479 9129
rect 5445 9163 5503 9169
rect 5445 9129 5457 9163
rect 5491 9160 5503 9163
rect 5534 9160 5540 9172
rect 5491 9132 5540 9160
rect 5491 9129 5503 9132
rect 5445 9123 5503 9129
rect 5534 9120 5540 9132
rect 5592 9120 5598 9172
rect 6546 9160 6552 9172
rect 6507 9132 6552 9160
rect 6546 9120 6552 9132
rect 6604 9120 6610 9172
rect 8018 9160 8024 9172
rect 7979 9132 8024 9160
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 8386 9160 8392 9172
rect 8347 9132 8392 9160
rect 8386 9120 8392 9132
rect 8444 9160 8450 9172
rect 8662 9160 8668 9172
rect 8444 9132 8668 9160
rect 8444 9120 8450 9132
rect 8662 9120 8668 9132
rect 8720 9120 8726 9172
rect 9677 9163 9735 9169
rect 9677 9129 9689 9163
rect 9723 9160 9735 9163
rect 9766 9160 9772 9172
rect 9723 9132 9772 9160
rect 9723 9129 9735 9132
rect 9677 9123 9735 9129
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 10134 9160 10140 9172
rect 10095 9132 10140 9160
rect 10134 9120 10140 9132
rect 10192 9120 10198 9172
rect 10778 9120 10784 9172
rect 10836 9160 10842 9172
rect 11609 9163 11667 9169
rect 11609 9160 11621 9163
rect 10836 9132 11621 9160
rect 10836 9120 10842 9132
rect 11609 9129 11621 9132
rect 11655 9160 11667 9163
rect 12066 9160 12072 9172
rect 11655 9132 12072 9160
rect 11655 9129 11667 9132
rect 11609 9123 11667 9129
rect 12066 9120 12072 9132
rect 12124 9120 12130 9172
rect 15657 9163 15715 9169
rect 15657 9129 15669 9163
rect 15703 9160 15715 9163
rect 17402 9160 17408 9172
rect 15703 9132 17408 9160
rect 15703 9129 15715 9132
rect 15657 9123 15715 9129
rect 17402 9120 17408 9132
rect 17460 9120 17466 9172
rect 18966 9160 18972 9172
rect 18927 9132 18972 9160
rect 18966 9120 18972 9132
rect 19024 9120 19030 9172
rect 19334 9160 19340 9172
rect 19295 9132 19340 9160
rect 19334 9120 19340 9132
rect 19392 9120 19398 9172
rect 2866 9052 2872 9104
rect 2924 9092 2930 9104
rect 4065 9095 4123 9101
rect 4065 9092 4077 9095
rect 2924 9064 4077 9092
rect 2924 9052 2930 9064
rect 4065 9061 4077 9064
rect 4111 9061 4123 9095
rect 4065 9055 4123 9061
rect 11054 9052 11060 9104
rect 11112 9092 11118 9104
rect 11149 9095 11207 9101
rect 11149 9092 11161 9095
rect 11112 9064 11161 9092
rect 11112 9052 11118 9064
rect 11149 9061 11161 9064
rect 11195 9061 11207 9095
rect 14918 9092 14924 9104
rect 14879 9064 14924 9092
rect 11149 9055 11207 9061
rect 14918 9052 14924 9064
rect 14976 9052 14982 9104
rect 15565 9095 15623 9101
rect 15565 9061 15577 9095
rect 15611 9092 15623 9095
rect 15930 9092 15936 9104
rect 15611 9064 15936 9092
rect 15611 9061 15623 9064
rect 15565 9055 15623 9061
rect 15930 9052 15936 9064
rect 15988 9092 15994 9104
rect 16485 9095 16543 9101
rect 16485 9092 16497 9095
rect 15988 9064 16497 9092
rect 15988 9052 15994 9064
rect 16485 9061 16497 9064
rect 16531 9092 16543 9095
rect 16758 9092 16764 9104
rect 16531 9064 16764 9092
rect 16531 9061 16543 9064
rect 16485 9055 16543 9061
rect 16758 9052 16764 9064
rect 16816 9052 16822 9104
rect 1486 9024 1492 9036
rect 1447 8996 1492 9024
rect 1486 8984 1492 8996
rect 1544 8984 1550 9036
rect 1756 9027 1814 9033
rect 1756 8993 1768 9027
rect 1802 9024 1814 9027
rect 4985 9027 5043 9033
rect 1802 8996 2728 9024
rect 1802 8993 1814 8996
rect 1756 8987 1814 8993
rect 2700 8956 2728 8996
rect 4985 8993 4997 9027
rect 5031 9024 5043 9027
rect 5353 9027 5411 9033
rect 5353 9024 5365 9027
rect 5031 8996 5365 9024
rect 5031 8993 5043 8996
rect 4985 8987 5043 8993
rect 5353 8993 5365 8996
rect 5399 9024 5411 9027
rect 5442 9024 5448 9036
rect 5399 8996 5448 9024
rect 5399 8993 5411 8996
rect 5353 8987 5411 8993
rect 5442 8984 5448 8996
rect 5500 8984 5506 9036
rect 5534 8984 5540 9036
rect 5592 9024 5598 9036
rect 5813 9027 5871 9033
rect 5813 9024 5825 9027
rect 5592 8996 5825 9024
rect 5592 8984 5598 8996
rect 5813 8993 5825 8996
rect 5859 8993 5871 9027
rect 5813 8987 5871 8993
rect 5905 9027 5963 9033
rect 5905 8993 5917 9027
rect 5951 9024 5963 9027
rect 6270 9024 6276 9036
rect 5951 8996 6276 9024
rect 5951 8993 5963 8996
rect 5905 8987 5963 8993
rect 6270 8984 6276 8996
rect 6328 8984 6334 9036
rect 8481 9027 8539 9033
rect 8481 8993 8493 9027
rect 8527 9024 8539 9027
rect 9582 9024 9588 9036
rect 8527 8996 9588 9024
rect 8527 8993 8539 8996
rect 8481 8987 8539 8993
rect 9582 8984 9588 8996
rect 9640 8984 9646 9036
rect 10042 9024 10048 9036
rect 10003 8996 10048 9024
rect 10042 8984 10048 8996
rect 10100 8984 10106 9036
rect 11330 8984 11336 9036
rect 11388 9024 11394 9036
rect 11882 9024 11888 9036
rect 11388 8996 11888 9024
rect 11388 8984 11394 8996
rect 11882 8984 11888 8996
rect 11940 9024 11946 9036
rect 12049 9027 12107 9033
rect 12049 9024 12061 9027
rect 11940 8996 12061 9024
rect 11940 8984 11946 8996
rect 12049 8993 12061 8996
rect 12095 8993 12107 9027
rect 12049 8987 12107 8993
rect 16022 8984 16028 9036
rect 16080 9024 16086 9036
rect 16666 9024 16672 9036
rect 16080 8996 16672 9024
rect 16080 8984 16086 8996
rect 16666 8984 16672 8996
rect 16724 8984 16730 9036
rect 16942 9033 16948 9036
rect 16936 9024 16948 9033
rect 16903 8996 16948 9024
rect 16936 8987 16948 8996
rect 16942 8984 16948 8987
rect 17000 8984 17006 9036
rect 3234 8956 3240 8968
rect 2700 8928 3240 8956
rect 3234 8916 3240 8928
rect 3292 8916 3298 8968
rect 5460 8956 5488 8984
rect 5997 8959 6055 8965
rect 5997 8956 6009 8959
rect 5460 8928 6009 8956
rect 5997 8925 6009 8928
rect 6043 8925 6055 8959
rect 5997 8919 6055 8925
rect 8573 8959 8631 8965
rect 8573 8925 8585 8959
rect 8619 8925 8631 8959
rect 8573 8919 8631 8925
rect 10321 8959 10379 8965
rect 10321 8925 10333 8959
rect 10367 8956 10379 8959
rect 10962 8956 10968 8968
rect 10367 8928 10968 8956
rect 10367 8925 10379 8928
rect 10321 8919 10379 8925
rect 2869 8891 2927 8897
rect 2869 8857 2881 8891
rect 2915 8888 2927 8891
rect 3142 8888 3148 8900
rect 2915 8860 3148 8888
rect 2915 8857 2927 8860
rect 2869 8851 2927 8857
rect 3142 8848 3148 8860
rect 3200 8848 3206 8900
rect 3252 8888 3280 8916
rect 3789 8891 3847 8897
rect 3789 8888 3801 8891
rect 3252 8860 3801 8888
rect 3789 8857 3801 8860
rect 3835 8888 3847 8891
rect 3878 8888 3884 8900
rect 3835 8860 3884 8888
rect 3835 8857 3847 8860
rect 3789 8851 3847 8857
rect 3878 8848 3884 8860
rect 3936 8888 3942 8900
rect 4525 8891 4583 8897
rect 4525 8888 4537 8891
rect 3936 8860 4537 8888
rect 3936 8848 3942 8860
rect 4525 8857 4537 8860
rect 4571 8857 4583 8891
rect 4525 8851 4583 8857
rect 8294 8848 8300 8900
rect 8352 8888 8358 8900
rect 8588 8888 8616 8919
rect 10962 8916 10968 8928
rect 11020 8916 11026 8968
rect 11422 8916 11428 8968
rect 11480 8956 11486 8968
rect 11793 8959 11851 8965
rect 11793 8956 11805 8959
rect 11480 8928 11805 8956
rect 11480 8916 11486 8928
rect 11793 8925 11805 8928
rect 11839 8925 11851 8959
rect 11793 8919 11851 8925
rect 13814 8916 13820 8968
rect 13872 8956 13878 8968
rect 14185 8959 14243 8965
rect 14185 8956 14197 8959
rect 13872 8928 14197 8956
rect 13872 8916 13878 8928
rect 14185 8925 14197 8928
rect 14231 8925 14243 8959
rect 14550 8956 14556 8968
rect 14511 8928 14556 8956
rect 14185 8919 14243 8925
rect 14550 8916 14556 8928
rect 14608 8916 14614 8968
rect 16209 8959 16267 8965
rect 16209 8925 16221 8959
rect 16255 8956 16267 8959
rect 16482 8956 16488 8968
rect 16255 8928 16488 8956
rect 16255 8925 16267 8928
rect 16209 8919 16267 8925
rect 16482 8916 16488 8928
rect 16540 8916 16546 8968
rect 9401 8891 9459 8897
rect 9401 8888 9413 8891
rect 8352 8860 8616 8888
rect 8680 8860 9413 8888
rect 8352 8848 8358 8860
rect 6914 8820 6920 8832
rect 6875 8792 6920 8820
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 7190 8820 7196 8832
rect 7151 8792 7196 8820
rect 7190 8780 7196 8792
rect 7248 8780 7254 8832
rect 7282 8780 7288 8832
rect 7340 8820 7346 8832
rect 7561 8823 7619 8829
rect 7561 8820 7573 8823
rect 7340 8792 7573 8820
rect 7340 8780 7346 8792
rect 7561 8789 7573 8792
rect 7607 8789 7619 8823
rect 7561 8783 7619 8789
rect 8202 8780 8208 8832
rect 8260 8820 8266 8832
rect 8680 8820 8708 8860
rect 9401 8857 9413 8860
rect 9447 8857 9459 8891
rect 9401 8851 9459 8857
rect 8260 8792 8708 8820
rect 8260 8780 8266 8792
rect 8938 8780 8944 8832
rect 8996 8820 9002 8832
rect 9033 8823 9091 8829
rect 9033 8820 9045 8823
rect 8996 8792 9045 8820
rect 8996 8780 9002 8792
rect 9033 8789 9045 8792
rect 9079 8789 9091 8823
rect 10870 8820 10876 8832
rect 10831 8792 10876 8820
rect 9033 8783 9091 8789
rect 10870 8780 10876 8792
rect 10928 8780 10934 8832
rect 13078 8780 13084 8832
rect 13136 8820 13142 8832
rect 13173 8823 13231 8829
rect 13173 8820 13185 8823
rect 13136 8792 13185 8820
rect 13136 8780 13142 8792
rect 13173 8789 13185 8792
rect 13219 8789 13231 8823
rect 13906 8820 13912 8832
rect 13867 8792 13912 8820
rect 13173 8783 13231 8789
rect 13906 8780 13912 8792
rect 13964 8780 13970 8832
rect 17954 8780 17960 8832
rect 18012 8820 18018 8832
rect 18049 8823 18107 8829
rect 18049 8820 18061 8823
rect 18012 8792 18061 8820
rect 18012 8780 18018 8792
rect 18049 8789 18061 8792
rect 18095 8789 18107 8823
rect 18598 8820 18604 8832
rect 18559 8792 18604 8820
rect 18049 8783 18107 8789
rect 18598 8780 18604 8792
rect 18656 8780 18662 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 2498 8576 2504 8628
rect 2556 8616 2562 8628
rect 2685 8619 2743 8625
rect 2685 8616 2697 8619
rect 2556 8588 2697 8616
rect 2556 8576 2562 8588
rect 2685 8585 2697 8588
rect 2731 8585 2743 8619
rect 2685 8579 2743 8585
rect 8294 8576 8300 8628
rect 8352 8616 8358 8628
rect 10045 8619 10103 8625
rect 10045 8616 10057 8619
rect 8352 8588 10057 8616
rect 8352 8576 8358 8588
rect 10045 8585 10057 8588
rect 10091 8585 10103 8619
rect 10045 8579 10103 8585
rect 10689 8619 10747 8625
rect 10689 8585 10701 8619
rect 10735 8616 10747 8619
rect 10962 8616 10968 8628
rect 10735 8588 10968 8616
rect 10735 8585 10747 8588
rect 10689 8579 10747 8585
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 11422 8576 11428 8628
rect 11480 8616 11486 8628
rect 11793 8619 11851 8625
rect 11793 8616 11805 8619
rect 11480 8588 11805 8616
rect 11480 8576 11486 8588
rect 11793 8585 11805 8588
rect 11839 8585 11851 8619
rect 11793 8579 11851 8585
rect 11808 8548 11836 8579
rect 11882 8576 11888 8628
rect 11940 8616 11946 8628
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 11940 8588 12173 8616
rect 11940 8576 11946 8588
rect 12161 8585 12173 8588
rect 12207 8585 12219 8619
rect 13630 8616 13636 8628
rect 12161 8579 12219 8585
rect 13004 8588 13636 8616
rect 12805 8551 12863 8557
rect 12805 8548 12817 8551
rect 11808 8520 12817 8548
rect 12805 8517 12817 8520
rect 12851 8548 12863 8551
rect 13004 8548 13032 8588
rect 13630 8576 13636 8588
rect 13688 8576 13694 8628
rect 13906 8576 13912 8628
rect 13964 8616 13970 8628
rect 14369 8619 14427 8625
rect 14369 8616 14381 8619
rect 13964 8588 14381 8616
rect 13964 8576 13970 8588
rect 14369 8585 14381 8588
rect 14415 8585 14427 8619
rect 14369 8579 14427 8585
rect 16666 8576 16672 8628
rect 16724 8616 16730 8628
rect 17129 8619 17187 8625
rect 17129 8616 17141 8619
rect 16724 8588 17141 8616
rect 16724 8576 16730 8588
rect 17129 8585 17141 8588
rect 17175 8585 17187 8619
rect 17129 8579 17187 8585
rect 17865 8619 17923 8625
rect 17865 8585 17877 8619
rect 17911 8616 17923 8619
rect 18046 8616 18052 8628
rect 17911 8588 18052 8616
rect 17911 8585 17923 8588
rect 17865 8579 17923 8585
rect 18046 8576 18052 8588
rect 18104 8616 18110 8628
rect 18104 8588 18552 8616
rect 18104 8576 18110 8588
rect 12851 8520 13032 8548
rect 12851 8517 12863 8520
rect 12805 8511 12863 8517
rect 1397 8483 1455 8489
rect 1397 8449 1409 8483
rect 1443 8480 1455 8483
rect 1762 8480 1768 8492
rect 1443 8452 1768 8480
rect 1443 8449 1455 8452
rect 1397 8443 1455 8449
rect 1762 8440 1768 8452
rect 1820 8440 1826 8492
rect 3142 8480 3148 8492
rect 3103 8452 3148 8480
rect 3142 8440 3148 8452
rect 3200 8440 3206 8492
rect 3234 8440 3240 8492
rect 3292 8480 3298 8492
rect 6638 8480 6644 8492
rect 3292 8452 3337 8480
rect 6599 8452 6644 8480
rect 3292 8440 3298 8452
rect 6638 8440 6644 8452
rect 6696 8480 6702 8492
rect 6696 8452 7144 8480
rect 6696 8440 6702 8452
rect 4522 8421 4528 8424
rect 3973 8415 4031 8421
rect 3973 8381 3985 8415
rect 4019 8412 4031 8415
rect 4249 8415 4307 8421
rect 4249 8412 4261 8415
rect 4019 8384 4261 8412
rect 4019 8381 4031 8384
rect 3973 8375 4031 8381
rect 4249 8381 4261 8384
rect 4295 8381 4307 8415
rect 4516 8412 4528 8421
rect 4249 8375 4307 8381
rect 4356 8384 4528 8412
rect 2590 8344 2596 8356
rect 2503 8316 2596 8344
rect 2590 8304 2596 8316
rect 2648 8344 2654 8356
rect 3053 8347 3111 8353
rect 3053 8344 3065 8347
rect 2648 8316 3065 8344
rect 2648 8304 2654 8316
rect 3053 8313 3065 8316
rect 3099 8313 3111 8347
rect 3053 8307 3111 8313
rect 3602 8304 3608 8356
rect 3660 8344 3666 8356
rect 3789 8347 3847 8353
rect 3789 8344 3801 8347
rect 3660 8316 3801 8344
rect 3660 8304 3666 8316
rect 3789 8313 3801 8316
rect 3835 8344 3847 8347
rect 4356 8344 4384 8384
rect 4516 8375 4528 8384
rect 4522 8372 4528 8375
rect 4580 8372 4586 8424
rect 6270 8412 6276 8424
rect 6183 8384 6276 8412
rect 6270 8372 6276 8384
rect 6328 8412 6334 8424
rect 6730 8412 6736 8424
rect 6328 8384 6736 8412
rect 6328 8372 6334 8384
rect 6730 8372 6736 8384
rect 6788 8372 6794 8424
rect 7116 8412 7144 8452
rect 7190 8440 7196 8492
rect 7248 8480 7254 8492
rect 7377 8483 7435 8489
rect 7377 8480 7389 8483
rect 7248 8452 7389 8480
rect 7248 8440 7254 8452
rect 7377 8449 7389 8452
rect 7423 8449 7435 8483
rect 7377 8443 7435 8449
rect 10870 8440 10876 8492
rect 10928 8480 10934 8492
rect 13004 8489 13032 8520
rect 15289 8551 15347 8557
rect 15289 8517 15301 8551
rect 15335 8548 15347 8551
rect 16117 8551 16175 8557
rect 16117 8548 16129 8551
rect 15335 8520 16129 8548
rect 15335 8517 15347 8520
rect 15289 8511 15347 8517
rect 16117 8517 16129 8520
rect 16163 8548 16175 8551
rect 16390 8548 16396 8560
rect 16163 8520 16396 8548
rect 16163 8517 16175 8520
rect 16117 8511 16175 8517
rect 16390 8508 16396 8520
rect 16448 8508 16454 8560
rect 11333 8483 11391 8489
rect 11333 8480 11345 8483
rect 10928 8452 11345 8480
rect 10928 8440 10934 8452
rect 11333 8449 11345 8452
rect 11379 8449 11391 8483
rect 11333 8443 11391 8449
rect 12989 8483 13047 8489
rect 12989 8449 13001 8483
rect 13035 8449 13047 8483
rect 12989 8443 13047 8449
rect 15838 8440 15844 8492
rect 15896 8480 15902 8492
rect 18524 8489 18552 8588
rect 16669 8483 16727 8489
rect 16669 8480 16681 8483
rect 15896 8452 16681 8480
rect 15896 8440 15902 8452
rect 16669 8449 16681 8452
rect 16715 8449 16727 8483
rect 16669 8443 16727 8449
rect 18509 8483 18567 8489
rect 18509 8449 18521 8483
rect 18555 8449 18567 8483
rect 18690 8480 18696 8492
rect 18651 8452 18696 8480
rect 18509 8443 18567 8449
rect 18690 8440 18696 8452
rect 18748 8440 18754 8492
rect 7285 8415 7343 8421
rect 7285 8412 7297 8415
rect 7116 8384 7297 8412
rect 7285 8381 7297 8384
rect 7331 8381 7343 8415
rect 7285 8375 7343 8381
rect 8573 8415 8631 8421
rect 8573 8381 8585 8415
rect 8619 8412 8631 8415
rect 8665 8415 8723 8421
rect 8665 8412 8677 8415
rect 8619 8384 8677 8412
rect 8619 8381 8631 8384
rect 8573 8375 8631 8381
rect 8665 8381 8677 8384
rect 8711 8412 8723 8415
rect 9490 8412 9496 8424
rect 8711 8384 9496 8412
rect 8711 8381 8723 8384
rect 8665 8375 8723 8381
rect 9490 8372 9496 8384
rect 9548 8372 9554 8424
rect 15930 8412 15936 8424
rect 15891 8384 15936 8412
rect 15930 8372 15936 8384
rect 15988 8412 15994 8424
rect 16577 8415 16635 8421
rect 16577 8412 16589 8415
rect 15988 8384 16589 8412
rect 15988 8372 15994 8384
rect 16577 8381 16589 8384
rect 16623 8412 16635 8415
rect 17770 8412 17776 8424
rect 16623 8384 17776 8412
rect 16623 8381 16635 8384
rect 16577 8375 16635 8381
rect 17770 8372 17776 8384
rect 17828 8372 17834 8424
rect 3835 8316 4384 8344
rect 5460 8316 6868 8344
rect 3835 8313 3847 8316
rect 3789 8307 3847 8313
rect 1949 8279 2007 8285
rect 1949 8245 1961 8279
rect 1995 8276 2007 8279
rect 2222 8276 2228 8288
rect 1995 8248 2228 8276
rect 1995 8245 2007 8248
rect 1949 8239 2007 8245
rect 2222 8236 2228 8248
rect 2280 8236 2286 8288
rect 2774 8236 2780 8288
rect 2832 8276 2838 8288
rect 3973 8279 4031 8285
rect 3973 8276 3985 8279
rect 2832 8248 3985 8276
rect 2832 8236 2838 8248
rect 3973 8245 3985 8248
rect 4019 8276 4031 8279
rect 4065 8279 4123 8285
rect 4065 8276 4077 8279
rect 4019 8248 4077 8276
rect 4019 8245 4031 8248
rect 3973 8239 4031 8245
rect 4065 8245 4077 8248
rect 4111 8245 4123 8279
rect 4065 8239 4123 8245
rect 4614 8236 4620 8288
rect 4672 8276 4678 8288
rect 5460 8276 5488 8316
rect 4672 8248 5488 8276
rect 5629 8279 5687 8285
rect 4672 8236 4678 8248
rect 5629 8245 5641 8279
rect 5675 8276 5687 8279
rect 6178 8276 6184 8288
rect 5675 8248 6184 8276
rect 5675 8245 5687 8248
rect 5629 8239 5687 8245
rect 6178 8236 6184 8248
rect 6236 8236 6242 8288
rect 6840 8285 6868 8316
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 7193 8347 7251 8353
rect 7193 8344 7205 8347
rect 6972 8316 7205 8344
rect 6972 8304 6978 8316
rect 7193 8313 7205 8316
rect 7239 8344 7251 8347
rect 7742 8344 7748 8356
rect 7239 8316 7748 8344
rect 7239 8313 7251 8316
rect 7193 8307 7251 8313
rect 7742 8304 7748 8316
rect 7800 8304 7806 8356
rect 8205 8347 8263 8353
rect 8205 8313 8217 8347
rect 8251 8344 8263 8347
rect 8932 8347 8990 8353
rect 8932 8344 8944 8347
rect 8251 8316 8944 8344
rect 8251 8313 8263 8316
rect 8205 8307 8263 8313
rect 8932 8313 8944 8316
rect 8978 8344 8990 8347
rect 9122 8344 9128 8356
rect 8978 8316 9128 8344
rect 8978 8313 8990 8316
rect 8932 8307 8990 8313
rect 9122 8304 9128 8316
rect 9180 8304 9186 8356
rect 13078 8304 13084 8356
rect 13136 8344 13142 8356
rect 13234 8347 13292 8353
rect 13234 8344 13246 8347
rect 13136 8316 13246 8344
rect 13136 8304 13142 8316
rect 13234 8313 13246 8316
rect 13280 8313 13292 8347
rect 16482 8344 16488 8356
rect 16443 8316 16488 8344
rect 13234 8307 13292 8313
rect 16482 8304 16488 8316
rect 16540 8304 16546 8356
rect 18414 8344 18420 8356
rect 18375 8316 18420 8344
rect 18414 8304 18420 8316
rect 18472 8344 18478 8356
rect 19061 8347 19119 8353
rect 19061 8344 19073 8347
rect 18472 8316 19073 8344
rect 18472 8304 18478 8316
rect 19061 8313 19073 8316
rect 19107 8313 19119 8347
rect 19061 8307 19119 8313
rect 6825 8279 6883 8285
rect 6825 8245 6837 8279
rect 6871 8245 6883 8279
rect 11146 8276 11152 8288
rect 11107 8248 11152 8276
rect 6825 8239 6883 8245
rect 11146 8236 11152 8248
rect 11204 8236 11210 8288
rect 15657 8279 15715 8285
rect 15657 8245 15669 8279
rect 15703 8276 15715 8279
rect 15838 8276 15844 8288
rect 15703 8248 15844 8276
rect 15703 8245 15715 8248
rect 15657 8239 15715 8245
rect 15838 8236 15844 8248
rect 15896 8236 15902 8288
rect 18046 8276 18052 8288
rect 18007 8248 18052 8276
rect 18046 8236 18052 8248
rect 18104 8236 18110 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1857 8075 1915 8081
rect 1857 8041 1869 8075
rect 1903 8072 1915 8075
rect 2038 8072 2044 8084
rect 1903 8044 2044 8072
rect 1903 8041 1915 8044
rect 1857 8035 1915 8041
rect 2038 8032 2044 8044
rect 2096 8032 2102 8084
rect 2777 8075 2835 8081
rect 2777 8041 2789 8075
rect 2823 8072 2835 8075
rect 3142 8072 3148 8084
rect 2823 8044 3148 8072
rect 2823 8041 2835 8044
rect 2777 8035 2835 8041
rect 3142 8032 3148 8044
rect 3200 8032 3206 8084
rect 4433 8075 4491 8081
rect 4433 8041 4445 8075
rect 4479 8072 4491 8075
rect 4614 8072 4620 8084
rect 4479 8044 4620 8072
rect 4479 8041 4491 8044
rect 4433 8035 4491 8041
rect 4614 8032 4620 8044
rect 4672 8032 4678 8084
rect 7466 8072 7472 8084
rect 7427 8044 7472 8072
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 8113 8075 8171 8081
rect 8113 8041 8125 8075
rect 8159 8072 8171 8075
rect 8294 8072 8300 8084
rect 8159 8044 8300 8072
rect 8159 8041 8171 8044
rect 8113 8035 8171 8041
rect 8294 8032 8300 8044
rect 8352 8032 8358 8084
rect 9766 8032 9772 8084
rect 9824 8072 9830 8084
rect 10873 8075 10931 8081
rect 9824 8044 10824 8072
rect 9824 8032 9830 8044
rect 9122 7964 9128 8016
rect 9180 8004 9186 8016
rect 10796 8004 10824 8044
rect 10873 8041 10885 8075
rect 10919 8072 10931 8075
rect 11330 8072 11336 8084
rect 10919 8044 11336 8072
rect 10919 8041 10931 8044
rect 10873 8035 10931 8041
rect 11330 8032 11336 8044
rect 11388 8032 11394 8084
rect 11698 8072 11704 8084
rect 11659 8044 11704 8072
rect 11698 8032 11704 8044
rect 11756 8032 11762 8084
rect 12066 8072 12072 8084
rect 12027 8044 12072 8072
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 13170 8032 13176 8084
rect 13228 8072 13234 8084
rect 13265 8075 13323 8081
rect 13265 8072 13277 8075
rect 13228 8044 13277 8072
rect 13228 8032 13234 8044
rect 13265 8041 13277 8044
rect 13311 8041 13323 8075
rect 13265 8035 13323 8041
rect 13633 8075 13691 8081
rect 13633 8041 13645 8075
rect 13679 8072 13691 8075
rect 13722 8072 13728 8084
rect 13679 8044 13728 8072
rect 13679 8041 13691 8044
rect 13633 8035 13691 8041
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 16390 8072 16396 8084
rect 16351 8044 16396 8072
rect 16390 8032 16396 8044
rect 16448 8032 16454 8084
rect 16942 8032 16948 8084
rect 17000 8072 17006 8084
rect 17037 8075 17095 8081
rect 17037 8072 17049 8075
rect 17000 8044 17049 8072
rect 17000 8032 17006 8044
rect 17037 8041 17049 8044
rect 17083 8041 17095 8075
rect 17586 8072 17592 8084
rect 17547 8044 17592 8072
rect 17037 8035 17095 8041
rect 17586 8032 17592 8044
rect 17644 8032 17650 8084
rect 17770 8004 17776 8016
rect 9180 7976 10272 8004
rect 10796 7976 17776 8004
rect 9180 7964 9186 7976
rect 1765 7939 1823 7945
rect 1765 7905 1777 7939
rect 1811 7936 1823 7939
rect 2222 7936 2228 7948
rect 1811 7908 2228 7936
rect 1811 7905 1823 7908
rect 1765 7899 1823 7905
rect 2222 7896 2228 7908
rect 2280 7896 2286 7948
rect 2774 7896 2780 7948
rect 2832 7936 2838 7948
rect 3053 7939 3111 7945
rect 3053 7936 3065 7939
rect 2832 7908 3065 7936
rect 2832 7896 2838 7908
rect 3053 7905 3065 7908
rect 3099 7905 3111 7939
rect 3053 7899 3111 7905
rect 5169 7939 5227 7945
rect 5169 7905 5181 7939
rect 5215 7936 5227 7939
rect 5994 7936 6000 7948
rect 5215 7908 6000 7936
rect 5215 7905 5227 7908
rect 5169 7899 5227 7905
rect 5994 7896 6000 7908
rect 6052 7936 6058 7948
rect 6345 7939 6403 7945
rect 6345 7936 6357 7939
rect 6052 7908 6357 7936
rect 6052 7896 6058 7908
rect 6345 7905 6357 7908
rect 6391 7905 6403 7939
rect 6345 7899 6403 7905
rect 7558 7896 7564 7948
rect 7616 7936 7622 7948
rect 9214 7936 9220 7948
rect 7616 7908 9220 7936
rect 7616 7896 7622 7908
rect 9214 7896 9220 7908
rect 9272 7896 9278 7948
rect 9766 7896 9772 7948
rect 9824 7936 9830 7948
rect 10045 7939 10103 7945
rect 10045 7936 10057 7939
rect 9824 7908 10057 7936
rect 9824 7896 9830 7908
rect 10045 7905 10057 7908
rect 10091 7905 10103 7939
rect 10045 7899 10103 7905
rect 2038 7868 2044 7880
rect 1999 7840 2044 7868
rect 2038 7828 2044 7840
rect 2096 7828 2102 7880
rect 4338 7828 4344 7880
rect 4396 7868 4402 7880
rect 4522 7868 4528 7880
rect 4396 7840 4528 7868
rect 4396 7828 4402 7840
rect 4522 7828 4528 7840
rect 4580 7828 4586 7880
rect 4709 7871 4767 7877
rect 4709 7837 4721 7871
rect 4755 7868 4767 7871
rect 4798 7868 4804 7880
rect 4755 7840 4804 7868
rect 4755 7837 4767 7840
rect 4709 7831 4767 7837
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 6089 7871 6147 7877
rect 6089 7837 6101 7871
rect 6135 7837 6147 7871
rect 8570 7868 8576 7880
rect 8531 7840 8576 7868
rect 6089 7831 6147 7837
rect 1397 7735 1455 7741
rect 1397 7701 1409 7735
rect 1443 7732 1455 7735
rect 1578 7732 1584 7744
rect 1443 7704 1584 7732
rect 1443 7701 1455 7704
rect 1397 7695 1455 7701
rect 1578 7692 1584 7704
rect 1636 7692 1642 7744
rect 3510 7732 3516 7744
rect 3423 7704 3516 7732
rect 3510 7692 3516 7704
rect 3568 7732 3574 7744
rect 3789 7735 3847 7741
rect 3789 7732 3801 7735
rect 3568 7704 3801 7732
rect 3568 7692 3574 7704
rect 3789 7701 3801 7704
rect 3835 7701 3847 7735
rect 3789 7695 3847 7701
rect 3970 7692 3976 7744
rect 4028 7732 4034 7744
rect 4065 7735 4123 7741
rect 4065 7732 4077 7735
rect 4028 7704 4077 7732
rect 4028 7692 4034 7704
rect 4065 7701 4077 7704
rect 4111 7701 4123 7735
rect 5534 7732 5540 7744
rect 5495 7704 5540 7732
rect 4065 7695 4123 7701
rect 5534 7692 5540 7704
rect 5592 7692 5598 7744
rect 5905 7735 5963 7741
rect 5905 7701 5917 7735
rect 5951 7732 5963 7735
rect 5994 7732 6000 7744
rect 5951 7704 6000 7732
rect 5951 7701 5963 7704
rect 5905 7695 5963 7701
rect 5994 7692 6000 7704
rect 6052 7692 6058 7744
rect 6104 7732 6132 7831
rect 8570 7828 8576 7840
rect 8628 7828 8634 7880
rect 10134 7868 10140 7880
rect 10095 7840 10140 7868
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 10244 7877 10272 7976
rect 17770 7964 17776 7976
rect 17828 7964 17834 8016
rect 13262 7896 13268 7948
rect 13320 7936 13326 7948
rect 13725 7939 13783 7945
rect 13725 7936 13737 7939
rect 13320 7908 13737 7936
rect 13320 7896 13326 7908
rect 13725 7905 13737 7908
rect 13771 7905 13783 7939
rect 17954 7936 17960 7948
rect 17915 7908 17960 7936
rect 13725 7899 13783 7905
rect 17954 7896 17960 7908
rect 18012 7896 18018 7948
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 11146 7828 11152 7880
rect 11204 7868 11210 7880
rect 12161 7871 12219 7877
rect 12161 7868 12173 7871
rect 11204 7840 12173 7868
rect 11204 7828 11210 7840
rect 12161 7837 12173 7840
rect 12207 7837 12219 7871
rect 12161 7831 12219 7837
rect 12250 7828 12256 7880
rect 12308 7868 12314 7880
rect 13078 7868 13084 7880
rect 12308 7840 13084 7868
rect 12308 7828 12314 7840
rect 13078 7828 13084 7840
rect 13136 7868 13142 7880
rect 13906 7868 13912 7880
rect 13136 7840 13912 7868
rect 13136 7828 13142 7840
rect 13906 7828 13912 7840
rect 13964 7828 13970 7880
rect 15105 7871 15163 7877
rect 15105 7837 15117 7871
rect 15151 7868 15163 7871
rect 15654 7868 15660 7880
rect 15151 7840 15660 7868
rect 15151 7837 15163 7840
rect 15105 7831 15163 7837
rect 15654 7828 15660 7840
rect 15712 7868 15718 7880
rect 16485 7871 16543 7877
rect 16485 7868 16497 7871
rect 15712 7840 16497 7868
rect 15712 7828 15718 7840
rect 16485 7837 16497 7840
rect 16531 7837 16543 7871
rect 16485 7831 16543 7837
rect 16669 7871 16727 7877
rect 16669 7837 16681 7871
rect 16715 7868 16727 7871
rect 16758 7868 16764 7880
rect 16715 7840 16764 7868
rect 16715 7837 16727 7840
rect 16669 7831 16727 7837
rect 16758 7828 16764 7840
rect 16816 7828 16822 7880
rect 17862 7828 17868 7880
rect 17920 7868 17926 7880
rect 18049 7871 18107 7877
rect 18049 7868 18061 7871
rect 17920 7840 18061 7868
rect 17920 7828 17926 7840
rect 18049 7837 18061 7840
rect 18095 7837 18107 7871
rect 18049 7831 18107 7837
rect 18233 7871 18291 7877
rect 18233 7837 18245 7871
rect 18279 7868 18291 7871
rect 18598 7868 18604 7880
rect 18279 7840 18604 7868
rect 18279 7837 18291 7840
rect 18233 7831 18291 7837
rect 18598 7828 18604 7840
rect 18656 7868 18662 7880
rect 18969 7871 19027 7877
rect 18969 7868 18981 7871
rect 18656 7840 18981 7868
rect 18656 7828 18662 7840
rect 18969 7837 18981 7840
rect 19015 7837 19027 7871
rect 18969 7831 19027 7837
rect 8754 7760 8760 7812
rect 8812 7800 8818 7812
rect 9401 7803 9459 7809
rect 9401 7800 9413 7803
rect 8812 7772 9413 7800
rect 8812 7760 8818 7772
rect 9401 7769 9413 7772
rect 9447 7769 9459 7803
rect 9674 7800 9680 7812
rect 9587 7772 9680 7800
rect 9401 7763 9459 7769
rect 9674 7760 9680 7772
rect 9732 7800 9738 7812
rect 10962 7800 10968 7812
rect 9732 7772 10968 7800
rect 9732 7760 9738 7772
rect 10962 7760 10968 7772
rect 11020 7760 11026 7812
rect 14737 7803 14795 7809
rect 14737 7769 14749 7803
rect 14783 7800 14795 7803
rect 14783 7772 16068 7800
rect 14783 7769 14795 7772
rect 14737 7763 14795 7769
rect 6362 7732 6368 7744
rect 6104 7704 6368 7732
rect 6362 7692 6368 7704
rect 6420 7692 6426 7744
rect 8386 7732 8392 7744
rect 8347 7704 8392 7732
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 8478 7692 8484 7744
rect 8536 7732 8542 7744
rect 9033 7735 9091 7741
rect 9033 7732 9045 7735
rect 8536 7704 9045 7732
rect 8536 7692 8542 7704
rect 9033 7701 9045 7704
rect 9079 7701 9091 7735
rect 11238 7732 11244 7744
rect 11199 7704 11244 7732
rect 9033 7695 9091 7701
rect 11238 7692 11244 7704
rect 11296 7692 11302 7744
rect 11422 7692 11428 7744
rect 11480 7732 11486 7744
rect 11517 7735 11575 7741
rect 11517 7732 11529 7735
rect 11480 7704 11529 7732
rect 11480 7692 11486 7704
rect 11517 7701 11529 7704
rect 11563 7701 11575 7735
rect 11517 7695 11575 7701
rect 14182 7692 14188 7744
rect 14240 7732 14246 7744
rect 14277 7735 14335 7741
rect 14277 7732 14289 7735
rect 14240 7704 14289 7732
rect 14240 7692 14246 7704
rect 14277 7701 14289 7704
rect 14323 7701 14335 7735
rect 15746 7732 15752 7744
rect 15707 7704 15752 7732
rect 14277 7695 14335 7701
rect 15746 7692 15752 7704
rect 15804 7692 15810 7744
rect 16040 7741 16068 7772
rect 16390 7760 16396 7812
rect 16448 7800 16454 7812
rect 17405 7803 17463 7809
rect 17405 7800 17417 7803
rect 16448 7772 17417 7800
rect 16448 7760 16454 7772
rect 17405 7769 17417 7772
rect 17451 7800 17463 7803
rect 18322 7800 18328 7812
rect 17451 7772 18328 7800
rect 17451 7769 17463 7772
rect 17405 7763 17463 7769
rect 18322 7760 18328 7772
rect 18380 7760 18386 7812
rect 16025 7735 16083 7741
rect 16025 7701 16037 7735
rect 16071 7732 16083 7735
rect 16574 7732 16580 7744
rect 16071 7704 16580 7732
rect 16071 7701 16083 7704
rect 16025 7695 16083 7701
rect 16574 7692 16580 7704
rect 16632 7692 16638 7744
rect 18598 7732 18604 7744
rect 18559 7704 18604 7732
rect 18598 7692 18604 7704
rect 18656 7692 18662 7744
rect 19705 7735 19763 7741
rect 19705 7701 19717 7735
rect 19751 7732 19763 7735
rect 20070 7732 20076 7744
rect 19751 7704 20076 7732
rect 19751 7701 19763 7704
rect 19705 7695 19763 7701
rect 20070 7692 20076 7704
rect 20128 7692 20134 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 2130 7488 2136 7540
rect 2188 7528 2194 7540
rect 2409 7531 2467 7537
rect 2409 7528 2421 7531
rect 2188 7500 2421 7528
rect 2188 7488 2194 7500
rect 2409 7497 2421 7500
rect 2455 7528 2467 7531
rect 2593 7531 2651 7537
rect 2593 7528 2605 7531
rect 2455 7500 2605 7528
rect 2455 7497 2467 7500
rect 2409 7491 2467 7497
rect 2593 7497 2605 7500
rect 2639 7497 2651 7531
rect 2958 7528 2964 7540
rect 2919 7500 2964 7528
rect 2593 7491 2651 7497
rect 2958 7488 2964 7500
rect 3016 7488 3022 7540
rect 8205 7531 8263 7537
rect 5092 7500 8156 7528
rect 566 7420 572 7472
rect 624 7460 630 7472
rect 5092 7460 5120 7500
rect 624 7432 5120 7460
rect 5169 7463 5227 7469
rect 624 7420 630 7432
rect 5169 7429 5181 7463
rect 5215 7429 5227 7463
rect 5169 7423 5227 7429
rect 6641 7463 6699 7469
rect 6641 7429 6653 7463
rect 6687 7460 6699 7463
rect 8128 7460 8156 7500
rect 8205 7497 8217 7531
rect 8251 7528 8263 7531
rect 8570 7528 8576 7540
rect 8251 7500 8576 7528
rect 8251 7497 8263 7500
rect 8205 7491 8263 7497
rect 8570 7488 8576 7500
rect 8628 7488 8634 7540
rect 8662 7488 8668 7540
rect 8720 7528 8726 7540
rect 10781 7531 10839 7537
rect 8720 7500 8765 7528
rect 8720 7488 8726 7500
rect 10781 7497 10793 7531
rect 10827 7528 10839 7531
rect 11146 7528 11152 7540
rect 10827 7500 11152 7528
rect 10827 7497 10839 7500
rect 10781 7491 10839 7497
rect 11146 7488 11152 7500
rect 11204 7488 11210 7540
rect 11885 7531 11943 7537
rect 11885 7497 11897 7531
rect 11931 7528 11943 7531
rect 12250 7528 12256 7540
rect 11931 7500 12256 7528
rect 11931 7497 11943 7500
rect 11885 7491 11943 7497
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 13633 7531 13691 7537
rect 13633 7497 13645 7531
rect 13679 7528 13691 7531
rect 13722 7528 13728 7540
rect 13679 7500 13728 7528
rect 13679 7497 13691 7500
rect 13633 7491 13691 7497
rect 13722 7488 13728 7500
rect 13780 7488 13786 7540
rect 13906 7488 13912 7540
rect 13964 7528 13970 7540
rect 14645 7531 14703 7537
rect 14645 7528 14657 7531
rect 13964 7500 14657 7528
rect 13964 7488 13970 7500
rect 14645 7497 14657 7500
rect 14691 7497 14703 7531
rect 15470 7528 15476 7540
rect 15431 7500 15476 7528
rect 14645 7491 14703 7497
rect 15470 7488 15476 7500
rect 15528 7488 15534 7540
rect 15654 7528 15660 7540
rect 15615 7500 15660 7528
rect 15654 7488 15660 7500
rect 15712 7488 15718 7540
rect 8389 7463 8447 7469
rect 8389 7460 8401 7463
rect 6687 7432 7512 7460
rect 8128 7432 8401 7460
rect 6687 7429 6699 7432
rect 6641 7423 6699 7429
rect 1670 7352 1676 7404
rect 1728 7392 1734 7404
rect 1857 7395 1915 7401
rect 1857 7392 1869 7395
rect 1728 7364 1869 7392
rect 1728 7352 1734 7364
rect 1857 7361 1869 7364
rect 1903 7361 1915 7395
rect 2038 7392 2044 7404
rect 1951 7364 2044 7392
rect 1857 7355 1915 7361
rect 2038 7352 2044 7364
rect 2096 7392 2102 7404
rect 2498 7392 2504 7404
rect 2096 7364 2504 7392
rect 2096 7352 2102 7364
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 3418 7392 3424 7404
rect 3379 7364 3424 7392
rect 3418 7352 3424 7364
rect 3476 7352 3482 7404
rect 3602 7392 3608 7404
rect 3563 7364 3608 7392
rect 3602 7352 3608 7364
rect 3660 7352 3666 7404
rect 3329 7327 3387 7333
rect 3329 7293 3341 7327
rect 3375 7324 3387 7327
rect 3694 7324 3700 7336
rect 3375 7296 3700 7324
rect 3375 7293 3387 7296
rect 3329 7287 3387 7293
rect 3694 7284 3700 7296
rect 3752 7284 3758 7336
rect 5184 7324 5212 7423
rect 7484 7404 7512 7432
rect 8389 7429 8401 7432
rect 8435 7460 8447 7463
rect 8481 7463 8539 7469
rect 8481 7460 8493 7463
rect 8435 7432 8493 7460
rect 8435 7429 8447 7432
rect 8389 7423 8447 7429
rect 8481 7429 8493 7432
rect 8527 7429 8539 7463
rect 8481 7423 8539 7429
rect 9122 7420 9128 7472
rect 9180 7460 9186 7472
rect 10134 7460 10140 7472
rect 9180 7432 9352 7460
rect 10047 7432 10140 7460
rect 9180 7420 9186 7432
rect 5810 7392 5816 7404
rect 5771 7364 5816 7392
rect 5810 7352 5816 7364
rect 5868 7352 5874 7404
rect 6914 7352 6920 7404
rect 6972 7392 6978 7404
rect 7282 7392 7288 7404
rect 6972 7364 7288 7392
rect 6972 7352 6978 7364
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 7466 7392 7472 7404
rect 7427 7364 7472 7392
rect 7466 7352 7472 7364
rect 7524 7352 7530 7404
rect 9324 7401 9352 7432
rect 10134 7420 10140 7432
rect 10192 7460 10198 7472
rect 12342 7460 12348 7472
rect 10192 7432 12348 7460
rect 10192 7420 10198 7432
rect 12342 7420 12348 7432
rect 12400 7420 12406 7472
rect 15286 7420 15292 7472
rect 15344 7460 15350 7472
rect 15344 7432 18092 7460
rect 15344 7420 15350 7432
rect 9309 7395 9367 7401
rect 9309 7361 9321 7395
rect 9355 7361 9367 7395
rect 9766 7392 9772 7404
rect 9679 7364 9772 7392
rect 9309 7355 9367 7361
rect 9766 7352 9772 7364
rect 9824 7392 9830 7404
rect 10962 7392 10968 7404
rect 9824 7364 10968 7392
rect 9824 7352 9830 7364
rect 10962 7352 10968 7364
rect 11020 7352 11026 7404
rect 11330 7392 11336 7404
rect 11291 7364 11336 7392
rect 11330 7352 11336 7364
rect 11388 7352 11394 7404
rect 12434 7352 12440 7404
rect 12492 7392 12498 7404
rect 13170 7392 13176 7404
rect 12492 7364 12537 7392
rect 13083 7364 13176 7392
rect 12492 7352 12498 7364
rect 13170 7352 13176 7364
rect 13228 7392 13234 7404
rect 14090 7392 14096 7404
rect 13228 7364 14096 7392
rect 13228 7352 13234 7364
rect 14090 7352 14096 7364
rect 14148 7352 14154 7404
rect 14274 7392 14280 7404
rect 14235 7364 14280 7392
rect 14274 7352 14280 7364
rect 14332 7352 14338 7404
rect 14458 7352 14464 7404
rect 14516 7392 14522 7404
rect 15102 7392 15108 7404
rect 14516 7364 15108 7392
rect 14516 7352 14522 7364
rect 15102 7352 15108 7364
rect 15160 7352 15166 7404
rect 15197 7395 15255 7401
rect 15197 7361 15209 7395
rect 15243 7392 15255 7395
rect 15838 7392 15844 7404
rect 15243 7364 15844 7392
rect 15243 7361 15255 7364
rect 15197 7355 15255 7361
rect 15838 7352 15844 7364
rect 15896 7392 15902 7404
rect 16298 7392 16304 7404
rect 15896 7364 16304 7392
rect 15896 7352 15902 7364
rect 16298 7352 16304 7364
rect 16356 7352 16362 7404
rect 7193 7327 7251 7333
rect 7193 7324 7205 7327
rect 5184 7296 7205 7324
rect 7193 7293 7205 7296
rect 7239 7324 7251 7327
rect 8478 7324 8484 7336
rect 7239 7296 8484 7324
rect 7239 7293 7251 7296
rect 7193 7287 7251 7293
rect 8478 7284 8484 7296
rect 8536 7284 8542 7336
rect 8570 7284 8576 7336
rect 8628 7324 8634 7336
rect 9033 7327 9091 7333
rect 9033 7324 9045 7327
rect 8628 7296 9045 7324
rect 8628 7284 8634 7296
rect 9033 7293 9045 7296
rect 9079 7293 9091 7327
rect 9033 7287 9091 7293
rect 10870 7284 10876 7336
rect 10928 7324 10934 7336
rect 11241 7327 11299 7333
rect 11241 7324 11253 7327
rect 10928 7296 11253 7324
rect 10928 7284 10934 7296
rect 11241 7293 11253 7296
rect 11287 7293 11299 7327
rect 11241 7287 11299 7293
rect 15470 7284 15476 7336
rect 15528 7324 15534 7336
rect 16025 7327 16083 7333
rect 16025 7324 16037 7327
rect 15528 7296 16037 7324
rect 15528 7284 15534 7296
rect 16025 7293 16037 7296
rect 16071 7324 16083 7327
rect 17589 7327 17647 7333
rect 17589 7324 17601 7327
rect 16071 7296 17601 7324
rect 16071 7293 16083 7296
rect 16025 7287 16083 7293
rect 17589 7293 17601 7296
rect 17635 7324 17647 7327
rect 17954 7324 17960 7336
rect 17635 7296 17960 7324
rect 17635 7293 17647 7296
rect 17589 7287 17647 7293
rect 17954 7284 17960 7296
rect 18012 7284 18018 7336
rect 18064 7324 18092 7432
rect 18322 7420 18328 7472
rect 18380 7460 18386 7472
rect 19613 7463 19671 7469
rect 18380 7432 18644 7460
rect 18380 7420 18386 7432
rect 18506 7392 18512 7404
rect 18419 7364 18512 7392
rect 18506 7352 18512 7364
rect 18564 7352 18570 7404
rect 18616 7401 18644 7432
rect 19613 7429 19625 7463
rect 19659 7460 19671 7463
rect 20530 7460 20536 7472
rect 19659 7432 20536 7460
rect 19659 7429 19671 7432
rect 19613 7423 19671 7429
rect 20530 7420 20536 7432
rect 20588 7420 20594 7472
rect 18601 7395 18659 7401
rect 18601 7361 18613 7395
rect 18647 7392 18659 7395
rect 18782 7392 18788 7404
rect 18647 7364 18788 7392
rect 18647 7361 18659 7364
rect 18601 7355 18659 7361
rect 18782 7352 18788 7364
rect 18840 7352 18846 7404
rect 19334 7352 19340 7404
rect 19392 7392 19398 7404
rect 19521 7395 19579 7401
rect 19521 7392 19533 7395
rect 19392 7364 19533 7392
rect 19392 7352 19398 7364
rect 19521 7361 19533 7364
rect 19567 7392 19579 7395
rect 20165 7395 20223 7401
rect 20165 7392 20177 7395
rect 19567 7364 20177 7392
rect 19567 7361 19579 7364
rect 19521 7355 19579 7361
rect 20165 7361 20177 7364
rect 20211 7361 20223 7395
rect 20165 7355 20223 7361
rect 18414 7324 18420 7336
rect 18064 7296 18420 7324
rect 18414 7284 18420 7296
rect 18472 7284 18478 7336
rect 18524 7324 18552 7352
rect 19061 7327 19119 7333
rect 19061 7324 19073 7327
rect 18524 7296 19073 7324
rect 19061 7293 19073 7296
rect 19107 7293 19119 7327
rect 19061 7287 19119 7293
rect 1762 7256 1768 7268
rect 1675 7228 1768 7256
rect 1762 7216 1768 7228
rect 1820 7256 1826 7268
rect 2777 7259 2835 7265
rect 2777 7256 2789 7259
rect 1820 7228 2789 7256
rect 1820 7216 1826 7228
rect 2777 7225 2789 7228
rect 2823 7225 2835 7259
rect 2777 7219 2835 7225
rect 5077 7259 5135 7265
rect 5077 7225 5089 7259
rect 5123 7256 5135 7259
rect 5123 7228 5580 7256
rect 5123 7225 5135 7228
rect 5077 7219 5135 7225
rect 5552 7200 5580 7228
rect 5626 7216 5632 7268
rect 5684 7256 5690 7268
rect 6086 7256 6092 7268
rect 5684 7228 6092 7256
rect 5684 7216 5690 7228
rect 6086 7216 6092 7228
rect 6144 7216 6150 7268
rect 8389 7259 8447 7265
rect 8389 7225 8401 7259
rect 8435 7256 8447 7259
rect 9125 7259 9183 7265
rect 9125 7256 9137 7259
rect 8435 7228 9137 7256
rect 8435 7225 8447 7228
rect 8389 7219 8447 7225
rect 9125 7225 9137 7228
rect 9171 7256 9183 7259
rect 9582 7256 9588 7268
rect 9171 7228 9588 7256
rect 9171 7225 9183 7228
rect 9125 7219 9183 7225
rect 9582 7216 9588 7228
rect 9640 7216 9646 7268
rect 11054 7216 11060 7268
rect 11112 7256 11118 7268
rect 12161 7259 12219 7265
rect 12161 7256 12173 7259
rect 11112 7228 12173 7256
rect 11112 7216 11118 7228
rect 12161 7225 12173 7228
rect 12207 7225 12219 7259
rect 12161 7219 12219 7225
rect 13541 7259 13599 7265
rect 13541 7225 13553 7259
rect 13587 7256 13599 7259
rect 13998 7256 14004 7268
rect 13587 7228 14004 7256
rect 13587 7225 13599 7228
rect 13541 7219 13599 7225
rect 13998 7216 14004 7228
rect 14056 7256 14062 7268
rect 14458 7256 14464 7268
rect 14056 7228 14464 7256
rect 14056 7216 14062 7228
rect 14458 7216 14464 7228
rect 14516 7216 14522 7268
rect 17221 7259 17279 7265
rect 17221 7256 17233 7259
rect 16132 7228 17233 7256
rect 1394 7188 1400 7200
rect 1355 7160 1400 7188
rect 1394 7148 1400 7160
rect 1452 7148 1458 7200
rect 2593 7191 2651 7197
rect 2593 7157 2605 7191
rect 2639 7188 2651 7191
rect 2866 7188 2872 7200
rect 2639 7160 2872 7188
rect 2639 7157 2651 7160
rect 2593 7151 2651 7157
rect 2866 7148 2872 7160
rect 2924 7148 2930 7200
rect 4065 7191 4123 7197
rect 4065 7157 4077 7191
rect 4111 7188 4123 7191
rect 4433 7191 4491 7197
rect 4433 7188 4445 7191
rect 4111 7160 4445 7188
rect 4111 7157 4123 7160
rect 4065 7151 4123 7157
rect 4433 7157 4445 7160
rect 4479 7188 4491 7191
rect 4798 7188 4804 7200
rect 4479 7160 4804 7188
rect 4479 7157 4491 7160
rect 4433 7151 4491 7157
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 5534 7188 5540 7200
rect 5495 7160 5540 7188
rect 5534 7148 5540 7160
rect 5592 7148 5598 7200
rect 5994 7148 6000 7200
rect 6052 7188 6058 7200
rect 6181 7191 6239 7197
rect 6181 7188 6193 7191
rect 6052 7160 6193 7188
rect 6052 7148 6058 7160
rect 6181 7157 6193 7160
rect 6227 7188 6239 7191
rect 6362 7188 6368 7200
rect 6227 7160 6368 7188
rect 6227 7157 6239 7160
rect 6181 7151 6239 7157
rect 6362 7148 6368 7160
rect 6420 7148 6426 7200
rect 6822 7188 6828 7200
rect 6783 7160 6828 7188
rect 6822 7148 6828 7160
rect 6880 7148 6886 7200
rect 9858 7148 9864 7200
rect 9916 7188 9922 7200
rect 10597 7191 10655 7197
rect 10597 7188 10609 7191
rect 9916 7160 10609 7188
rect 9916 7148 9922 7160
rect 10597 7157 10609 7160
rect 10643 7188 10655 7191
rect 11149 7191 11207 7197
rect 11149 7188 11161 7191
rect 10643 7160 11161 7188
rect 10643 7157 10655 7160
rect 10597 7151 10655 7157
rect 11149 7157 11161 7160
rect 11195 7188 11207 7191
rect 11330 7188 11336 7200
rect 11195 7160 11336 7188
rect 11195 7157 11207 7160
rect 11149 7151 11207 7157
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 14090 7148 14096 7200
rect 14148 7188 14154 7200
rect 14366 7188 14372 7200
rect 14148 7160 14372 7188
rect 14148 7148 14154 7160
rect 14366 7148 14372 7160
rect 14424 7148 14430 7200
rect 15746 7148 15752 7200
rect 15804 7188 15810 7200
rect 16132 7197 16160 7228
rect 17221 7225 17233 7228
rect 17267 7256 17279 7259
rect 17862 7256 17868 7268
rect 17267 7228 17868 7256
rect 17267 7225 17279 7228
rect 17221 7219 17279 7225
rect 17862 7216 17868 7228
rect 17920 7216 17926 7268
rect 18506 7256 18512 7268
rect 18064 7228 18512 7256
rect 16117 7191 16175 7197
rect 16117 7188 16129 7191
rect 15804 7160 16129 7188
rect 15804 7148 15810 7160
rect 16117 7157 16129 7160
rect 16163 7157 16175 7191
rect 16758 7188 16764 7200
rect 16719 7160 16764 7188
rect 16117 7151 16175 7157
rect 16758 7148 16764 7160
rect 16816 7148 16822 7200
rect 18064 7197 18092 7228
rect 18506 7216 18512 7228
rect 18564 7216 18570 7268
rect 18049 7191 18107 7197
rect 18049 7157 18061 7191
rect 18095 7157 18107 7191
rect 19978 7188 19984 7200
rect 19939 7160 19984 7188
rect 18049 7151 18107 7157
rect 19978 7148 19984 7160
rect 20036 7148 20042 7200
rect 20070 7148 20076 7200
rect 20128 7188 20134 7200
rect 20622 7188 20628 7200
rect 20128 7160 20628 7188
rect 20128 7148 20134 7160
rect 20622 7148 20628 7160
rect 20680 7148 20686 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1397 6987 1455 6993
rect 1397 6953 1409 6987
rect 1443 6984 1455 6987
rect 1762 6984 1768 6996
rect 1443 6956 1768 6984
rect 1443 6953 1455 6956
rect 1397 6947 1455 6953
rect 1762 6944 1768 6956
rect 1820 6944 1826 6996
rect 3513 6987 3571 6993
rect 3513 6953 3525 6987
rect 3559 6984 3571 6987
rect 3602 6984 3608 6996
rect 3559 6956 3608 6984
rect 3559 6953 3571 6956
rect 3513 6947 3571 6953
rect 3602 6944 3608 6956
rect 3660 6944 3666 6996
rect 7374 6944 7380 6996
rect 7432 6984 7438 6996
rect 8662 6984 8668 6996
rect 7432 6956 8668 6984
rect 7432 6944 7438 6956
rect 8662 6944 8668 6956
rect 8720 6944 8726 6996
rect 9033 6987 9091 6993
rect 9033 6953 9045 6987
rect 9079 6984 9091 6987
rect 9122 6984 9128 6996
rect 9079 6956 9128 6984
rect 9079 6953 9091 6956
rect 9033 6947 9091 6953
rect 9122 6944 9128 6956
rect 9180 6984 9186 6996
rect 9401 6987 9459 6993
rect 9401 6984 9413 6987
rect 9180 6956 9413 6984
rect 9180 6944 9186 6956
rect 9401 6953 9413 6956
rect 9447 6953 9459 6987
rect 9674 6984 9680 6996
rect 9635 6956 9680 6984
rect 9401 6947 9459 6953
rect 9674 6944 9680 6956
rect 9732 6944 9738 6996
rect 10045 6987 10103 6993
rect 10045 6953 10057 6987
rect 10091 6984 10103 6987
rect 10778 6984 10784 6996
rect 10091 6956 10784 6984
rect 10091 6953 10103 6956
rect 10045 6947 10103 6953
rect 1670 6876 1676 6928
rect 1728 6916 1734 6928
rect 1857 6919 1915 6925
rect 1857 6916 1869 6919
rect 1728 6888 1869 6916
rect 1728 6876 1734 6888
rect 1857 6885 1869 6888
rect 1903 6885 1915 6919
rect 1857 6879 1915 6885
rect 2869 6919 2927 6925
rect 2869 6885 2881 6919
rect 2915 6916 2927 6919
rect 3970 6916 3976 6928
rect 2915 6888 3976 6916
rect 2915 6885 2927 6888
rect 2869 6879 2927 6885
rect 3970 6876 3976 6888
rect 4028 6876 4034 6928
rect 5810 6876 5816 6928
rect 5868 6916 5874 6928
rect 10060 6916 10088 6947
rect 10778 6944 10784 6956
rect 10836 6944 10842 6996
rect 13909 6987 13967 6993
rect 13909 6953 13921 6987
rect 13955 6984 13967 6987
rect 14274 6984 14280 6996
rect 13955 6956 14280 6984
rect 13955 6953 13967 6956
rect 13909 6947 13967 6953
rect 14274 6944 14280 6956
rect 14332 6944 14338 6996
rect 16758 6944 16764 6996
rect 16816 6984 16822 6996
rect 17773 6987 17831 6993
rect 17773 6984 17785 6987
rect 16816 6956 17785 6984
rect 16816 6944 16822 6956
rect 17773 6953 17785 6956
rect 17819 6953 17831 6987
rect 18414 6984 18420 6996
rect 18375 6956 18420 6984
rect 17773 6947 17831 6953
rect 18414 6944 18420 6956
rect 18472 6944 18478 6996
rect 19242 6984 19248 6996
rect 19203 6956 19248 6984
rect 19242 6944 19248 6956
rect 19300 6944 19306 6996
rect 5868 6888 6868 6916
rect 5868 6876 5874 6888
rect 2777 6851 2835 6857
rect 2777 6817 2789 6851
rect 2823 6848 2835 6851
rect 4062 6848 4068 6860
rect 2823 6820 4068 6848
rect 2823 6817 2835 6820
rect 2777 6811 2835 6817
rect 4062 6808 4068 6820
rect 4120 6808 4126 6860
rect 4433 6851 4491 6857
rect 4433 6817 4445 6851
rect 4479 6848 4491 6851
rect 4614 6848 4620 6860
rect 4479 6820 4620 6848
rect 4479 6817 4491 6820
rect 4433 6811 4491 6817
rect 4614 6808 4620 6820
rect 4672 6808 4678 6860
rect 6253 6851 6311 6857
rect 6253 6848 6265 6851
rect 5920 6820 6265 6848
rect 3050 6780 3056 6792
rect 2963 6752 3056 6780
rect 3050 6740 3056 6752
rect 3108 6780 3114 6792
rect 3510 6780 3516 6792
rect 3108 6752 3516 6780
rect 3108 6740 3114 6752
rect 3510 6740 3516 6752
rect 3568 6740 3574 6792
rect 4246 6740 4252 6792
rect 4304 6780 4310 6792
rect 4525 6783 4583 6789
rect 4525 6780 4537 6783
rect 4304 6752 4537 6780
rect 4304 6740 4310 6752
rect 4525 6749 4537 6752
rect 4571 6749 4583 6783
rect 4525 6743 4583 6749
rect 4709 6783 4767 6789
rect 4709 6749 4721 6783
rect 4755 6780 4767 6783
rect 4798 6780 4804 6792
rect 4755 6752 4804 6780
rect 4755 6749 4767 6752
rect 4709 6743 4767 6749
rect 2498 6672 2504 6724
rect 2556 6712 2562 6724
rect 3881 6715 3939 6721
rect 3881 6712 3893 6715
rect 2556 6684 3893 6712
rect 2556 6672 2562 6684
rect 3881 6681 3893 6684
rect 3927 6712 3939 6715
rect 4724 6712 4752 6743
rect 4798 6740 4804 6752
rect 4856 6740 4862 6792
rect 5718 6712 5724 6724
rect 3927 6684 4752 6712
rect 5184 6684 5724 6712
rect 3927 6681 3939 6684
rect 3881 6675 3939 6681
rect 5184 6656 5212 6684
rect 5718 6672 5724 6684
rect 5776 6672 5782 6724
rect 2222 6644 2228 6656
rect 2183 6616 2228 6644
rect 2222 6604 2228 6616
rect 2280 6604 2286 6656
rect 2409 6647 2467 6653
rect 2409 6613 2421 6647
rect 2455 6644 2467 6647
rect 2682 6644 2688 6656
rect 2455 6616 2688 6644
rect 2455 6613 2467 6616
rect 2409 6607 2467 6613
rect 2682 6604 2688 6616
rect 2740 6604 2746 6656
rect 4062 6644 4068 6656
rect 4023 6616 4068 6644
rect 4062 6604 4068 6616
rect 4120 6604 4126 6656
rect 5166 6644 5172 6656
rect 5127 6616 5172 6644
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 5629 6647 5687 6653
rect 5629 6613 5641 6647
rect 5675 6644 5687 6647
rect 5920 6644 5948 6820
rect 6253 6817 6265 6820
rect 6299 6817 6311 6851
rect 6840 6848 6868 6888
rect 9600 6888 10088 6916
rect 13173 6919 13231 6925
rect 7374 6848 7380 6860
rect 6840 6820 7380 6848
rect 6253 6811 6311 6817
rect 7374 6808 7380 6820
rect 7432 6808 7438 6860
rect 8478 6848 8484 6860
rect 8439 6820 8484 6848
rect 8478 6808 8484 6820
rect 8536 6808 8542 6860
rect 9398 6808 9404 6860
rect 9456 6848 9462 6860
rect 9600 6848 9628 6888
rect 13173 6885 13185 6919
rect 13219 6916 13231 6919
rect 13219 6888 13860 6916
rect 13219 6885 13231 6888
rect 13173 6879 13231 6885
rect 11606 6848 11612 6860
rect 9456 6820 9628 6848
rect 11567 6820 11612 6848
rect 9456 6808 9462 6820
rect 11606 6808 11612 6820
rect 11664 6848 11670 6860
rect 13832 6848 13860 6888
rect 16298 6876 16304 6928
rect 16356 6916 16362 6928
rect 16356 6888 16620 6916
rect 16356 6876 16362 6888
rect 14274 6848 14280 6860
rect 11664 6820 13584 6848
rect 13832 6820 14280 6848
rect 11664 6808 11670 6820
rect 5994 6740 6000 6792
rect 6052 6780 6058 6792
rect 6052 6752 6097 6780
rect 6052 6740 6058 6752
rect 9030 6740 9036 6792
rect 9088 6780 9094 6792
rect 10042 6780 10048 6792
rect 9088 6752 10048 6780
rect 9088 6740 9094 6752
rect 10042 6740 10048 6752
rect 10100 6780 10106 6792
rect 10137 6783 10195 6789
rect 10137 6780 10149 6783
rect 10100 6752 10149 6780
rect 10100 6740 10106 6752
rect 10137 6749 10149 6752
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 10226 6740 10232 6792
rect 10284 6780 10290 6792
rect 10284 6752 10329 6780
rect 10284 6740 10290 6752
rect 10778 6740 10784 6792
rect 10836 6780 10842 6792
rect 11422 6780 11428 6792
rect 10836 6752 11428 6780
rect 10836 6740 10842 6752
rect 11422 6740 11428 6752
rect 11480 6780 11486 6792
rect 11701 6783 11759 6789
rect 11701 6780 11713 6783
rect 11480 6752 11713 6780
rect 11480 6740 11486 6752
rect 11701 6749 11713 6752
rect 11747 6749 11759 6783
rect 11882 6780 11888 6792
rect 11843 6752 11888 6780
rect 11701 6743 11759 6749
rect 11882 6740 11888 6752
rect 11940 6740 11946 6792
rect 13262 6780 13268 6792
rect 13223 6752 13268 6780
rect 13262 6740 13268 6752
rect 13320 6740 13326 6792
rect 13446 6780 13452 6792
rect 13407 6752 13452 6780
rect 13446 6740 13452 6752
rect 13504 6740 13510 6792
rect 13556 6780 13584 6820
rect 14274 6808 14280 6820
rect 14332 6808 14338 6860
rect 15381 6851 15439 6857
rect 15381 6817 15393 6851
rect 15427 6848 15439 6851
rect 16482 6848 16488 6860
rect 15427 6820 16488 6848
rect 15427 6817 15439 6820
rect 15381 6811 15439 6817
rect 16482 6808 16488 6820
rect 16540 6808 16546 6860
rect 16592 6848 16620 6888
rect 16666 6857 16672 6860
rect 16660 6848 16672 6857
rect 16592 6820 16672 6848
rect 16660 6811 16672 6820
rect 16666 6808 16672 6811
rect 16724 6808 16730 6860
rect 14553 6783 14611 6789
rect 14553 6780 14565 6783
rect 13556 6752 14565 6780
rect 14553 6749 14565 6752
rect 14599 6749 14611 6783
rect 14553 6743 14611 6749
rect 16022 6740 16028 6792
rect 16080 6780 16086 6792
rect 16393 6783 16451 6789
rect 16393 6780 16405 6783
rect 16080 6752 16405 6780
rect 16080 6740 16086 6752
rect 16393 6749 16405 6752
rect 16439 6749 16451 6783
rect 19334 6780 19340 6792
rect 19295 6752 19340 6780
rect 16393 6743 16451 6749
rect 19334 6740 19340 6752
rect 19392 6740 19398 6792
rect 19426 6740 19432 6792
rect 19484 6780 19490 6792
rect 19484 6752 19529 6780
rect 19484 6740 19490 6752
rect 12802 6712 12808 6724
rect 12763 6684 12808 6712
rect 12802 6672 12808 6684
rect 12860 6672 12866 6724
rect 18877 6715 18935 6721
rect 18877 6681 18889 6715
rect 18923 6712 18935 6715
rect 20533 6715 20591 6721
rect 20533 6712 20545 6715
rect 18923 6684 20545 6712
rect 18923 6681 18935 6684
rect 18877 6675 18935 6681
rect 20533 6681 20545 6684
rect 20579 6712 20591 6715
rect 20990 6712 20996 6724
rect 20579 6684 20996 6712
rect 20579 6681 20591 6684
rect 20533 6675 20591 6681
rect 20990 6672 20996 6684
rect 21048 6672 21054 6724
rect 5994 6644 6000 6656
rect 5675 6616 6000 6644
rect 5675 6613 5687 6616
rect 5629 6607 5687 6613
rect 5994 6604 6000 6616
rect 6052 6604 6058 6656
rect 7374 6644 7380 6656
rect 7335 6616 7380 6644
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 7926 6644 7932 6656
rect 7887 6616 7932 6644
rect 7926 6604 7932 6616
rect 7984 6604 7990 6656
rect 8294 6644 8300 6656
rect 8255 6616 8300 6644
rect 8294 6604 8300 6616
rect 8352 6604 8358 6656
rect 9766 6604 9772 6656
rect 9824 6644 9830 6656
rect 10781 6647 10839 6653
rect 10781 6644 10793 6647
rect 9824 6616 10793 6644
rect 9824 6604 9830 6616
rect 10781 6613 10793 6616
rect 10827 6644 10839 6647
rect 10870 6644 10876 6656
rect 10827 6616 10876 6644
rect 10827 6613 10839 6616
rect 10781 6607 10839 6613
rect 10870 6604 10876 6616
rect 10928 6604 10934 6656
rect 11238 6644 11244 6656
rect 11199 6616 11244 6644
rect 11238 6604 11244 6616
rect 11296 6604 11302 6656
rect 12526 6644 12532 6656
rect 12487 6616 12532 6644
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 14274 6644 14280 6656
rect 14235 6616 14280 6644
rect 14274 6604 14280 6616
rect 14332 6604 14338 6656
rect 14734 6604 14740 6656
rect 14792 6644 14798 6656
rect 15013 6647 15071 6653
rect 15013 6644 15025 6647
rect 14792 6616 15025 6644
rect 14792 6604 14798 6616
rect 15013 6613 15025 6616
rect 15059 6613 15071 6647
rect 16206 6644 16212 6656
rect 16167 6616 16212 6644
rect 15013 6607 15071 6613
rect 16206 6604 16212 6616
rect 16264 6604 16270 6656
rect 18690 6644 18696 6656
rect 18651 6616 18696 6644
rect 18690 6604 18696 6616
rect 18748 6604 18754 6656
rect 19978 6644 19984 6656
rect 19939 6616 19984 6644
rect 19978 6604 19984 6616
rect 20036 6604 20042 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 4982 6440 4988 6452
rect 4943 6412 4988 6440
rect 4982 6400 4988 6412
rect 5040 6400 5046 6452
rect 5169 6443 5227 6449
rect 5169 6409 5181 6443
rect 5215 6440 5227 6443
rect 5442 6440 5448 6452
rect 5215 6412 5448 6440
rect 5215 6409 5227 6412
rect 5169 6403 5227 6409
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 6822 6440 6828 6452
rect 6783 6412 6828 6440
rect 6822 6400 6828 6412
rect 6880 6400 6886 6452
rect 8297 6443 8355 6449
rect 8297 6409 8309 6443
rect 8343 6440 8355 6443
rect 8386 6440 8392 6452
rect 8343 6412 8392 6440
rect 8343 6409 8355 6412
rect 8297 6403 8355 6409
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 9030 6440 9036 6452
rect 8991 6412 9036 6440
rect 9030 6400 9036 6412
rect 9088 6400 9094 6452
rect 9398 6440 9404 6452
rect 9359 6412 9404 6440
rect 9398 6400 9404 6412
rect 9456 6400 9462 6452
rect 10226 6400 10232 6452
rect 10284 6440 10290 6452
rect 11425 6443 11483 6449
rect 11425 6440 11437 6443
rect 10284 6412 11437 6440
rect 10284 6400 10290 6412
rect 11425 6409 11437 6412
rect 11471 6409 11483 6443
rect 11882 6440 11888 6452
rect 11843 6412 11888 6440
rect 11425 6403 11483 6409
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 14185 6443 14243 6449
rect 14185 6409 14197 6443
rect 14231 6440 14243 6443
rect 16022 6440 16028 6452
rect 14231 6412 16028 6440
rect 14231 6409 14243 6412
rect 14185 6403 14243 6409
rect 6086 6332 6092 6384
rect 6144 6372 6150 6384
rect 8573 6375 8631 6381
rect 8573 6372 8585 6375
rect 6144 6344 8585 6372
rect 6144 6332 6150 6344
rect 8573 6341 8585 6344
rect 8619 6372 8631 6375
rect 9122 6372 9128 6384
rect 8619 6344 9128 6372
rect 8619 6341 8631 6344
rect 8573 6335 8631 6341
rect 9122 6332 9128 6344
rect 9180 6372 9186 6384
rect 9180 6344 9536 6372
rect 9180 6332 9186 6344
rect 4154 6264 4160 6316
rect 4212 6304 4218 6316
rect 5166 6304 5172 6316
rect 4212 6276 5172 6304
rect 4212 6264 4218 6276
rect 5166 6264 5172 6276
rect 5224 6304 5230 6316
rect 5629 6307 5687 6313
rect 5629 6304 5641 6307
rect 5224 6276 5641 6304
rect 5224 6264 5230 6276
rect 5629 6273 5641 6276
rect 5675 6273 5687 6307
rect 5629 6267 5687 6273
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6304 5871 6307
rect 5994 6304 6000 6316
rect 5859 6276 6000 6304
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 5994 6264 6000 6276
rect 6052 6304 6058 6316
rect 6454 6304 6460 6316
rect 6052 6276 6460 6304
rect 6052 6264 6058 6276
rect 6454 6264 6460 6276
rect 6512 6264 6518 6316
rect 7374 6264 7380 6316
rect 7432 6304 7438 6316
rect 9508 6313 9536 6344
rect 7469 6307 7527 6313
rect 7469 6304 7481 6307
rect 7432 6276 7481 6304
rect 7432 6264 7438 6276
rect 7469 6273 7481 6276
rect 7515 6304 7527 6307
rect 7837 6307 7895 6313
rect 7837 6304 7849 6307
rect 7515 6276 7849 6304
rect 7515 6273 7527 6276
rect 7469 6267 7527 6273
rect 7837 6273 7849 6276
rect 7883 6273 7895 6307
rect 7837 6267 7895 6273
rect 9493 6307 9551 6313
rect 9493 6273 9505 6307
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 12526 6264 12532 6316
rect 12584 6304 12590 6316
rect 12989 6307 13047 6313
rect 12989 6304 13001 6307
rect 12584 6276 13001 6304
rect 12584 6264 12590 6276
rect 12989 6273 13001 6276
rect 13035 6273 13047 6307
rect 12989 6267 13047 6273
rect 13814 6264 13820 6316
rect 13872 6304 13878 6316
rect 14292 6313 14320 6412
rect 16022 6400 16028 6412
rect 16080 6440 16086 6452
rect 16393 6443 16451 6449
rect 16393 6440 16405 6443
rect 16080 6412 16405 6440
rect 16080 6400 16086 6412
rect 16393 6409 16405 6412
rect 16439 6440 16451 6443
rect 16482 6440 16488 6452
rect 16439 6412 16488 6440
rect 16439 6409 16451 6412
rect 16393 6403 16451 6409
rect 16482 6400 16488 6412
rect 16540 6440 16546 6452
rect 17773 6443 17831 6449
rect 17773 6440 17785 6443
rect 16540 6412 17785 6440
rect 16540 6400 16546 6412
rect 17773 6409 17785 6412
rect 17819 6409 17831 6443
rect 17773 6403 17831 6409
rect 14277 6307 14335 6313
rect 14277 6304 14289 6307
rect 13872 6276 14289 6304
rect 13872 6264 13878 6276
rect 14277 6273 14289 6276
rect 14323 6273 14335 6307
rect 17788 6304 17816 6403
rect 19978 6400 19984 6452
rect 20036 6440 20042 6452
rect 20533 6443 20591 6449
rect 20533 6440 20545 6443
rect 20036 6412 20545 6440
rect 20036 6400 20042 6412
rect 20533 6409 20545 6412
rect 20579 6409 20591 6443
rect 20533 6403 20591 6409
rect 19426 6372 19432 6384
rect 19387 6344 19432 6372
rect 19426 6332 19432 6344
rect 19484 6372 19490 6384
rect 20349 6375 20407 6381
rect 20349 6372 20361 6375
rect 19484 6344 20361 6372
rect 19484 6332 19490 6344
rect 20349 6341 20361 6344
rect 20395 6341 20407 6375
rect 20349 6335 20407 6341
rect 18049 6307 18107 6313
rect 18049 6304 18061 6307
rect 17788 6276 18061 6304
rect 14277 6267 14335 6273
rect 18049 6273 18061 6276
rect 18095 6273 18107 6307
rect 20990 6304 20996 6316
rect 20951 6276 20996 6304
rect 18049 6267 18107 6273
rect 20990 6264 20996 6276
rect 21048 6264 21054 6316
rect 21177 6307 21235 6313
rect 21177 6273 21189 6307
rect 21223 6304 21235 6307
rect 21450 6304 21456 6316
rect 21223 6276 21456 6304
rect 21223 6273 21235 6276
rect 21177 6267 21235 6273
rect 21450 6264 21456 6276
rect 21508 6264 21514 6316
rect 2225 6239 2283 6245
rect 2225 6205 2237 6239
rect 2271 6236 2283 6239
rect 2492 6239 2550 6245
rect 2271 6208 2305 6236
rect 2271 6205 2283 6208
rect 2225 6199 2283 6205
rect 2492 6205 2504 6239
rect 2538 6236 2550 6239
rect 3050 6236 3056 6248
rect 2538 6208 3056 6236
rect 2538 6205 2550 6208
rect 2492 6199 2550 6205
rect 2133 6171 2191 6177
rect 2133 6137 2145 6171
rect 2179 6168 2191 6171
rect 2240 6168 2268 6199
rect 3050 6196 3056 6208
rect 3108 6196 3114 6248
rect 4982 6196 4988 6248
rect 5040 6236 5046 6248
rect 5537 6239 5595 6245
rect 5537 6236 5549 6239
rect 5040 6208 5549 6236
rect 5040 6196 5046 6208
rect 5537 6205 5549 6208
rect 5583 6205 5595 6239
rect 5537 6199 5595 6205
rect 7098 6196 7104 6248
rect 7156 6236 7162 6248
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 7156 6208 7297 6236
rect 7156 6196 7162 6208
rect 7285 6205 7297 6208
rect 7331 6236 7343 6239
rect 7926 6236 7932 6248
rect 7331 6208 7932 6236
rect 7331 6205 7343 6208
rect 7285 6199 7343 6205
rect 7926 6196 7932 6208
rect 7984 6196 7990 6248
rect 16850 6236 16856 6248
rect 16811 6208 16856 6236
rect 16850 6196 16856 6208
rect 16908 6236 16914 6248
rect 17405 6239 17463 6245
rect 17405 6236 17417 6239
rect 16908 6208 17417 6236
rect 16908 6196 16914 6208
rect 17405 6205 17417 6208
rect 17451 6205 17463 6239
rect 17405 6199 17463 6205
rect 18138 6196 18144 6248
rect 18196 6236 18202 6248
rect 18316 6239 18374 6245
rect 18316 6236 18328 6239
rect 18196 6208 18328 6236
rect 18196 6196 18202 6208
rect 18316 6205 18328 6208
rect 18362 6236 18374 6239
rect 18690 6236 18696 6248
rect 18362 6208 18696 6236
rect 18362 6205 18374 6208
rect 18316 6199 18374 6205
rect 18690 6196 18696 6208
rect 18748 6196 18754 6248
rect 20898 6236 20904 6248
rect 20859 6208 20904 6236
rect 20898 6196 20904 6208
rect 20956 6236 20962 6248
rect 21545 6239 21603 6245
rect 21545 6236 21557 6239
rect 20956 6208 21557 6236
rect 20956 6196 20962 6208
rect 21545 6205 21557 6208
rect 21591 6205 21603 6239
rect 22278 6236 22284 6248
rect 22239 6208 22284 6236
rect 21545 6199 21603 6205
rect 22278 6196 22284 6208
rect 22336 6236 22342 6248
rect 22741 6239 22799 6245
rect 22741 6236 22753 6239
rect 22336 6208 22753 6236
rect 22336 6196 22342 6208
rect 22741 6205 22753 6208
rect 22787 6205 22799 6239
rect 22741 6199 22799 6205
rect 2774 6168 2780 6180
rect 2179 6140 2780 6168
rect 2179 6137 2191 6140
rect 2133 6131 2191 6137
rect 2774 6128 2780 6140
rect 2832 6128 2838 6180
rect 7190 6168 7196 6180
rect 7103 6140 7196 6168
rect 7190 6128 7196 6140
rect 7248 6168 7254 6180
rect 8294 6168 8300 6180
rect 7248 6140 8300 6168
rect 7248 6128 7254 6140
rect 8294 6128 8300 6140
rect 8352 6128 8358 6180
rect 9766 6177 9772 6180
rect 9760 6168 9772 6177
rect 9727 6140 9772 6168
rect 9760 6131 9772 6140
rect 9766 6128 9772 6131
rect 9824 6128 9830 6180
rect 12805 6171 12863 6177
rect 12805 6168 12817 6171
rect 12176 6140 12817 6168
rect 12176 6112 12204 6140
rect 12805 6137 12817 6140
rect 12851 6137 12863 6171
rect 12805 6131 12863 6137
rect 14544 6171 14602 6177
rect 14544 6137 14556 6171
rect 14590 6168 14602 6171
rect 14642 6168 14648 6180
rect 14590 6140 14648 6168
rect 14590 6137 14602 6140
rect 14544 6131 14602 6137
rect 14642 6128 14648 6140
rect 14700 6128 14706 6180
rect 17310 6128 17316 6180
rect 17368 6168 17374 6180
rect 19334 6168 19340 6180
rect 17368 6140 19340 6168
rect 17368 6128 17374 6140
rect 19334 6128 19340 6140
rect 19392 6168 19398 6180
rect 19981 6171 20039 6177
rect 19981 6168 19993 6171
rect 19392 6140 19993 6168
rect 19392 6128 19398 6140
rect 19981 6137 19993 6140
rect 20027 6137 20039 6171
rect 19981 6131 20039 6137
rect 1670 6100 1676 6112
rect 1631 6072 1676 6100
rect 1670 6060 1676 6072
rect 1728 6060 1734 6112
rect 3605 6103 3663 6109
rect 3605 6069 3617 6103
rect 3651 6100 3663 6103
rect 3786 6100 3792 6112
rect 3651 6072 3792 6100
rect 3651 6069 3663 6072
rect 3605 6063 3663 6069
rect 3786 6060 3792 6072
rect 3844 6060 3850 6112
rect 4246 6100 4252 6112
rect 4207 6072 4252 6100
rect 4246 6060 4252 6072
rect 4304 6060 4310 6112
rect 4614 6100 4620 6112
rect 4527 6072 4620 6100
rect 4614 6060 4620 6072
rect 4672 6100 4678 6112
rect 5442 6100 5448 6112
rect 4672 6072 5448 6100
rect 4672 6060 4678 6072
rect 5442 6060 5448 6072
rect 5500 6060 5506 6112
rect 6086 6060 6092 6112
rect 6144 6100 6150 6112
rect 6181 6103 6239 6109
rect 6181 6100 6193 6103
rect 6144 6072 6193 6100
rect 6144 6060 6150 6072
rect 6181 6069 6193 6072
rect 6227 6069 6239 6103
rect 6181 6063 6239 6069
rect 6454 6060 6460 6112
rect 6512 6100 6518 6112
rect 6641 6103 6699 6109
rect 6641 6100 6653 6103
rect 6512 6072 6653 6100
rect 6512 6060 6518 6072
rect 6641 6069 6653 6072
rect 6687 6100 6699 6103
rect 7282 6100 7288 6112
rect 6687 6072 7288 6100
rect 6687 6069 6699 6072
rect 6641 6063 6699 6069
rect 7282 6060 7288 6072
rect 7340 6060 7346 6112
rect 9858 6060 9864 6112
rect 9916 6100 9922 6112
rect 10873 6103 10931 6109
rect 10873 6100 10885 6103
rect 9916 6072 10885 6100
rect 9916 6060 9922 6072
rect 10873 6069 10885 6072
rect 10919 6069 10931 6103
rect 12158 6100 12164 6112
rect 12119 6072 12164 6100
rect 10873 6063 10931 6069
rect 12158 6060 12164 6072
rect 12216 6060 12222 6112
rect 12434 6060 12440 6112
rect 12492 6100 12498 6112
rect 12894 6100 12900 6112
rect 12492 6072 12537 6100
rect 12855 6072 12900 6100
rect 12492 6060 12498 6072
rect 12894 6060 12900 6072
rect 12952 6060 12958 6112
rect 13446 6100 13452 6112
rect 13407 6072 13452 6100
rect 13446 6060 13452 6072
rect 13504 6060 13510 6112
rect 15194 6060 15200 6112
rect 15252 6100 15258 6112
rect 15657 6103 15715 6109
rect 15657 6100 15669 6103
rect 15252 6072 15669 6100
rect 15252 6060 15258 6072
rect 15657 6069 15669 6072
rect 15703 6100 15715 6103
rect 16298 6100 16304 6112
rect 15703 6072 16304 6100
rect 15703 6069 15715 6072
rect 15657 6063 15715 6069
rect 16298 6060 16304 6072
rect 16356 6060 16362 6112
rect 17034 6100 17040 6112
rect 16995 6072 17040 6100
rect 17034 6060 17040 6072
rect 17092 6060 17098 6112
rect 22462 6100 22468 6112
rect 22423 6072 22468 6100
rect 22462 6060 22468 6072
rect 22520 6060 22526 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 2777 5899 2835 5905
rect 2777 5865 2789 5899
rect 2823 5896 2835 5899
rect 3050 5896 3056 5908
rect 2823 5868 3056 5896
rect 2823 5865 2835 5868
rect 2777 5859 2835 5865
rect 3050 5856 3056 5868
rect 3108 5856 3114 5908
rect 4798 5856 4804 5908
rect 4856 5896 4862 5908
rect 5445 5899 5503 5905
rect 5445 5896 5457 5899
rect 4856 5868 5457 5896
rect 4856 5856 4862 5868
rect 5445 5865 5457 5868
rect 5491 5865 5503 5899
rect 5445 5859 5503 5865
rect 6089 5899 6147 5905
rect 6089 5865 6101 5899
rect 6135 5896 6147 5899
rect 6178 5896 6184 5908
rect 6135 5868 6184 5896
rect 6135 5865 6147 5868
rect 6089 5859 6147 5865
rect 6178 5856 6184 5868
rect 6236 5856 6242 5908
rect 6454 5896 6460 5908
rect 6415 5868 6460 5896
rect 6454 5856 6460 5868
rect 6512 5856 6518 5908
rect 6549 5899 6607 5905
rect 6549 5865 6561 5899
rect 6595 5896 6607 5899
rect 7190 5896 7196 5908
rect 6595 5868 7196 5896
rect 6595 5865 6607 5868
rect 6549 5859 6607 5865
rect 7190 5856 7196 5868
rect 7248 5856 7254 5908
rect 7926 5896 7932 5908
rect 7887 5868 7932 5896
rect 7926 5856 7932 5868
rect 7984 5856 7990 5908
rect 9493 5899 9551 5905
rect 9493 5865 9505 5899
rect 9539 5896 9551 5899
rect 9766 5896 9772 5908
rect 9539 5868 9772 5896
rect 9539 5865 9551 5868
rect 9493 5859 9551 5865
rect 9766 5856 9772 5868
rect 9824 5896 9830 5908
rect 11057 5899 11115 5905
rect 11057 5896 11069 5899
rect 9824 5868 11069 5896
rect 9824 5856 9830 5868
rect 11057 5865 11069 5868
rect 11103 5896 11115 5899
rect 13446 5896 13452 5908
rect 11103 5868 13452 5896
rect 11103 5865 11115 5868
rect 11057 5859 11115 5865
rect 13446 5856 13452 5868
rect 13504 5856 13510 5908
rect 14369 5899 14427 5905
rect 14369 5865 14381 5899
rect 14415 5896 14427 5899
rect 14642 5896 14648 5908
rect 14415 5868 14648 5896
rect 14415 5865 14427 5868
rect 14369 5859 14427 5865
rect 14642 5856 14648 5868
rect 14700 5856 14706 5908
rect 18138 5896 18144 5908
rect 18099 5868 18144 5896
rect 18138 5856 18144 5868
rect 18196 5856 18202 5908
rect 18969 5899 19027 5905
rect 18969 5865 18981 5899
rect 19015 5896 19027 5899
rect 19242 5896 19248 5908
rect 19015 5868 19248 5896
rect 19015 5865 19027 5868
rect 18969 5859 19027 5865
rect 19242 5856 19248 5868
rect 19300 5856 19306 5908
rect 19518 5856 19524 5908
rect 19576 5896 19582 5908
rect 19705 5899 19763 5905
rect 19705 5896 19717 5899
rect 19576 5868 19717 5896
rect 19576 5856 19582 5868
rect 19705 5865 19717 5868
rect 19751 5865 19763 5899
rect 19705 5859 19763 5865
rect 20714 5856 20720 5908
rect 20772 5896 20778 5908
rect 20901 5899 20959 5905
rect 20901 5896 20913 5899
rect 20772 5868 20913 5896
rect 20772 5856 20778 5868
rect 20901 5865 20913 5868
rect 20947 5865 20959 5899
rect 20901 5859 20959 5865
rect 1762 5828 1768 5840
rect 1412 5800 1768 5828
rect 1412 5769 1440 5800
rect 1762 5788 1768 5800
rect 1820 5828 1826 5840
rect 11701 5831 11759 5837
rect 1820 5800 2820 5828
rect 1820 5788 1826 5800
rect 2792 5772 2820 5800
rect 9692 5800 11652 5828
rect 1670 5769 1676 5772
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5729 1455 5763
rect 1664 5760 1676 5769
rect 1583 5732 1676 5760
rect 1397 5723 1455 5729
rect 1664 5723 1676 5732
rect 1728 5760 1734 5772
rect 2406 5760 2412 5772
rect 1728 5732 2412 5760
rect 1670 5720 1676 5723
rect 1728 5720 1734 5732
rect 2406 5720 2412 5732
rect 2464 5720 2470 5772
rect 2774 5720 2780 5772
rect 2832 5760 2838 5772
rect 4065 5763 4123 5769
rect 4065 5760 4077 5763
rect 2832 5732 4077 5760
rect 2832 5720 2838 5732
rect 4065 5729 4077 5732
rect 4111 5760 4123 5763
rect 4154 5760 4160 5772
rect 4111 5732 4160 5760
rect 4111 5729 4123 5732
rect 4065 5723 4123 5729
rect 4154 5720 4160 5732
rect 4212 5720 4218 5772
rect 4338 5769 4344 5772
rect 4332 5760 4344 5769
rect 4299 5732 4344 5760
rect 4332 5723 4344 5732
rect 4338 5720 4344 5723
rect 4396 5720 4402 5772
rect 6914 5760 6920 5772
rect 6875 5732 6920 5760
rect 6914 5720 6920 5732
rect 6972 5720 6978 5772
rect 8294 5760 8300 5772
rect 8255 5732 8300 5760
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 9122 5720 9128 5772
rect 9180 5760 9186 5772
rect 9692 5769 9720 5800
rect 9677 5763 9735 5769
rect 9677 5760 9689 5763
rect 9180 5732 9689 5760
rect 9180 5720 9186 5732
rect 9677 5729 9689 5732
rect 9723 5729 9735 5763
rect 9677 5723 9735 5729
rect 9944 5763 10002 5769
rect 9944 5729 9956 5763
rect 9990 5760 10002 5763
rect 10686 5760 10692 5772
rect 9990 5732 10692 5760
rect 9990 5729 10002 5732
rect 9944 5723 10002 5729
rect 10686 5720 10692 5732
rect 10744 5720 10750 5772
rect 11624 5760 11652 5800
rect 11701 5797 11713 5831
rect 11747 5828 11759 5831
rect 12342 5828 12348 5840
rect 11747 5800 12348 5828
rect 11747 5797 11759 5800
rect 11701 5791 11759 5797
rect 12342 5788 12348 5800
rect 12400 5788 12406 5840
rect 15565 5831 15623 5837
rect 15565 5797 15577 5831
rect 15611 5828 15623 5831
rect 16114 5828 16120 5840
rect 15611 5800 16120 5828
rect 15611 5797 15623 5800
rect 15565 5791 15623 5797
rect 16114 5788 16120 5800
rect 16172 5828 16178 5840
rect 16758 5828 16764 5840
rect 16172 5800 16764 5828
rect 16172 5788 16178 5800
rect 16758 5788 16764 5800
rect 16816 5828 16822 5840
rect 17006 5831 17064 5837
rect 17006 5828 17018 5831
rect 16816 5800 17018 5828
rect 16816 5788 16822 5800
rect 17006 5797 17018 5800
rect 17052 5797 17064 5831
rect 17006 5791 17064 5797
rect 19426 5788 19432 5840
rect 19484 5828 19490 5840
rect 20533 5831 20591 5837
rect 20533 5828 20545 5831
rect 19484 5800 20545 5828
rect 19484 5788 19490 5800
rect 20533 5797 20545 5800
rect 20579 5828 20591 5831
rect 21450 5828 21456 5840
rect 20579 5800 21456 5828
rect 20579 5797 20591 5800
rect 20533 5791 20591 5797
rect 21450 5788 21456 5800
rect 21508 5788 21514 5840
rect 12066 5760 12072 5772
rect 11624 5732 12072 5760
rect 12066 5720 12072 5732
rect 12124 5760 12130 5772
rect 12161 5763 12219 5769
rect 12161 5760 12173 5763
rect 12124 5732 12173 5760
rect 12124 5720 12130 5732
rect 12161 5729 12173 5732
rect 12207 5729 12219 5763
rect 12161 5723 12219 5729
rect 12428 5763 12486 5769
rect 12428 5729 12440 5763
rect 12474 5760 12486 5763
rect 12986 5760 12992 5772
rect 12474 5732 12992 5760
rect 12474 5729 12486 5732
rect 12428 5723 12486 5729
rect 12986 5720 12992 5732
rect 13044 5720 13050 5772
rect 15654 5760 15660 5772
rect 15615 5732 15660 5760
rect 15654 5720 15660 5732
rect 15712 5720 15718 5772
rect 19613 5763 19671 5769
rect 19613 5729 19625 5763
rect 19659 5760 19671 5763
rect 19978 5760 19984 5772
rect 19659 5732 19984 5760
rect 19659 5729 19671 5732
rect 19613 5723 19671 5729
rect 19978 5720 19984 5732
rect 20036 5720 20042 5772
rect 20714 5720 20720 5772
rect 20772 5760 20778 5772
rect 21269 5763 21327 5769
rect 21269 5760 21281 5763
rect 20772 5732 21281 5760
rect 20772 5720 20778 5732
rect 21269 5729 21281 5732
rect 21315 5760 21327 5763
rect 22002 5760 22008 5772
rect 21315 5732 22008 5760
rect 21315 5729 21327 5732
rect 21269 5723 21327 5729
rect 22002 5720 22008 5732
rect 22060 5720 22066 5772
rect 22462 5720 22468 5772
rect 22520 5760 22526 5772
rect 23290 5760 23296 5772
rect 22520 5732 23296 5760
rect 22520 5720 22526 5732
rect 23290 5720 23296 5732
rect 23348 5720 23354 5772
rect 7009 5695 7067 5701
rect 7009 5661 7021 5695
rect 7055 5661 7067 5695
rect 7009 5655 7067 5661
rect 7193 5695 7251 5701
rect 7193 5661 7205 5695
rect 7239 5692 7251 5695
rect 7282 5692 7288 5704
rect 7239 5664 7288 5692
rect 7239 5661 7251 5664
rect 7193 5655 7251 5661
rect 3142 5584 3148 5636
rect 3200 5624 3206 5636
rect 3200 5596 3832 5624
rect 3200 5584 3206 5596
rect 3804 5568 3832 5596
rect 6914 5584 6920 5636
rect 6972 5624 6978 5636
rect 7024 5624 7052 5655
rect 7282 5652 7288 5664
rect 7340 5652 7346 5704
rect 8570 5692 8576 5704
rect 8531 5664 8576 5692
rect 8570 5652 8576 5664
rect 8628 5652 8634 5704
rect 10870 5652 10876 5704
rect 10928 5692 10934 5704
rect 11606 5692 11612 5704
rect 10928 5664 11612 5692
rect 10928 5652 10934 5664
rect 11606 5652 11612 5664
rect 11664 5652 11670 5704
rect 16482 5652 16488 5704
rect 16540 5692 16546 5704
rect 16761 5695 16819 5701
rect 16761 5692 16773 5695
rect 16540 5664 16773 5692
rect 16540 5652 16546 5664
rect 16761 5661 16773 5664
rect 16807 5661 16819 5695
rect 16761 5655 16819 5661
rect 19334 5652 19340 5704
rect 19392 5692 19398 5704
rect 19794 5692 19800 5704
rect 19392 5664 19800 5692
rect 19392 5652 19398 5664
rect 19794 5652 19800 5664
rect 19852 5652 19858 5704
rect 21361 5695 21419 5701
rect 21361 5661 21373 5695
rect 21407 5661 21419 5695
rect 21361 5655 21419 5661
rect 9030 5624 9036 5636
rect 6972 5596 7052 5624
rect 8991 5596 9036 5624
rect 6972 5584 6978 5596
rect 9030 5584 9036 5596
rect 9088 5584 9094 5636
rect 13722 5584 13728 5636
rect 13780 5624 13786 5636
rect 14645 5627 14703 5633
rect 14645 5624 14657 5627
rect 13780 5596 14657 5624
rect 13780 5584 13786 5596
rect 14645 5593 14657 5596
rect 14691 5593 14703 5627
rect 15838 5624 15844 5636
rect 15799 5596 15844 5624
rect 14645 5587 14703 5593
rect 15838 5584 15844 5596
rect 15896 5584 15902 5636
rect 19245 5627 19303 5633
rect 19245 5593 19257 5627
rect 19291 5624 19303 5627
rect 21376 5624 21404 5655
rect 21450 5652 21456 5704
rect 21508 5692 21514 5704
rect 21508 5664 21553 5692
rect 21508 5652 21514 5664
rect 21542 5624 21548 5636
rect 19291 5596 21548 5624
rect 19291 5593 19303 5596
rect 19245 5587 19303 5593
rect 21542 5584 21548 5596
rect 21600 5584 21606 5636
rect 3694 5556 3700 5568
rect 3655 5528 3700 5556
rect 3694 5516 3700 5528
rect 3752 5516 3758 5568
rect 3786 5516 3792 5568
rect 3844 5556 3850 5568
rect 7558 5556 7564 5568
rect 3844 5528 7564 5556
rect 3844 5516 3850 5528
rect 7558 5516 7564 5528
rect 7616 5516 7622 5568
rect 9398 5516 9404 5568
rect 9456 5556 9462 5568
rect 9858 5556 9864 5568
rect 9456 5528 9864 5556
rect 9456 5516 9462 5528
rect 9858 5516 9864 5528
rect 9916 5516 9922 5568
rect 12069 5559 12127 5565
rect 12069 5525 12081 5559
rect 12115 5556 12127 5559
rect 13262 5556 13268 5568
rect 12115 5528 13268 5556
rect 12115 5525 12127 5528
rect 12069 5519 12127 5525
rect 13262 5516 13268 5528
rect 13320 5556 13326 5568
rect 13446 5556 13452 5568
rect 13320 5528 13452 5556
rect 13320 5516 13326 5528
rect 13446 5516 13452 5528
rect 13504 5516 13510 5568
rect 13541 5559 13599 5565
rect 13541 5525 13553 5559
rect 13587 5556 13599 5559
rect 13630 5556 13636 5568
rect 13587 5528 13636 5556
rect 13587 5525 13599 5528
rect 13541 5519 13599 5525
rect 13630 5516 13636 5528
rect 13688 5516 13694 5568
rect 15105 5559 15163 5565
rect 15105 5525 15117 5559
rect 15151 5556 15163 5559
rect 15378 5556 15384 5568
rect 15151 5528 15384 5556
rect 15151 5525 15163 5528
rect 15105 5519 15163 5525
rect 15378 5516 15384 5528
rect 15436 5516 15442 5568
rect 16485 5559 16543 5565
rect 16485 5525 16497 5559
rect 16531 5556 16543 5559
rect 16666 5556 16672 5568
rect 16531 5528 16672 5556
rect 16531 5525 16543 5528
rect 16485 5519 16543 5525
rect 16666 5516 16672 5528
rect 16724 5516 16730 5568
rect 23474 5556 23480 5568
rect 23435 5528 23480 5556
rect 23474 5516 23480 5528
rect 23532 5516 23538 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 2406 5352 2412 5364
rect 2367 5324 2412 5352
rect 2406 5312 2412 5324
rect 2464 5312 2470 5364
rect 2869 5355 2927 5361
rect 2869 5321 2881 5355
rect 2915 5352 2927 5355
rect 3050 5352 3056 5364
rect 2915 5324 3056 5352
rect 2915 5321 2927 5324
rect 2869 5315 2927 5321
rect 1397 5287 1455 5293
rect 1397 5253 1409 5287
rect 1443 5284 1455 5287
rect 2774 5284 2780 5296
rect 1443 5256 2780 5284
rect 1443 5253 1455 5256
rect 1397 5247 1455 5253
rect 2774 5244 2780 5256
rect 2832 5244 2838 5296
rect 1578 5176 1584 5228
rect 1636 5216 1642 5228
rect 1857 5219 1915 5225
rect 1857 5216 1869 5219
rect 1636 5188 1869 5216
rect 1636 5176 1642 5188
rect 1857 5185 1869 5188
rect 1903 5185 1915 5219
rect 1857 5179 1915 5185
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5216 2099 5219
rect 2884 5216 2912 5315
rect 3050 5312 3056 5324
rect 3108 5312 3114 5364
rect 3786 5312 3792 5364
rect 3844 5352 3850 5364
rect 4154 5352 4160 5364
rect 3844 5324 4160 5352
rect 3844 5312 3850 5324
rect 4154 5312 4160 5324
rect 4212 5352 4218 5364
rect 4617 5355 4675 5361
rect 4617 5352 4629 5355
rect 4212 5324 4629 5352
rect 4212 5312 4218 5324
rect 4617 5321 4629 5324
rect 4663 5352 4675 5355
rect 6086 5352 6092 5364
rect 4663 5324 6092 5352
rect 4663 5321 4675 5324
rect 4617 5315 4675 5321
rect 6086 5312 6092 5324
rect 6144 5312 6150 5364
rect 9122 5352 9128 5364
rect 9083 5324 9128 5352
rect 9122 5312 9128 5324
rect 9180 5312 9186 5364
rect 12986 5352 12992 5364
rect 12947 5324 12992 5352
rect 12986 5312 12992 5324
rect 13044 5312 13050 5364
rect 14642 5312 14648 5364
rect 14700 5352 14706 5364
rect 14921 5355 14979 5361
rect 14921 5352 14933 5355
rect 14700 5324 14933 5352
rect 14700 5312 14706 5324
rect 14921 5321 14933 5324
rect 14967 5321 14979 5355
rect 14921 5315 14979 5321
rect 16482 5312 16488 5364
rect 16540 5352 16546 5364
rect 17402 5352 17408 5364
rect 16540 5324 17408 5352
rect 16540 5312 16546 5324
rect 17402 5312 17408 5324
rect 17460 5312 17466 5364
rect 18049 5355 18107 5361
rect 18049 5321 18061 5355
rect 18095 5352 18107 5355
rect 18230 5352 18236 5364
rect 18095 5324 18236 5352
rect 18095 5321 18107 5324
rect 18049 5315 18107 5321
rect 18230 5312 18236 5324
rect 18288 5312 18294 5364
rect 19613 5355 19671 5361
rect 19613 5321 19625 5355
rect 19659 5352 19671 5355
rect 20714 5352 20720 5364
rect 19659 5324 20720 5352
rect 19659 5321 19671 5324
rect 19613 5315 19671 5321
rect 20714 5312 20720 5324
rect 20772 5312 20778 5364
rect 21450 5312 21456 5364
rect 21508 5352 21514 5364
rect 21637 5355 21695 5361
rect 21637 5352 21649 5355
rect 21508 5324 21649 5352
rect 21508 5312 21514 5324
rect 21637 5321 21649 5324
rect 21683 5321 21695 5355
rect 21637 5315 21695 5321
rect 22094 5312 22100 5364
rect 22152 5352 22158 5364
rect 23290 5352 23296 5364
rect 22152 5324 22197 5352
rect 23251 5324 23296 5352
rect 22152 5312 22158 5324
rect 23290 5312 23296 5324
rect 23348 5312 23354 5364
rect 6178 5284 6184 5296
rect 5828 5256 6184 5284
rect 2087 5188 2912 5216
rect 2087 5185 2099 5188
rect 2041 5179 2099 5185
rect 3694 5176 3700 5228
rect 3752 5216 3758 5228
rect 5828 5225 5856 5256
rect 6178 5244 6184 5256
rect 6236 5284 6242 5296
rect 6362 5284 6368 5296
rect 6236 5256 6368 5284
rect 6236 5244 6242 5256
rect 6362 5244 6368 5256
rect 6420 5244 6426 5296
rect 6822 5284 6828 5296
rect 6564 5256 6828 5284
rect 4249 5219 4307 5225
rect 4249 5216 4261 5219
rect 3752 5188 4261 5216
rect 3752 5176 3758 5188
rect 4249 5185 4261 5188
rect 4295 5216 4307 5219
rect 5813 5219 5871 5225
rect 5813 5216 5825 5219
rect 4295 5188 5825 5216
rect 4295 5185 4307 5188
rect 4249 5179 4307 5185
rect 5813 5185 5825 5188
rect 5859 5185 5871 5219
rect 5813 5179 5871 5185
rect 1394 5108 1400 5160
rect 1452 5148 1458 5160
rect 1765 5151 1823 5157
rect 1765 5148 1777 5151
rect 1452 5120 1777 5148
rect 1452 5108 1458 5120
rect 1765 5117 1777 5120
rect 1811 5117 1823 5151
rect 1765 5111 1823 5117
rect 4065 5151 4123 5157
rect 4065 5117 4077 5151
rect 4111 5148 4123 5151
rect 4154 5148 4160 5160
rect 4111 5120 4160 5148
rect 4111 5117 4123 5120
rect 4065 5111 4123 5117
rect 4154 5108 4160 5120
rect 4212 5108 4218 5160
rect 5442 5108 5448 5160
rect 5500 5148 5506 5160
rect 6178 5148 6184 5160
rect 5500 5120 6184 5148
rect 5500 5108 5506 5120
rect 6178 5108 6184 5120
rect 6236 5148 6242 5160
rect 6564 5157 6592 5256
rect 6822 5244 6828 5256
rect 6880 5244 6886 5296
rect 12066 5244 12072 5296
rect 12124 5284 12130 5296
rect 12161 5287 12219 5293
rect 12161 5284 12173 5287
rect 12124 5256 12173 5284
rect 12124 5244 12130 5256
rect 12161 5253 12173 5256
rect 12207 5253 12219 5287
rect 12161 5247 12219 5253
rect 16301 5287 16359 5293
rect 16301 5253 16313 5287
rect 16347 5284 16359 5287
rect 18138 5284 18144 5296
rect 16347 5256 18144 5284
rect 16347 5253 16359 5256
rect 16301 5247 16359 5253
rect 8849 5219 8907 5225
rect 8849 5185 8861 5219
rect 8895 5216 8907 5219
rect 8895 5188 9444 5216
rect 8895 5185 8907 5188
rect 8849 5179 8907 5185
rect 6549 5151 6607 5157
rect 6549 5148 6561 5151
rect 6236 5120 6561 5148
rect 6236 5108 6242 5120
rect 6549 5117 6561 5120
rect 6595 5117 6607 5151
rect 6822 5148 6828 5160
rect 6783 5120 6828 5148
rect 6549 5111 6607 5117
rect 6822 5108 6828 5120
rect 6880 5108 6886 5160
rect 7092 5151 7150 5157
rect 7092 5117 7104 5151
rect 7138 5148 7150 5151
rect 7558 5148 7564 5160
rect 7138 5120 7564 5148
rect 7138 5117 7150 5120
rect 7092 5111 7150 5117
rect 7558 5108 7564 5120
rect 7616 5108 7622 5160
rect 9122 5108 9128 5160
rect 9180 5148 9186 5160
rect 9309 5151 9367 5157
rect 9309 5148 9321 5151
rect 9180 5120 9321 5148
rect 9180 5108 9186 5120
rect 9309 5117 9321 5120
rect 9355 5117 9367 5151
rect 9416 5148 9444 5188
rect 9582 5157 9588 5160
rect 9576 5148 9588 5157
rect 9416 5120 9588 5148
rect 9309 5111 9367 5117
rect 9576 5111 9588 5120
rect 9582 5108 9588 5111
rect 9640 5108 9646 5160
rect 3513 5083 3571 5089
rect 3513 5049 3525 5083
rect 3559 5080 3571 5083
rect 5077 5083 5135 5089
rect 3559 5052 3924 5080
rect 3559 5049 3571 5052
rect 3513 5043 3571 5049
rect 3896 5024 3924 5052
rect 5077 5049 5089 5083
rect 5123 5080 5135 5083
rect 6730 5080 6736 5092
rect 5123 5052 5580 5080
rect 5123 5049 5135 5052
rect 5077 5043 5135 5049
rect 5552 5024 5580 5052
rect 6288 5052 6736 5080
rect 6288 5024 6316 5052
rect 6730 5040 6736 5052
rect 6788 5040 6794 5092
rect 9950 5040 9956 5092
rect 10008 5080 10014 5092
rect 11241 5083 11299 5089
rect 11241 5080 11253 5083
rect 10008 5052 11253 5080
rect 10008 5040 10014 5052
rect 11241 5049 11253 5052
rect 11287 5049 11299 5083
rect 12176 5080 12204 5247
rect 17052 5225 17080 5256
rect 18138 5244 18144 5256
rect 18196 5244 18202 5296
rect 19518 5244 19524 5296
rect 19576 5284 19582 5296
rect 20625 5287 20683 5293
rect 20625 5284 20637 5287
rect 19576 5256 20637 5284
rect 19576 5244 19582 5256
rect 20625 5253 20637 5256
rect 20671 5253 20683 5287
rect 22370 5284 22376 5296
rect 22331 5256 22376 5284
rect 20625 5247 20683 5253
rect 22370 5244 22376 5256
rect 22428 5244 22434 5296
rect 17037 5219 17095 5225
rect 17037 5185 17049 5219
rect 17083 5185 17095 5219
rect 17770 5216 17776 5228
rect 17731 5188 17776 5216
rect 17037 5179 17095 5185
rect 17770 5176 17776 5188
rect 17828 5216 17834 5228
rect 18598 5216 18604 5228
rect 17828 5188 18460 5216
rect 18559 5188 18604 5216
rect 17828 5176 17834 5188
rect 12342 5108 12348 5160
rect 12400 5148 12406 5160
rect 12526 5148 12532 5160
rect 12400 5120 12532 5148
rect 12400 5108 12406 5120
rect 12526 5108 12532 5120
rect 12584 5108 12590 5160
rect 13541 5151 13599 5157
rect 13541 5117 13553 5151
rect 13587 5117 13599 5151
rect 15654 5148 15660 5160
rect 15615 5120 15660 5148
rect 13541 5111 13599 5117
rect 13357 5083 13415 5089
rect 13357 5080 13369 5083
rect 12176 5052 13369 5080
rect 11241 5043 11299 5049
rect 13357 5049 13369 5052
rect 13403 5080 13415 5083
rect 13556 5080 13584 5111
rect 15654 5108 15660 5120
rect 15712 5108 15718 5160
rect 16574 5108 16580 5160
rect 16632 5148 16638 5160
rect 18432 5157 18460 5188
rect 18598 5176 18604 5188
rect 18656 5176 18662 5228
rect 19794 5176 19800 5228
rect 19852 5216 19858 5228
rect 20165 5219 20223 5225
rect 20165 5216 20177 5219
rect 19852 5188 20177 5216
rect 19852 5176 19858 5188
rect 20165 5185 20177 5188
rect 20211 5216 20223 5219
rect 20254 5216 20260 5228
rect 20211 5188 20260 5216
rect 20211 5185 20223 5188
rect 20165 5179 20223 5185
rect 20254 5176 20260 5188
rect 20312 5216 20318 5228
rect 20993 5219 21051 5225
rect 20993 5216 21005 5219
rect 20312 5188 21005 5216
rect 20312 5176 20318 5188
rect 20993 5185 21005 5188
rect 21039 5185 21051 5219
rect 20993 5179 21051 5185
rect 16761 5151 16819 5157
rect 16761 5148 16773 5151
rect 16632 5120 16773 5148
rect 16632 5108 16638 5120
rect 16761 5117 16773 5120
rect 16807 5117 16819 5151
rect 16761 5111 16819 5117
rect 18417 5151 18475 5157
rect 18417 5117 18429 5151
rect 18463 5117 18475 5151
rect 18417 5111 18475 5117
rect 18506 5108 18512 5160
rect 18564 5148 18570 5160
rect 18564 5120 18609 5148
rect 18564 5108 18570 5120
rect 20714 5108 20720 5160
rect 20772 5148 20778 5160
rect 21177 5151 21235 5157
rect 21177 5148 21189 5151
rect 20772 5120 21189 5148
rect 20772 5108 20778 5120
rect 21177 5117 21189 5120
rect 21223 5148 21235 5151
rect 21818 5148 21824 5160
rect 21223 5120 21824 5148
rect 21223 5117 21235 5120
rect 21177 5111 21235 5117
rect 21818 5108 21824 5120
rect 21876 5108 21882 5160
rect 22738 5148 22744 5160
rect 22699 5120 22744 5148
rect 22738 5108 22744 5120
rect 22796 5108 22802 5160
rect 13403 5052 13584 5080
rect 13403 5049 13415 5052
rect 13357 5043 13415 5049
rect 13630 5040 13636 5092
rect 13688 5080 13694 5092
rect 13786 5083 13844 5089
rect 13786 5080 13798 5083
rect 13688 5052 13798 5080
rect 13688 5040 13694 5052
rect 13786 5049 13798 5052
rect 13832 5049 13844 5083
rect 13786 5043 13844 5049
rect 16482 5040 16488 5092
rect 16540 5080 16546 5092
rect 16850 5080 16856 5092
rect 16540 5052 16856 5080
rect 16540 5040 16546 5052
rect 16850 5040 16856 5052
rect 16908 5040 16914 5092
rect 19981 5083 20039 5089
rect 19981 5080 19993 5083
rect 19076 5052 19993 5080
rect 3602 5012 3608 5024
rect 3563 4984 3608 5012
rect 3602 4972 3608 4984
rect 3660 4972 3666 5024
rect 3878 4972 3884 5024
rect 3936 5012 3942 5024
rect 3973 5015 4031 5021
rect 3973 5012 3985 5015
rect 3936 4984 3985 5012
rect 3936 4972 3942 4984
rect 3973 4981 3985 4984
rect 4019 4981 4031 5015
rect 5166 5012 5172 5024
rect 5127 4984 5172 5012
rect 3973 4975 4031 4981
rect 5166 4972 5172 4984
rect 5224 4972 5230 5024
rect 5534 5012 5540 5024
rect 5495 4984 5540 5012
rect 5534 4972 5540 4984
rect 5592 4972 5598 5024
rect 5626 4972 5632 5024
rect 5684 5012 5690 5024
rect 6270 5012 6276 5024
rect 5684 4984 5729 5012
rect 6231 4984 6276 5012
rect 5684 4972 5690 4984
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 8018 4972 8024 5024
rect 8076 5012 8082 5024
rect 8205 5015 8263 5021
rect 8205 5012 8217 5015
rect 8076 4984 8217 5012
rect 8076 4972 8082 4984
rect 8205 4981 8217 4984
rect 8251 4981 8263 5015
rect 10686 5012 10692 5024
rect 10647 4984 10692 5012
rect 8205 4975 8263 4981
rect 10686 4972 10692 4984
rect 10744 4972 10750 5024
rect 11146 4972 11152 5024
rect 11204 5012 11210 5024
rect 11609 5015 11667 5021
rect 11609 5012 11621 5015
rect 11204 4984 11621 5012
rect 11204 4972 11210 4984
rect 11609 4981 11621 4984
rect 11655 4981 11667 5015
rect 12710 5012 12716 5024
rect 12671 4984 12716 5012
rect 11609 4975 11667 4981
rect 12710 4972 12716 4984
rect 12768 4972 12774 5024
rect 12802 4972 12808 5024
rect 12860 5012 12866 5024
rect 13078 5012 13084 5024
rect 12860 4984 13084 5012
rect 12860 4972 12866 4984
rect 13078 4972 13084 4984
rect 13136 4972 13142 5024
rect 16390 5012 16396 5024
rect 16351 4984 16396 5012
rect 16390 4972 16396 4984
rect 16448 4972 16454 5024
rect 18966 4972 18972 5024
rect 19024 5012 19030 5024
rect 19076 5021 19104 5052
rect 19981 5049 19993 5052
rect 20027 5049 20039 5083
rect 19981 5043 20039 5049
rect 19061 5015 19119 5021
rect 19061 5012 19073 5015
rect 19024 4984 19073 5012
rect 19024 4972 19030 4984
rect 19061 4981 19073 4984
rect 19107 4981 19119 5015
rect 19061 4975 19119 4981
rect 19334 4972 19340 5024
rect 19392 5012 19398 5024
rect 19521 5015 19579 5021
rect 19521 5012 19533 5015
rect 19392 4984 19533 5012
rect 19392 4972 19398 4984
rect 19521 4981 19533 4984
rect 19567 5012 19579 5015
rect 20073 5015 20131 5021
rect 20073 5012 20085 5015
rect 19567 4984 20085 5012
rect 19567 4981 19579 4984
rect 19521 4975 19579 4981
rect 20073 4981 20085 4984
rect 20119 4981 20131 5015
rect 21358 5012 21364 5024
rect 21319 4984 21364 5012
rect 20073 4975 20131 4981
rect 21358 4972 21364 4984
rect 21416 4972 21422 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1673 4811 1731 4817
rect 1673 4777 1685 4811
rect 1719 4808 1731 4811
rect 1762 4808 1768 4820
rect 1719 4780 1768 4808
rect 1719 4777 1731 4780
rect 1673 4771 1731 4777
rect 1762 4768 1768 4780
rect 1820 4768 1826 4820
rect 2869 4811 2927 4817
rect 2869 4777 2881 4811
rect 2915 4808 2927 4811
rect 2958 4808 2964 4820
rect 2915 4780 2964 4808
rect 2915 4777 2927 4780
rect 2869 4771 2927 4777
rect 2958 4768 2964 4780
rect 3016 4768 3022 4820
rect 3697 4811 3755 4817
rect 3697 4777 3709 4811
rect 3743 4808 3755 4811
rect 4154 4808 4160 4820
rect 3743 4780 4160 4808
rect 3743 4777 3755 4780
rect 3697 4771 3755 4777
rect 4154 4768 4160 4780
rect 4212 4768 4218 4820
rect 4338 4808 4344 4820
rect 4299 4780 4344 4808
rect 4338 4768 4344 4780
rect 4396 4768 4402 4820
rect 5166 4768 5172 4820
rect 5224 4808 5230 4820
rect 5905 4811 5963 4817
rect 5905 4808 5917 4811
rect 5224 4780 5917 4808
rect 5224 4768 5230 4780
rect 5905 4777 5917 4780
rect 5951 4777 5963 4811
rect 5905 4771 5963 4777
rect 5994 4768 6000 4820
rect 6052 4808 6058 4820
rect 6052 4780 6097 4808
rect 6052 4768 6058 4780
rect 6822 4768 6828 4820
rect 6880 4768 6886 4820
rect 7098 4808 7104 4820
rect 7059 4780 7104 4808
rect 7098 4768 7104 4780
rect 7156 4768 7162 4820
rect 9122 4768 9128 4820
rect 9180 4808 9186 4820
rect 9309 4811 9367 4817
rect 9309 4808 9321 4811
rect 9180 4780 9321 4808
rect 9180 4768 9186 4780
rect 9309 4777 9321 4780
rect 9355 4777 9367 4811
rect 10962 4808 10968 4820
rect 10923 4780 10968 4808
rect 9309 4771 9367 4777
rect 10962 4768 10968 4780
rect 11020 4768 11026 4820
rect 11330 4768 11336 4820
rect 11388 4808 11394 4820
rect 11425 4811 11483 4817
rect 11425 4808 11437 4811
rect 11388 4780 11437 4808
rect 11388 4768 11394 4780
rect 11425 4777 11437 4780
rect 11471 4777 11483 4811
rect 11425 4771 11483 4777
rect 11882 4768 11888 4820
rect 11940 4808 11946 4820
rect 11977 4811 12035 4817
rect 11977 4808 11989 4811
rect 11940 4780 11989 4808
rect 11940 4768 11946 4780
rect 11977 4777 11989 4780
rect 12023 4777 12035 4811
rect 11977 4771 12035 4777
rect 2774 4700 2780 4752
rect 2832 4740 2838 4752
rect 2832 4712 2877 4740
rect 2832 4700 2838 4712
rect 4430 4700 4436 4752
rect 4488 4740 4494 4752
rect 5350 4740 5356 4752
rect 4488 4712 5356 4740
rect 4488 4700 4494 4712
rect 5350 4700 5356 4712
rect 5408 4700 5414 4752
rect 6086 4700 6092 4752
rect 6144 4740 6150 4752
rect 6840 4740 6868 4768
rect 6917 4743 6975 4749
rect 6917 4740 6929 4743
rect 6144 4712 6929 4740
rect 6144 4700 6150 4712
rect 6917 4709 6929 4712
rect 6963 4709 6975 4743
rect 10502 4740 10508 4752
rect 10463 4712 10508 4740
rect 6917 4703 6975 4709
rect 10502 4700 10508 4712
rect 10560 4740 10566 4752
rect 10686 4740 10692 4752
rect 10560 4712 10692 4740
rect 10560 4700 10566 4712
rect 10686 4700 10692 4712
rect 10744 4700 10750 4752
rect 5534 4632 5540 4684
rect 5592 4672 5598 4684
rect 6822 4672 6828 4684
rect 5592 4644 6828 4672
rect 5592 4632 5598 4644
rect 6822 4632 6828 4644
rect 6880 4632 6886 4684
rect 7190 4632 7196 4684
rect 7248 4672 7254 4684
rect 7469 4675 7527 4681
rect 7469 4672 7481 4675
rect 7248 4644 7481 4672
rect 7248 4632 7254 4644
rect 7469 4641 7481 4644
rect 7515 4672 7527 4675
rect 7742 4672 7748 4684
rect 7515 4644 7748 4672
rect 7515 4641 7527 4644
rect 7469 4635 7527 4641
rect 7742 4632 7748 4644
rect 7800 4632 7806 4684
rect 9950 4672 9956 4684
rect 9911 4644 9956 4672
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 10042 4632 10048 4684
rect 10100 4672 10106 4684
rect 10781 4675 10839 4681
rect 10781 4672 10793 4675
rect 10100 4644 10793 4672
rect 10100 4632 10106 4644
rect 10781 4641 10793 4644
rect 10827 4641 10839 4675
rect 10781 4635 10839 4641
rect 11333 4675 11391 4681
rect 11333 4641 11345 4675
rect 11379 4672 11391 4675
rect 11698 4672 11704 4684
rect 11379 4644 11704 4672
rect 11379 4641 11391 4644
rect 11333 4635 11391 4641
rect 11698 4632 11704 4644
rect 11756 4632 11762 4684
rect 11992 4672 12020 4771
rect 12434 4768 12440 4820
rect 12492 4808 12498 4820
rect 12897 4811 12955 4817
rect 12897 4808 12909 4811
rect 12492 4780 12909 4808
rect 12492 4768 12498 4780
rect 12897 4777 12909 4780
rect 12943 4808 12955 4811
rect 13909 4811 13967 4817
rect 13909 4808 13921 4811
rect 12943 4780 13921 4808
rect 12943 4777 12955 4780
rect 12897 4771 12955 4777
rect 13909 4777 13921 4780
rect 13955 4777 13967 4811
rect 16114 4808 16120 4820
rect 16075 4780 16120 4808
rect 13909 4771 13967 4777
rect 16114 4768 16120 4780
rect 16172 4768 16178 4820
rect 16206 4768 16212 4820
rect 16264 4808 16270 4820
rect 16485 4811 16543 4817
rect 16485 4808 16497 4811
rect 16264 4780 16497 4808
rect 16264 4768 16270 4780
rect 16485 4777 16497 4780
rect 16531 4777 16543 4811
rect 16942 4808 16948 4820
rect 16903 4780 16948 4808
rect 16485 4771 16543 4777
rect 16942 4768 16948 4780
rect 17000 4808 17006 4820
rect 18138 4808 18144 4820
rect 17000 4780 18144 4808
rect 17000 4768 17006 4780
rect 18138 4768 18144 4780
rect 18196 4768 18202 4820
rect 20254 4808 20260 4820
rect 20215 4780 20260 4808
rect 20254 4768 20260 4780
rect 20312 4768 20318 4820
rect 21542 4808 21548 4820
rect 21503 4780 21548 4808
rect 21542 4768 21548 4780
rect 21600 4768 21606 4820
rect 21818 4808 21824 4820
rect 21779 4780 21824 4808
rect 21818 4768 21824 4780
rect 21876 4768 21882 4820
rect 12986 4740 12992 4752
rect 12899 4712 12992 4740
rect 12986 4700 12992 4712
rect 13044 4740 13050 4752
rect 13722 4740 13728 4752
rect 13044 4712 13728 4740
rect 13044 4700 13050 4712
rect 13722 4700 13728 4712
rect 13780 4700 13786 4752
rect 19337 4743 19395 4749
rect 19337 4740 19349 4743
rect 15304 4712 19349 4740
rect 15304 4684 15332 4712
rect 19337 4709 19349 4712
rect 19383 4740 19395 4743
rect 19978 4740 19984 4752
rect 19383 4712 19984 4740
rect 19383 4709 19395 4712
rect 19337 4703 19395 4709
rect 19978 4700 19984 4712
rect 20036 4700 20042 4752
rect 11992 4644 12664 4672
rect 2958 4604 2964 4616
rect 2919 4576 2964 4604
rect 2958 4564 2964 4576
rect 3016 4564 3022 4616
rect 6086 4604 6092 4616
rect 6047 4576 6092 4604
rect 6086 4564 6092 4576
rect 6144 4564 6150 4616
rect 7558 4604 7564 4616
rect 7519 4576 7564 4604
rect 7558 4564 7564 4576
rect 7616 4564 7622 4616
rect 7653 4607 7711 4613
rect 7653 4573 7665 4607
rect 7699 4573 7711 4607
rect 7653 4567 7711 4573
rect 2406 4536 2412 4548
rect 2367 4508 2412 4536
rect 2406 4496 2412 4508
rect 2464 4496 2470 4548
rect 2317 4471 2375 4477
rect 2317 4437 2329 4471
rect 2363 4468 2375 4471
rect 2976 4468 3004 4564
rect 5261 4539 5319 4545
rect 5261 4505 5273 4539
rect 5307 4536 5319 4539
rect 5626 4536 5632 4548
rect 5307 4508 5632 4536
rect 5307 4505 5319 4508
rect 5261 4499 5319 4505
rect 5626 4496 5632 4508
rect 5684 4536 5690 4548
rect 6730 4536 6736 4548
rect 5684 4508 6736 4536
rect 5684 4496 5690 4508
rect 6730 4496 6736 4508
rect 6788 4496 6794 4548
rect 7282 4496 7288 4548
rect 7340 4536 7346 4548
rect 7668 4536 7696 4567
rect 10134 4564 10140 4616
rect 10192 4604 10198 4616
rect 10686 4604 10692 4616
rect 10192 4576 10692 4604
rect 10192 4564 10198 4576
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 11606 4604 11612 4616
rect 11519 4576 11612 4604
rect 11606 4564 11612 4576
rect 11664 4604 11670 4616
rect 12636 4604 12664 4644
rect 12710 4632 12716 4684
rect 12768 4672 12774 4684
rect 14093 4675 14151 4681
rect 14093 4672 14105 4675
rect 12768 4644 14105 4672
rect 12768 4632 12774 4644
rect 14093 4641 14105 4644
rect 14139 4672 14151 4675
rect 14642 4672 14648 4684
rect 14139 4644 14648 4672
rect 14139 4641 14151 4644
rect 14093 4635 14151 4641
rect 14642 4632 14648 4644
rect 14700 4632 14706 4684
rect 15286 4672 15292 4684
rect 15247 4644 15292 4672
rect 15286 4632 15292 4644
rect 15344 4632 15350 4684
rect 16850 4672 16856 4684
rect 16811 4644 16856 4672
rect 16850 4632 16856 4644
rect 16908 4632 16914 4684
rect 17494 4672 17500 4684
rect 17455 4644 17500 4672
rect 17494 4632 17500 4644
rect 17552 4672 17558 4684
rect 17865 4675 17923 4681
rect 17865 4672 17877 4675
rect 17552 4644 17877 4672
rect 17552 4632 17558 4644
rect 17865 4641 17877 4644
rect 17911 4641 17923 4675
rect 17865 4635 17923 4641
rect 13078 4604 13084 4616
rect 11664 4576 12480 4604
rect 12636 4576 13084 4604
rect 11664 4564 11670 4576
rect 7340 4508 7696 4536
rect 7340 4496 7346 4508
rect 4614 4468 4620 4480
rect 2363 4440 3004 4468
rect 4575 4440 4620 4468
rect 2363 4437 2375 4440
rect 2317 4431 2375 4437
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 5534 4468 5540 4480
rect 5495 4440 5540 4468
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 8110 4468 8116 4480
rect 8071 4440 8116 4468
rect 8110 4428 8116 4440
rect 8168 4428 8174 4480
rect 8294 4428 8300 4480
rect 8352 4468 8358 4480
rect 8481 4471 8539 4477
rect 8481 4468 8493 4471
rect 8352 4440 8493 4468
rect 8352 4428 8358 4440
rect 8481 4437 8493 4440
rect 8527 4437 8539 4471
rect 8846 4468 8852 4480
rect 8807 4440 8852 4468
rect 8481 4431 8539 4437
rect 8846 4428 8852 4440
rect 8904 4428 8910 4480
rect 10137 4471 10195 4477
rect 10137 4437 10149 4471
rect 10183 4468 10195 4471
rect 10962 4468 10968 4480
rect 10183 4440 10968 4468
rect 10183 4437 10195 4440
rect 10137 4431 10195 4437
rect 10962 4428 10968 4440
rect 11020 4428 11026 4480
rect 12452 4477 12480 4576
rect 13078 4564 13084 4576
rect 13136 4564 13142 4616
rect 13630 4604 13636 4616
rect 13591 4576 13636 4604
rect 13630 4564 13636 4576
rect 13688 4564 13694 4616
rect 13722 4564 13728 4616
rect 13780 4604 13786 4616
rect 15013 4607 15071 4613
rect 15013 4604 15025 4607
rect 13780 4576 15025 4604
rect 13780 4564 13786 4576
rect 15013 4573 15025 4576
rect 15059 4573 15071 4607
rect 15013 4567 15071 4573
rect 16574 4564 16580 4616
rect 16632 4604 16638 4616
rect 17129 4607 17187 4613
rect 17129 4604 17141 4607
rect 16632 4576 17141 4604
rect 16632 4564 16638 4576
rect 17129 4573 17141 4576
rect 17175 4604 17187 4607
rect 17678 4604 17684 4616
rect 17175 4576 17684 4604
rect 17175 4573 17187 4576
rect 17129 4567 17187 4573
rect 17678 4564 17684 4576
rect 17736 4564 17742 4616
rect 12529 4539 12587 4545
rect 12529 4505 12541 4539
rect 12575 4536 12587 4539
rect 14366 4536 14372 4548
rect 12575 4508 14372 4536
rect 12575 4505 12587 4508
rect 12529 4499 12587 4505
rect 14366 4496 14372 4508
rect 14424 4536 14430 4548
rect 14645 4539 14703 4545
rect 14645 4536 14657 4539
rect 14424 4508 14657 4536
rect 14424 4496 14430 4508
rect 14645 4505 14657 4508
rect 14691 4505 14703 4539
rect 15470 4536 15476 4548
rect 15431 4508 15476 4536
rect 14645 4499 14703 4505
rect 15470 4496 15476 4508
rect 15528 4496 15534 4548
rect 17880 4536 17908 4635
rect 18046 4632 18052 4684
rect 18104 4672 18110 4684
rect 18417 4675 18475 4681
rect 18417 4672 18429 4675
rect 18104 4644 18429 4672
rect 18104 4632 18110 4644
rect 18417 4641 18429 4644
rect 18463 4641 18475 4675
rect 18417 4635 18475 4641
rect 19518 4632 19524 4684
rect 19576 4672 19582 4684
rect 19613 4675 19671 4681
rect 19613 4672 19625 4675
rect 19576 4644 19625 4672
rect 19576 4632 19582 4644
rect 19613 4641 19625 4644
rect 19659 4641 19671 4675
rect 19613 4635 19671 4641
rect 20901 4675 20959 4681
rect 20901 4641 20913 4675
rect 20947 4672 20959 4675
rect 21358 4672 21364 4684
rect 20947 4644 21364 4672
rect 20947 4641 20959 4644
rect 20901 4635 20959 4641
rect 21358 4632 21364 4644
rect 21416 4632 21422 4684
rect 18506 4604 18512 4616
rect 18467 4576 18512 4604
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 18598 4564 18604 4616
rect 18656 4604 18662 4616
rect 18656 4576 18749 4604
rect 18656 4564 18662 4576
rect 18616 4536 18644 4564
rect 17880 4508 18644 4536
rect 19797 4539 19855 4545
rect 19797 4505 19809 4539
rect 19843 4536 19855 4539
rect 21266 4536 21272 4548
rect 19843 4508 21272 4536
rect 19843 4505 19855 4508
rect 19797 4499 19855 4505
rect 21266 4496 21272 4508
rect 21324 4496 21330 4548
rect 12437 4471 12495 4477
rect 12437 4437 12449 4471
rect 12483 4468 12495 4471
rect 13262 4468 13268 4480
rect 12483 4440 13268 4468
rect 12483 4437 12495 4440
rect 12437 4431 12495 4437
rect 13262 4428 13268 4440
rect 13320 4428 13326 4480
rect 14277 4471 14335 4477
rect 14277 4437 14289 4471
rect 14323 4468 14335 4471
rect 17494 4468 17500 4480
rect 14323 4440 17500 4468
rect 14323 4437 14335 4440
rect 14277 4431 14335 4437
rect 17494 4428 17500 4440
rect 17552 4428 17558 4480
rect 18049 4471 18107 4477
rect 18049 4437 18061 4471
rect 18095 4468 18107 4471
rect 18322 4468 18328 4480
rect 18095 4440 18328 4468
rect 18095 4437 18107 4440
rect 18049 4431 18107 4437
rect 18322 4428 18328 4440
rect 18380 4428 18386 4480
rect 20530 4468 20536 4480
rect 20491 4440 20536 4468
rect 20530 4428 20536 4440
rect 20588 4428 20594 4480
rect 20806 4428 20812 4480
rect 20864 4468 20870 4480
rect 21085 4471 21143 4477
rect 21085 4468 21097 4471
rect 20864 4440 21097 4468
rect 20864 4428 20870 4440
rect 21085 4437 21097 4440
rect 21131 4437 21143 4471
rect 21085 4431 21143 4437
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 3786 4264 3792 4276
rect 3747 4236 3792 4264
rect 3786 4224 3792 4236
rect 3844 4224 3850 4276
rect 5994 4224 6000 4276
rect 6052 4264 6058 4276
rect 6181 4267 6239 4273
rect 6181 4264 6193 4267
rect 6052 4236 6193 4264
rect 6052 4224 6058 4236
rect 6181 4233 6193 4236
rect 6227 4233 6239 4267
rect 7558 4264 7564 4276
rect 7519 4236 7564 4264
rect 6181 4227 6239 4233
rect 7558 4224 7564 4236
rect 7616 4224 7622 4276
rect 9950 4264 9956 4276
rect 9863 4236 9956 4264
rect 2958 4128 2964 4140
rect 2919 4100 2964 4128
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 3804 4128 3832 4224
rect 7282 4196 7288 4208
rect 6932 4168 7288 4196
rect 3881 4131 3939 4137
rect 3881 4128 3893 4131
rect 3804 4100 3893 4128
rect 3881 4097 3893 4100
rect 3927 4097 3939 4131
rect 3881 4091 3939 4097
rect 6641 4131 6699 4137
rect 6641 4097 6653 4131
rect 6687 4128 6699 4131
rect 6932 4128 6960 4168
rect 7282 4156 7288 4168
rect 7340 4156 7346 4208
rect 8110 4156 8116 4208
rect 8168 4196 8174 4208
rect 8168 4168 8248 4196
rect 8168 4156 8174 4168
rect 6687 4100 6960 4128
rect 8220 4128 8248 4168
rect 8297 4131 8355 4137
rect 8297 4128 8309 4131
rect 8220 4100 8309 4128
rect 6687 4097 6699 4100
rect 6641 4091 6699 4097
rect 8297 4097 8309 4100
rect 8343 4128 8355 4131
rect 9766 4128 9772 4140
rect 8343 4100 9772 4128
rect 8343 4097 8355 4100
rect 8297 4091 8355 4097
rect 9766 4088 9772 4100
rect 9824 4088 9830 4140
rect 9876 4137 9904 4236
rect 9950 4224 9956 4236
rect 10008 4264 10014 4276
rect 10689 4267 10747 4273
rect 10689 4264 10701 4267
rect 10008 4236 10701 4264
rect 10008 4224 10014 4236
rect 10689 4233 10701 4236
rect 10735 4264 10747 4267
rect 11606 4264 11612 4276
rect 10735 4236 11612 4264
rect 10735 4233 10747 4236
rect 10689 4227 10747 4233
rect 11606 4224 11612 4236
rect 11664 4224 11670 4276
rect 11698 4224 11704 4276
rect 11756 4264 11762 4276
rect 11756 4236 11801 4264
rect 11756 4224 11762 4236
rect 12526 4224 12532 4276
rect 12584 4264 12590 4276
rect 14001 4267 14059 4273
rect 14001 4264 14013 4267
rect 12584 4236 14013 4264
rect 12584 4224 12590 4236
rect 14001 4233 14013 4236
rect 14047 4233 14059 4267
rect 15286 4264 15292 4276
rect 15247 4236 15292 4264
rect 14001 4227 14059 4233
rect 15286 4224 15292 4236
rect 15344 4224 15350 4276
rect 16114 4224 16120 4276
rect 16172 4264 16178 4276
rect 16172 4236 16712 4264
rect 16172 4224 16178 4236
rect 11146 4156 11152 4208
rect 11204 4196 11210 4208
rect 12437 4199 12495 4205
rect 12437 4196 12449 4199
rect 11204 4168 12449 4196
rect 11204 4156 11210 4168
rect 12437 4165 12449 4168
rect 12483 4165 12495 4199
rect 12437 4159 12495 4165
rect 16206 4156 16212 4208
rect 16264 4196 16270 4208
rect 16264 4168 16528 4196
rect 16264 4156 16270 4168
rect 9861 4131 9919 4137
rect 9861 4097 9873 4131
rect 9907 4097 9919 4131
rect 9861 4091 9919 4097
rect 11241 4131 11299 4137
rect 11241 4097 11253 4131
rect 11287 4128 11299 4131
rect 12158 4128 12164 4140
rect 11287 4100 12164 4128
rect 11287 4097 11299 4100
rect 11241 4091 11299 4097
rect 3421 4063 3479 4069
rect 3421 4029 3433 4063
rect 3467 4060 3479 4063
rect 3467 4032 3832 4060
rect 3467 4029 3479 4032
rect 3421 4023 3479 4029
rect 1857 3995 1915 4001
rect 1857 3961 1869 3995
rect 1903 3992 1915 3995
rect 2225 3995 2283 4001
rect 2225 3992 2237 3995
rect 1903 3964 2237 3992
rect 1903 3961 1915 3964
rect 1857 3955 1915 3961
rect 2225 3961 2237 3964
rect 2271 3992 2283 3995
rect 2406 3992 2412 4004
rect 2271 3964 2412 3992
rect 2271 3961 2283 3964
rect 2225 3955 2283 3961
rect 2406 3952 2412 3964
rect 2464 3952 2470 4004
rect 2777 3995 2835 4001
rect 2777 3961 2789 3995
rect 2823 3992 2835 3995
rect 3602 3992 3608 4004
rect 2823 3964 3608 3992
rect 2823 3961 2835 3964
rect 2777 3955 2835 3961
rect 3602 3952 3608 3964
rect 3660 3952 3666 4004
rect 3804 3992 3832 4032
rect 5994 4020 6000 4072
rect 6052 4060 6058 4072
rect 7466 4060 7472 4072
rect 6052 4032 7472 4060
rect 6052 4020 6058 4032
rect 7466 4020 7472 4032
rect 7524 4020 7530 4072
rect 8113 4063 8171 4069
rect 8113 4029 8125 4063
rect 8159 4060 8171 4063
rect 8202 4060 8208 4072
rect 8159 4032 8208 4060
rect 8159 4029 8171 4032
rect 8113 4023 8171 4029
rect 8202 4020 8208 4032
rect 8260 4020 8266 4072
rect 8570 4020 8576 4072
rect 8628 4060 8634 4072
rect 8757 4063 8815 4069
rect 8757 4060 8769 4063
rect 8628 4032 8769 4060
rect 8628 4020 8634 4032
rect 8757 4029 8769 4032
rect 8803 4060 8815 4063
rect 9876 4060 9904 4091
rect 12158 4088 12164 4100
rect 12216 4088 12222 4140
rect 12802 4088 12808 4140
rect 12860 4128 12866 4140
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 12860 4100 12909 4128
rect 12860 4088 12866 4100
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 12897 4091 12955 4097
rect 13081 4131 13139 4137
rect 13081 4097 13093 4131
rect 13127 4128 13139 4131
rect 13262 4128 13268 4140
rect 13127 4100 13268 4128
rect 13127 4097 13139 4100
rect 13081 4091 13139 4097
rect 8803 4032 9904 4060
rect 11057 4063 11115 4069
rect 8803 4029 8815 4032
rect 8757 4023 8815 4029
rect 11057 4029 11069 4063
rect 11103 4060 11115 4063
rect 11330 4060 11336 4072
rect 11103 4032 11336 4060
rect 11103 4029 11115 4032
rect 11057 4023 11115 4029
rect 11330 4020 11336 4032
rect 11388 4020 11394 4072
rect 12912 4060 12940 4091
rect 13262 4088 13268 4100
rect 13320 4088 13326 4140
rect 13909 4131 13967 4137
rect 13909 4097 13921 4131
rect 13955 4128 13967 4131
rect 13998 4128 14004 4140
rect 13955 4100 14004 4128
rect 13955 4097 13967 4100
rect 13909 4091 13967 4097
rect 13998 4088 14004 4100
rect 14056 4128 14062 4140
rect 14553 4131 14611 4137
rect 14553 4128 14565 4131
rect 14056 4100 14565 4128
rect 14056 4088 14062 4100
rect 14553 4097 14565 4100
rect 14599 4097 14611 4131
rect 16500 4128 16528 4168
rect 16684 4137 16712 4236
rect 18506 4224 18512 4276
rect 18564 4264 18570 4276
rect 19613 4267 19671 4273
rect 19613 4264 19625 4267
rect 18564 4236 19625 4264
rect 18564 4224 18570 4236
rect 19613 4233 19625 4236
rect 19659 4264 19671 4267
rect 20530 4264 20536 4276
rect 19659 4236 20536 4264
rect 19659 4233 19671 4236
rect 19613 4227 19671 4233
rect 20530 4224 20536 4236
rect 20588 4224 20594 4276
rect 21085 4267 21143 4273
rect 21085 4233 21097 4267
rect 21131 4264 21143 4267
rect 21358 4264 21364 4276
rect 21131 4236 21364 4264
rect 21131 4233 21143 4236
rect 21085 4227 21143 4233
rect 21358 4224 21364 4236
rect 21416 4224 21422 4276
rect 19518 4196 19524 4208
rect 19352 4168 19524 4196
rect 16577 4131 16635 4137
rect 16577 4128 16589 4131
rect 16500 4100 16589 4128
rect 14553 4091 14611 4097
rect 16577 4097 16589 4100
rect 16623 4097 16635 4131
rect 16577 4091 16635 4097
rect 16669 4131 16727 4137
rect 16669 4097 16681 4131
rect 16715 4097 16727 4131
rect 16669 4091 16727 4097
rect 18693 4131 18751 4137
rect 18693 4097 18705 4131
rect 18739 4128 18751 4131
rect 18782 4128 18788 4140
rect 18739 4100 18788 4128
rect 18739 4097 18751 4100
rect 18693 4091 18751 4097
rect 18782 4088 18788 4100
rect 18840 4088 18846 4140
rect 19153 4131 19211 4137
rect 19153 4097 19165 4131
rect 19199 4128 19211 4131
rect 19352 4128 19380 4168
rect 19518 4156 19524 4168
rect 19576 4156 19582 4208
rect 20254 4128 20260 4140
rect 19199 4100 19380 4128
rect 20215 4100 20260 4128
rect 19199 4097 19211 4100
rect 19153 4091 19211 4097
rect 20254 4088 20260 4100
rect 20312 4088 20318 4140
rect 13449 4063 13507 4069
rect 13449 4060 13461 4063
rect 12912 4032 13461 4060
rect 13449 4029 13461 4032
rect 13495 4060 13507 4063
rect 13538 4060 13544 4072
rect 13495 4032 13544 4060
rect 13495 4029 13507 4032
rect 13449 4023 13507 4029
rect 13538 4020 13544 4032
rect 13596 4020 13602 4072
rect 14366 4060 14372 4072
rect 14327 4032 14372 4060
rect 14366 4020 14372 4032
rect 14424 4020 14430 4072
rect 14734 4020 14740 4072
rect 14792 4060 14798 4072
rect 15470 4060 15476 4072
rect 14792 4032 15476 4060
rect 14792 4020 14798 4032
rect 15470 4020 15476 4032
rect 15528 4060 15534 4072
rect 16485 4063 16543 4069
rect 16485 4060 16497 4063
rect 15528 4032 16497 4060
rect 15528 4020 15534 4032
rect 16485 4029 16497 4032
rect 16531 4029 16543 4063
rect 18417 4063 18475 4069
rect 18417 4060 18429 4063
rect 16485 4023 16543 4029
rect 17420 4032 18429 4060
rect 4148 3995 4206 4001
rect 4148 3992 4160 3995
rect 3804 3964 4160 3992
rect 4148 3961 4160 3964
rect 4194 3992 4206 3995
rect 4246 3992 4252 4004
rect 4194 3964 4252 3992
rect 4194 3961 4206 3964
rect 4148 3955 4206 3961
rect 4246 3952 4252 3964
rect 4304 3952 4310 4004
rect 4890 3952 4896 4004
rect 4948 3992 4954 4004
rect 5813 3995 5871 4001
rect 5813 3992 5825 3995
rect 4948 3964 5825 3992
rect 4948 3952 4954 3964
rect 5813 3961 5825 3964
rect 5859 3992 5871 3995
rect 6086 3992 6092 4004
rect 5859 3964 6092 3992
rect 5859 3961 5871 3964
rect 5813 3955 5871 3961
rect 6086 3952 6092 3964
rect 6144 3952 6150 4004
rect 8846 3992 8852 4004
rect 8220 3964 8852 3992
rect 2314 3924 2320 3936
rect 2275 3896 2320 3924
rect 2314 3884 2320 3896
rect 2372 3884 2378 3936
rect 2682 3924 2688 3936
rect 2643 3896 2688 3924
rect 2682 3884 2688 3896
rect 2740 3884 2746 3936
rect 4338 3884 4344 3936
rect 4396 3924 4402 3936
rect 5261 3927 5319 3933
rect 5261 3924 5273 3927
rect 4396 3896 5273 3924
rect 4396 3884 4402 3896
rect 5261 3893 5273 3896
rect 5307 3893 5319 3927
rect 7190 3924 7196 3936
rect 7151 3896 7196 3924
rect 5261 3887 5319 3893
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 7742 3924 7748 3936
rect 7703 3896 7748 3924
rect 7742 3884 7748 3896
rect 7800 3884 7806 3936
rect 7834 3884 7840 3936
rect 7892 3924 7898 3936
rect 8220 3933 8248 3964
rect 8846 3952 8852 3964
rect 8904 3952 8910 4004
rect 9769 3995 9827 4001
rect 9769 3992 9781 3995
rect 9140 3964 9781 3992
rect 8205 3927 8263 3933
rect 8205 3924 8217 3927
rect 7892 3896 8217 3924
rect 7892 3884 7898 3896
rect 8205 3893 8217 3896
rect 8251 3893 8263 3927
rect 8205 3887 8263 3893
rect 8938 3884 8944 3936
rect 8996 3924 9002 3936
rect 9140 3933 9168 3964
rect 9769 3961 9781 3964
rect 9815 3961 9827 3995
rect 11238 3992 11244 4004
rect 9769 3955 9827 3961
rect 9876 3964 11244 3992
rect 9125 3927 9183 3933
rect 9125 3924 9137 3927
rect 8996 3896 9137 3924
rect 8996 3884 9002 3896
rect 9125 3893 9137 3896
rect 9171 3893 9183 3927
rect 9306 3924 9312 3936
rect 9267 3896 9312 3924
rect 9125 3887 9183 3893
rect 9306 3884 9312 3896
rect 9364 3884 9370 3936
rect 9490 3884 9496 3936
rect 9548 3924 9554 3936
rect 9677 3927 9735 3933
rect 9677 3924 9689 3927
rect 9548 3896 9689 3924
rect 9548 3884 9554 3896
rect 9677 3893 9689 3896
rect 9723 3924 9735 3927
rect 9876 3924 9904 3964
rect 11238 3952 11244 3964
rect 11296 3952 11302 4004
rect 13906 3952 13912 4004
rect 13964 3992 13970 4004
rect 14461 3995 14519 4001
rect 14461 3992 14473 3995
rect 13964 3964 14473 3992
rect 13964 3952 13970 3964
rect 14461 3961 14473 3964
rect 14507 3961 14519 3995
rect 14461 3955 14519 3961
rect 15930 3952 15936 4004
rect 15988 3992 15994 4004
rect 16025 3995 16083 4001
rect 16025 3992 16037 3995
rect 15988 3964 16037 3992
rect 15988 3952 15994 3964
rect 16025 3961 16037 3964
rect 16071 3992 16083 3995
rect 16574 3992 16580 4004
rect 16071 3964 16580 3992
rect 16071 3961 16083 3964
rect 16025 3955 16083 3961
rect 16574 3952 16580 3964
rect 16632 3952 16638 4004
rect 17420 3936 17448 4032
rect 18417 4029 18429 4032
rect 18463 4029 18475 4063
rect 18417 4023 18475 4029
rect 20073 4063 20131 4069
rect 20073 4029 20085 4063
rect 20119 4060 20131 4063
rect 20162 4060 20168 4072
rect 20119 4032 20168 4060
rect 20119 4029 20131 4032
rect 20073 4023 20131 4029
rect 20162 4020 20168 4032
rect 20220 4060 20226 4072
rect 20625 4063 20683 4069
rect 20625 4060 20637 4063
rect 20220 4032 20637 4060
rect 20220 4020 20226 4032
rect 20625 4029 20637 4032
rect 20671 4060 20683 4063
rect 20990 4060 20996 4072
rect 20671 4032 20996 4060
rect 20671 4029 20683 4032
rect 20625 4023 20683 4029
rect 20990 4020 20996 4032
rect 21048 4020 21054 4072
rect 21174 4060 21180 4072
rect 21135 4032 21180 4060
rect 21174 4020 21180 4032
rect 21232 4060 21238 4072
rect 21729 4063 21787 4069
rect 21729 4060 21741 4063
rect 21232 4032 21741 4060
rect 21232 4020 21238 4032
rect 21729 4029 21741 4032
rect 21775 4029 21787 4063
rect 21729 4023 21787 4029
rect 22094 4020 22100 4072
rect 22152 4060 22158 4072
rect 22278 4060 22284 4072
rect 22152 4032 22197 4060
rect 22239 4032 22284 4060
rect 22152 4020 22158 4032
rect 22278 4020 22284 4032
rect 22336 4060 22342 4072
rect 22741 4063 22799 4069
rect 22741 4060 22753 4063
rect 22336 4032 22753 4060
rect 22336 4020 22342 4032
rect 22741 4029 22753 4032
rect 22787 4029 22799 4063
rect 22741 4023 22799 4029
rect 18509 3995 18567 4001
rect 18509 3992 18521 3995
rect 17788 3964 18521 3992
rect 17788 3936 17816 3964
rect 18509 3961 18521 3964
rect 18555 3961 18567 3995
rect 22370 3992 22376 4004
rect 18509 3955 18567 3961
rect 21376 3964 22376 3992
rect 9723 3896 9904 3924
rect 9723 3893 9735 3896
rect 9677 3887 9735 3893
rect 11974 3884 11980 3936
rect 12032 3924 12038 3936
rect 12161 3927 12219 3933
rect 12161 3924 12173 3927
rect 12032 3896 12173 3924
rect 12032 3884 12038 3896
rect 12161 3893 12173 3896
rect 12207 3924 12219 3927
rect 12805 3927 12863 3933
rect 12805 3924 12817 3927
rect 12207 3896 12817 3924
rect 12207 3893 12219 3896
rect 12161 3887 12219 3893
rect 12805 3893 12817 3896
rect 12851 3924 12863 3927
rect 13446 3924 13452 3936
rect 12851 3896 13452 3924
rect 12851 3893 12863 3896
rect 12805 3887 12863 3893
rect 13446 3884 13452 3896
rect 13504 3884 13510 3936
rect 16117 3927 16175 3933
rect 16117 3893 16129 3927
rect 16163 3924 16175 3927
rect 16482 3924 16488 3936
rect 16163 3896 16488 3924
rect 16163 3893 16175 3896
rect 16117 3887 16175 3893
rect 16482 3884 16488 3896
rect 16540 3884 16546 3936
rect 17402 3924 17408 3936
rect 17363 3896 17408 3924
rect 17402 3884 17408 3896
rect 17460 3884 17466 3936
rect 17770 3924 17776 3936
rect 17731 3896 17776 3924
rect 17770 3884 17776 3896
rect 17828 3884 17834 3936
rect 18046 3924 18052 3936
rect 18007 3896 18052 3924
rect 18046 3884 18052 3896
rect 18104 3884 18110 3936
rect 19426 3924 19432 3936
rect 19387 3896 19432 3924
rect 19426 3884 19432 3896
rect 19484 3924 19490 3936
rect 21376 3933 21404 3964
rect 22370 3952 22376 3964
rect 22428 3952 22434 4004
rect 19981 3927 20039 3933
rect 19981 3924 19993 3927
rect 19484 3896 19993 3924
rect 19484 3884 19490 3896
rect 19981 3893 19993 3896
rect 20027 3893 20039 3927
rect 19981 3887 20039 3893
rect 21361 3927 21419 3933
rect 21361 3893 21373 3927
rect 21407 3893 21419 3927
rect 21361 3887 21419 3893
rect 22094 3884 22100 3936
rect 22152 3924 22158 3936
rect 22465 3927 22523 3933
rect 22465 3924 22477 3927
rect 22152 3896 22477 3924
rect 22152 3884 22158 3896
rect 22465 3893 22477 3896
rect 22511 3893 22523 3927
rect 22465 3887 22523 3893
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1486 3680 1492 3732
rect 1544 3720 1550 3732
rect 1581 3723 1639 3729
rect 1581 3720 1593 3723
rect 1544 3692 1593 3720
rect 1544 3680 1550 3692
rect 1581 3689 1593 3692
rect 1627 3689 1639 3723
rect 1581 3683 1639 3689
rect 1596 3652 1624 3683
rect 1854 3680 1860 3732
rect 1912 3720 1918 3732
rect 2225 3723 2283 3729
rect 2225 3720 2237 3723
rect 1912 3692 2237 3720
rect 1912 3680 1918 3692
rect 2225 3689 2237 3692
rect 2271 3720 2283 3723
rect 2590 3720 2596 3732
rect 2271 3692 2596 3720
rect 2271 3689 2283 3692
rect 2225 3683 2283 3689
rect 2590 3680 2596 3692
rect 2648 3680 2654 3732
rect 2958 3680 2964 3732
rect 3016 3720 3022 3732
rect 3145 3723 3203 3729
rect 3145 3720 3157 3723
rect 3016 3692 3157 3720
rect 3016 3680 3022 3692
rect 3145 3689 3157 3692
rect 3191 3720 3203 3723
rect 3510 3720 3516 3732
rect 3191 3692 3516 3720
rect 3191 3689 3203 3692
rect 3145 3683 3203 3689
rect 3510 3680 3516 3692
rect 3568 3680 3574 3732
rect 3602 3680 3608 3732
rect 3660 3720 3666 3732
rect 3660 3692 3705 3720
rect 3660 3680 3666 3692
rect 5166 3680 5172 3732
rect 5224 3720 5230 3732
rect 5353 3723 5411 3729
rect 5353 3720 5365 3723
rect 5224 3692 5365 3720
rect 5224 3680 5230 3692
rect 5353 3689 5365 3692
rect 5399 3689 5411 3723
rect 5353 3683 5411 3689
rect 6086 3680 6092 3732
rect 6144 3720 6150 3732
rect 6917 3723 6975 3729
rect 6917 3720 6929 3723
rect 6144 3692 6929 3720
rect 6144 3680 6150 3692
rect 6917 3689 6929 3692
rect 6963 3720 6975 3723
rect 7926 3720 7932 3732
rect 6963 3692 7932 3720
rect 6963 3689 6975 3692
rect 6917 3683 6975 3689
rect 7926 3680 7932 3692
rect 7984 3680 7990 3732
rect 8021 3723 8079 3729
rect 8021 3689 8033 3723
rect 8067 3720 8079 3723
rect 8754 3720 8760 3732
rect 8067 3692 8760 3720
rect 8067 3689 8079 3692
rect 8021 3683 8079 3689
rect 8754 3680 8760 3692
rect 8812 3680 8818 3732
rect 9401 3723 9459 3729
rect 9401 3689 9413 3723
rect 9447 3720 9459 3723
rect 9490 3720 9496 3732
rect 9447 3692 9496 3720
rect 9447 3689 9459 3692
rect 9401 3683 9459 3689
rect 9490 3680 9496 3692
rect 9548 3680 9554 3732
rect 10137 3723 10195 3729
rect 10137 3689 10149 3723
rect 10183 3720 10195 3723
rect 10778 3720 10784 3732
rect 10183 3692 10784 3720
rect 10183 3689 10195 3692
rect 10137 3683 10195 3689
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 11054 3680 11060 3732
rect 11112 3720 11118 3732
rect 11241 3723 11299 3729
rect 11241 3720 11253 3723
rect 11112 3692 11253 3720
rect 11112 3680 11118 3692
rect 11241 3689 11253 3692
rect 11287 3689 11299 3723
rect 12618 3720 12624 3732
rect 11241 3683 11299 3689
rect 11992 3692 12624 3720
rect 2133 3655 2191 3661
rect 2133 3652 2145 3655
rect 1596 3624 2145 3652
rect 2133 3621 2145 3624
rect 2179 3621 2191 3655
rect 2133 3615 2191 3621
rect 2869 3655 2927 3661
rect 2869 3621 2881 3655
rect 2915 3652 2927 3655
rect 3786 3652 3792 3664
rect 2915 3624 3792 3652
rect 2915 3621 2927 3624
rect 2869 3615 2927 3621
rect 2222 3544 2228 3596
rect 2280 3584 2286 3596
rect 2884 3584 2912 3615
rect 3786 3612 3792 3624
rect 3844 3652 3850 3664
rect 5804 3655 5862 3661
rect 3844 3624 5580 3652
rect 3844 3612 3850 3624
rect 5552 3593 5580 3624
rect 5804 3621 5816 3655
rect 5850 3652 5862 3655
rect 6362 3652 6368 3664
rect 5850 3624 6368 3652
rect 5850 3621 5862 3624
rect 5804 3615 5862 3621
rect 6362 3612 6368 3624
rect 6420 3612 6426 3664
rect 7006 3612 7012 3664
rect 7064 3652 7070 3664
rect 8202 3652 8208 3664
rect 7064 3624 8208 3652
rect 7064 3612 7070 3624
rect 8202 3612 8208 3624
rect 8260 3612 8266 3664
rect 10597 3655 10655 3661
rect 10597 3621 10609 3655
rect 10643 3652 10655 3655
rect 11146 3652 11152 3664
rect 10643 3624 11152 3652
rect 10643 3621 10655 3624
rect 10597 3615 10655 3621
rect 11146 3612 11152 3624
rect 11204 3612 11210 3664
rect 11330 3612 11336 3664
rect 11388 3652 11394 3664
rect 11992 3661 12020 3692
rect 12618 3680 12624 3692
rect 12676 3680 12682 3732
rect 13078 3720 13084 3732
rect 13039 3692 13084 3720
rect 13078 3680 13084 3692
rect 13136 3720 13142 3732
rect 13633 3723 13691 3729
rect 13633 3720 13645 3723
rect 13136 3692 13645 3720
rect 13136 3680 13142 3692
rect 13633 3689 13645 3692
rect 13679 3689 13691 3723
rect 13633 3683 13691 3689
rect 13906 3680 13912 3732
rect 13964 3720 13970 3732
rect 14001 3723 14059 3729
rect 14001 3720 14013 3723
rect 13964 3692 14013 3720
rect 13964 3680 13970 3692
rect 14001 3689 14013 3692
rect 14047 3689 14059 3723
rect 14366 3720 14372 3732
rect 14327 3692 14372 3720
rect 14001 3683 14059 3689
rect 14366 3680 14372 3692
rect 14424 3680 14430 3732
rect 14642 3720 14648 3732
rect 14603 3692 14648 3720
rect 14642 3680 14648 3692
rect 14700 3680 14706 3732
rect 15930 3720 15936 3732
rect 15891 3692 15936 3720
rect 15930 3680 15936 3692
rect 15988 3680 15994 3732
rect 16577 3723 16635 3729
rect 16577 3689 16589 3723
rect 16623 3720 16635 3723
rect 16666 3720 16672 3732
rect 16623 3692 16672 3720
rect 16623 3689 16635 3692
rect 16577 3683 16635 3689
rect 16666 3680 16672 3692
rect 16724 3720 16730 3732
rect 16850 3720 16856 3732
rect 16724 3692 16856 3720
rect 16724 3680 16730 3692
rect 16850 3680 16856 3692
rect 16908 3680 16914 3732
rect 17678 3680 17684 3732
rect 17736 3720 17742 3732
rect 18049 3723 18107 3729
rect 18049 3720 18061 3723
rect 17736 3692 18061 3720
rect 17736 3680 17742 3692
rect 18049 3689 18061 3692
rect 18095 3689 18107 3723
rect 18690 3720 18696 3732
rect 18651 3692 18696 3720
rect 18049 3683 18107 3689
rect 18690 3680 18696 3692
rect 18748 3720 18754 3732
rect 20165 3723 20223 3729
rect 20165 3720 20177 3723
rect 18748 3692 20177 3720
rect 18748 3680 18754 3692
rect 20165 3689 20177 3692
rect 20211 3720 20223 3723
rect 20254 3720 20260 3732
rect 20211 3692 20260 3720
rect 20211 3689 20223 3692
rect 20165 3683 20223 3689
rect 20254 3680 20260 3692
rect 20312 3680 20318 3732
rect 11968 3655 12026 3661
rect 11968 3652 11980 3655
rect 11388 3624 11980 3652
rect 11388 3612 11394 3624
rect 11968 3621 11980 3624
rect 12014 3621 12026 3655
rect 13814 3652 13820 3664
rect 11968 3615 12026 3621
rect 13372 3624 13820 3652
rect 2280 3556 2912 3584
rect 5537 3587 5595 3593
rect 2280 3544 2286 3556
rect 5537 3553 5549 3587
rect 5583 3553 5595 3587
rect 5537 3547 5595 3553
rect 2406 3516 2412 3528
rect 2367 3488 2412 3516
rect 2406 3476 2412 3488
rect 2464 3476 2470 3528
rect 1762 3380 1768 3392
rect 1723 3352 1768 3380
rect 1762 3340 1768 3352
rect 1820 3340 1826 3392
rect 3418 3340 3424 3392
rect 3476 3380 3482 3392
rect 4430 3380 4436 3392
rect 3476 3352 4436 3380
rect 3476 3340 3482 3352
rect 4430 3340 4436 3352
rect 4488 3380 4494 3392
rect 4525 3383 4583 3389
rect 4525 3380 4537 3383
rect 4488 3352 4537 3380
rect 4488 3340 4494 3352
rect 4525 3349 4537 3352
rect 4571 3349 4583 3383
rect 4890 3380 4896 3392
rect 4851 3352 4896 3380
rect 4525 3343 4583 3349
rect 4890 3340 4896 3352
rect 4948 3340 4954 3392
rect 5552 3380 5580 3547
rect 7190 3544 7196 3596
rect 7248 3584 7254 3596
rect 7926 3584 7932 3596
rect 7248 3556 7932 3584
rect 7248 3544 7254 3556
rect 7926 3544 7932 3556
rect 7984 3584 7990 3596
rect 8389 3587 8447 3593
rect 8389 3584 8401 3587
rect 7984 3556 8401 3584
rect 7984 3544 7990 3556
rect 8389 3553 8401 3556
rect 8435 3553 8447 3587
rect 9950 3584 9956 3596
rect 9911 3556 9956 3584
rect 8389 3547 8447 3553
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 10505 3587 10563 3593
rect 10505 3553 10517 3587
rect 10551 3553 10563 3587
rect 11698 3584 11704 3596
rect 11611 3556 11704 3584
rect 10505 3547 10563 3553
rect 6914 3476 6920 3528
rect 6972 3516 6978 3528
rect 8478 3516 8484 3528
rect 6972 3488 8484 3516
rect 6972 3476 6978 3488
rect 8478 3476 8484 3488
rect 8536 3476 8542 3528
rect 8570 3476 8576 3528
rect 8628 3516 8634 3528
rect 8628 3488 8673 3516
rect 8628 3476 8634 3488
rect 7466 3408 7472 3460
rect 7524 3448 7530 3460
rect 7561 3451 7619 3457
rect 7561 3448 7573 3451
rect 7524 3420 7573 3448
rect 7524 3408 7530 3420
rect 7561 3417 7573 3420
rect 7607 3448 7619 3451
rect 8588 3448 8616 3476
rect 7607 3420 8616 3448
rect 7607 3417 7619 3420
rect 7561 3411 7619 3417
rect 7742 3380 7748 3392
rect 5552 3352 7748 3380
rect 7742 3340 7748 3352
rect 7800 3380 7806 3392
rect 7837 3383 7895 3389
rect 7837 3380 7849 3383
rect 7800 3352 7849 3380
rect 7800 3340 7806 3352
rect 7837 3349 7849 3352
rect 7883 3349 7895 3383
rect 10520 3380 10548 3547
rect 11698 3544 11704 3556
rect 11756 3584 11762 3596
rect 13372 3584 13400 3624
rect 13814 3612 13820 3624
rect 13872 3612 13878 3664
rect 14550 3612 14556 3664
rect 14608 3652 14614 3664
rect 19426 3652 19432 3664
rect 14608 3624 19432 3652
rect 14608 3612 14614 3624
rect 19426 3612 19432 3624
rect 19484 3612 19490 3664
rect 20990 3612 20996 3664
rect 21048 3652 21054 3664
rect 21048 3624 22232 3652
rect 21048 3612 21054 3624
rect 11756 3556 13400 3584
rect 11756 3544 11762 3556
rect 13446 3544 13452 3596
rect 13504 3584 13510 3596
rect 13630 3584 13636 3596
rect 13504 3556 13636 3584
rect 13504 3544 13510 3556
rect 13630 3544 13636 3556
rect 13688 3544 13694 3596
rect 14182 3584 14188 3596
rect 14143 3556 14188 3584
rect 14182 3544 14188 3556
rect 14240 3544 14246 3596
rect 15289 3587 15347 3593
rect 15289 3584 15301 3587
rect 15028 3556 15301 3584
rect 10781 3519 10839 3525
rect 10781 3485 10793 3519
rect 10827 3516 10839 3519
rect 11330 3516 11336 3528
rect 10827 3488 11336 3516
rect 10827 3485 10839 3488
rect 10781 3479 10839 3485
rect 11330 3476 11336 3488
rect 11388 3476 11394 3528
rect 13722 3380 13728 3392
rect 10520 3352 13728 3380
rect 7837 3343 7895 3349
rect 13722 3340 13728 3352
rect 13780 3340 13786 3392
rect 14734 3340 14740 3392
rect 14792 3380 14798 3392
rect 15028 3389 15056 3556
rect 15289 3553 15301 3556
rect 15335 3553 15347 3587
rect 15289 3547 15347 3553
rect 16482 3544 16488 3596
rect 16540 3584 16546 3596
rect 16936 3587 16994 3593
rect 16936 3584 16948 3587
rect 16540 3556 16948 3584
rect 16540 3544 16546 3556
rect 16936 3553 16948 3556
rect 16982 3584 16994 3587
rect 18966 3584 18972 3596
rect 16982 3556 18972 3584
rect 16982 3553 16994 3556
rect 16936 3547 16994 3553
rect 18966 3544 18972 3556
rect 19024 3544 19030 3596
rect 19518 3584 19524 3596
rect 19479 3556 19524 3584
rect 19518 3544 19524 3556
rect 19576 3544 19582 3596
rect 19613 3587 19671 3593
rect 19613 3553 19625 3587
rect 19659 3584 19671 3587
rect 20533 3587 20591 3593
rect 20533 3584 20545 3587
rect 19659 3556 20545 3584
rect 19659 3553 19671 3556
rect 19613 3547 19671 3553
rect 20533 3553 20545 3556
rect 20579 3553 20591 3587
rect 20533 3547 20591 3553
rect 21085 3587 21143 3593
rect 21085 3553 21097 3587
rect 21131 3584 21143 3587
rect 22094 3584 22100 3596
rect 21131 3556 22100 3584
rect 21131 3553 21143 3556
rect 21085 3547 21143 3553
rect 16298 3476 16304 3528
rect 16356 3516 16362 3528
rect 16669 3519 16727 3525
rect 16669 3516 16681 3519
rect 16356 3488 16681 3516
rect 16356 3476 16362 3488
rect 16669 3485 16681 3488
rect 16715 3485 16727 3519
rect 16669 3479 16727 3485
rect 18782 3476 18788 3528
rect 18840 3516 18846 3528
rect 18840 3488 19380 3516
rect 18840 3476 18846 3488
rect 15473 3451 15531 3457
rect 15473 3417 15485 3451
rect 15519 3448 15531 3451
rect 16206 3448 16212 3460
rect 15519 3420 16212 3448
rect 15519 3417 15531 3420
rect 15473 3411 15531 3417
rect 16206 3408 16212 3420
rect 16264 3408 16270 3460
rect 19150 3448 19156 3460
rect 19111 3420 19156 3448
rect 19150 3408 19156 3420
rect 19208 3408 19214 3460
rect 19352 3448 19380 3488
rect 19426 3476 19432 3528
rect 19484 3516 19490 3528
rect 19628 3516 19656 3547
rect 21468 3528 21496 3556
rect 22094 3544 22100 3556
rect 22152 3544 22158 3596
rect 22204 3593 22232 3624
rect 22189 3587 22247 3593
rect 22189 3553 22201 3587
rect 22235 3584 22247 3587
rect 22554 3584 22560 3596
rect 22235 3556 22560 3584
rect 22235 3553 22247 3556
rect 22189 3547 22247 3553
rect 22554 3544 22560 3556
rect 22612 3544 22618 3596
rect 19484 3488 19656 3516
rect 19705 3519 19763 3525
rect 19484 3476 19490 3488
rect 19705 3485 19717 3519
rect 19751 3485 19763 3519
rect 19705 3479 19763 3485
rect 19720 3448 19748 3479
rect 21450 3476 21456 3528
rect 21508 3476 21514 3528
rect 19352 3420 19748 3448
rect 15013 3383 15071 3389
rect 15013 3380 15025 3383
rect 14792 3352 15025 3380
rect 14792 3340 14798 3352
rect 15013 3349 15025 3352
rect 15059 3349 15071 3383
rect 18966 3380 18972 3392
rect 18927 3352 18972 3380
rect 15013 3343 15071 3349
rect 18966 3340 18972 3352
rect 19024 3340 19030 3392
rect 21266 3380 21272 3392
rect 21227 3352 21272 3380
rect 21266 3340 21272 3352
rect 21324 3340 21330 3392
rect 21910 3340 21916 3392
rect 21968 3380 21974 3392
rect 22373 3383 22431 3389
rect 22373 3380 22385 3383
rect 21968 3352 22385 3380
rect 21968 3340 21974 3352
rect 22373 3349 22385 3352
rect 22419 3349 22431 3383
rect 22373 3343 22431 3349
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1854 3176 1860 3188
rect 1815 3148 1860 3176
rect 1854 3136 1860 3148
rect 1912 3136 1918 3188
rect 3510 3176 3516 3188
rect 3471 3148 3516 3176
rect 3510 3136 3516 3148
rect 3568 3176 3574 3188
rect 4065 3179 4123 3185
rect 4065 3176 4077 3179
rect 3568 3148 4077 3176
rect 3568 3136 3574 3148
rect 4065 3145 4077 3148
rect 4111 3176 4123 3179
rect 4154 3176 4160 3188
rect 4111 3148 4160 3176
rect 4111 3145 4123 3148
rect 4065 3139 4123 3145
rect 4154 3136 4160 3148
rect 4212 3136 4218 3188
rect 4522 3136 4528 3188
rect 4580 3176 4586 3188
rect 4893 3179 4951 3185
rect 4893 3176 4905 3179
rect 4580 3148 4905 3176
rect 4580 3136 4586 3148
rect 4893 3145 4905 3148
rect 4939 3145 4951 3179
rect 4893 3139 4951 3145
rect 6825 3179 6883 3185
rect 6825 3145 6837 3179
rect 6871 3176 6883 3179
rect 7834 3176 7840 3188
rect 6871 3148 7840 3176
rect 6871 3145 6883 3148
rect 6825 3139 6883 3145
rect 7834 3136 7840 3148
rect 7892 3136 7898 3188
rect 8113 3179 8171 3185
rect 8113 3145 8125 3179
rect 8159 3176 8171 3179
rect 8386 3176 8392 3188
rect 8159 3148 8392 3176
rect 8159 3145 8171 3148
rect 8113 3139 8171 3145
rect 8386 3136 8392 3148
rect 8444 3136 8450 3188
rect 9769 3179 9827 3185
rect 9769 3145 9781 3179
rect 9815 3176 9827 3179
rect 9858 3176 9864 3188
rect 9815 3148 9864 3176
rect 9815 3145 9827 3148
rect 9769 3139 9827 3145
rect 9858 3136 9864 3148
rect 9916 3176 9922 3188
rect 10778 3176 10784 3188
rect 9916 3148 10784 3176
rect 9916 3136 9922 3148
rect 10778 3136 10784 3148
rect 10836 3176 10842 3188
rect 11149 3179 11207 3185
rect 11149 3176 11161 3179
rect 10836 3148 11161 3176
rect 10836 3136 10842 3148
rect 11149 3145 11161 3148
rect 11195 3176 11207 3179
rect 11330 3176 11336 3188
rect 11195 3148 11336 3176
rect 11195 3145 11207 3148
rect 11149 3139 11207 3145
rect 11330 3136 11336 3148
rect 11388 3136 11394 3188
rect 11698 3136 11704 3188
rect 11756 3176 11762 3188
rect 11793 3179 11851 3185
rect 11793 3176 11805 3179
rect 11756 3148 11805 3176
rect 11756 3136 11762 3148
rect 11793 3145 11805 3148
rect 11839 3176 11851 3179
rect 12161 3179 12219 3185
rect 12161 3176 12173 3179
rect 11839 3148 12173 3176
rect 11839 3145 11851 3148
rect 11793 3139 11851 3145
rect 12161 3145 12173 3148
rect 12207 3145 12219 3179
rect 13998 3176 14004 3188
rect 13959 3148 14004 3176
rect 12161 3139 12219 3145
rect 4430 3000 4436 3052
rect 4488 3040 4494 3052
rect 5353 3043 5411 3049
rect 5353 3040 5365 3043
rect 4488 3012 5365 3040
rect 4488 3000 4494 3012
rect 5353 3009 5365 3012
rect 5399 3009 5411 3043
rect 5353 3003 5411 3009
rect 5445 3043 5503 3049
rect 5445 3009 5457 3043
rect 5491 3009 5503 3043
rect 7466 3040 7472 3052
rect 7427 3012 7472 3040
rect 5445 3003 5503 3009
rect 2133 2975 2191 2981
rect 2133 2941 2145 2975
rect 2179 2972 2191 2975
rect 2222 2972 2228 2984
rect 2179 2944 2228 2972
rect 2179 2941 2191 2944
rect 2133 2935 2191 2941
rect 2222 2932 2228 2944
rect 2280 2932 2286 2984
rect 2406 2981 2412 2984
rect 2400 2972 2412 2981
rect 2367 2944 2412 2972
rect 2400 2935 2412 2944
rect 2406 2932 2412 2935
rect 2464 2932 2470 2984
rect 4890 2932 4896 2984
rect 4948 2972 4954 2984
rect 5460 2972 5488 3003
rect 7466 3000 7472 3012
rect 7524 3000 7530 3052
rect 7742 3000 7748 3052
rect 7800 3040 7806 3052
rect 8389 3043 8447 3049
rect 8389 3040 8401 3043
rect 7800 3012 8401 3040
rect 7800 3000 7806 3012
rect 8389 3009 8401 3012
rect 8435 3009 8447 3043
rect 12176 3040 12204 3139
rect 13998 3136 14004 3148
rect 14056 3176 14062 3188
rect 14553 3179 14611 3185
rect 14553 3176 14565 3179
rect 14056 3148 14565 3176
rect 14056 3136 14062 3148
rect 14553 3145 14565 3148
rect 14599 3145 14611 3179
rect 14553 3139 14611 3145
rect 15013 3179 15071 3185
rect 15013 3145 15025 3179
rect 15059 3176 15071 3179
rect 16298 3176 16304 3188
rect 15059 3148 16304 3176
rect 15059 3145 15071 3148
rect 15013 3139 15071 3145
rect 12621 3043 12679 3049
rect 12621 3040 12633 3043
rect 12176 3012 12633 3040
rect 8389 3003 8447 3009
rect 12621 3009 12633 3012
rect 12667 3009 12679 3043
rect 14568 3040 14596 3139
rect 15120 3120 15148 3148
rect 16298 3136 16304 3148
rect 16356 3136 16362 3188
rect 16482 3176 16488 3188
rect 16443 3148 16488 3176
rect 16482 3136 16488 3148
rect 16540 3136 16546 3188
rect 17218 3136 17224 3188
rect 17276 3176 17282 3188
rect 17405 3179 17463 3185
rect 17405 3176 17417 3179
rect 17276 3148 17417 3176
rect 17276 3136 17282 3148
rect 17405 3145 17417 3148
rect 17451 3145 17463 3179
rect 17405 3139 17463 3145
rect 15102 3068 15108 3120
rect 15160 3068 15166 3120
rect 16316 3108 16344 3136
rect 17037 3111 17095 3117
rect 17037 3108 17049 3111
rect 16316 3080 17049 3108
rect 17037 3077 17049 3080
rect 17083 3077 17095 3111
rect 17037 3071 17095 3077
rect 14568 3012 15240 3040
rect 12621 3003 12679 3009
rect 4948 2944 5488 2972
rect 4948 2932 4954 2944
rect 11054 2932 11060 2984
rect 11112 2972 11118 2984
rect 11241 2975 11299 2981
rect 11241 2972 11253 2975
rect 11112 2944 11253 2972
rect 11112 2932 11118 2944
rect 11241 2941 11253 2944
rect 11287 2941 11299 2975
rect 15102 2972 15108 2984
rect 15063 2944 15108 2972
rect 11241 2935 11299 2941
rect 15102 2932 15108 2944
rect 15160 2932 15166 2984
rect 15212 2972 15240 3012
rect 15361 2975 15419 2981
rect 15361 2972 15373 2975
rect 15212 2944 15373 2972
rect 15361 2941 15373 2944
rect 15407 2941 15419 2975
rect 15361 2935 15419 2941
rect 4246 2864 4252 2916
rect 4304 2904 4310 2916
rect 4801 2907 4859 2913
rect 4801 2904 4813 2907
rect 4304 2876 4813 2904
rect 4304 2864 4310 2876
rect 4801 2873 4813 2876
rect 4847 2904 4859 2907
rect 5258 2904 5264 2916
rect 4847 2876 5264 2904
rect 4847 2873 4859 2876
rect 4801 2867 4859 2873
rect 5258 2864 5264 2876
rect 5316 2864 5322 2916
rect 6641 2907 6699 2913
rect 6641 2873 6653 2907
rect 6687 2904 6699 2907
rect 7282 2904 7288 2916
rect 6687 2876 7288 2904
rect 6687 2873 6699 2876
rect 6641 2867 6699 2873
rect 7282 2864 7288 2876
rect 7340 2864 7346 2916
rect 8656 2907 8714 2913
rect 8656 2873 8668 2907
rect 8702 2904 8714 2907
rect 9950 2904 9956 2916
rect 8702 2876 9956 2904
rect 8702 2873 8714 2876
rect 8656 2867 8714 2873
rect 9600 2848 9628 2876
rect 9950 2864 9956 2876
rect 10008 2904 10014 2916
rect 10321 2907 10379 2913
rect 10321 2904 10333 2907
rect 10008 2876 10333 2904
rect 10008 2864 10014 2876
rect 10321 2873 10333 2876
rect 10367 2873 10379 2907
rect 10321 2867 10379 2873
rect 12888 2907 12946 2913
rect 12888 2873 12900 2907
rect 12934 2904 12946 2907
rect 13078 2904 13084 2916
rect 12934 2876 13084 2904
rect 12934 2873 12946 2876
rect 12888 2867 12946 2873
rect 13078 2864 13084 2876
rect 13136 2864 13142 2916
rect 17420 2904 17448 3139
rect 17586 3136 17592 3188
rect 17644 3176 17650 3188
rect 17773 3179 17831 3185
rect 17773 3176 17785 3179
rect 17644 3148 17785 3176
rect 17644 3136 17650 3148
rect 17773 3145 17785 3148
rect 17819 3145 17831 3179
rect 17773 3139 17831 3145
rect 18049 3179 18107 3185
rect 18049 3145 18061 3179
rect 18095 3176 18107 3179
rect 18138 3176 18144 3188
rect 18095 3148 18144 3176
rect 18095 3145 18107 3148
rect 18049 3139 18107 3145
rect 17788 2972 17816 3139
rect 18138 3136 18144 3148
rect 18196 3136 18202 3188
rect 18782 3136 18788 3188
rect 18840 3176 18846 3188
rect 19153 3179 19211 3185
rect 19153 3176 19165 3179
rect 18840 3148 19165 3176
rect 18840 3136 18846 3148
rect 19153 3145 19165 3148
rect 19199 3145 19211 3179
rect 19153 3139 19211 3145
rect 19518 3136 19524 3188
rect 19576 3176 19582 3188
rect 19613 3179 19671 3185
rect 19613 3176 19625 3179
rect 19576 3148 19625 3176
rect 19576 3136 19582 3148
rect 19613 3145 19625 3148
rect 19659 3176 19671 3179
rect 20622 3176 20628 3188
rect 19659 3148 20628 3176
rect 19659 3145 19671 3148
rect 19613 3139 19671 3145
rect 20622 3136 20628 3148
rect 20680 3136 20686 3188
rect 22554 3176 22560 3188
rect 22515 3148 22560 3176
rect 22554 3136 22560 3148
rect 22612 3136 22618 3188
rect 23842 3176 23848 3188
rect 23803 3148 23848 3176
rect 23842 3136 23848 3148
rect 23900 3136 23906 3188
rect 18693 3043 18751 3049
rect 18693 3009 18705 3043
rect 18739 3040 18751 3043
rect 18966 3040 18972 3052
rect 18739 3012 18972 3040
rect 18739 3009 18751 3012
rect 18693 3003 18751 3009
rect 18966 3000 18972 3012
rect 19024 3000 19030 3052
rect 20162 3000 20168 3052
rect 20220 3040 20226 3052
rect 20257 3043 20315 3049
rect 20257 3040 20269 3043
rect 20220 3012 20269 3040
rect 20220 3000 20226 3012
rect 20257 3009 20269 3012
rect 20303 3040 20315 3043
rect 20625 3043 20683 3049
rect 20625 3040 20637 3043
rect 20303 3012 20637 3040
rect 20303 3009 20315 3012
rect 20257 3003 20315 3009
rect 20625 3009 20637 3012
rect 20671 3009 20683 3043
rect 20625 3003 20683 3009
rect 18417 2975 18475 2981
rect 18417 2972 18429 2975
rect 17788 2944 18429 2972
rect 18417 2941 18429 2944
rect 18463 2972 18475 2975
rect 19150 2972 19156 2984
rect 18463 2944 19156 2972
rect 18463 2941 18475 2944
rect 18417 2935 18475 2941
rect 19150 2932 19156 2944
rect 19208 2932 19214 2984
rect 19242 2932 19248 2984
rect 19300 2972 19306 2984
rect 19981 2975 20039 2981
rect 19981 2972 19993 2975
rect 19300 2944 19993 2972
rect 19300 2932 19306 2944
rect 19981 2941 19993 2944
rect 20027 2972 20039 2975
rect 21361 2975 21419 2981
rect 21361 2972 21373 2975
rect 20027 2944 21373 2972
rect 20027 2941 20039 2944
rect 19981 2935 20039 2941
rect 21361 2941 21373 2944
rect 21407 2941 21419 2975
rect 21634 2972 21640 2984
rect 21595 2944 21640 2972
rect 21361 2935 21419 2941
rect 21634 2932 21640 2944
rect 21692 2972 21698 2984
rect 22189 2975 22247 2981
rect 22189 2972 22201 2975
rect 21692 2944 22201 2972
rect 21692 2932 21698 2944
rect 22189 2941 22201 2944
rect 22235 2941 22247 2975
rect 23658 2972 23664 2984
rect 23619 2944 23664 2972
rect 22189 2935 22247 2941
rect 23658 2932 23664 2944
rect 23716 2972 23722 2984
rect 24213 2975 24271 2981
rect 24213 2972 24225 2975
rect 23716 2944 24225 2972
rect 23716 2932 23722 2944
rect 24213 2941 24225 2944
rect 24259 2941 24271 2975
rect 24213 2935 24271 2941
rect 18509 2907 18567 2913
rect 18509 2904 18521 2907
rect 17420 2876 18521 2904
rect 18509 2873 18521 2876
rect 18555 2904 18567 2907
rect 18966 2904 18972 2916
rect 18555 2876 18972 2904
rect 18555 2873 18567 2876
rect 18509 2867 18567 2873
rect 18966 2864 18972 2876
rect 19024 2864 19030 2916
rect 19518 2864 19524 2916
rect 19576 2904 19582 2916
rect 19576 2876 20116 2904
rect 19576 2864 19582 2876
rect 6178 2836 6184 2848
rect 6139 2808 6184 2836
rect 6178 2796 6184 2808
rect 6236 2836 6242 2848
rect 7193 2839 7251 2845
rect 7193 2836 7205 2839
rect 6236 2808 7205 2836
rect 6236 2796 6242 2808
rect 7193 2805 7205 2808
rect 7239 2805 7251 2839
rect 7193 2799 7251 2805
rect 9582 2796 9588 2848
rect 9640 2796 9646 2848
rect 11422 2836 11428 2848
rect 11383 2808 11428 2836
rect 11422 2796 11428 2808
rect 11480 2796 11486 2848
rect 20088 2845 20116 2876
rect 20073 2839 20131 2845
rect 20073 2805 20085 2839
rect 20119 2836 20131 2839
rect 20993 2839 21051 2845
rect 20993 2836 21005 2839
rect 20119 2808 21005 2836
rect 20119 2805 20131 2808
rect 20073 2799 20131 2805
rect 20993 2805 21005 2808
rect 21039 2805 21051 2839
rect 21818 2836 21824 2848
rect 21779 2808 21824 2836
rect 20993 2799 21051 2805
rect 21818 2796 21824 2808
rect 21876 2796 21882 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 2409 2635 2467 2641
rect 2409 2601 2421 2635
rect 2455 2632 2467 2635
rect 3418 2632 3424 2644
rect 2455 2604 3424 2632
rect 2455 2601 2467 2604
rect 2409 2595 2467 2601
rect 3418 2592 3424 2604
rect 3476 2592 3482 2644
rect 3513 2635 3571 2641
rect 3513 2601 3525 2635
rect 3559 2632 3571 2635
rect 3694 2632 3700 2644
rect 3559 2604 3700 2632
rect 3559 2601 3571 2604
rect 3513 2595 3571 2601
rect 1949 2567 2007 2573
rect 1949 2533 1961 2567
rect 1995 2564 2007 2567
rect 2777 2567 2835 2573
rect 2777 2564 2789 2567
rect 1995 2536 2789 2564
rect 1995 2533 2007 2536
rect 1949 2527 2007 2533
rect 2777 2533 2789 2536
rect 2823 2564 2835 2567
rect 2866 2564 2872 2576
rect 2823 2536 2872 2564
rect 2823 2533 2835 2536
rect 2777 2527 2835 2533
rect 2866 2524 2872 2536
rect 2924 2524 2930 2576
rect 1397 2431 1455 2437
rect 1397 2397 1409 2431
rect 1443 2428 1455 2431
rect 2038 2428 2044 2440
rect 1443 2400 2044 2428
rect 1443 2397 1455 2400
rect 1397 2391 1455 2397
rect 2038 2388 2044 2400
rect 2096 2388 2102 2440
rect 2317 2431 2375 2437
rect 2317 2397 2329 2431
rect 2363 2428 2375 2431
rect 2869 2431 2927 2437
rect 2869 2428 2881 2431
rect 2363 2400 2881 2428
rect 2363 2397 2375 2400
rect 2317 2391 2375 2397
rect 2869 2397 2881 2400
rect 2915 2397 2927 2431
rect 2869 2391 2927 2397
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2428 3111 2431
rect 3528 2428 3556 2595
rect 3694 2592 3700 2604
rect 3752 2592 3758 2644
rect 3878 2632 3884 2644
rect 3839 2604 3884 2632
rect 3878 2592 3884 2604
rect 3936 2592 3942 2644
rect 5442 2632 5448 2644
rect 5403 2604 5448 2632
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 6362 2632 6368 2644
rect 6323 2604 6368 2632
rect 6362 2592 6368 2604
rect 6420 2592 6426 2644
rect 7926 2632 7932 2644
rect 7887 2604 7932 2632
rect 7926 2592 7932 2604
rect 7984 2592 7990 2644
rect 8110 2632 8116 2644
rect 8071 2604 8116 2632
rect 8110 2592 8116 2604
rect 8168 2592 8174 2644
rect 9582 2632 9588 2644
rect 9543 2604 9588 2632
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 10042 2592 10048 2644
rect 10100 2632 10106 2644
rect 10137 2635 10195 2641
rect 10137 2632 10149 2635
rect 10100 2604 10149 2632
rect 10100 2592 10106 2604
rect 10137 2601 10149 2604
rect 10183 2601 10195 2635
rect 10778 2632 10784 2644
rect 10739 2604 10784 2632
rect 10137 2595 10195 2601
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 11333 2635 11391 2641
rect 11333 2601 11345 2635
rect 11379 2632 11391 2635
rect 11974 2632 11980 2644
rect 11379 2604 11980 2632
rect 11379 2601 11391 2604
rect 11333 2595 11391 2601
rect 3896 2496 3924 2592
rect 4154 2524 4160 2576
rect 4212 2564 4218 2576
rect 4310 2567 4368 2573
rect 4310 2564 4322 2567
rect 4212 2536 4322 2564
rect 4212 2524 4218 2536
rect 4310 2533 4322 2536
rect 4356 2533 4368 2567
rect 4310 2527 4368 2533
rect 9766 2524 9772 2576
rect 9824 2564 9830 2576
rect 10229 2567 10287 2573
rect 10229 2564 10241 2567
rect 9824 2536 10241 2564
rect 9824 2524 9830 2536
rect 10229 2533 10241 2536
rect 10275 2533 10287 2567
rect 10229 2527 10287 2533
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 3896 2468 4077 2496
rect 4065 2465 4077 2468
rect 4111 2496 4123 2499
rect 5997 2499 6055 2505
rect 5997 2496 6009 2499
rect 4111 2468 6009 2496
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 5997 2465 6009 2468
rect 6043 2465 6055 2499
rect 5997 2459 6055 2465
rect 7101 2499 7159 2505
rect 7101 2465 7113 2499
rect 7147 2496 7159 2499
rect 8294 2496 8300 2508
rect 7147 2468 8300 2496
rect 7147 2465 7159 2468
rect 7101 2459 7159 2465
rect 8294 2456 8300 2468
rect 8352 2456 8358 2508
rect 8478 2496 8484 2508
rect 8439 2468 8484 2496
rect 8478 2456 8484 2468
rect 8536 2496 8542 2508
rect 9125 2499 9183 2505
rect 9125 2496 9137 2499
rect 8536 2468 9137 2496
rect 8536 2456 8542 2468
rect 9125 2465 9137 2468
rect 9171 2496 9183 2499
rect 9490 2496 9496 2508
rect 9171 2468 9496 2496
rect 9171 2465 9183 2468
rect 9125 2459 9183 2465
rect 9490 2456 9496 2468
rect 9548 2456 9554 2508
rect 11440 2505 11468 2604
rect 11974 2592 11980 2604
rect 12032 2592 12038 2644
rect 12437 2635 12495 2641
rect 12437 2601 12449 2635
rect 12483 2632 12495 2635
rect 12989 2635 13047 2641
rect 12989 2632 13001 2635
rect 12483 2604 13001 2632
rect 12483 2601 12495 2604
rect 12437 2595 12495 2601
rect 12989 2601 13001 2604
rect 13035 2632 13047 2635
rect 13446 2632 13452 2644
rect 13035 2604 13452 2632
rect 13035 2601 13047 2604
rect 12989 2595 13047 2601
rect 13446 2592 13452 2604
rect 13504 2592 13510 2644
rect 14182 2632 14188 2644
rect 14143 2604 14188 2632
rect 14182 2592 14188 2604
rect 14240 2592 14246 2644
rect 14458 2592 14464 2644
rect 14516 2632 14522 2644
rect 14734 2632 14740 2644
rect 14516 2604 14740 2632
rect 14516 2592 14522 2604
rect 14734 2592 14740 2604
rect 14792 2592 14798 2644
rect 15470 2632 15476 2644
rect 15431 2604 15476 2632
rect 15470 2592 15476 2604
rect 15528 2592 15534 2644
rect 16482 2592 16488 2644
rect 16540 2632 16546 2644
rect 16669 2635 16727 2641
rect 16669 2632 16681 2635
rect 16540 2604 16681 2632
rect 16540 2592 16546 2604
rect 16669 2601 16681 2604
rect 16715 2601 16727 2635
rect 16669 2595 16727 2601
rect 17862 2592 17868 2644
rect 17920 2632 17926 2644
rect 18049 2635 18107 2641
rect 18049 2632 18061 2635
rect 17920 2604 18061 2632
rect 17920 2592 17926 2604
rect 18049 2601 18061 2604
rect 18095 2601 18107 2635
rect 18049 2595 18107 2601
rect 18325 2635 18383 2641
rect 18325 2601 18337 2635
rect 18371 2632 18383 2635
rect 19242 2632 19248 2644
rect 18371 2604 19248 2632
rect 18371 2601 18383 2604
rect 18325 2595 18383 2601
rect 11425 2499 11483 2505
rect 11425 2465 11437 2499
rect 11471 2465 11483 2499
rect 11425 2459 11483 2465
rect 13081 2499 13139 2505
rect 13081 2465 13093 2499
rect 13127 2496 13139 2499
rect 14200 2496 14228 2592
rect 15286 2524 15292 2576
rect 15344 2564 15350 2576
rect 15933 2567 15991 2573
rect 15933 2564 15945 2567
rect 15344 2536 15945 2564
rect 15344 2524 15350 2536
rect 15933 2533 15945 2536
rect 15979 2533 15991 2567
rect 18064 2564 18092 2595
rect 19242 2592 19248 2604
rect 19300 2592 19306 2644
rect 20622 2592 20628 2644
rect 20680 2632 20686 2644
rect 20809 2635 20867 2641
rect 20809 2632 20821 2635
rect 20680 2604 20821 2632
rect 20680 2592 20686 2604
rect 20809 2601 20821 2604
rect 20855 2601 20867 2635
rect 21450 2632 21456 2644
rect 21411 2604 21456 2632
rect 20809 2595 20867 2601
rect 21450 2592 21456 2604
rect 21508 2592 21514 2644
rect 18785 2567 18843 2573
rect 18785 2564 18797 2567
rect 18064 2536 18797 2564
rect 15933 2527 15991 2533
rect 18785 2533 18797 2536
rect 18831 2533 18843 2567
rect 19429 2567 19487 2573
rect 19429 2564 19441 2567
rect 18785 2527 18843 2533
rect 18892 2536 19441 2564
rect 14277 2499 14335 2505
rect 14277 2496 14289 2499
rect 13127 2468 13768 2496
rect 14200 2468 14289 2496
rect 13127 2465 13139 2468
rect 13081 2459 13139 2465
rect 3099 2400 3556 2428
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 2884 2360 2912 2391
rect 6914 2388 6920 2440
rect 6972 2428 6978 2440
rect 7653 2431 7711 2437
rect 7653 2428 7665 2431
rect 6972 2400 7665 2428
rect 6972 2388 6978 2400
rect 7653 2397 7665 2400
rect 7699 2428 7711 2431
rect 8573 2431 8631 2437
rect 8573 2428 8585 2431
rect 7699 2400 8585 2428
rect 7699 2397 7711 2400
rect 7653 2391 7711 2397
rect 8573 2397 8585 2400
rect 8619 2428 8631 2431
rect 8662 2428 8668 2440
rect 8619 2400 8668 2428
rect 8619 2397 8631 2400
rect 8573 2391 8631 2397
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2428 8815 2431
rect 9582 2428 9588 2440
rect 8803 2400 9588 2428
rect 8803 2397 8815 2400
rect 8757 2391 8815 2397
rect 9582 2388 9588 2400
rect 9640 2388 9646 2440
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2428 10471 2431
rect 10778 2428 10784 2440
rect 10459 2400 10784 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 10778 2388 10784 2400
rect 10836 2388 10842 2440
rect 11974 2428 11980 2440
rect 11935 2400 11980 2428
rect 11974 2388 11980 2400
rect 12032 2428 12038 2440
rect 13096 2428 13124 2459
rect 13262 2428 13268 2440
rect 12032 2400 13124 2428
rect 13175 2400 13268 2428
rect 12032 2388 12038 2400
rect 13262 2388 13268 2400
rect 13320 2428 13326 2440
rect 13633 2431 13691 2437
rect 13633 2428 13645 2431
rect 13320 2400 13645 2428
rect 13320 2388 13326 2400
rect 13633 2397 13645 2400
rect 13679 2397 13691 2431
rect 13740 2428 13768 2468
rect 14277 2465 14289 2468
rect 14323 2465 14335 2499
rect 14277 2459 14335 2465
rect 14734 2456 14740 2508
rect 14792 2496 14798 2508
rect 14829 2499 14887 2505
rect 14829 2496 14841 2499
rect 14792 2468 14841 2496
rect 14792 2456 14798 2468
rect 14829 2465 14841 2468
rect 14875 2496 14887 2499
rect 15841 2499 15899 2505
rect 15841 2496 15853 2499
rect 14875 2468 15853 2496
rect 14875 2465 14887 2468
rect 14829 2459 14887 2465
rect 15841 2465 15853 2468
rect 15887 2465 15899 2499
rect 17126 2496 17132 2508
rect 17087 2468 17132 2496
rect 15841 2459 15899 2465
rect 17126 2456 17132 2468
rect 17184 2496 17190 2508
rect 17681 2499 17739 2505
rect 17681 2496 17693 2499
rect 17184 2468 17693 2496
rect 17184 2456 17190 2468
rect 17681 2465 17693 2468
rect 17727 2465 17739 2499
rect 18690 2496 18696 2508
rect 18651 2468 18696 2496
rect 17681 2459 17739 2465
rect 18690 2456 18696 2468
rect 18748 2496 18754 2508
rect 18892 2496 18920 2536
rect 19429 2533 19441 2536
rect 19475 2533 19487 2567
rect 19429 2527 19487 2533
rect 18748 2468 18920 2496
rect 18748 2456 18754 2468
rect 19334 2456 19340 2508
rect 19392 2496 19398 2508
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 19392 2468 19901 2496
rect 19392 2456 19398 2468
rect 19889 2465 19901 2468
rect 19935 2496 19947 2499
rect 20441 2499 20499 2505
rect 20441 2496 20453 2499
rect 19935 2468 20453 2496
rect 19935 2465 19947 2468
rect 19889 2459 19947 2465
rect 20441 2465 20453 2468
rect 20487 2465 20499 2499
rect 22186 2496 22192 2508
rect 22099 2468 22192 2496
rect 20441 2459 20499 2465
rect 22186 2456 22192 2468
rect 22244 2496 22250 2508
rect 22741 2499 22799 2505
rect 22741 2496 22753 2499
rect 22244 2468 22753 2496
rect 22244 2456 22250 2468
rect 22741 2465 22753 2468
rect 22787 2465 22799 2499
rect 24026 2496 24032 2508
rect 23987 2468 24032 2496
rect 22741 2459 22799 2465
rect 24026 2456 24032 2468
rect 24084 2496 24090 2508
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 24084 2468 24593 2496
rect 24084 2456 24090 2468
rect 24581 2465 24593 2468
rect 24627 2465 24639 2499
rect 24581 2459 24639 2465
rect 14918 2428 14924 2440
rect 13740 2400 14924 2428
rect 13633 2391 13691 2397
rect 14918 2388 14924 2400
rect 14976 2388 14982 2440
rect 15930 2388 15936 2440
rect 15988 2428 15994 2440
rect 16025 2431 16083 2437
rect 16025 2428 16037 2431
rect 15988 2400 16037 2428
rect 15988 2388 15994 2400
rect 16025 2397 16037 2400
rect 16071 2397 16083 2431
rect 18874 2428 18880 2440
rect 18835 2400 18880 2428
rect 16025 2391 16083 2397
rect 18874 2388 18880 2400
rect 18932 2428 18938 2440
rect 19705 2431 19763 2437
rect 19705 2428 19717 2431
rect 18932 2400 19717 2428
rect 18932 2388 18938 2400
rect 19705 2397 19717 2400
rect 19751 2397 19763 2431
rect 19705 2391 19763 2397
rect 3326 2360 3332 2372
rect 2884 2332 3332 2360
rect 3326 2320 3332 2332
rect 3384 2320 3390 2372
rect 9769 2363 9827 2369
rect 9769 2329 9781 2363
rect 9815 2360 9827 2363
rect 10870 2360 10876 2372
rect 9815 2332 10876 2360
rect 9815 2329 9827 2332
rect 9769 2323 9827 2329
rect 10870 2320 10876 2332
rect 10928 2320 10934 2372
rect 11606 2360 11612 2372
rect 11567 2332 11612 2360
rect 11606 2320 11612 2332
rect 11664 2320 11670 2372
rect 12621 2363 12679 2369
rect 12621 2329 12633 2363
rect 12667 2360 12679 2363
rect 13722 2360 13728 2372
rect 12667 2332 13728 2360
rect 12667 2329 12679 2332
rect 12621 2323 12679 2329
rect 13722 2320 13728 2332
rect 13780 2320 13786 2372
rect 14461 2363 14519 2369
rect 14461 2329 14473 2363
rect 14507 2360 14519 2363
rect 15470 2360 15476 2372
rect 14507 2332 15476 2360
rect 14507 2329 14519 2332
rect 14461 2323 14519 2329
rect 15470 2320 15476 2332
rect 15528 2320 15534 2372
rect 7282 2292 7288 2304
rect 7243 2264 7288 2292
rect 7282 2252 7288 2264
rect 7340 2252 7346 2304
rect 15286 2292 15292 2304
rect 15247 2264 15292 2292
rect 15286 2252 15292 2264
rect 15344 2252 15350 2304
rect 17310 2292 17316 2304
rect 17271 2264 17316 2292
rect 17310 2252 17316 2264
rect 17368 2252 17374 2304
rect 20070 2292 20076 2304
rect 20031 2264 20076 2292
rect 20070 2252 20076 2264
rect 20128 2252 20134 2304
rect 22373 2295 22431 2301
rect 22373 2261 22385 2295
rect 22419 2292 22431 2295
rect 24118 2292 24124 2304
rect 22419 2264 24124 2292
rect 22419 2261 22431 2264
rect 22373 2255 22431 2261
rect 24118 2252 24124 2264
rect 24176 2252 24182 2304
rect 24210 2252 24216 2304
rect 24268 2292 24274 2304
rect 24268 2264 24313 2292
rect 24268 2252 24274 2264
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 14642 1980 14648 2032
rect 14700 2020 14706 2032
rect 15746 2020 15752 2032
rect 14700 1992 15752 2020
rect 14700 1980 14706 1992
rect 15746 1980 15752 1992
rect 15804 1980 15810 2032
rect 14366 1844 14372 1896
rect 14424 1884 14430 1896
rect 18690 1884 18696 1896
rect 14424 1856 18696 1884
rect 14424 1844 14430 1856
rect 18690 1844 18696 1856
rect 18748 1844 18754 1896
<< via1 >>
rect 7564 27412 7616 27464
rect 7656 27412 7708 27464
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 1952 25304 2004 25356
rect 2412 25304 2464 25356
rect 5356 25304 5408 25356
rect 2964 25168 3016 25220
rect 2136 25100 2188 25152
rect 2320 25143 2372 25152
rect 2320 25109 2329 25143
rect 2329 25109 2363 25143
rect 2363 25109 2372 25143
rect 2320 25100 2372 25109
rect 2872 25100 2924 25152
rect 3056 25143 3108 25152
rect 3056 25109 3065 25143
rect 3065 25109 3099 25143
rect 3099 25109 3108 25143
rect 3056 25100 3108 25109
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 2412 24939 2464 24948
rect 2412 24905 2421 24939
rect 2421 24905 2455 24939
rect 2455 24905 2464 24939
rect 2412 24896 2464 24905
rect 4068 24828 4120 24880
rect 6184 24828 6236 24880
rect 2044 24803 2096 24812
rect 2044 24769 2053 24803
rect 2053 24769 2087 24803
rect 2087 24769 2096 24803
rect 2044 24760 2096 24769
rect 3056 24735 3108 24744
rect 3056 24701 3065 24735
rect 3065 24701 3099 24735
rect 3099 24701 3108 24735
rect 3056 24692 3108 24701
rect 3332 24692 3384 24744
rect 3608 24735 3660 24744
rect 3608 24701 3617 24735
rect 3617 24701 3651 24735
rect 3651 24701 3660 24735
rect 3608 24692 3660 24701
rect 12348 24692 12400 24744
rect 1400 24556 1452 24608
rect 2596 24599 2648 24608
rect 2596 24565 2605 24599
rect 2605 24565 2639 24599
rect 2639 24565 2648 24599
rect 2596 24556 2648 24565
rect 3424 24556 3476 24608
rect 6920 24556 6972 24608
rect 7840 24556 7892 24608
rect 16120 24599 16172 24608
rect 16120 24565 16129 24599
rect 16129 24565 16163 24599
rect 16163 24565 16172 24599
rect 16120 24556 16172 24565
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 1952 24395 2004 24404
rect 1952 24361 1961 24395
rect 1961 24361 1995 24395
rect 1995 24361 2004 24395
rect 1952 24352 2004 24361
rect 2780 24352 2832 24404
rect 4804 24352 4856 24404
rect 6000 24352 6052 24404
rect 7840 24395 7892 24404
rect 7840 24361 7849 24395
rect 7849 24361 7883 24395
rect 7883 24361 7892 24395
rect 7840 24352 7892 24361
rect 14280 24395 14332 24404
rect 14280 24361 14289 24395
rect 14289 24361 14323 24395
rect 14323 24361 14332 24395
rect 14280 24352 14332 24361
rect 15476 24395 15528 24404
rect 15476 24361 15485 24395
rect 15485 24361 15519 24395
rect 15519 24361 15528 24395
rect 15476 24352 15528 24361
rect 18512 24352 18564 24404
rect 18880 24395 18932 24404
rect 18880 24361 18889 24395
rect 18889 24361 18923 24395
rect 18923 24361 18932 24395
rect 18880 24352 18932 24361
rect 22468 24352 22520 24404
rect 6092 24284 6144 24336
rect 2044 24216 2096 24268
rect 3608 24216 3660 24268
rect 11796 24216 11848 24268
rect 13636 24216 13688 24268
rect 15292 24259 15344 24268
rect 15292 24225 15301 24259
rect 15301 24225 15335 24259
rect 15335 24225 15344 24259
rect 15292 24216 15344 24225
rect 16856 24216 16908 24268
rect 17408 24216 17460 24268
rect 18972 24216 19024 24268
rect 20812 24216 20864 24268
rect 3332 24148 3384 24200
rect 4528 24191 4580 24200
rect 4528 24157 4537 24191
rect 4537 24157 4571 24191
rect 4571 24157 4580 24191
rect 4528 24148 4580 24157
rect 2504 24080 2556 24132
rect 7380 24148 7432 24200
rect 8116 24191 8168 24200
rect 1676 24012 1728 24064
rect 2688 24012 2740 24064
rect 3332 24012 3384 24064
rect 5356 24080 5408 24132
rect 8116 24157 8125 24191
rect 8125 24157 8159 24191
rect 8159 24157 8168 24191
rect 8116 24148 8168 24157
rect 9036 24080 9088 24132
rect 12256 24123 12308 24132
rect 12256 24089 12265 24123
rect 12265 24089 12299 24123
rect 12299 24089 12308 24123
rect 12256 24080 12308 24089
rect 17776 24123 17828 24132
rect 17776 24089 17785 24123
rect 17785 24089 17819 24123
rect 17819 24089 17828 24123
rect 17776 24080 17828 24089
rect 4068 24055 4120 24064
rect 4068 24021 4077 24055
rect 4077 24021 4111 24055
rect 4111 24021 4120 24055
rect 4068 24012 4120 24021
rect 5448 24012 5500 24064
rect 6920 24055 6972 24064
rect 6920 24021 6929 24055
rect 6929 24021 6963 24055
rect 6963 24021 6972 24055
rect 6920 24012 6972 24021
rect 7380 24055 7432 24064
rect 7380 24021 7389 24055
rect 7389 24021 7423 24055
rect 7423 24021 7432 24055
rect 7380 24012 7432 24021
rect 7472 24055 7524 24064
rect 7472 24021 7481 24055
rect 7481 24021 7515 24055
rect 7515 24021 7524 24055
rect 7472 24012 7524 24021
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 2044 23851 2096 23860
rect 2044 23817 2053 23851
rect 2053 23817 2087 23851
rect 2087 23817 2096 23851
rect 2044 23808 2096 23817
rect 2320 23808 2372 23860
rect 2780 23808 2832 23860
rect 3148 23851 3200 23860
rect 3148 23817 3157 23851
rect 3157 23817 3191 23851
rect 3191 23817 3200 23851
rect 3148 23808 3200 23817
rect 3240 23808 3292 23860
rect 3608 23851 3660 23860
rect 3608 23817 3617 23851
rect 3617 23817 3651 23851
rect 3651 23817 3660 23851
rect 3608 23808 3660 23817
rect 5356 23808 5408 23860
rect 6000 23851 6052 23860
rect 6000 23817 6009 23851
rect 6009 23817 6043 23851
rect 6043 23817 6052 23851
rect 6000 23808 6052 23817
rect 6092 23808 6144 23860
rect 6276 23808 6328 23860
rect 9036 23808 9088 23860
rect 10784 23808 10836 23860
rect 12624 23851 12676 23860
rect 12624 23817 12633 23851
rect 12633 23817 12667 23851
rect 12667 23817 12676 23851
rect 12624 23808 12676 23817
rect 2688 23715 2740 23724
rect 2688 23681 2697 23715
rect 2697 23681 2731 23715
rect 2731 23681 2740 23715
rect 2688 23672 2740 23681
rect 2504 23647 2556 23656
rect 2504 23613 2513 23647
rect 2513 23613 2547 23647
rect 2547 23613 2556 23647
rect 2504 23604 2556 23613
rect 2596 23647 2648 23656
rect 2596 23613 2605 23647
rect 2605 23613 2639 23647
rect 2639 23613 2648 23647
rect 2596 23604 2648 23613
rect 4160 23604 4212 23656
rect 6368 23604 6420 23656
rect 6920 23604 6972 23656
rect 9864 23604 9916 23656
rect 10784 23604 10836 23656
rect 13360 23808 13412 23860
rect 14004 23783 14056 23792
rect 14004 23749 14013 23783
rect 14013 23749 14047 23783
rect 14047 23749 14056 23783
rect 14004 23740 14056 23749
rect 15660 23808 15712 23860
rect 17040 23851 17092 23860
rect 17040 23817 17049 23851
rect 17049 23817 17083 23851
rect 17083 23817 17092 23851
rect 17040 23808 17092 23817
rect 18236 23851 18288 23860
rect 18236 23817 18245 23851
rect 18245 23817 18279 23851
rect 18279 23817 18288 23851
rect 18236 23808 18288 23817
rect 19708 23808 19760 23860
rect 21364 23851 21416 23860
rect 21364 23817 21373 23851
rect 21373 23817 21407 23851
rect 21407 23817 21416 23851
rect 21364 23808 21416 23817
rect 25320 23808 25372 23860
rect 15108 23783 15160 23792
rect 15108 23749 15117 23783
rect 15117 23749 15151 23783
rect 15151 23749 15160 23783
rect 15108 23740 15160 23749
rect 3976 23579 4028 23588
rect 3976 23545 3985 23579
rect 3985 23545 4019 23579
rect 4019 23545 4028 23579
rect 3976 23536 4028 23545
rect 4896 23536 4948 23588
rect 7380 23536 7432 23588
rect 7564 23536 7616 23588
rect 7932 23536 7984 23588
rect 3332 23468 3384 23520
rect 6828 23468 6880 23520
rect 8116 23468 8168 23520
rect 11428 23511 11480 23520
rect 11428 23477 11437 23511
rect 11437 23477 11471 23511
rect 11471 23477 11480 23511
rect 11428 23468 11480 23477
rect 11796 23468 11848 23520
rect 13636 23511 13688 23520
rect 13636 23477 13645 23511
rect 13645 23477 13679 23511
rect 13679 23477 13688 23511
rect 13636 23468 13688 23477
rect 14556 23468 14608 23520
rect 17408 23604 17460 23656
rect 19432 23647 19484 23656
rect 15292 23468 15344 23520
rect 16856 23468 16908 23520
rect 19432 23613 19441 23647
rect 19441 23613 19475 23647
rect 19475 23613 19484 23647
rect 19432 23604 19484 23613
rect 21088 23604 21140 23656
rect 23480 23604 23532 23656
rect 17592 23468 17644 23520
rect 18604 23511 18656 23520
rect 18604 23477 18613 23511
rect 18613 23477 18647 23511
rect 18647 23477 18656 23511
rect 18604 23468 18656 23477
rect 18972 23511 19024 23520
rect 18972 23477 18981 23511
rect 18981 23477 19015 23511
rect 19015 23477 19024 23511
rect 18972 23468 19024 23477
rect 20812 23468 20864 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 2320 23264 2372 23316
rect 2780 23264 2832 23316
rect 3976 23264 4028 23316
rect 5264 23307 5316 23316
rect 5264 23273 5273 23307
rect 5273 23273 5307 23307
rect 5307 23273 5316 23307
rect 5264 23264 5316 23273
rect 9864 23307 9916 23316
rect 9864 23273 9873 23307
rect 9873 23273 9907 23307
rect 9907 23273 9916 23307
rect 9864 23264 9916 23273
rect 13636 23264 13688 23316
rect 14832 23264 14884 23316
rect 17224 23307 17276 23316
rect 17224 23273 17233 23307
rect 17233 23273 17267 23307
rect 17267 23273 17276 23307
rect 17224 23264 17276 23273
rect 18972 23264 19024 23316
rect 21088 23307 21140 23316
rect 21088 23273 21097 23307
rect 21097 23273 21131 23307
rect 21131 23273 21140 23307
rect 21088 23264 21140 23273
rect 23480 23264 23532 23316
rect 2228 23196 2280 23248
rect 2596 23196 2648 23248
rect 3608 23196 3660 23248
rect 4160 23196 4212 23248
rect 6368 23196 6420 23248
rect 6828 23196 6880 23248
rect 5172 23171 5224 23180
rect 5172 23137 5181 23171
rect 5181 23137 5215 23171
rect 5215 23137 5224 23171
rect 5172 23128 5224 23137
rect 7380 23128 7432 23180
rect 9772 23128 9824 23180
rect 12164 23128 12216 23180
rect 15384 23128 15436 23180
rect 17040 23171 17092 23180
rect 17040 23137 17049 23171
rect 17049 23137 17083 23171
rect 17083 23137 17092 23171
rect 17040 23128 17092 23137
rect 18236 23128 18288 23180
rect 20904 23171 20956 23180
rect 20904 23137 20913 23171
rect 20913 23137 20947 23171
rect 20947 23137 20956 23171
rect 20904 23128 20956 23137
rect 22192 23171 22244 23180
rect 22192 23137 22201 23171
rect 22201 23137 22235 23171
rect 22235 23137 22244 23171
rect 22192 23128 22244 23137
rect 2044 23060 2096 23112
rect 2688 23060 2740 23112
rect 4160 23060 4212 23112
rect 4436 23060 4488 23112
rect 6368 23103 6420 23112
rect 4896 22992 4948 23044
rect 6368 23069 6377 23103
rect 6377 23069 6411 23103
rect 6411 23069 6420 23103
rect 6368 23060 6420 23069
rect 13544 23103 13596 23112
rect 13544 23069 13553 23103
rect 13553 23069 13587 23103
rect 13587 23069 13596 23103
rect 13544 23060 13596 23069
rect 1860 22924 1912 22976
rect 2872 22967 2924 22976
rect 2872 22933 2881 22967
rect 2881 22933 2915 22967
rect 2915 22933 2924 22967
rect 2872 22924 2924 22933
rect 3332 22924 3384 22976
rect 4804 22967 4856 22976
rect 4804 22933 4813 22967
rect 4813 22933 4847 22967
rect 4847 22933 4856 22967
rect 4804 22924 4856 22933
rect 8484 22967 8536 22976
rect 8484 22933 8493 22967
rect 8493 22933 8527 22967
rect 8527 22933 8536 22967
rect 8484 22924 8536 22933
rect 14464 22967 14516 22976
rect 14464 22933 14473 22967
rect 14473 22933 14507 22967
rect 14507 22933 14516 22967
rect 14464 22924 14516 22933
rect 15476 22967 15528 22976
rect 15476 22933 15485 22967
rect 15485 22933 15519 22967
rect 15519 22933 15528 22967
rect 15476 22924 15528 22933
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 2136 22720 2188 22772
rect 2228 22584 2280 22636
rect 3608 22720 3660 22772
rect 4896 22763 4948 22772
rect 4896 22729 4905 22763
rect 4905 22729 4939 22763
rect 4939 22729 4948 22763
rect 4896 22720 4948 22729
rect 6184 22763 6236 22772
rect 6184 22729 6193 22763
rect 6193 22729 6227 22763
rect 6227 22729 6236 22763
rect 6184 22720 6236 22729
rect 6368 22720 6420 22772
rect 7472 22720 7524 22772
rect 16396 22720 16448 22772
rect 16856 22763 16908 22772
rect 16856 22729 16865 22763
rect 16865 22729 16899 22763
rect 16899 22729 16908 22763
rect 16856 22720 16908 22729
rect 17040 22720 17092 22772
rect 20904 22763 20956 22772
rect 20904 22729 20913 22763
rect 20913 22729 20947 22763
rect 20947 22729 20956 22763
rect 20904 22720 20956 22729
rect 8392 22695 8444 22704
rect 8392 22661 8401 22695
rect 8401 22661 8435 22695
rect 8435 22661 8444 22695
rect 8392 22652 8444 22661
rect 12900 22695 12952 22704
rect 12900 22661 12909 22695
rect 12909 22661 12943 22695
rect 12943 22661 12952 22695
rect 12900 22652 12952 22661
rect 5632 22627 5684 22636
rect 5632 22593 5641 22627
rect 5641 22593 5675 22627
rect 5675 22593 5684 22627
rect 5632 22584 5684 22593
rect 5540 22559 5592 22568
rect 1584 22423 1636 22432
rect 1584 22389 1593 22423
rect 1593 22389 1627 22423
rect 1627 22389 1636 22423
rect 1584 22380 1636 22389
rect 2872 22380 2924 22432
rect 5540 22525 5549 22559
rect 5549 22525 5583 22559
rect 5583 22525 5592 22559
rect 5540 22516 5592 22525
rect 7380 22584 7432 22636
rect 8484 22584 8536 22636
rect 14464 22584 14516 22636
rect 6828 22516 6880 22568
rect 12164 22559 12216 22568
rect 12164 22525 12173 22559
rect 12173 22525 12207 22559
rect 12207 22525 12216 22559
rect 12164 22516 12216 22525
rect 12900 22516 12952 22568
rect 15476 22516 15528 22568
rect 6368 22448 6420 22500
rect 3792 22380 3844 22432
rect 5172 22423 5224 22432
rect 5172 22389 5181 22423
rect 5181 22389 5215 22423
rect 5215 22389 5224 22423
rect 5172 22380 5224 22389
rect 6184 22380 6236 22432
rect 7472 22380 7524 22432
rect 8116 22380 8168 22432
rect 14556 22448 14608 22500
rect 14832 22448 14884 22500
rect 19340 22516 19392 22568
rect 22192 22559 22244 22568
rect 22192 22525 22201 22559
rect 22201 22525 22235 22559
rect 22235 22525 22244 22559
rect 22192 22516 22244 22525
rect 18512 22448 18564 22500
rect 8484 22380 8536 22432
rect 9772 22423 9824 22432
rect 9772 22389 9781 22423
rect 9781 22389 9815 22423
rect 9815 22389 9824 22423
rect 9772 22380 9824 22389
rect 9864 22380 9916 22432
rect 14004 22423 14056 22432
rect 14004 22389 14013 22423
rect 14013 22389 14047 22423
rect 14047 22389 14056 22423
rect 14004 22380 14056 22389
rect 14740 22380 14792 22432
rect 15384 22423 15436 22432
rect 15384 22389 15393 22423
rect 15393 22389 15427 22423
rect 15427 22389 15436 22423
rect 15384 22380 15436 22389
rect 18236 22423 18288 22432
rect 18236 22389 18245 22423
rect 18245 22389 18279 22423
rect 18279 22389 18288 22423
rect 18236 22380 18288 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 1952 22176 2004 22228
rect 2228 22108 2280 22160
rect 5172 22176 5224 22228
rect 5632 22219 5684 22228
rect 5632 22185 5641 22219
rect 5641 22185 5675 22219
rect 5675 22185 5684 22219
rect 5632 22176 5684 22185
rect 4436 22151 4488 22160
rect 1676 22083 1728 22092
rect 1676 22049 1710 22083
rect 1710 22049 1728 22083
rect 1676 22040 1728 22049
rect 2412 22040 2464 22092
rect 3976 22040 4028 22092
rect 4436 22117 4445 22151
rect 4445 22117 4479 22151
rect 4479 22117 4488 22151
rect 4436 22108 4488 22117
rect 5540 22108 5592 22160
rect 4528 22083 4580 22092
rect 1768 21836 1820 21888
rect 2688 21904 2740 21956
rect 4528 22049 4537 22083
rect 4537 22049 4571 22083
rect 4571 22049 4580 22083
rect 4528 22040 4580 22049
rect 6828 22176 6880 22228
rect 8484 22219 8536 22228
rect 8484 22185 8493 22219
rect 8493 22185 8527 22219
rect 8527 22185 8536 22219
rect 8484 22176 8536 22185
rect 13820 22219 13872 22228
rect 13820 22185 13829 22219
rect 13829 22185 13863 22219
rect 13863 22185 13872 22219
rect 13820 22176 13872 22185
rect 14004 22176 14056 22228
rect 14372 22176 14424 22228
rect 14740 22176 14792 22228
rect 6644 22040 6696 22092
rect 6828 22083 6880 22092
rect 6828 22049 6837 22083
rect 6837 22049 6871 22083
rect 6871 22049 6880 22083
rect 6828 22040 6880 22049
rect 8760 22040 8812 22092
rect 10876 22083 10928 22092
rect 10876 22049 10885 22083
rect 10885 22049 10919 22083
rect 10919 22049 10928 22083
rect 10876 22040 10928 22049
rect 13268 22040 13320 22092
rect 14464 22040 14516 22092
rect 15568 22083 15620 22092
rect 15568 22049 15591 22083
rect 15591 22049 15620 22083
rect 15568 22040 15620 22049
rect 4620 22015 4672 22024
rect 4620 21981 4629 22015
rect 4629 21981 4663 22015
rect 4663 21981 4672 22015
rect 4620 21972 4672 21981
rect 10968 22015 11020 22024
rect 6736 21904 6788 21956
rect 10968 21981 10977 22015
rect 10977 21981 11011 22015
rect 11011 21981 11020 22015
rect 10968 21972 11020 21981
rect 11060 21972 11112 22024
rect 13636 21972 13688 22024
rect 14096 21972 14148 22024
rect 9680 21904 9732 21956
rect 13728 21904 13780 21956
rect 16672 21947 16724 21956
rect 16672 21913 16681 21947
rect 16681 21913 16715 21947
rect 16715 21913 16724 21947
rect 16672 21904 16724 21913
rect 7380 21879 7432 21888
rect 7380 21845 7389 21879
rect 7389 21845 7423 21879
rect 7423 21845 7432 21879
rect 7380 21836 7432 21845
rect 7656 21836 7708 21888
rect 9496 21836 9548 21888
rect 11060 21836 11112 21888
rect 11152 21836 11204 21888
rect 13268 21879 13320 21888
rect 13268 21845 13277 21879
rect 13277 21845 13311 21879
rect 13311 21845 13320 21879
rect 13268 21836 13320 21845
rect 13360 21879 13412 21888
rect 13360 21845 13369 21879
rect 13369 21845 13403 21879
rect 13403 21845 13412 21879
rect 13360 21836 13412 21845
rect 14556 21836 14608 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 4712 21675 4764 21684
rect 4712 21641 4721 21675
rect 4721 21641 4755 21675
rect 4755 21641 4764 21675
rect 4712 21632 4764 21641
rect 6828 21632 6880 21684
rect 10876 21632 10928 21684
rect 13636 21632 13688 21684
rect 15568 21675 15620 21684
rect 15568 21641 15577 21675
rect 15577 21641 15611 21675
rect 15611 21641 15620 21675
rect 15568 21632 15620 21641
rect 10968 21564 11020 21616
rect 2228 21539 2280 21548
rect 2228 21505 2237 21539
rect 2237 21505 2271 21539
rect 2271 21505 2280 21539
rect 2228 21496 2280 21505
rect 5172 21496 5224 21548
rect 8208 21496 8260 21548
rect 9496 21539 9548 21548
rect 9496 21505 9505 21539
rect 9505 21505 9539 21539
rect 9539 21505 9548 21539
rect 9496 21496 9548 21505
rect 11428 21539 11480 21548
rect 11428 21505 11437 21539
rect 11437 21505 11471 21539
rect 11471 21505 11480 21539
rect 11428 21496 11480 21505
rect 12992 21539 13044 21548
rect 12992 21505 13001 21539
rect 13001 21505 13035 21539
rect 13035 21505 13044 21539
rect 12992 21496 13044 21505
rect 5356 21428 5408 21480
rect 2320 21360 2372 21412
rect 2688 21360 2740 21412
rect 4712 21360 4764 21412
rect 8116 21428 8168 21480
rect 11244 21471 11296 21480
rect 11244 21437 11253 21471
rect 11253 21437 11287 21471
rect 11287 21437 11296 21471
rect 11244 21428 11296 21437
rect 3608 21335 3660 21344
rect 3608 21301 3617 21335
rect 3617 21301 3651 21335
rect 3651 21301 3660 21335
rect 3608 21292 3660 21301
rect 4988 21292 5040 21344
rect 6000 21360 6052 21412
rect 6644 21360 6696 21412
rect 6828 21360 6880 21412
rect 7564 21360 7616 21412
rect 8852 21403 8904 21412
rect 8852 21369 8861 21403
rect 8861 21369 8895 21403
rect 8895 21369 8904 21403
rect 8852 21360 8904 21369
rect 13084 21360 13136 21412
rect 14556 21360 14608 21412
rect 7012 21335 7064 21344
rect 7012 21301 7021 21335
rect 7021 21301 7055 21335
rect 7055 21301 7064 21335
rect 7012 21292 7064 21301
rect 7656 21292 7708 21344
rect 8944 21335 8996 21344
rect 8944 21301 8953 21335
rect 8953 21301 8987 21335
rect 8987 21301 8996 21335
rect 8944 21292 8996 21301
rect 9036 21292 9088 21344
rect 10968 21292 11020 21344
rect 11152 21335 11204 21344
rect 11152 21301 11161 21335
rect 11161 21301 11195 21335
rect 11195 21301 11204 21335
rect 11152 21292 11204 21301
rect 12164 21292 12216 21344
rect 13636 21292 13688 21344
rect 14096 21335 14148 21344
rect 14096 21301 14105 21335
rect 14105 21301 14139 21335
rect 14139 21301 14148 21335
rect 14096 21292 14148 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 2320 21131 2372 21140
rect 2320 21097 2329 21131
rect 2329 21097 2363 21131
rect 2363 21097 2372 21131
rect 2320 21088 2372 21097
rect 4528 21088 4580 21140
rect 5540 21088 5592 21140
rect 2872 21063 2924 21072
rect 2872 21029 2881 21063
rect 2881 21029 2915 21063
rect 2915 21029 2924 21063
rect 2872 21020 2924 21029
rect 3792 21063 3844 21072
rect 3792 21029 3801 21063
rect 3801 21029 3835 21063
rect 3835 21029 3844 21063
rect 3792 21020 3844 21029
rect 6184 21088 6236 21140
rect 7564 21088 7616 21140
rect 7840 21131 7892 21140
rect 7840 21097 7849 21131
rect 7849 21097 7883 21131
rect 7883 21097 7892 21131
rect 7840 21088 7892 21097
rect 9036 21131 9088 21140
rect 9036 21097 9045 21131
rect 9045 21097 9079 21131
rect 9079 21097 9088 21131
rect 9036 21088 9088 21097
rect 11428 21088 11480 21140
rect 12992 21088 13044 21140
rect 13268 21088 13320 21140
rect 15568 21131 15620 21140
rect 15568 21097 15577 21131
rect 15577 21097 15611 21131
rect 15611 21097 15620 21131
rect 15568 21088 15620 21097
rect 6000 21020 6052 21072
rect 9496 21020 9548 21072
rect 13728 21020 13780 21072
rect 14004 21020 14056 21072
rect 1400 20995 1452 21004
rect 1400 20961 1409 20995
rect 1409 20961 1443 20995
rect 1443 20961 1452 20995
rect 1400 20952 1452 20961
rect 2780 20995 2832 21004
rect 2780 20961 2789 20995
rect 2789 20961 2823 20995
rect 2823 20961 2832 20995
rect 2780 20952 2832 20961
rect 4988 20952 5040 21004
rect 5448 20952 5500 21004
rect 2964 20927 3016 20936
rect 2964 20893 2973 20927
rect 2973 20893 3007 20927
rect 3007 20893 3016 20927
rect 2964 20884 3016 20893
rect 3608 20884 3660 20936
rect 4896 20927 4948 20936
rect 1676 20816 1728 20868
rect 3792 20816 3844 20868
rect 1584 20791 1636 20800
rect 1584 20757 1593 20791
rect 1593 20757 1627 20791
rect 1627 20757 1636 20791
rect 1584 20748 1636 20757
rect 4160 20748 4212 20800
rect 4896 20893 4905 20927
rect 4905 20893 4939 20927
rect 4939 20893 4948 20927
rect 4896 20884 4948 20893
rect 6368 20927 6420 20936
rect 6368 20893 6377 20927
rect 6377 20893 6411 20927
rect 6411 20893 6420 20927
rect 6368 20884 6420 20893
rect 6092 20816 6144 20868
rect 7196 20884 7248 20936
rect 13360 20952 13412 21004
rect 14740 20952 14792 21004
rect 14004 20927 14056 20936
rect 5172 20748 5224 20800
rect 5540 20748 5592 20800
rect 7380 20748 7432 20800
rect 8116 20748 8168 20800
rect 8392 20748 8444 20800
rect 14004 20893 14013 20927
rect 14013 20893 14047 20927
rect 14047 20893 14056 20927
rect 14004 20884 14056 20893
rect 14464 20884 14516 20936
rect 9864 20748 9916 20800
rect 10876 20748 10928 20800
rect 12348 20791 12400 20800
rect 12348 20757 12357 20791
rect 12357 20757 12391 20791
rect 12391 20757 12400 20791
rect 12348 20748 12400 20757
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 2964 20544 3016 20596
rect 5540 20587 5592 20596
rect 5540 20553 5549 20587
rect 5549 20553 5583 20587
rect 5583 20553 5592 20587
rect 5540 20544 5592 20553
rect 6184 20544 6236 20596
rect 7196 20587 7248 20596
rect 7196 20553 7205 20587
rect 7205 20553 7239 20587
rect 7239 20553 7248 20587
rect 7196 20544 7248 20553
rect 8300 20544 8352 20596
rect 11060 20544 11112 20596
rect 14004 20544 14056 20596
rect 14740 20587 14792 20596
rect 14740 20553 14749 20587
rect 14749 20553 14783 20587
rect 14783 20553 14792 20587
rect 14740 20544 14792 20553
rect 15568 20544 15620 20596
rect 2412 20340 2464 20392
rect 2688 20340 2740 20392
rect 4068 20340 4120 20392
rect 7380 20383 7432 20392
rect 7380 20349 7389 20383
rect 7389 20349 7423 20383
rect 7423 20349 7432 20383
rect 7380 20340 7432 20349
rect 2872 20315 2924 20324
rect 2872 20281 2881 20315
rect 2881 20281 2915 20315
rect 2915 20281 2924 20315
rect 2872 20272 2924 20281
rect 3608 20272 3660 20324
rect 8392 20272 8444 20324
rect 12532 20340 12584 20392
rect 12992 20340 13044 20392
rect 1400 20204 1452 20256
rect 2964 20204 3016 20256
rect 3240 20204 3292 20256
rect 3792 20204 3844 20256
rect 4436 20204 4488 20256
rect 4896 20204 4948 20256
rect 6184 20204 6236 20256
rect 6368 20204 6420 20256
rect 9864 20204 9916 20256
rect 11888 20247 11940 20256
rect 11888 20213 11897 20247
rect 11897 20213 11931 20247
rect 11931 20213 11940 20247
rect 11888 20204 11940 20213
rect 12716 20204 12768 20256
rect 13544 20204 13596 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 1952 20043 2004 20052
rect 1952 20009 1961 20043
rect 1961 20009 1995 20043
rect 1995 20009 2004 20043
rect 1952 20000 2004 20009
rect 2412 20043 2464 20052
rect 2412 20009 2421 20043
rect 2421 20009 2455 20043
rect 2455 20009 2464 20043
rect 2412 20000 2464 20009
rect 3608 20000 3660 20052
rect 6000 20043 6052 20052
rect 6000 20009 6009 20043
rect 6009 20009 6043 20043
rect 6043 20009 6052 20043
rect 6000 20000 6052 20009
rect 6920 20043 6972 20052
rect 6920 20009 6929 20043
rect 6929 20009 6963 20043
rect 6963 20009 6972 20043
rect 6920 20000 6972 20009
rect 9036 20000 9088 20052
rect 9680 20000 9732 20052
rect 11060 20000 11112 20052
rect 11888 20000 11940 20052
rect 12992 20000 13044 20052
rect 4436 19932 4488 19984
rect 10876 19932 10928 19984
rect 12532 19975 12584 19984
rect 12532 19941 12541 19975
rect 12541 19941 12575 19975
rect 12575 19941 12584 19975
rect 12532 19932 12584 19941
rect 14740 19932 14792 19984
rect 15292 19932 15344 19984
rect 2320 19864 2372 19916
rect 4068 19907 4120 19916
rect 4068 19873 4084 19907
rect 4084 19873 4118 19907
rect 4118 19873 4120 19907
rect 4068 19864 4120 19873
rect 15108 19864 15160 19916
rect 7012 19839 7064 19848
rect 7012 19805 7021 19839
rect 7021 19805 7055 19839
rect 7055 19805 7064 19839
rect 7012 19796 7064 19805
rect 3056 19771 3108 19780
rect 3056 19737 3065 19771
rect 3065 19737 3099 19771
rect 3099 19737 3108 19771
rect 3056 19728 3108 19737
rect 6092 19728 6144 19780
rect 6644 19728 6696 19780
rect 7380 19796 7432 19848
rect 9864 19796 9916 19848
rect 10508 19839 10560 19848
rect 10508 19805 10517 19839
rect 10517 19805 10551 19839
rect 10551 19805 10560 19839
rect 10508 19796 10560 19805
rect 13820 19796 13872 19848
rect 12532 19728 12584 19780
rect 14464 19728 14516 19780
rect 1584 19703 1636 19712
rect 1584 19669 1593 19703
rect 1593 19669 1627 19703
rect 1627 19669 1636 19703
rect 1584 19660 1636 19669
rect 3792 19703 3844 19712
rect 3792 19669 3801 19703
rect 3801 19669 3835 19703
rect 3835 19669 3844 19703
rect 3792 19660 3844 19669
rect 4436 19660 4488 19712
rect 5540 19660 5592 19712
rect 7932 19660 7984 19712
rect 8392 19703 8444 19712
rect 8392 19669 8401 19703
rect 8401 19669 8435 19703
rect 8435 19669 8444 19703
rect 8392 19660 8444 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 2320 19499 2372 19508
rect 2320 19465 2329 19499
rect 2329 19465 2363 19499
rect 2363 19465 2372 19499
rect 2320 19456 2372 19465
rect 6092 19456 6144 19508
rect 6920 19456 6972 19508
rect 7196 19456 7248 19508
rect 7656 19499 7708 19508
rect 7656 19465 7665 19499
rect 7665 19465 7699 19499
rect 7699 19465 7708 19499
rect 7656 19456 7708 19465
rect 9956 19456 10008 19508
rect 10508 19456 10560 19508
rect 12624 19499 12676 19508
rect 7472 19388 7524 19440
rect 7840 19388 7892 19440
rect 12624 19465 12633 19499
rect 12633 19465 12667 19499
rect 12667 19465 12676 19499
rect 12624 19456 12676 19465
rect 12716 19388 12768 19440
rect 1308 19320 1360 19372
rect 2320 19320 2372 19372
rect 4436 19363 4488 19372
rect 2964 19252 3016 19304
rect 1492 19116 1544 19168
rect 2044 19159 2096 19168
rect 2044 19125 2053 19159
rect 2053 19125 2087 19159
rect 2087 19125 2096 19159
rect 2044 19116 2096 19125
rect 2688 19159 2740 19168
rect 2688 19125 2697 19159
rect 2697 19125 2731 19159
rect 2731 19125 2740 19159
rect 2688 19116 2740 19125
rect 4436 19329 4445 19363
rect 4445 19329 4479 19363
rect 4479 19329 4488 19363
rect 4436 19320 4488 19329
rect 4160 19295 4212 19304
rect 4160 19261 4169 19295
rect 4169 19261 4203 19295
rect 4203 19261 4212 19295
rect 4160 19252 4212 19261
rect 5356 19295 5408 19304
rect 5356 19261 5365 19295
rect 5365 19261 5399 19295
rect 5399 19261 5408 19295
rect 5356 19252 5408 19261
rect 5448 19252 5500 19304
rect 7012 19320 7064 19372
rect 7564 19320 7616 19372
rect 8392 19320 8444 19372
rect 8944 19252 8996 19304
rect 9680 19295 9732 19304
rect 9680 19261 9689 19295
rect 9689 19261 9723 19295
rect 9723 19261 9732 19295
rect 9680 19252 9732 19261
rect 4896 19227 4948 19236
rect 4896 19193 4905 19227
rect 4905 19193 4939 19227
rect 4939 19193 4948 19227
rect 4896 19184 4948 19193
rect 7012 19184 7064 19236
rect 7932 19184 7984 19236
rect 10876 19320 10928 19372
rect 11428 19363 11480 19372
rect 11428 19329 11437 19363
rect 11437 19329 11471 19363
rect 11471 19329 11480 19363
rect 11428 19320 11480 19329
rect 14556 19456 14608 19508
rect 11060 19252 11112 19304
rect 12164 19252 12216 19304
rect 12992 19295 13044 19304
rect 12992 19261 13001 19295
rect 13001 19261 13035 19295
rect 13035 19261 13044 19295
rect 12992 19252 13044 19261
rect 14096 19295 14148 19304
rect 12716 19184 12768 19236
rect 14096 19261 14105 19295
rect 14105 19261 14139 19295
rect 14139 19261 14148 19295
rect 14096 19252 14148 19261
rect 14464 19295 14516 19304
rect 14464 19261 14498 19295
rect 14498 19261 14516 19295
rect 14464 19252 14516 19261
rect 3240 19116 3292 19168
rect 3884 19116 3936 19168
rect 4252 19159 4304 19168
rect 4252 19125 4261 19159
rect 4261 19125 4295 19159
rect 4295 19125 4304 19159
rect 4252 19116 4304 19125
rect 5080 19116 5132 19168
rect 8208 19116 8260 19168
rect 8392 19116 8444 19168
rect 9220 19159 9272 19168
rect 9220 19125 9229 19159
rect 9229 19125 9263 19159
rect 9263 19125 9272 19159
rect 9220 19116 9272 19125
rect 10784 19159 10836 19168
rect 10784 19125 10793 19159
rect 10793 19125 10827 19159
rect 10827 19125 10836 19159
rect 10784 19116 10836 19125
rect 13084 19159 13136 19168
rect 13084 19125 13093 19159
rect 13093 19125 13127 19159
rect 13127 19125 13136 19159
rect 13084 19116 13136 19125
rect 13820 19116 13872 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 4252 18912 4304 18964
rect 5172 18912 5224 18964
rect 7012 18912 7064 18964
rect 7380 18912 7432 18964
rect 8024 18912 8076 18964
rect 8944 18912 8996 18964
rect 10876 18912 10928 18964
rect 11152 18912 11204 18964
rect 14464 18912 14516 18964
rect 15292 18955 15344 18964
rect 15292 18921 15301 18955
rect 15301 18921 15335 18955
rect 15335 18921 15344 18955
rect 15292 18912 15344 18921
rect 4160 18844 4212 18896
rect 4436 18844 4488 18896
rect 1676 18776 1728 18828
rect 3976 18776 4028 18828
rect 5448 18844 5500 18896
rect 9496 18844 9548 18896
rect 9956 18844 10008 18896
rect 11060 18844 11112 18896
rect 13084 18844 13136 18896
rect 6460 18819 6512 18828
rect 6460 18785 6469 18819
rect 6469 18785 6503 18819
rect 6503 18785 6512 18819
rect 6460 18776 6512 18785
rect 6736 18776 6788 18828
rect 7472 18776 7524 18828
rect 10048 18819 10100 18828
rect 3792 18708 3844 18760
rect 5080 18751 5132 18760
rect 5080 18717 5089 18751
rect 5089 18717 5123 18751
rect 5123 18717 5132 18751
rect 5080 18708 5132 18717
rect 6644 18751 6696 18760
rect 6644 18717 6653 18751
rect 6653 18717 6687 18751
rect 6687 18717 6696 18751
rect 6644 18708 6696 18717
rect 7840 18708 7892 18760
rect 6920 18640 6972 18692
rect 10048 18785 10057 18819
rect 10057 18785 10091 18819
rect 10091 18785 10100 18819
rect 10048 18776 10100 18785
rect 11428 18776 11480 18828
rect 12808 18776 12860 18828
rect 13544 18776 13596 18828
rect 8208 18751 8260 18760
rect 8208 18717 8217 18751
rect 8217 18717 8251 18751
rect 8251 18717 8260 18751
rect 8208 18708 8260 18717
rect 9956 18708 10008 18760
rect 10140 18751 10192 18760
rect 10140 18717 10149 18751
rect 10149 18717 10183 18751
rect 10183 18717 10192 18751
rect 10140 18708 10192 18717
rect 10416 18708 10468 18760
rect 12716 18751 12768 18760
rect 12716 18717 12725 18751
rect 12725 18717 12759 18751
rect 12759 18717 12768 18751
rect 12716 18708 12768 18717
rect 11060 18640 11112 18692
rect 1400 18572 1452 18624
rect 2044 18615 2096 18624
rect 2044 18581 2053 18615
rect 2053 18581 2087 18615
rect 2087 18581 2096 18615
rect 2044 18572 2096 18581
rect 2688 18615 2740 18624
rect 2688 18581 2697 18615
rect 2697 18581 2731 18615
rect 2731 18581 2740 18615
rect 2688 18572 2740 18581
rect 3240 18572 3292 18624
rect 6368 18572 6420 18624
rect 7656 18615 7708 18624
rect 7656 18581 7665 18615
rect 7665 18581 7699 18615
rect 7699 18581 7708 18615
rect 7656 18572 7708 18581
rect 9404 18615 9456 18624
rect 9404 18581 9413 18615
rect 9413 18581 9447 18615
rect 9447 18581 9456 18615
rect 9404 18572 9456 18581
rect 9864 18572 9916 18624
rect 12532 18615 12584 18624
rect 12532 18581 12541 18615
rect 12541 18581 12575 18615
rect 12575 18581 12584 18615
rect 12532 18572 12584 18581
rect 15384 18572 15436 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 3792 18411 3844 18420
rect 3792 18377 3801 18411
rect 3801 18377 3835 18411
rect 3835 18377 3844 18411
rect 3792 18368 3844 18377
rect 8392 18411 8444 18420
rect 8392 18377 8401 18411
rect 8401 18377 8435 18411
rect 8435 18377 8444 18411
rect 8392 18368 8444 18377
rect 9312 18368 9364 18420
rect 10416 18368 10468 18420
rect 13084 18368 13136 18420
rect 2596 18300 2648 18352
rect 8024 18300 8076 18352
rect 12716 18300 12768 18352
rect 3240 18275 3292 18284
rect 3240 18241 3249 18275
rect 3249 18241 3283 18275
rect 3283 18241 3292 18275
rect 3240 18232 3292 18241
rect 7012 18275 7064 18284
rect 7012 18241 7021 18275
rect 7021 18241 7055 18275
rect 7055 18241 7064 18275
rect 7012 18232 7064 18241
rect 2044 18164 2096 18216
rect 2964 18164 3016 18216
rect 3148 18207 3200 18216
rect 3148 18173 3157 18207
rect 3157 18173 3191 18207
rect 3191 18173 3200 18207
rect 3148 18164 3200 18173
rect 4068 18164 4120 18216
rect 4896 18164 4948 18216
rect 9496 18207 9548 18216
rect 9496 18173 9505 18207
rect 9505 18173 9539 18207
rect 9539 18173 9548 18207
rect 9496 18164 9548 18173
rect 13728 18232 13780 18284
rect 14464 18232 14516 18284
rect 10048 18164 10100 18216
rect 11060 18164 11112 18216
rect 12532 18164 12584 18216
rect 4436 18096 4488 18148
rect 5080 18096 5132 18148
rect 6460 18096 6512 18148
rect 7380 18096 7432 18148
rect 9404 18096 9456 18148
rect 12256 18139 12308 18148
rect 12256 18105 12265 18139
rect 12265 18105 12299 18139
rect 12299 18105 12308 18139
rect 12256 18096 12308 18105
rect 14188 18096 14240 18148
rect 14648 18096 14700 18148
rect 1584 18071 1636 18080
rect 1584 18037 1593 18071
rect 1593 18037 1627 18071
rect 1627 18037 1636 18071
rect 1584 18028 1636 18037
rect 2964 18028 3016 18080
rect 3424 18028 3476 18080
rect 5540 18028 5592 18080
rect 6736 18028 6788 18080
rect 7104 18028 7156 18080
rect 10876 18071 10928 18080
rect 10876 18037 10885 18071
rect 10885 18037 10919 18071
rect 10919 18037 10928 18071
rect 10876 18028 10928 18037
rect 11520 18028 11572 18080
rect 14004 18028 14056 18080
rect 14740 18028 14792 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 1676 17824 1728 17876
rect 3424 17824 3476 17876
rect 4620 17824 4672 17876
rect 5172 17867 5224 17876
rect 5172 17833 5181 17867
rect 5181 17833 5215 17867
rect 5215 17833 5224 17867
rect 5172 17824 5224 17833
rect 6828 17824 6880 17876
rect 9036 17824 9088 17876
rect 9496 17867 9548 17876
rect 9496 17833 9505 17867
rect 9505 17833 9539 17867
rect 9539 17833 9548 17867
rect 9496 17824 9548 17833
rect 14464 17867 14516 17876
rect 14464 17833 14473 17867
rect 14473 17833 14507 17867
rect 14507 17833 14516 17867
rect 14464 17824 14516 17833
rect 3976 17756 4028 17808
rect 6644 17756 6696 17808
rect 9956 17799 10008 17808
rect 9956 17765 9965 17799
rect 9965 17765 9999 17799
rect 9999 17765 10008 17799
rect 9956 17756 10008 17765
rect 5172 17688 5224 17740
rect 6736 17688 6788 17740
rect 8208 17688 8260 17740
rect 10784 17688 10836 17740
rect 11428 17731 11480 17740
rect 11428 17697 11462 17731
rect 11462 17697 11480 17731
rect 11428 17688 11480 17697
rect 2596 17620 2648 17672
rect 3056 17663 3108 17672
rect 3056 17629 3065 17663
rect 3065 17629 3099 17663
rect 3099 17629 3108 17663
rect 3056 17620 3108 17629
rect 4896 17620 4948 17672
rect 5540 17620 5592 17672
rect 2228 17552 2280 17604
rect 1952 17527 2004 17536
rect 1952 17493 1961 17527
rect 1961 17493 1995 17527
rect 1995 17493 2004 17527
rect 1952 17484 2004 17493
rect 2688 17484 2740 17536
rect 3608 17484 3660 17536
rect 6184 17484 6236 17536
rect 6460 17527 6512 17536
rect 6460 17493 6469 17527
rect 6469 17493 6503 17527
rect 6503 17493 6512 17527
rect 6460 17484 6512 17493
rect 7840 17620 7892 17672
rect 9496 17620 9548 17672
rect 11152 17663 11204 17672
rect 11152 17629 11161 17663
rect 11161 17629 11195 17663
rect 11195 17629 11204 17663
rect 11152 17620 11204 17629
rect 10324 17595 10376 17604
rect 10324 17561 10333 17595
rect 10333 17561 10367 17595
rect 10367 17561 10376 17595
rect 10324 17552 10376 17561
rect 6828 17484 6880 17536
rect 7380 17484 7432 17536
rect 12532 17527 12584 17536
rect 12532 17493 12541 17527
rect 12541 17493 12575 17527
rect 12575 17493 12584 17527
rect 12532 17484 12584 17493
rect 13176 17484 13228 17536
rect 14188 17484 14240 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 2228 17280 2280 17332
rect 4620 17280 4672 17332
rect 5172 17280 5224 17332
rect 6460 17280 6512 17332
rect 6828 17280 6880 17332
rect 8576 17323 8628 17332
rect 8576 17289 8585 17323
rect 8585 17289 8619 17323
rect 8619 17289 8628 17323
rect 8576 17280 8628 17289
rect 10784 17280 10836 17332
rect 12808 17323 12860 17332
rect 12808 17289 12817 17323
rect 12817 17289 12851 17323
rect 12851 17289 12860 17323
rect 12808 17280 12860 17289
rect 13912 17280 13964 17332
rect 5632 17255 5684 17264
rect 5632 17221 5641 17255
rect 5641 17221 5675 17255
rect 5675 17221 5684 17255
rect 5632 17212 5684 17221
rect 11152 17212 11204 17264
rect 11796 17212 11848 17264
rect 12716 17212 12768 17264
rect 7380 17187 7432 17196
rect 7380 17153 7389 17187
rect 7389 17153 7423 17187
rect 7423 17153 7432 17187
rect 7380 17144 7432 17153
rect 8208 17144 8260 17196
rect 9496 17144 9548 17196
rect 10876 17144 10928 17196
rect 12348 17144 12400 17196
rect 1952 17076 2004 17128
rect 2872 17119 2924 17128
rect 2872 17085 2881 17119
rect 2881 17085 2915 17119
rect 2915 17085 2924 17119
rect 2872 17076 2924 17085
rect 4068 17076 4120 17128
rect 5540 17076 5592 17128
rect 6460 17076 6512 17128
rect 8668 17076 8720 17128
rect 9220 17076 9272 17128
rect 10048 17076 10100 17128
rect 3240 17051 3292 17060
rect 3240 17017 3274 17051
rect 3274 17017 3292 17051
rect 3240 17008 3292 17017
rect 7656 17008 7708 17060
rect 8208 17008 8260 17060
rect 9956 17008 10008 17060
rect 13176 17008 13228 17060
rect 1492 16940 1544 16992
rect 3056 16940 3108 16992
rect 4712 16940 4764 16992
rect 6828 16983 6880 16992
rect 6828 16949 6837 16983
rect 6837 16949 6871 16983
rect 6871 16949 6880 16983
rect 6828 16940 6880 16949
rect 11428 16940 11480 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1676 16736 1728 16788
rect 2596 16736 2648 16788
rect 3424 16779 3476 16788
rect 3424 16745 3433 16779
rect 3433 16745 3467 16779
rect 3467 16745 3476 16779
rect 3424 16736 3476 16745
rect 3976 16736 4028 16788
rect 6736 16779 6788 16788
rect 6736 16745 6745 16779
rect 6745 16745 6779 16779
rect 6779 16745 6788 16779
rect 6736 16736 6788 16745
rect 8208 16779 8260 16788
rect 5172 16668 5224 16720
rect 8208 16745 8217 16779
rect 8217 16745 8251 16779
rect 8251 16745 8260 16779
rect 8208 16736 8260 16745
rect 8668 16779 8720 16788
rect 8668 16745 8677 16779
rect 8677 16745 8711 16779
rect 8711 16745 8720 16779
rect 8668 16736 8720 16745
rect 9496 16779 9548 16788
rect 9496 16745 9505 16779
rect 9505 16745 9539 16779
rect 9539 16745 9548 16779
rect 9496 16736 9548 16745
rect 9956 16779 10008 16788
rect 9956 16745 9965 16779
rect 9965 16745 9999 16779
rect 9999 16745 10008 16779
rect 9956 16736 10008 16745
rect 10048 16736 10100 16788
rect 10692 16736 10744 16788
rect 7472 16668 7524 16720
rect 7748 16668 7800 16720
rect 2228 16600 2280 16652
rect 2044 16532 2096 16584
rect 3240 16600 3292 16652
rect 4712 16575 4764 16584
rect 4712 16541 4721 16575
rect 4721 16541 4755 16575
rect 4755 16541 4764 16575
rect 4712 16532 4764 16541
rect 2412 16464 2464 16516
rect 2596 16464 2648 16516
rect 4896 16600 4948 16652
rect 4988 16600 5040 16652
rect 5540 16643 5592 16652
rect 5540 16609 5549 16643
rect 5549 16609 5583 16643
rect 5583 16609 5592 16643
rect 5540 16600 5592 16609
rect 6000 16643 6052 16652
rect 6000 16609 6009 16643
rect 6009 16609 6043 16643
rect 6043 16609 6052 16643
rect 6000 16600 6052 16609
rect 7840 16600 7892 16652
rect 11704 16736 11756 16788
rect 13084 16779 13136 16788
rect 13084 16745 13093 16779
rect 13093 16745 13127 16779
rect 13127 16745 13136 16779
rect 13084 16736 13136 16745
rect 15752 16779 15804 16788
rect 15752 16745 15761 16779
rect 15761 16745 15795 16779
rect 15795 16745 15804 16779
rect 15752 16736 15804 16745
rect 6092 16575 6144 16584
rect 6092 16541 6101 16575
rect 6101 16541 6135 16575
rect 6135 16541 6144 16575
rect 6092 16532 6144 16541
rect 7748 16575 7800 16584
rect 5356 16464 5408 16516
rect 7748 16541 7757 16575
rect 7757 16541 7791 16575
rect 7791 16541 7800 16575
rect 7748 16532 7800 16541
rect 10232 16532 10284 16584
rect 12532 16668 12584 16720
rect 11796 16600 11848 16652
rect 11980 16643 12032 16652
rect 11980 16609 12014 16643
rect 12014 16609 12032 16643
rect 11980 16600 12032 16609
rect 15660 16643 15712 16652
rect 15660 16609 15669 16643
rect 15669 16609 15703 16643
rect 15703 16609 15712 16643
rect 15660 16600 15712 16609
rect 15936 16575 15988 16584
rect 9404 16464 9456 16516
rect 15936 16541 15945 16575
rect 15945 16541 15979 16575
rect 15979 16541 15988 16575
rect 15936 16532 15988 16541
rect 1768 16396 1820 16448
rect 2780 16396 2832 16448
rect 4068 16439 4120 16448
rect 4068 16405 4077 16439
rect 4077 16405 4111 16439
rect 4111 16405 4120 16439
rect 4068 16396 4120 16405
rect 6920 16396 6972 16448
rect 10140 16396 10192 16448
rect 10692 16396 10744 16448
rect 15292 16439 15344 16448
rect 15292 16405 15301 16439
rect 15301 16405 15335 16439
rect 15335 16405 15344 16439
rect 15292 16396 15344 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 1860 16192 1912 16244
rect 4712 16235 4764 16244
rect 4712 16201 4721 16235
rect 4721 16201 4755 16235
rect 4755 16201 4764 16235
rect 4712 16192 4764 16201
rect 5356 16192 5408 16244
rect 6092 16192 6144 16244
rect 6644 16235 6696 16244
rect 6644 16201 6653 16235
rect 6653 16201 6687 16235
rect 6687 16201 6696 16235
rect 6644 16192 6696 16201
rect 9312 16192 9364 16244
rect 10048 16192 10100 16244
rect 11796 16235 11848 16244
rect 11796 16201 11805 16235
rect 11805 16201 11839 16235
rect 11839 16201 11848 16235
rect 11796 16192 11848 16201
rect 15936 16192 15988 16244
rect 6736 16124 6788 16176
rect 15752 16124 15804 16176
rect 16120 16124 16172 16176
rect 2320 16099 2372 16108
rect 2320 16065 2329 16099
rect 2329 16065 2363 16099
rect 2363 16065 2372 16099
rect 2320 16056 2372 16065
rect 1768 15988 1820 16040
rect 9036 16056 9088 16108
rect 6644 15988 6696 16040
rect 7932 15988 7984 16040
rect 8576 15988 8628 16040
rect 15660 16031 15712 16040
rect 1584 15895 1636 15904
rect 1584 15861 1593 15895
rect 1593 15861 1627 15895
rect 1627 15861 1636 15895
rect 1584 15852 1636 15861
rect 2872 15920 2924 15972
rect 6092 15920 6144 15972
rect 6920 15920 6972 15972
rect 10140 15963 10192 15972
rect 10140 15929 10174 15963
rect 10174 15929 10192 15963
rect 10140 15920 10192 15929
rect 11796 15920 11848 15972
rect 15660 15997 15669 16031
rect 15669 15997 15703 16031
rect 15703 15997 15712 16031
rect 15660 15988 15712 15997
rect 13912 15920 13964 15972
rect 4528 15852 4580 15904
rect 5724 15895 5776 15904
rect 5724 15861 5733 15895
rect 5733 15861 5767 15895
rect 5767 15861 5776 15895
rect 5724 15852 5776 15861
rect 7840 15852 7892 15904
rect 11336 15852 11388 15904
rect 11980 15852 12032 15904
rect 15108 15895 15160 15904
rect 15108 15861 15117 15895
rect 15117 15861 15151 15895
rect 15151 15861 15160 15895
rect 15108 15852 15160 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2044 15648 2096 15700
rect 2228 15691 2280 15700
rect 2228 15657 2237 15691
rect 2237 15657 2271 15691
rect 2271 15657 2280 15691
rect 2228 15648 2280 15657
rect 2412 15691 2464 15700
rect 2412 15657 2421 15691
rect 2421 15657 2455 15691
rect 2455 15657 2464 15691
rect 2412 15648 2464 15657
rect 4068 15648 4120 15700
rect 4252 15691 4304 15700
rect 4252 15657 4261 15691
rect 4261 15657 4295 15691
rect 4295 15657 4304 15691
rect 4252 15648 4304 15657
rect 5172 15648 5224 15700
rect 5540 15648 5592 15700
rect 5724 15648 5776 15700
rect 7748 15648 7800 15700
rect 9404 15691 9456 15700
rect 9404 15657 9413 15691
rect 9413 15657 9447 15691
rect 9447 15657 9456 15691
rect 9404 15648 9456 15657
rect 10140 15648 10192 15700
rect 10784 15691 10836 15700
rect 10784 15657 10793 15691
rect 10793 15657 10827 15691
rect 10827 15657 10836 15691
rect 10784 15648 10836 15657
rect 11244 15691 11296 15700
rect 11244 15657 11253 15691
rect 11253 15657 11287 15691
rect 11287 15657 11296 15691
rect 11244 15648 11296 15657
rect 12440 15648 12492 15700
rect 12808 15691 12860 15700
rect 12808 15657 12817 15691
rect 12817 15657 12851 15691
rect 12851 15657 12860 15691
rect 12808 15648 12860 15657
rect 3976 15580 4028 15632
rect 6000 15580 6052 15632
rect 7932 15580 7984 15632
rect 11520 15580 11572 15632
rect 13912 15648 13964 15700
rect 14556 15648 14608 15700
rect 15752 15623 15804 15632
rect 2044 15512 2096 15564
rect 2688 15512 2740 15564
rect 3792 15512 3844 15564
rect 4068 15555 4120 15564
rect 4068 15521 4077 15555
rect 4077 15521 4111 15555
rect 4111 15521 4120 15555
rect 4068 15512 4120 15521
rect 6644 15512 6696 15564
rect 12716 15555 12768 15564
rect 12716 15521 12725 15555
rect 12725 15521 12759 15555
rect 12759 15521 12768 15555
rect 12716 15512 12768 15521
rect 2596 15444 2648 15496
rect 4528 15444 4580 15496
rect 9864 15444 9916 15496
rect 10968 15444 11020 15496
rect 11428 15487 11480 15496
rect 11428 15453 11437 15487
rect 11437 15453 11471 15487
rect 11471 15453 11480 15487
rect 11428 15444 11480 15453
rect 13084 15444 13136 15496
rect 15752 15589 15761 15623
rect 15761 15589 15795 15623
rect 15795 15589 15804 15623
rect 15752 15580 15804 15589
rect 13820 15512 13872 15564
rect 15936 15512 15988 15564
rect 15844 15487 15896 15496
rect 15844 15453 15853 15487
rect 15853 15453 15887 15487
rect 15887 15453 15896 15487
rect 15844 15444 15896 15453
rect 3240 15376 3292 15428
rect 5448 15308 5500 15360
rect 10048 15419 10100 15428
rect 10048 15385 10057 15419
rect 10057 15385 10091 15419
rect 10091 15385 10100 15419
rect 10048 15376 10100 15385
rect 6920 15308 6972 15360
rect 14464 15308 14516 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2596 15104 2648 15156
rect 4068 15104 4120 15156
rect 6092 15104 6144 15156
rect 6920 15104 6972 15156
rect 8576 15147 8628 15156
rect 8576 15113 8585 15147
rect 8585 15113 8619 15147
rect 8619 15113 8628 15147
rect 8576 15104 8628 15113
rect 10140 15147 10192 15156
rect 10140 15113 10149 15147
rect 10149 15113 10183 15147
rect 10183 15113 10192 15147
rect 10140 15104 10192 15113
rect 10968 15104 11020 15156
rect 11244 15147 11296 15156
rect 11244 15113 11253 15147
rect 11253 15113 11287 15147
rect 11287 15113 11296 15147
rect 11244 15104 11296 15113
rect 11520 15147 11572 15156
rect 11520 15113 11529 15147
rect 11529 15113 11563 15147
rect 11563 15113 11572 15147
rect 11520 15104 11572 15113
rect 12348 15104 12400 15156
rect 13084 15147 13136 15156
rect 13084 15113 13093 15147
rect 13093 15113 13127 15147
rect 13127 15113 13136 15147
rect 13084 15104 13136 15113
rect 3976 15036 4028 15088
rect 6644 15036 6696 15088
rect 2872 15011 2924 15020
rect 2872 14977 2881 15011
rect 2881 14977 2915 15011
rect 2915 14977 2924 15011
rect 2872 14968 2924 14977
rect 3516 14968 3568 15020
rect 6000 14968 6052 15020
rect 7932 14968 7984 15020
rect 1400 14943 1452 14952
rect 1400 14909 1409 14943
rect 1409 14909 1443 14943
rect 1443 14909 1452 14943
rect 1400 14900 1452 14909
rect 3976 14943 4028 14952
rect 3976 14909 3985 14943
rect 3985 14909 4019 14943
rect 4019 14909 4028 14943
rect 3976 14900 4028 14909
rect 5540 14943 5592 14952
rect 5540 14909 5549 14943
rect 5549 14909 5583 14943
rect 5583 14909 5592 14943
rect 5540 14900 5592 14909
rect 2780 14875 2832 14884
rect 2780 14841 2789 14875
rect 2789 14841 2823 14875
rect 2823 14841 2832 14875
rect 2780 14832 2832 14841
rect 6460 14900 6512 14952
rect 7196 14943 7248 14952
rect 7196 14909 7205 14943
rect 7205 14909 7239 14943
rect 7239 14909 7248 14943
rect 7196 14900 7248 14909
rect 8576 14900 8628 14952
rect 9312 14900 9364 14952
rect 12808 14900 12860 14952
rect 12716 14875 12768 14884
rect 12716 14841 12725 14875
rect 12725 14841 12759 14875
rect 12759 14841 12768 14875
rect 12716 14832 12768 14841
rect 13268 14832 13320 14884
rect 13452 14875 13504 14884
rect 13452 14841 13461 14875
rect 13461 14841 13495 14875
rect 13495 14841 13504 14875
rect 13452 14832 13504 14841
rect 14096 14832 14148 14884
rect 3148 14764 3200 14816
rect 3516 14807 3568 14816
rect 3516 14773 3525 14807
rect 3525 14773 3559 14807
rect 3559 14773 3568 14807
rect 3516 14764 3568 14773
rect 4160 14807 4212 14816
rect 4160 14773 4169 14807
rect 4169 14773 4203 14807
rect 4203 14773 4212 14807
rect 4160 14764 4212 14773
rect 5448 14764 5500 14816
rect 6828 14807 6880 14816
rect 6828 14773 6837 14807
rect 6837 14773 6871 14807
rect 6871 14773 6880 14807
rect 6828 14764 6880 14773
rect 7288 14807 7340 14816
rect 7288 14773 7297 14807
rect 7297 14773 7331 14807
rect 7331 14773 7340 14807
rect 7288 14764 7340 14773
rect 14924 14764 14976 14816
rect 15384 14764 15436 14816
rect 15752 14764 15804 14816
rect 15936 14764 15988 14816
rect 16672 14807 16724 14816
rect 16672 14773 16681 14807
rect 16681 14773 16715 14807
rect 16715 14773 16724 14807
rect 16672 14764 16724 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2228 14560 2280 14612
rect 3792 14603 3844 14612
rect 3792 14569 3801 14603
rect 3801 14569 3835 14603
rect 3835 14569 3844 14603
rect 3792 14560 3844 14569
rect 6000 14603 6052 14612
rect 6000 14569 6009 14603
rect 6009 14569 6043 14603
rect 6043 14569 6052 14603
rect 6000 14560 6052 14569
rect 7932 14603 7984 14612
rect 7932 14569 7941 14603
rect 7941 14569 7975 14603
rect 7975 14569 7984 14603
rect 7932 14560 7984 14569
rect 9680 14603 9732 14612
rect 9680 14569 9689 14603
rect 9689 14569 9723 14603
rect 9723 14569 9732 14603
rect 9680 14560 9732 14569
rect 14096 14603 14148 14612
rect 14096 14569 14105 14603
rect 14105 14569 14139 14603
rect 14139 14569 14148 14603
rect 14096 14560 14148 14569
rect 14924 14603 14976 14612
rect 14924 14569 14933 14603
rect 14933 14569 14967 14603
rect 14967 14569 14976 14603
rect 14924 14560 14976 14569
rect 2872 14535 2924 14544
rect 2872 14501 2881 14535
rect 2881 14501 2915 14535
rect 2915 14501 2924 14535
rect 2872 14492 2924 14501
rect 4528 14492 4580 14544
rect 15568 14492 15620 14544
rect 15844 14492 15896 14544
rect 2412 14424 2464 14476
rect 2504 14356 2556 14408
rect 3240 14424 3292 14476
rect 4068 14467 4120 14476
rect 4068 14433 4077 14467
rect 4077 14433 4111 14467
rect 4111 14433 4120 14467
rect 4068 14424 4120 14433
rect 3516 14399 3568 14408
rect 3516 14365 3525 14399
rect 3525 14365 3559 14399
rect 3559 14365 3568 14399
rect 3516 14356 3568 14365
rect 3792 14356 3844 14408
rect 6184 14424 6236 14476
rect 10324 14424 10376 14476
rect 12256 14424 12308 14476
rect 13544 14424 13596 14476
rect 15660 14467 15712 14476
rect 15660 14433 15669 14467
rect 15669 14433 15703 14467
rect 15703 14433 15712 14467
rect 15660 14424 15712 14433
rect 6460 14356 6512 14408
rect 9680 14356 9732 14408
rect 11336 14356 11388 14408
rect 12716 14399 12768 14408
rect 12716 14365 12725 14399
rect 12725 14365 12759 14399
rect 12759 14365 12768 14399
rect 12716 14356 12768 14365
rect 13912 14356 13964 14408
rect 16672 14356 16724 14408
rect 12440 14288 12492 14340
rect 1952 14263 2004 14272
rect 1952 14229 1961 14263
rect 1961 14229 1995 14263
rect 1995 14229 2004 14263
rect 1952 14220 2004 14229
rect 2228 14263 2280 14272
rect 2228 14229 2237 14263
rect 2237 14229 2271 14263
rect 2271 14229 2280 14263
rect 2228 14220 2280 14229
rect 2964 14220 3016 14272
rect 5540 14220 5592 14272
rect 7288 14220 7340 14272
rect 8852 14263 8904 14272
rect 8852 14229 8861 14263
rect 8861 14229 8895 14263
rect 8895 14229 8904 14263
rect 8852 14220 8904 14229
rect 12164 14220 12216 14272
rect 12532 14263 12584 14272
rect 12532 14229 12541 14263
rect 12541 14229 12575 14263
rect 12575 14229 12584 14263
rect 12532 14220 12584 14229
rect 15476 14220 15528 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 3332 14016 3384 14068
rect 4068 14016 4120 14068
rect 4528 14059 4580 14068
rect 4528 14025 4537 14059
rect 4537 14025 4571 14059
rect 4571 14025 4580 14059
rect 4528 14016 4580 14025
rect 5172 14059 5224 14068
rect 5172 14025 5181 14059
rect 5181 14025 5215 14059
rect 5215 14025 5224 14059
rect 5172 14016 5224 14025
rect 5540 14016 5592 14068
rect 6184 14059 6236 14068
rect 6184 14025 6193 14059
rect 6193 14025 6227 14059
rect 6227 14025 6236 14059
rect 6184 14016 6236 14025
rect 6460 14016 6512 14068
rect 6644 14059 6696 14068
rect 6644 14025 6653 14059
rect 6653 14025 6687 14059
rect 6687 14025 6696 14059
rect 6644 14016 6696 14025
rect 7288 14016 7340 14068
rect 8484 14016 8536 14068
rect 9864 14059 9916 14068
rect 9864 14025 9873 14059
rect 9873 14025 9907 14059
rect 9907 14025 9916 14059
rect 9864 14016 9916 14025
rect 10048 14016 10100 14068
rect 10324 14059 10376 14068
rect 10324 14025 10333 14059
rect 10333 14025 10367 14059
rect 10367 14025 10376 14059
rect 10324 14016 10376 14025
rect 11336 14059 11388 14068
rect 11336 14025 11345 14059
rect 11345 14025 11379 14059
rect 11379 14025 11388 14059
rect 11336 14016 11388 14025
rect 12256 14059 12308 14068
rect 12256 14025 12265 14059
rect 12265 14025 12299 14059
rect 12299 14025 12308 14059
rect 12256 14016 12308 14025
rect 12716 14059 12768 14068
rect 12716 14025 12725 14059
rect 12725 14025 12759 14059
rect 12759 14025 12768 14059
rect 12716 14016 12768 14025
rect 13820 14016 13872 14068
rect 13912 14016 13964 14068
rect 2228 13923 2280 13932
rect 2228 13889 2237 13923
rect 2237 13889 2271 13923
rect 2271 13889 2280 13923
rect 2228 13880 2280 13889
rect 3700 13923 3752 13932
rect 3700 13889 3709 13923
rect 3709 13889 3743 13923
rect 3743 13889 3752 13923
rect 3700 13880 3752 13889
rect 2044 13855 2096 13864
rect 2044 13821 2053 13855
rect 2053 13821 2087 13855
rect 2087 13821 2096 13855
rect 2044 13812 2096 13821
rect 3056 13855 3108 13864
rect 3056 13821 3065 13855
rect 3065 13821 3099 13855
rect 3099 13821 3108 13855
rect 3608 13855 3660 13864
rect 3056 13812 3108 13821
rect 3608 13821 3617 13855
rect 3617 13821 3651 13855
rect 3651 13821 3660 13855
rect 3608 13812 3660 13821
rect 3516 13787 3568 13796
rect 3516 13753 3525 13787
rect 3525 13753 3559 13787
rect 3559 13753 3568 13787
rect 3516 13744 3568 13753
rect 6092 13880 6144 13932
rect 8760 13948 8812 14000
rect 9312 13948 9364 14000
rect 7564 13880 7616 13932
rect 9404 13923 9456 13932
rect 9404 13889 9413 13923
rect 9413 13889 9447 13923
rect 9447 13889 9456 13923
rect 9404 13880 9456 13889
rect 10140 13880 10192 13932
rect 10692 13880 10744 13932
rect 5908 13812 5960 13864
rect 6828 13812 6880 13864
rect 7932 13812 7984 13864
rect 8852 13812 8904 13864
rect 10048 13812 10100 13864
rect 15384 13812 15436 13864
rect 15568 13812 15620 13864
rect 4896 13744 4948 13796
rect 5540 13787 5592 13796
rect 5540 13753 5549 13787
rect 5549 13753 5583 13787
rect 5583 13753 5592 13787
rect 5540 13744 5592 13753
rect 8484 13744 8536 13796
rect 9220 13787 9272 13796
rect 9220 13753 9229 13787
rect 9229 13753 9263 13787
rect 9263 13753 9272 13787
rect 9220 13744 9272 13753
rect 9864 13744 9916 13796
rect 11152 13744 11204 13796
rect 12532 13744 12584 13796
rect 2044 13676 2096 13728
rect 7380 13676 7432 13728
rect 8300 13719 8352 13728
rect 8300 13685 8309 13719
rect 8309 13685 8343 13719
rect 8343 13685 8352 13719
rect 8300 13676 8352 13685
rect 8760 13719 8812 13728
rect 8760 13685 8769 13719
rect 8769 13685 8803 13719
rect 8803 13685 8812 13719
rect 8760 13676 8812 13685
rect 13728 13719 13780 13728
rect 13728 13685 13737 13719
rect 13737 13685 13771 13719
rect 13771 13685 13780 13719
rect 16212 13719 16264 13728
rect 13728 13676 13780 13685
rect 16212 13685 16221 13719
rect 16221 13685 16255 13719
rect 16255 13685 16264 13719
rect 16212 13676 16264 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 3056 13472 3108 13524
rect 3516 13515 3568 13524
rect 3516 13481 3525 13515
rect 3525 13481 3559 13515
rect 3559 13481 3568 13515
rect 3516 13472 3568 13481
rect 3700 13472 3752 13524
rect 3976 13472 4028 13524
rect 4344 13472 4396 13524
rect 4620 13472 4672 13524
rect 5540 13515 5592 13524
rect 5540 13481 5549 13515
rect 5549 13481 5583 13515
rect 5583 13481 5592 13515
rect 5540 13472 5592 13481
rect 5908 13515 5960 13524
rect 5908 13481 5917 13515
rect 5917 13481 5951 13515
rect 5951 13481 5960 13515
rect 5908 13472 5960 13481
rect 6552 13472 6604 13524
rect 7564 13515 7616 13524
rect 7564 13481 7573 13515
rect 7573 13481 7607 13515
rect 7607 13481 7616 13515
rect 7564 13472 7616 13481
rect 8392 13472 8444 13524
rect 8944 13472 8996 13524
rect 9680 13515 9732 13524
rect 9680 13481 9689 13515
rect 9689 13481 9723 13515
rect 9723 13481 9732 13515
rect 9680 13472 9732 13481
rect 9956 13472 10008 13524
rect 10692 13515 10744 13524
rect 10692 13481 10701 13515
rect 10701 13481 10735 13515
rect 10735 13481 10744 13515
rect 10692 13472 10744 13481
rect 13728 13472 13780 13524
rect 14004 13472 14056 13524
rect 15476 13472 15528 13524
rect 15660 13472 15712 13524
rect 16672 13515 16724 13524
rect 16672 13481 16681 13515
rect 16681 13481 16715 13515
rect 16715 13481 16724 13515
rect 16672 13472 16724 13481
rect 17316 13515 17368 13524
rect 17316 13481 17325 13515
rect 17325 13481 17359 13515
rect 17359 13481 17368 13515
rect 17316 13472 17368 13481
rect 1400 13379 1452 13388
rect 1400 13345 1409 13379
rect 1409 13345 1443 13379
rect 1443 13345 1452 13379
rect 1400 13336 1452 13345
rect 2688 13336 2740 13388
rect 3700 13336 3752 13388
rect 5356 13336 5408 13388
rect 6368 13379 6420 13388
rect 6368 13345 6377 13379
rect 6377 13345 6411 13379
rect 6411 13345 6420 13379
rect 6368 13336 6420 13345
rect 7932 13404 7984 13456
rect 11060 13447 11112 13456
rect 11060 13413 11069 13447
rect 11069 13413 11103 13447
rect 11103 13413 11112 13447
rect 11060 13404 11112 13413
rect 12164 13447 12216 13456
rect 12164 13413 12173 13447
rect 12173 13413 12207 13447
rect 12207 13413 12216 13447
rect 12164 13404 12216 13413
rect 12808 13404 12860 13456
rect 17408 13404 17460 13456
rect 8392 13379 8444 13388
rect 8392 13345 8401 13379
rect 8401 13345 8435 13379
rect 8435 13345 8444 13379
rect 8392 13336 8444 13345
rect 9036 13336 9088 13388
rect 11520 13336 11572 13388
rect 13728 13379 13780 13388
rect 13728 13345 13737 13379
rect 13737 13345 13771 13379
rect 13771 13345 13780 13379
rect 13728 13336 13780 13345
rect 14556 13336 14608 13388
rect 15568 13336 15620 13388
rect 15752 13379 15804 13388
rect 15752 13345 15761 13379
rect 15761 13345 15795 13379
rect 15795 13345 15804 13379
rect 15752 13336 15804 13345
rect 1768 13200 1820 13252
rect 2044 13200 2096 13252
rect 3240 13200 3292 13252
rect 5540 13268 5592 13320
rect 6460 13311 6512 13320
rect 6460 13277 6469 13311
rect 6469 13277 6503 13311
rect 6503 13277 6512 13311
rect 6460 13268 6512 13277
rect 6552 13311 6604 13320
rect 6552 13277 6561 13311
rect 6561 13277 6595 13311
rect 6595 13277 6604 13311
rect 6552 13268 6604 13277
rect 6736 13268 6788 13320
rect 7932 13268 7984 13320
rect 8484 13311 8536 13320
rect 8484 13277 8493 13311
rect 8493 13277 8527 13311
rect 8527 13277 8536 13311
rect 8484 13268 8536 13277
rect 8208 13200 8260 13252
rect 2412 13175 2464 13184
rect 2412 13141 2421 13175
rect 2421 13141 2455 13175
rect 2455 13141 2464 13175
rect 2412 13132 2464 13141
rect 4436 13175 4488 13184
rect 4436 13141 4445 13175
rect 4445 13141 4479 13175
rect 4479 13141 4488 13175
rect 4436 13132 4488 13141
rect 8024 13175 8076 13184
rect 8024 13141 8033 13175
rect 8033 13141 8067 13175
rect 8067 13141 8076 13175
rect 8024 13132 8076 13141
rect 10692 13268 10744 13320
rect 11152 13268 11204 13320
rect 13452 13268 13504 13320
rect 13544 13268 13596 13320
rect 14740 13268 14792 13320
rect 16212 13268 16264 13320
rect 16672 13268 16724 13320
rect 17684 13268 17736 13320
rect 12164 13200 12216 13252
rect 15568 13200 15620 13252
rect 16028 13200 16080 13252
rect 9404 13132 9456 13184
rect 11428 13175 11480 13184
rect 11428 13141 11437 13175
rect 11437 13141 11471 13175
rect 11471 13141 11480 13175
rect 11428 13132 11480 13141
rect 12900 13175 12952 13184
rect 12900 13141 12909 13175
rect 12909 13141 12943 13175
rect 12943 13141 12952 13175
rect 12900 13132 12952 13141
rect 15844 13132 15896 13184
rect 16764 13132 16816 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2044 12928 2096 12980
rect 2320 12928 2372 12980
rect 3700 12928 3752 12980
rect 6552 12928 6604 12980
rect 7932 12928 7984 12980
rect 8392 12971 8444 12980
rect 8392 12937 8401 12971
rect 8401 12937 8435 12971
rect 8435 12937 8444 12971
rect 8392 12928 8444 12937
rect 9036 12971 9088 12980
rect 9036 12937 9045 12971
rect 9045 12937 9079 12971
rect 9079 12937 9088 12971
rect 9036 12928 9088 12937
rect 10692 12928 10744 12980
rect 12532 12971 12584 12980
rect 12532 12937 12541 12971
rect 12541 12937 12575 12971
rect 12575 12937 12584 12971
rect 12532 12928 12584 12937
rect 13544 12971 13596 12980
rect 13544 12937 13553 12971
rect 13553 12937 13587 12971
rect 13587 12937 13596 12971
rect 13544 12928 13596 12937
rect 14004 12971 14056 12980
rect 14004 12937 14013 12971
rect 14013 12937 14047 12971
rect 14047 12937 14056 12971
rect 14004 12928 14056 12937
rect 14556 12971 14608 12980
rect 14556 12937 14565 12971
rect 14565 12937 14599 12971
rect 14599 12937 14608 12971
rect 14556 12928 14608 12937
rect 14740 12928 14792 12980
rect 17408 12971 17460 12980
rect 17408 12937 17417 12971
rect 17417 12937 17451 12971
rect 17451 12937 17460 12971
rect 17408 12928 17460 12937
rect 4068 12903 4120 12912
rect 4068 12869 4077 12903
rect 4077 12869 4111 12903
rect 4111 12869 4120 12903
rect 4068 12860 4120 12869
rect 6460 12860 6512 12912
rect 4988 12835 5040 12844
rect 4988 12801 4997 12835
rect 4997 12801 5031 12835
rect 5031 12801 5040 12835
rect 4988 12792 5040 12801
rect 5172 12835 5224 12844
rect 5172 12801 5181 12835
rect 5181 12801 5215 12835
rect 5215 12801 5224 12835
rect 5172 12792 5224 12801
rect 6736 12792 6788 12844
rect 8668 12792 8720 12844
rect 9128 12835 9180 12844
rect 9128 12801 9137 12835
rect 9137 12801 9171 12835
rect 9171 12801 9180 12835
rect 9128 12792 9180 12801
rect 4896 12767 4948 12776
rect 4896 12733 4905 12767
rect 4905 12733 4939 12767
rect 4939 12733 4948 12767
rect 4896 12724 4948 12733
rect 9404 12767 9456 12776
rect 9404 12733 9438 12767
rect 9438 12733 9456 12767
rect 9404 12724 9456 12733
rect 9956 12724 10008 12776
rect 2688 12656 2740 12708
rect 12440 12792 12492 12844
rect 13452 12792 13504 12844
rect 15200 12792 15252 12844
rect 12900 12767 12952 12776
rect 12900 12733 12909 12767
rect 12909 12733 12943 12767
rect 12943 12733 12952 12767
rect 12900 12724 12952 12733
rect 16212 12724 16264 12776
rect 18052 12767 18104 12776
rect 18052 12733 18061 12767
rect 18061 12733 18095 12767
rect 18095 12733 18104 12767
rect 18052 12724 18104 12733
rect 18328 12767 18380 12776
rect 18328 12733 18362 12767
rect 18362 12733 18380 12767
rect 18328 12724 18380 12733
rect 16488 12656 16540 12708
rect 1860 12631 1912 12640
rect 1860 12597 1869 12631
rect 1869 12597 1903 12631
rect 1903 12597 1912 12631
rect 1860 12588 1912 12597
rect 3424 12631 3476 12640
rect 3424 12597 3433 12631
rect 3433 12597 3467 12631
rect 3467 12597 3476 12631
rect 3424 12588 3476 12597
rect 4528 12631 4580 12640
rect 4528 12597 4537 12631
rect 4537 12597 4571 12631
rect 4571 12597 4580 12631
rect 4528 12588 4580 12597
rect 5632 12631 5684 12640
rect 5632 12597 5641 12631
rect 5641 12597 5675 12631
rect 5675 12597 5684 12631
rect 5632 12588 5684 12597
rect 7196 12631 7248 12640
rect 7196 12597 7205 12631
rect 7205 12597 7239 12631
rect 7239 12597 7248 12631
rect 7196 12588 7248 12597
rect 7288 12631 7340 12640
rect 7288 12597 7297 12631
rect 7297 12597 7331 12631
rect 7331 12597 7340 12631
rect 7288 12588 7340 12597
rect 10784 12588 10836 12640
rect 14096 12631 14148 12640
rect 14096 12597 14105 12631
rect 14105 12597 14139 12631
rect 14139 12597 14148 12631
rect 14096 12588 14148 12597
rect 16856 12631 16908 12640
rect 16856 12597 16865 12631
rect 16865 12597 16899 12631
rect 16899 12597 16908 12631
rect 16856 12588 16908 12597
rect 19432 12631 19484 12640
rect 19432 12597 19441 12631
rect 19441 12597 19475 12631
rect 19475 12597 19484 12631
rect 19432 12588 19484 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1676 12384 1728 12436
rect 1952 12384 2004 12436
rect 2320 12384 2372 12436
rect 2596 12384 2648 12436
rect 2688 12384 2740 12436
rect 5172 12384 5224 12436
rect 6736 12427 6788 12436
rect 6736 12393 6745 12427
rect 6745 12393 6779 12427
rect 6779 12393 6788 12427
rect 6736 12384 6788 12393
rect 7288 12427 7340 12436
rect 7288 12393 7297 12427
rect 7297 12393 7331 12427
rect 7331 12393 7340 12427
rect 7288 12384 7340 12393
rect 8208 12384 8260 12436
rect 9128 12427 9180 12436
rect 9128 12393 9137 12427
rect 9137 12393 9171 12427
rect 9171 12393 9180 12427
rect 9128 12384 9180 12393
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 10140 12427 10192 12436
rect 10140 12393 10149 12427
rect 10149 12393 10183 12427
rect 10183 12393 10192 12427
rect 10140 12384 10192 12393
rect 12900 12384 12952 12436
rect 14464 12384 14516 12436
rect 15108 12384 15160 12436
rect 15844 12427 15896 12436
rect 15844 12393 15853 12427
rect 15853 12393 15887 12427
rect 15887 12393 15896 12427
rect 15844 12384 15896 12393
rect 17408 12384 17460 12436
rect 17592 12384 17644 12436
rect 18052 12427 18104 12436
rect 18052 12393 18061 12427
rect 18061 12393 18095 12427
rect 18095 12393 18104 12427
rect 18052 12384 18104 12393
rect 9496 12316 9548 12368
rect 13084 12316 13136 12368
rect 13728 12316 13780 12368
rect 1952 12248 2004 12300
rect 4068 12291 4120 12300
rect 1400 12223 1452 12232
rect 1400 12189 1409 12223
rect 1409 12189 1443 12223
rect 1443 12189 1452 12223
rect 1400 12180 1452 12189
rect 4068 12257 4077 12291
rect 4077 12257 4111 12291
rect 4111 12257 4120 12291
rect 4068 12248 4120 12257
rect 4436 12248 4488 12300
rect 5080 12248 5132 12300
rect 6000 12248 6052 12300
rect 7472 12248 7524 12300
rect 8024 12248 8076 12300
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 10048 12248 10100 12257
rect 10876 12248 10928 12300
rect 11612 12291 11664 12300
rect 11612 12257 11621 12291
rect 11621 12257 11655 12291
rect 11655 12257 11664 12291
rect 11612 12248 11664 12257
rect 11704 12291 11756 12300
rect 11704 12257 11713 12291
rect 11713 12257 11747 12291
rect 11747 12257 11756 12291
rect 11704 12248 11756 12257
rect 14096 12248 14148 12300
rect 15752 12291 15804 12300
rect 15752 12257 15761 12291
rect 15761 12257 15795 12291
rect 15795 12257 15804 12291
rect 15752 12248 15804 12257
rect 17040 12248 17092 12300
rect 3516 12180 3568 12232
rect 8300 12223 8352 12232
rect 3148 12044 3200 12096
rect 3608 12044 3660 12096
rect 4252 12087 4304 12096
rect 4252 12053 4261 12087
rect 4261 12053 4295 12087
rect 4295 12053 4304 12087
rect 4252 12044 4304 12053
rect 4620 12044 4672 12096
rect 4896 12044 4948 12096
rect 8300 12189 8309 12223
rect 8309 12189 8343 12223
rect 8343 12189 8352 12223
rect 8300 12180 8352 12189
rect 8484 12223 8536 12232
rect 8484 12189 8493 12223
rect 8493 12189 8527 12223
rect 8527 12189 8536 12223
rect 8484 12180 8536 12189
rect 10324 12223 10376 12232
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 10784 12180 10836 12232
rect 11888 12223 11940 12232
rect 11888 12189 11897 12223
rect 11897 12189 11931 12223
rect 11931 12189 11940 12223
rect 11888 12180 11940 12189
rect 13452 12223 13504 12232
rect 13452 12189 13461 12223
rect 13461 12189 13495 12223
rect 13495 12189 13504 12223
rect 16028 12223 16080 12232
rect 13452 12180 13504 12189
rect 13728 12112 13780 12164
rect 16028 12189 16037 12223
rect 16037 12189 16071 12223
rect 16071 12189 16080 12223
rect 16028 12180 16080 12189
rect 16856 12180 16908 12232
rect 17316 12180 17368 12232
rect 17592 12223 17644 12232
rect 17040 12112 17092 12164
rect 17592 12189 17601 12223
rect 17601 12189 17635 12223
rect 17635 12189 17644 12223
rect 17592 12180 17644 12189
rect 5540 12044 5592 12096
rect 10784 12087 10836 12096
rect 10784 12053 10793 12087
rect 10793 12053 10827 12087
rect 10827 12053 10836 12087
rect 10784 12044 10836 12053
rect 11244 12044 11296 12096
rect 13820 12087 13872 12096
rect 13820 12053 13829 12087
rect 13829 12053 13863 12087
rect 13863 12053 13872 12087
rect 13820 12044 13872 12053
rect 14740 12044 14792 12096
rect 15292 12044 15344 12096
rect 16396 12087 16448 12096
rect 16396 12053 16405 12087
rect 16405 12053 16439 12087
rect 16439 12053 16448 12087
rect 16396 12044 16448 12053
rect 16948 12087 17000 12096
rect 16948 12053 16957 12087
rect 16957 12053 16991 12087
rect 16991 12053 17000 12087
rect 16948 12044 17000 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1584 11883 1636 11892
rect 1584 11849 1593 11883
rect 1593 11849 1627 11883
rect 1627 11849 1636 11883
rect 1584 11840 1636 11849
rect 4068 11840 4120 11892
rect 6552 11840 6604 11892
rect 8300 11840 8352 11892
rect 8760 11840 8812 11892
rect 10048 11840 10100 11892
rect 1400 11772 1452 11824
rect 1860 11772 1912 11824
rect 1400 11679 1452 11688
rect 1400 11645 1409 11679
rect 1409 11645 1443 11679
rect 1443 11645 1452 11679
rect 1400 11636 1452 11645
rect 8484 11772 8536 11824
rect 10324 11840 10376 11892
rect 10968 11840 11020 11892
rect 11612 11840 11664 11892
rect 12532 11840 12584 11892
rect 12808 11840 12860 11892
rect 14096 11840 14148 11892
rect 14648 11840 14700 11892
rect 15844 11840 15896 11892
rect 11704 11772 11756 11824
rect 15752 11772 15804 11824
rect 10784 11704 10836 11756
rect 14740 11704 14792 11756
rect 15384 11704 15436 11756
rect 2780 11636 2832 11688
rect 3424 11636 3476 11688
rect 6644 11636 6696 11688
rect 6920 11636 6972 11688
rect 11244 11679 11296 11688
rect 11244 11645 11253 11679
rect 11253 11645 11287 11679
rect 11287 11645 11296 11679
rect 11244 11636 11296 11645
rect 11428 11636 11480 11688
rect 12624 11636 12676 11688
rect 13084 11636 13136 11688
rect 17316 11636 17368 11688
rect 2964 11568 3016 11620
rect 2780 11543 2832 11552
rect 2780 11509 2789 11543
rect 2789 11509 2823 11543
rect 2823 11509 2832 11543
rect 2780 11500 2832 11509
rect 3424 11500 3476 11552
rect 5540 11568 5592 11620
rect 6000 11568 6052 11620
rect 8484 11568 8536 11620
rect 11152 11611 11204 11620
rect 11152 11577 11161 11611
rect 11161 11577 11195 11611
rect 11195 11577 11204 11611
rect 11152 11568 11204 11577
rect 12716 11568 12768 11620
rect 5632 11500 5684 11552
rect 6644 11543 6696 11552
rect 6644 11509 6653 11543
rect 6653 11509 6687 11543
rect 6687 11509 6696 11543
rect 6644 11500 6696 11509
rect 8208 11543 8260 11552
rect 8208 11509 8217 11543
rect 8217 11509 8251 11543
rect 8251 11509 8260 11543
rect 8208 11500 8260 11509
rect 13452 11500 13504 11552
rect 13820 11500 13872 11552
rect 14832 11543 14884 11552
rect 14832 11509 14841 11543
rect 14841 11509 14875 11543
rect 14875 11509 14884 11543
rect 14832 11500 14884 11509
rect 15476 11543 15528 11552
rect 15476 11509 15485 11543
rect 15485 11509 15519 11543
rect 15519 11509 15528 11543
rect 15476 11500 15528 11509
rect 17040 11500 17092 11552
rect 17592 11500 17644 11552
rect 18604 11500 18656 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1400 11296 1452 11348
rect 1952 11339 2004 11348
rect 1952 11305 1961 11339
rect 1961 11305 1995 11339
rect 1995 11305 2004 11339
rect 1952 11296 2004 11305
rect 2044 11296 2096 11348
rect 4068 11296 4120 11348
rect 5448 11296 5500 11348
rect 5632 11296 5684 11348
rect 6920 11296 6972 11348
rect 7472 11339 7524 11348
rect 7472 11305 7481 11339
rect 7481 11305 7515 11339
rect 7515 11305 7524 11339
rect 7472 11296 7524 11305
rect 8208 11296 8260 11348
rect 8300 11296 8352 11348
rect 8944 11339 8996 11348
rect 3148 11228 3200 11280
rect 3424 11271 3476 11280
rect 3424 11237 3433 11271
rect 3433 11237 3467 11271
rect 3467 11237 3476 11271
rect 3424 11228 3476 11237
rect 2136 11160 2188 11212
rect 2780 11203 2832 11212
rect 2780 11169 2789 11203
rect 2789 11169 2823 11203
rect 2823 11169 2832 11203
rect 2780 11160 2832 11169
rect 4344 11160 4396 11212
rect 4804 11160 4856 11212
rect 6000 11228 6052 11280
rect 6736 11228 6788 11280
rect 8944 11305 8953 11339
rect 8953 11305 8987 11339
rect 8987 11305 8996 11339
rect 8944 11296 8996 11305
rect 10140 11296 10192 11348
rect 12440 11296 12492 11348
rect 13268 11339 13320 11348
rect 13268 11305 13277 11339
rect 13277 11305 13311 11339
rect 13311 11305 13320 11339
rect 13268 11296 13320 11305
rect 13728 11296 13780 11348
rect 14280 11339 14332 11348
rect 7748 11160 7800 11212
rect 8300 11203 8352 11212
rect 8300 11169 8309 11203
rect 8309 11169 8343 11203
rect 8343 11169 8352 11203
rect 8300 11160 8352 11169
rect 9588 11228 9640 11280
rect 10048 11228 10100 11280
rect 11336 11228 11388 11280
rect 13912 11271 13964 11280
rect 2964 11135 3016 11144
rect 2964 11101 2973 11135
rect 2973 11101 3007 11135
rect 3007 11101 3016 11135
rect 4620 11135 4672 11144
rect 2964 11092 3016 11101
rect 4620 11101 4629 11135
rect 4629 11101 4663 11135
rect 4663 11101 4672 11135
rect 4620 11092 4672 11101
rect 8392 11135 8444 11144
rect 8392 11101 8401 11135
rect 8401 11101 8435 11135
rect 8435 11101 8444 11135
rect 8392 11092 8444 11101
rect 10968 11160 11020 11212
rect 13912 11237 13921 11271
rect 13921 11237 13955 11271
rect 13955 11237 13964 11271
rect 13912 11228 13964 11237
rect 14280 11305 14289 11339
rect 14289 11305 14323 11339
rect 14323 11305 14332 11339
rect 14280 11296 14332 11305
rect 14924 11296 14976 11348
rect 16396 11296 16448 11348
rect 17132 11271 17184 11280
rect 17132 11237 17141 11271
rect 17141 11237 17175 11271
rect 17175 11237 17184 11271
rect 17132 11228 17184 11237
rect 15476 11160 15528 11212
rect 15752 11160 15804 11212
rect 16028 11160 16080 11212
rect 4068 11024 4120 11076
rect 4896 11024 4948 11076
rect 6920 11024 6972 11076
rect 10232 11024 10284 11076
rect 8576 10956 8628 11008
rect 9956 10999 10008 11008
rect 9956 10965 9965 10999
rect 9965 10965 9999 10999
rect 9999 10965 10008 10999
rect 9956 10956 10008 10965
rect 10324 10999 10376 11008
rect 10324 10965 10333 10999
rect 10333 10965 10367 10999
rect 10367 10965 10376 10999
rect 10324 10956 10376 10965
rect 12716 11024 12768 11076
rect 13452 11135 13504 11144
rect 13452 11101 13461 11135
rect 13461 11101 13495 11135
rect 13495 11101 13504 11135
rect 13452 11092 13504 11101
rect 15292 11092 15344 11144
rect 16304 11135 16356 11144
rect 16304 11101 16313 11135
rect 16313 11101 16347 11135
rect 16347 11101 16356 11135
rect 16304 11092 16356 11101
rect 17408 11160 17460 11212
rect 17868 11135 17920 11144
rect 17868 11101 17877 11135
rect 17877 11101 17911 11135
rect 17911 11101 17920 11135
rect 17868 11092 17920 11101
rect 15660 11067 15712 11076
rect 11428 10956 11480 11008
rect 13084 10956 13136 11008
rect 15660 11033 15669 11067
rect 15669 11033 15703 11067
rect 15703 11033 15712 11067
rect 15660 11024 15712 11033
rect 14648 10956 14700 11008
rect 18604 10956 18656 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 2688 10752 2740 10804
rect 3056 10752 3108 10804
rect 4344 10795 4396 10804
rect 4344 10761 4353 10795
rect 4353 10761 4387 10795
rect 4387 10761 4396 10795
rect 4344 10752 4396 10761
rect 5356 10752 5408 10804
rect 7196 10752 7248 10804
rect 8392 10752 8444 10804
rect 9680 10795 9732 10804
rect 9680 10761 9689 10795
rect 9689 10761 9723 10795
rect 9723 10761 9732 10795
rect 9680 10752 9732 10761
rect 11428 10752 11480 10804
rect 13452 10795 13504 10804
rect 13452 10761 13461 10795
rect 13461 10761 13495 10795
rect 13495 10761 13504 10795
rect 13452 10752 13504 10761
rect 14648 10795 14700 10804
rect 14648 10761 14657 10795
rect 14657 10761 14691 10795
rect 14691 10761 14700 10795
rect 14648 10752 14700 10761
rect 14740 10752 14792 10804
rect 2044 10659 2096 10668
rect 2044 10625 2053 10659
rect 2053 10625 2087 10659
rect 2087 10625 2096 10659
rect 2044 10616 2096 10625
rect 2320 10616 2372 10668
rect 1400 10548 1452 10600
rect 3424 10616 3476 10668
rect 3884 10616 3936 10668
rect 7748 10684 7800 10736
rect 8760 10684 8812 10736
rect 11060 10684 11112 10736
rect 6000 10616 6052 10668
rect 9956 10616 10008 10668
rect 13084 10659 13136 10668
rect 13084 10625 13093 10659
rect 13093 10625 13127 10659
rect 13127 10625 13136 10659
rect 13084 10616 13136 10625
rect 15844 10752 15896 10804
rect 16488 10752 16540 10804
rect 18052 10795 18104 10804
rect 18052 10761 18061 10795
rect 18061 10761 18095 10795
rect 18095 10761 18104 10795
rect 18052 10752 18104 10761
rect 18604 10659 18656 10668
rect 18604 10625 18613 10659
rect 18613 10625 18647 10659
rect 18647 10625 18656 10659
rect 18604 10616 18656 10625
rect 5540 10548 5592 10600
rect 6644 10548 6696 10600
rect 7104 10548 7156 10600
rect 9680 10548 9732 10600
rect 10232 10548 10284 10600
rect 10324 10548 10376 10600
rect 12624 10548 12676 10600
rect 1860 10523 1912 10532
rect 1860 10489 1869 10523
rect 1869 10489 1903 10523
rect 1903 10489 1912 10523
rect 1860 10480 1912 10489
rect 4068 10480 4120 10532
rect 8208 10480 8260 10532
rect 9312 10480 9364 10532
rect 9496 10480 9548 10532
rect 13176 10548 13228 10600
rect 13820 10591 13872 10600
rect 13820 10557 13829 10591
rect 13829 10557 13863 10591
rect 13863 10557 13872 10591
rect 13820 10548 13872 10557
rect 15752 10523 15804 10532
rect 15752 10489 15786 10523
rect 15786 10489 15804 10523
rect 15752 10480 15804 10489
rect 18236 10480 18288 10532
rect 5632 10412 5684 10464
rect 9128 10455 9180 10464
rect 9128 10421 9137 10455
rect 9137 10421 9171 10455
rect 9171 10421 9180 10455
rect 9128 10412 9180 10421
rect 9956 10412 10008 10464
rect 11612 10455 11664 10464
rect 11612 10421 11621 10455
rect 11621 10421 11655 10455
rect 11655 10421 11664 10455
rect 11612 10412 11664 10421
rect 12716 10412 12768 10464
rect 13912 10412 13964 10464
rect 16764 10412 16816 10464
rect 17408 10455 17460 10464
rect 17408 10421 17417 10455
rect 17417 10421 17451 10455
rect 17451 10421 17460 10455
rect 17408 10412 17460 10421
rect 18052 10412 18104 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2044 10208 2096 10260
rect 2596 10208 2648 10260
rect 3792 10251 3844 10260
rect 3792 10217 3801 10251
rect 3801 10217 3835 10251
rect 3835 10217 3844 10251
rect 3792 10208 3844 10217
rect 5632 10208 5684 10260
rect 10968 10208 11020 10260
rect 11612 10208 11664 10260
rect 12624 10208 12676 10260
rect 13820 10251 13872 10260
rect 13820 10217 13829 10251
rect 13829 10217 13863 10251
rect 13863 10217 13872 10251
rect 13820 10208 13872 10217
rect 15108 10251 15160 10260
rect 15108 10217 15117 10251
rect 15117 10217 15151 10251
rect 15151 10217 15160 10251
rect 15108 10208 15160 10217
rect 15752 10208 15804 10260
rect 18052 10251 18104 10260
rect 18052 10217 18061 10251
rect 18061 10217 18095 10251
rect 18095 10217 18104 10251
rect 18052 10208 18104 10217
rect 18512 10251 18564 10260
rect 18512 10217 18521 10251
rect 18521 10217 18555 10251
rect 18555 10217 18564 10251
rect 18512 10208 18564 10217
rect 18972 10251 19024 10260
rect 18972 10217 18981 10251
rect 18981 10217 19015 10251
rect 19015 10217 19024 10251
rect 18972 10208 19024 10217
rect 19432 10208 19484 10260
rect 6920 10183 6972 10192
rect 6920 10149 6929 10183
rect 6929 10149 6963 10183
rect 6963 10149 6972 10183
rect 6920 10140 6972 10149
rect 8208 10140 8260 10192
rect 8576 10140 8628 10192
rect 14188 10183 14240 10192
rect 14188 10149 14197 10183
rect 14197 10149 14231 10183
rect 14231 10149 14240 10183
rect 14188 10140 14240 10149
rect 1768 10115 1820 10124
rect 1768 10081 1777 10115
rect 1777 10081 1811 10115
rect 1811 10081 1820 10115
rect 1768 10072 1820 10081
rect 5264 10115 5316 10124
rect 5264 10081 5273 10115
rect 5273 10081 5307 10115
rect 5307 10081 5316 10115
rect 5264 10072 5316 10081
rect 6828 10115 6880 10124
rect 6828 10081 6837 10115
rect 6837 10081 6871 10115
rect 6871 10081 6880 10115
rect 6828 10072 6880 10081
rect 8760 10072 8812 10124
rect 1676 10004 1728 10056
rect 1952 10047 2004 10056
rect 1952 10013 1961 10047
rect 1961 10013 1995 10047
rect 1995 10013 2004 10047
rect 1952 10004 2004 10013
rect 4988 10004 5040 10056
rect 5448 10047 5500 10056
rect 5448 10013 5457 10047
rect 5457 10013 5491 10047
rect 5491 10013 5500 10047
rect 5448 10004 5500 10013
rect 1400 9979 1452 9988
rect 1400 9945 1409 9979
rect 1409 9945 1443 9979
rect 1443 9945 1452 9979
rect 1400 9936 1452 9945
rect 6552 9936 6604 9988
rect 8300 10004 8352 10056
rect 12440 10072 12492 10124
rect 15936 10072 15988 10124
rect 16304 10115 16356 10124
rect 16304 10081 16327 10115
rect 16327 10081 16356 10115
rect 18880 10115 18932 10124
rect 16304 10072 16356 10081
rect 18880 10081 18889 10115
rect 18889 10081 18923 10115
rect 18923 10081 18932 10115
rect 18880 10072 18932 10081
rect 9680 10047 9732 10056
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 12624 10004 12676 10056
rect 13268 10047 13320 10056
rect 13268 10013 13277 10047
rect 13277 10013 13311 10047
rect 13311 10013 13320 10047
rect 13268 10004 13320 10013
rect 13452 10047 13504 10056
rect 13452 10013 13461 10047
rect 13461 10013 13495 10047
rect 13495 10013 13504 10047
rect 13452 10004 13504 10013
rect 15844 10004 15896 10056
rect 16028 10047 16080 10056
rect 16028 10013 16037 10047
rect 16037 10013 16071 10047
rect 16071 10013 16080 10047
rect 16028 10004 16080 10013
rect 19064 10047 19116 10056
rect 9128 9936 9180 9988
rect 2780 9868 2832 9920
rect 4344 9911 4396 9920
rect 4344 9877 4353 9911
rect 4353 9877 4387 9911
rect 4387 9877 4396 9911
rect 4344 9868 4396 9877
rect 4620 9911 4672 9920
rect 4620 9877 4629 9911
rect 4629 9877 4663 9911
rect 4663 9877 4672 9911
rect 4620 9868 4672 9877
rect 5540 9868 5592 9920
rect 7472 9911 7524 9920
rect 7472 9877 7481 9911
rect 7481 9877 7515 9911
rect 7515 9877 7524 9911
rect 7472 9868 7524 9877
rect 8024 9911 8076 9920
rect 8024 9877 8033 9911
rect 8033 9877 8067 9911
rect 8067 9877 8076 9911
rect 8024 9868 8076 9877
rect 9864 9868 9916 9920
rect 11796 9936 11848 9988
rect 13636 9936 13688 9988
rect 11152 9868 11204 9920
rect 11980 9911 12032 9920
rect 11980 9877 11989 9911
rect 11989 9877 12023 9911
rect 12023 9877 12032 9911
rect 11980 9868 12032 9877
rect 14556 9911 14608 9920
rect 14556 9877 14565 9911
rect 14565 9877 14599 9911
rect 14599 9877 14608 9911
rect 14556 9868 14608 9877
rect 15936 9911 15988 9920
rect 15936 9877 15945 9911
rect 15945 9877 15979 9911
rect 15979 9877 15988 9911
rect 15936 9868 15988 9877
rect 16948 9868 17000 9920
rect 19064 10013 19073 10047
rect 19073 10013 19107 10047
rect 19107 10013 19116 10047
rect 19064 10004 19116 10013
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 1860 9664 1912 9716
rect 5264 9664 5316 9716
rect 1676 9596 1728 9648
rect 1952 9571 2004 9580
rect 1952 9537 1961 9571
rect 1961 9537 1995 9571
rect 1995 9537 2004 9571
rect 1952 9528 2004 9537
rect 2964 9528 3016 9580
rect 6736 9664 6788 9716
rect 1492 9460 1544 9512
rect 2780 9460 2832 9512
rect 3148 9460 3200 9512
rect 3792 9460 3844 9512
rect 7104 9664 7156 9716
rect 9680 9707 9732 9716
rect 9680 9673 9689 9707
rect 9689 9673 9723 9707
rect 9723 9673 9732 9707
rect 9680 9664 9732 9673
rect 8116 9596 8168 9648
rect 12624 9664 12676 9716
rect 12716 9664 12768 9716
rect 13268 9707 13320 9716
rect 13268 9673 13277 9707
rect 13277 9673 13311 9707
rect 13311 9673 13320 9707
rect 13268 9664 13320 9673
rect 19064 9707 19116 9716
rect 19064 9673 19073 9707
rect 19073 9673 19107 9707
rect 19107 9673 19116 9707
rect 19064 9664 19116 9673
rect 19340 9664 19392 9716
rect 20168 9664 20220 9716
rect 15384 9596 15436 9648
rect 16304 9639 16356 9648
rect 16304 9605 16313 9639
rect 16313 9605 16347 9639
rect 16347 9605 16356 9639
rect 16304 9596 16356 9605
rect 7932 9528 7984 9580
rect 9588 9528 9640 9580
rect 11336 9571 11388 9580
rect 11336 9537 11345 9571
rect 11345 9537 11379 9571
rect 11379 9537 11388 9571
rect 11336 9528 11388 9537
rect 2044 9392 2096 9444
rect 2228 9324 2280 9376
rect 4528 9324 4580 9376
rect 4988 9367 5040 9376
rect 4988 9333 4997 9367
rect 4997 9333 5031 9367
rect 5031 9333 5040 9367
rect 4988 9324 5040 9333
rect 6460 9324 6512 9376
rect 7472 9460 7524 9512
rect 13636 9460 13688 9512
rect 16028 9503 16080 9512
rect 16028 9469 16037 9503
rect 16037 9469 16071 9503
rect 16071 9469 16080 9503
rect 16028 9460 16080 9469
rect 18972 9596 19024 9648
rect 19432 9596 19484 9648
rect 16764 9528 16816 9580
rect 17960 9528 18012 9580
rect 18604 9571 18656 9580
rect 18604 9537 18613 9571
rect 18613 9537 18647 9571
rect 18647 9537 18656 9571
rect 18604 9528 18656 9537
rect 8300 9324 8352 9376
rect 10048 9324 10100 9376
rect 11612 9392 11664 9444
rect 13452 9392 13504 9444
rect 13912 9392 13964 9444
rect 17592 9460 17644 9512
rect 10784 9367 10836 9376
rect 10784 9333 10793 9367
rect 10793 9333 10827 9367
rect 10827 9333 10836 9367
rect 10784 9324 10836 9333
rect 10876 9324 10928 9376
rect 11704 9324 11756 9376
rect 12348 9324 12400 9376
rect 13636 9367 13688 9376
rect 13636 9333 13645 9367
rect 13645 9333 13679 9367
rect 13679 9333 13688 9367
rect 13636 9324 13688 9333
rect 17408 9367 17460 9376
rect 17408 9333 17417 9367
rect 17417 9333 17451 9367
rect 17451 9333 17460 9367
rect 17408 9324 17460 9333
rect 17776 9367 17828 9376
rect 17776 9333 17785 9367
rect 17785 9333 17819 9367
rect 17819 9333 17828 9367
rect 17776 9324 17828 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2964 9120 3016 9172
rect 5540 9120 5592 9172
rect 6552 9163 6604 9172
rect 6552 9129 6561 9163
rect 6561 9129 6595 9163
rect 6595 9129 6604 9163
rect 6552 9120 6604 9129
rect 8024 9163 8076 9172
rect 8024 9129 8033 9163
rect 8033 9129 8067 9163
rect 8067 9129 8076 9163
rect 8024 9120 8076 9129
rect 8392 9163 8444 9172
rect 8392 9129 8401 9163
rect 8401 9129 8435 9163
rect 8435 9129 8444 9163
rect 8392 9120 8444 9129
rect 8668 9120 8720 9172
rect 9772 9120 9824 9172
rect 10140 9163 10192 9172
rect 10140 9129 10149 9163
rect 10149 9129 10183 9163
rect 10183 9129 10192 9163
rect 10140 9120 10192 9129
rect 10784 9120 10836 9172
rect 12072 9120 12124 9172
rect 17408 9120 17460 9172
rect 18972 9163 19024 9172
rect 18972 9129 18981 9163
rect 18981 9129 19015 9163
rect 19015 9129 19024 9163
rect 18972 9120 19024 9129
rect 19340 9163 19392 9172
rect 19340 9129 19349 9163
rect 19349 9129 19383 9163
rect 19383 9129 19392 9163
rect 19340 9120 19392 9129
rect 2872 9052 2924 9104
rect 11060 9052 11112 9104
rect 14924 9095 14976 9104
rect 14924 9061 14933 9095
rect 14933 9061 14967 9095
rect 14967 9061 14976 9095
rect 14924 9052 14976 9061
rect 15936 9052 15988 9104
rect 16764 9052 16816 9104
rect 1492 9027 1544 9036
rect 1492 8993 1501 9027
rect 1501 8993 1535 9027
rect 1535 8993 1544 9027
rect 1492 8984 1544 8993
rect 5448 8984 5500 9036
rect 5540 8984 5592 9036
rect 6276 8984 6328 9036
rect 9588 8984 9640 9036
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 11336 8984 11388 9036
rect 11888 8984 11940 9036
rect 16028 8984 16080 9036
rect 16672 9027 16724 9036
rect 16672 8993 16681 9027
rect 16681 8993 16715 9027
rect 16715 8993 16724 9027
rect 16672 8984 16724 8993
rect 16948 9027 17000 9036
rect 16948 8993 16982 9027
rect 16982 8993 17000 9027
rect 16948 8984 17000 8993
rect 3240 8916 3292 8968
rect 3148 8848 3200 8900
rect 3884 8848 3936 8900
rect 8300 8848 8352 8900
rect 10968 8916 11020 8968
rect 11428 8916 11480 8968
rect 13820 8916 13872 8968
rect 14556 8959 14608 8968
rect 14556 8925 14565 8959
rect 14565 8925 14599 8959
rect 14599 8925 14608 8959
rect 14556 8916 14608 8925
rect 16488 8916 16540 8968
rect 6920 8823 6972 8832
rect 6920 8789 6929 8823
rect 6929 8789 6963 8823
rect 6963 8789 6972 8823
rect 6920 8780 6972 8789
rect 7196 8823 7248 8832
rect 7196 8789 7205 8823
rect 7205 8789 7239 8823
rect 7239 8789 7248 8823
rect 7196 8780 7248 8789
rect 7288 8780 7340 8832
rect 8208 8780 8260 8832
rect 8944 8780 8996 8832
rect 10876 8823 10928 8832
rect 10876 8789 10885 8823
rect 10885 8789 10919 8823
rect 10919 8789 10928 8823
rect 10876 8780 10928 8789
rect 13084 8780 13136 8832
rect 13912 8823 13964 8832
rect 13912 8789 13921 8823
rect 13921 8789 13955 8823
rect 13955 8789 13964 8823
rect 13912 8780 13964 8789
rect 17960 8780 18012 8832
rect 18604 8823 18656 8832
rect 18604 8789 18613 8823
rect 18613 8789 18647 8823
rect 18647 8789 18656 8823
rect 18604 8780 18656 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2504 8576 2556 8628
rect 8300 8576 8352 8628
rect 10968 8576 11020 8628
rect 11428 8576 11480 8628
rect 11888 8576 11940 8628
rect 13636 8576 13688 8628
rect 13912 8576 13964 8628
rect 16672 8576 16724 8628
rect 18052 8576 18104 8628
rect 1768 8440 1820 8492
rect 3148 8483 3200 8492
rect 3148 8449 3157 8483
rect 3157 8449 3191 8483
rect 3191 8449 3200 8483
rect 3148 8440 3200 8449
rect 3240 8483 3292 8492
rect 3240 8449 3249 8483
rect 3249 8449 3283 8483
rect 3283 8449 3292 8483
rect 6644 8483 6696 8492
rect 3240 8440 3292 8449
rect 6644 8449 6653 8483
rect 6653 8449 6687 8483
rect 6687 8449 6696 8483
rect 6644 8440 6696 8449
rect 4528 8415 4580 8424
rect 2596 8347 2648 8356
rect 2596 8313 2605 8347
rect 2605 8313 2639 8347
rect 2639 8313 2648 8347
rect 2596 8304 2648 8313
rect 3608 8304 3660 8356
rect 4528 8381 4562 8415
rect 4562 8381 4580 8415
rect 4528 8372 4580 8381
rect 6276 8415 6328 8424
rect 6276 8381 6285 8415
rect 6285 8381 6319 8415
rect 6319 8381 6328 8415
rect 6276 8372 6328 8381
rect 6736 8372 6788 8424
rect 7196 8440 7248 8492
rect 10876 8440 10928 8492
rect 16396 8508 16448 8560
rect 15844 8440 15896 8492
rect 18696 8483 18748 8492
rect 18696 8449 18705 8483
rect 18705 8449 18739 8483
rect 18739 8449 18748 8483
rect 18696 8440 18748 8449
rect 9496 8372 9548 8424
rect 15936 8415 15988 8424
rect 15936 8381 15945 8415
rect 15945 8381 15979 8415
rect 15979 8381 15988 8415
rect 15936 8372 15988 8381
rect 17776 8372 17828 8424
rect 2228 8236 2280 8288
rect 2780 8236 2832 8288
rect 4620 8236 4672 8288
rect 6184 8236 6236 8288
rect 6920 8304 6972 8356
rect 7748 8304 7800 8356
rect 9128 8304 9180 8356
rect 13084 8304 13136 8356
rect 16488 8347 16540 8356
rect 16488 8313 16497 8347
rect 16497 8313 16531 8347
rect 16531 8313 16540 8347
rect 16488 8304 16540 8313
rect 18420 8347 18472 8356
rect 18420 8313 18429 8347
rect 18429 8313 18463 8347
rect 18463 8313 18472 8347
rect 18420 8304 18472 8313
rect 11152 8279 11204 8288
rect 11152 8245 11161 8279
rect 11161 8245 11195 8279
rect 11195 8245 11204 8279
rect 11152 8236 11204 8245
rect 15844 8236 15896 8288
rect 18052 8279 18104 8288
rect 18052 8245 18061 8279
rect 18061 8245 18095 8279
rect 18095 8245 18104 8279
rect 18052 8236 18104 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 2044 8032 2096 8084
rect 3148 8032 3200 8084
rect 4620 8032 4672 8084
rect 7472 8075 7524 8084
rect 7472 8041 7481 8075
rect 7481 8041 7515 8075
rect 7515 8041 7524 8075
rect 7472 8032 7524 8041
rect 8300 8032 8352 8084
rect 9772 8032 9824 8084
rect 9128 7964 9180 8016
rect 11336 8032 11388 8084
rect 11704 8075 11756 8084
rect 11704 8041 11713 8075
rect 11713 8041 11747 8075
rect 11747 8041 11756 8075
rect 11704 8032 11756 8041
rect 12072 8075 12124 8084
rect 12072 8041 12081 8075
rect 12081 8041 12115 8075
rect 12115 8041 12124 8075
rect 12072 8032 12124 8041
rect 13176 8032 13228 8084
rect 13728 8032 13780 8084
rect 16396 8075 16448 8084
rect 16396 8041 16405 8075
rect 16405 8041 16439 8075
rect 16439 8041 16448 8075
rect 16396 8032 16448 8041
rect 16948 8032 17000 8084
rect 17592 8075 17644 8084
rect 17592 8041 17601 8075
rect 17601 8041 17635 8075
rect 17635 8041 17644 8075
rect 17592 8032 17644 8041
rect 2228 7896 2280 7948
rect 2780 7896 2832 7948
rect 6000 7896 6052 7948
rect 7564 7896 7616 7948
rect 9220 7896 9272 7948
rect 9772 7896 9824 7948
rect 2044 7871 2096 7880
rect 2044 7837 2053 7871
rect 2053 7837 2087 7871
rect 2087 7837 2096 7871
rect 2044 7828 2096 7837
rect 4344 7828 4396 7880
rect 4528 7871 4580 7880
rect 4528 7837 4537 7871
rect 4537 7837 4571 7871
rect 4571 7837 4580 7871
rect 4528 7828 4580 7837
rect 4804 7828 4856 7880
rect 8576 7871 8628 7880
rect 1584 7692 1636 7744
rect 3516 7735 3568 7744
rect 3516 7701 3525 7735
rect 3525 7701 3559 7735
rect 3559 7701 3568 7735
rect 3516 7692 3568 7701
rect 3976 7692 4028 7744
rect 5540 7735 5592 7744
rect 5540 7701 5549 7735
rect 5549 7701 5583 7735
rect 5583 7701 5592 7735
rect 5540 7692 5592 7701
rect 6000 7692 6052 7744
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 8576 7828 8628 7837
rect 10140 7871 10192 7880
rect 10140 7837 10149 7871
rect 10149 7837 10183 7871
rect 10183 7837 10192 7871
rect 10140 7828 10192 7837
rect 17776 7964 17828 8016
rect 13268 7896 13320 7948
rect 17960 7939 18012 7948
rect 17960 7905 17969 7939
rect 17969 7905 18003 7939
rect 18003 7905 18012 7939
rect 17960 7896 18012 7905
rect 11152 7828 11204 7880
rect 12256 7871 12308 7880
rect 12256 7837 12265 7871
rect 12265 7837 12299 7871
rect 12299 7837 12308 7871
rect 13084 7871 13136 7880
rect 12256 7828 12308 7837
rect 13084 7837 13093 7871
rect 13093 7837 13127 7871
rect 13127 7837 13136 7871
rect 13912 7871 13964 7880
rect 13084 7828 13136 7837
rect 13912 7837 13921 7871
rect 13921 7837 13955 7871
rect 13955 7837 13964 7871
rect 13912 7828 13964 7837
rect 15660 7828 15712 7880
rect 16764 7828 16816 7880
rect 17868 7828 17920 7880
rect 18604 7828 18656 7880
rect 8760 7760 8812 7812
rect 9680 7803 9732 7812
rect 9680 7769 9689 7803
rect 9689 7769 9723 7803
rect 9723 7769 9732 7803
rect 9680 7760 9732 7769
rect 10968 7760 11020 7812
rect 6368 7692 6420 7744
rect 8392 7735 8444 7744
rect 8392 7701 8401 7735
rect 8401 7701 8435 7735
rect 8435 7701 8444 7735
rect 8392 7692 8444 7701
rect 8484 7692 8536 7744
rect 11244 7735 11296 7744
rect 11244 7701 11253 7735
rect 11253 7701 11287 7735
rect 11287 7701 11296 7735
rect 11244 7692 11296 7701
rect 11428 7692 11480 7744
rect 14188 7692 14240 7744
rect 15752 7735 15804 7744
rect 15752 7701 15761 7735
rect 15761 7701 15795 7735
rect 15795 7701 15804 7735
rect 15752 7692 15804 7701
rect 16396 7760 16448 7812
rect 18328 7760 18380 7812
rect 16580 7692 16632 7744
rect 18604 7735 18656 7744
rect 18604 7701 18613 7735
rect 18613 7701 18647 7735
rect 18647 7701 18656 7735
rect 18604 7692 18656 7701
rect 20076 7692 20128 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 2136 7488 2188 7540
rect 2964 7531 3016 7540
rect 2964 7497 2973 7531
rect 2973 7497 3007 7531
rect 3007 7497 3016 7531
rect 2964 7488 3016 7497
rect 572 7420 624 7472
rect 8576 7488 8628 7540
rect 8668 7531 8720 7540
rect 8668 7497 8677 7531
rect 8677 7497 8711 7531
rect 8711 7497 8720 7531
rect 8668 7488 8720 7497
rect 11152 7488 11204 7540
rect 12256 7488 12308 7540
rect 13728 7488 13780 7540
rect 13912 7488 13964 7540
rect 15476 7531 15528 7540
rect 15476 7497 15485 7531
rect 15485 7497 15519 7531
rect 15519 7497 15528 7531
rect 15476 7488 15528 7497
rect 15660 7531 15712 7540
rect 15660 7497 15669 7531
rect 15669 7497 15703 7531
rect 15703 7497 15712 7531
rect 15660 7488 15712 7497
rect 1676 7352 1728 7404
rect 2044 7395 2096 7404
rect 2044 7361 2053 7395
rect 2053 7361 2087 7395
rect 2087 7361 2096 7395
rect 2044 7352 2096 7361
rect 2504 7352 2556 7404
rect 3424 7395 3476 7404
rect 3424 7361 3433 7395
rect 3433 7361 3467 7395
rect 3467 7361 3476 7395
rect 3424 7352 3476 7361
rect 3608 7395 3660 7404
rect 3608 7361 3617 7395
rect 3617 7361 3651 7395
rect 3651 7361 3660 7395
rect 3608 7352 3660 7361
rect 3700 7284 3752 7336
rect 9128 7420 9180 7472
rect 10140 7463 10192 7472
rect 5816 7395 5868 7404
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 6920 7352 6972 7404
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 7472 7395 7524 7404
rect 7472 7361 7481 7395
rect 7481 7361 7515 7395
rect 7515 7361 7524 7395
rect 7472 7352 7524 7361
rect 10140 7429 10149 7463
rect 10149 7429 10183 7463
rect 10183 7429 10192 7463
rect 10140 7420 10192 7429
rect 12348 7420 12400 7472
rect 15292 7420 15344 7472
rect 9772 7395 9824 7404
rect 9772 7361 9781 7395
rect 9781 7361 9815 7395
rect 9815 7361 9824 7395
rect 9772 7352 9824 7361
rect 10968 7352 11020 7404
rect 11336 7395 11388 7404
rect 11336 7361 11345 7395
rect 11345 7361 11379 7395
rect 11379 7361 11388 7395
rect 11336 7352 11388 7361
rect 12440 7395 12492 7404
rect 12440 7361 12449 7395
rect 12449 7361 12483 7395
rect 12483 7361 12492 7395
rect 13176 7395 13228 7404
rect 12440 7352 12492 7361
rect 13176 7361 13185 7395
rect 13185 7361 13219 7395
rect 13219 7361 13228 7395
rect 14096 7395 14148 7404
rect 13176 7352 13228 7361
rect 14096 7361 14105 7395
rect 14105 7361 14139 7395
rect 14139 7361 14148 7395
rect 14096 7352 14148 7361
rect 14280 7395 14332 7404
rect 14280 7361 14289 7395
rect 14289 7361 14323 7395
rect 14323 7361 14332 7395
rect 14280 7352 14332 7361
rect 14464 7352 14516 7404
rect 15108 7352 15160 7404
rect 15844 7352 15896 7404
rect 16304 7395 16356 7404
rect 16304 7361 16313 7395
rect 16313 7361 16347 7395
rect 16347 7361 16356 7395
rect 16304 7352 16356 7361
rect 8484 7284 8536 7336
rect 8576 7284 8628 7336
rect 10876 7284 10928 7336
rect 15476 7284 15528 7336
rect 17960 7284 18012 7336
rect 18328 7420 18380 7472
rect 18512 7395 18564 7404
rect 18512 7361 18521 7395
rect 18521 7361 18555 7395
rect 18555 7361 18564 7395
rect 18512 7352 18564 7361
rect 20536 7420 20588 7472
rect 18788 7352 18840 7404
rect 19340 7352 19392 7404
rect 18420 7327 18472 7336
rect 18420 7293 18429 7327
rect 18429 7293 18463 7327
rect 18463 7293 18472 7327
rect 18420 7284 18472 7293
rect 1768 7259 1820 7268
rect 1768 7225 1777 7259
rect 1777 7225 1811 7259
rect 1811 7225 1820 7259
rect 1768 7216 1820 7225
rect 5632 7259 5684 7268
rect 5632 7225 5641 7259
rect 5641 7225 5675 7259
rect 5675 7225 5684 7259
rect 5632 7216 5684 7225
rect 6092 7216 6144 7268
rect 9588 7216 9640 7268
rect 11060 7216 11112 7268
rect 14004 7259 14056 7268
rect 14004 7225 14013 7259
rect 14013 7225 14047 7259
rect 14047 7225 14056 7259
rect 14004 7216 14056 7225
rect 14464 7216 14516 7268
rect 1400 7191 1452 7200
rect 1400 7157 1409 7191
rect 1409 7157 1443 7191
rect 1443 7157 1452 7191
rect 1400 7148 1452 7157
rect 2872 7148 2924 7200
rect 4804 7148 4856 7200
rect 5540 7191 5592 7200
rect 5540 7157 5549 7191
rect 5549 7157 5583 7191
rect 5583 7157 5592 7191
rect 5540 7148 5592 7157
rect 6000 7148 6052 7200
rect 6368 7148 6420 7200
rect 6828 7191 6880 7200
rect 6828 7157 6837 7191
rect 6837 7157 6871 7191
rect 6871 7157 6880 7191
rect 6828 7148 6880 7157
rect 9864 7148 9916 7200
rect 11336 7148 11388 7200
rect 14096 7148 14148 7200
rect 14372 7148 14424 7200
rect 15752 7148 15804 7200
rect 17868 7216 17920 7268
rect 16764 7191 16816 7200
rect 16764 7157 16773 7191
rect 16773 7157 16807 7191
rect 16807 7157 16816 7191
rect 16764 7148 16816 7157
rect 18512 7216 18564 7268
rect 19984 7191 20036 7200
rect 19984 7157 19993 7191
rect 19993 7157 20027 7191
rect 20027 7157 20036 7191
rect 19984 7148 20036 7157
rect 20076 7191 20128 7200
rect 20076 7157 20085 7191
rect 20085 7157 20119 7191
rect 20119 7157 20128 7191
rect 20076 7148 20128 7157
rect 20628 7148 20680 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 1768 6944 1820 6996
rect 3608 6944 3660 6996
rect 7380 6944 7432 6996
rect 8668 6944 8720 6996
rect 9128 6944 9180 6996
rect 9680 6987 9732 6996
rect 9680 6953 9689 6987
rect 9689 6953 9723 6987
rect 9723 6953 9732 6987
rect 9680 6944 9732 6953
rect 1676 6876 1728 6928
rect 3976 6876 4028 6928
rect 5816 6876 5868 6928
rect 10784 6944 10836 6996
rect 14280 6944 14332 6996
rect 16764 6944 16816 6996
rect 18420 6987 18472 6996
rect 18420 6953 18429 6987
rect 18429 6953 18463 6987
rect 18463 6953 18472 6987
rect 18420 6944 18472 6953
rect 19248 6987 19300 6996
rect 19248 6953 19257 6987
rect 19257 6953 19291 6987
rect 19291 6953 19300 6987
rect 19248 6944 19300 6953
rect 4068 6808 4120 6860
rect 4620 6808 4672 6860
rect 3056 6783 3108 6792
rect 3056 6749 3065 6783
rect 3065 6749 3099 6783
rect 3099 6749 3108 6783
rect 3056 6740 3108 6749
rect 3516 6740 3568 6792
rect 4252 6740 4304 6792
rect 2504 6672 2556 6724
rect 4804 6740 4856 6792
rect 5724 6672 5776 6724
rect 2228 6647 2280 6656
rect 2228 6613 2237 6647
rect 2237 6613 2271 6647
rect 2271 6613 2280 6647
rect 2228 6604 2280 6613
rect 2688 6604 2740 6656
rect 4068 6647 4120 6656
rect 4068 6613 4077 6647
rect 4077 6613 4111 6647
rect 4111 6613 4120 6647
rect 4068 6604 4120 6613
rect 5172 6647 5224 6656
rect 5172 6613 5181 6647
rect 5181 6613 5215 6647
rect 5215 6613 5224 6647
rect 5172 6604 5224 6613
rect 7380 6808 7432 6860
rect 8484 6851 8536 6860
rect 8484 6817 8493 6851
rect 8493 6817 8527 6851
rect 8527 6817 8536 6851
rect 8484 6808 8536 6817
rect 9404 6808 9456 6860
rect 11612 6851 11664 6860
rect 11612 6817 11621 6851
rect 11621 6817 11655 6851
rect 11655 6817 11664 6851
rect 16304 6876 16356 6928
rect 11612 6808 11664 6817
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 9036 6740 9088 6792
rect 10048 6740 10100 6792
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 10232 6740 10284 6749
rect 10784 6740 10836 6792
rect 11428 6740 11480 6792
rect 11888 6783 11940 6792
rect 11888 6749 11897 6783
rect 11897 6749 11931 6783
rect 11931 6749 11940 6783
rect 11888 6740 11940 6749
rect 13268 6783 13320 6792
rect 13268 6749 13277 6783
rect 13277 6749 13311 6783
rect 13311 6749 13320 6783
rect 13268 6740 13320 6749
rect 13452 6783 13504 6792
rect 13452 6749 13461 6783
rect 13461 6749 13495 6783
rect 13495 6749 13504 6783
rect 13452 6740 13504 6749
rect 14280 6808 14332 6860
rect 16488 6808 16540 6860
rect 16672 6851 16724 6860
rect 16672 6817 16706 6851
rect 16706 6817 16724 6851
rect 16672 6808 16724 6817
rect 16028 6740 16080 6792
rect 19340 6783 19392 6792
rect 19340 6749 19349 6783
rect 19349 6749 19383 6783
rect 19383 6749 19392 6783
rect 19340 6740 19392 6749
rect 19432 6783 19484 6792
rect 19432 6749 19441 6783
rect 19441 6749 19475 6783
rect 19475 6749 19484 6783
rect 19432 6740 19484 6749
rect 12808 6715 12860 6724
rect 12808 6681 12817 6715
rect 12817 6681 12851 6715
rect 12851 6681 12860 6715
rect 12808 6672 12860 6681
rect 20996 6672 21048 6724
rect 6000 6604 6052 6656
rect 7380 6647 7432 6656
rect 7380 6613 7389 6647
rect 7389 6613 7423 6647
rect 7423 6613 7432 6647
rect 7380 6604 7432 6613
rect 7932 6647 7984 6656
rect 7932 6613 7941 6647
rect 7941 6613 7975 6647
rect 7975 6613 7984 6647
rect 7932 6604 7984 6613
rect 8300 6647 8352 6656
rect 8300 6613 8309 6647
rect 8309 6613 8343 6647
rect 8343 6613 8352 6647
rect 8300 6604 8352 6613
rect 9772 6604 9824 6656
rect 10876 6604 10928 6656
rect 11244 6647 11296 6656
rect 11244 6613 11253 6647
rect 11253 6613 11287 6647
rect 11287 6613 11296 6647
rect 11244 6604 11296 6613
rect 12532 6647 12584 6656
rect 12532 6613 12541 6647
rect 12541 6613 12575 6647
rect 12575 6613 12584 6647
rect 12532 6604 12584 6613
rect 14280 6647 14332 6656
rect 14280 6613 14289 6647
rect 14289 6613 14323 6647
rect 14323 6613 14332 6647
rect 14280 6604 14332 6613
rect 14740 6604 14792 6656
rect 16212 6647 16264 6656
rect 16212 6613 16221 6647
rect 16221 6613 16255 6647
rect 16255 6613 16264 6647
rect 16212 6604 16264 6613
rect 18696 6647 18748 6656
rect 18696 6613 18705 6647
rect 18705 6613 18739 6647
rect 18739 6613 18748 6647
rect 18696 6604 18748 6613
rect 19984 6647 20036 6656
rect 19984 6613 19993 6647
rect 19993 6613 20027 6647
rect 20027 6613 20036 6647
rect 19984 6604 20036 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 4988 6443 5040 6452
rect 4988 6409 4997 6443
rect 4997 6409 5031 6443
rect 5031 6409 5040 6443
rect 4988 6400 5040 6409
rect 5448 6400 5500 6452
rect 6828 6443 6880 6452
rect 6828 6409 6837 6443
rect 6837 6409 6871 6443
rect 6871 6409 6880 6443
rect 6828 6400 6880 6409
rect 8392 6400 8444 6452
rect 9036 6443 9088 6452
rect 9036 6409 9045 6443
rect 9045 6409 9079 6443
rect 9079 6409 9088 6443
rect 9036 6400 9088 6409
rect 9404 6443 9456 6452
rect 9404 6409 9413 6443
rect 9413 6409 9447 6443
rect 9447 6409 9456 6443
rect 9404 6400 9456 6409
rect 10232 6400 10284 6452
rect 11888 6443 11940 6452
rect 11888 6409 11897 6443
rect 11897 6409 11931 6443
rect 11931 6409 11940 6443
rect 11888 6400 11940 6409
rect 6092 6332 6144 6384
rect 9128 6332 9180 6384
rect 4160 6264 4212 6316
rect 5172 6264 5224 6316
rect 6000 6264 6052 6316
rect 6460 6264 6512 6316
rect 7380 6264 7432 6316
rect 12532 6264 12584 6316
rect 13820 6264 13872 6316
rect 16028 6400 16080 6452
rect 16488 6400 16540 6452
rect 19984 6400 20036 6452
rect 19432 6375 19484 6384
rect 19432 6341 19441 6375
rect 19441 6341 19475 6375
rect 19475 6341 19484 6375
rect 19432 6332 19484 6341
rect 20996 6307 21048 6316
rect 20996 6273 21005 6307
rect 21005 6273 21039 6307
rect 21039 6273 21048 6307
rect 20996 6264 21048 6273
rect 21456 6264 21508 6316
rect 3056 6196 3108 6248
rect 4988 6196 5040 6248
rect 7104 6196 7156 6248
rect 7932 6196 7984 6248
rect 16856 6239 16908 6248
rect 16856 6205 16865 6239
rect 16865 6205 16899 6239
rect 16899 6205 16908 6239
rect 16856 6196 16908 6205
rect 18144 6196 18196 6248
rect 18696 6196 18748 6248
rect 20904 6239 20956 6248
rect 20904 6205 20913 6239
rect 20913 6205 20947 6239
rect 20947 6205 20956 6239
rect 20904 6196 20956 6205
rect 22284 6239 22336 6248
rect 22284 6205 22293 6239
rect 22293 6205 22327 6239
rect 22327 6205 22336 6239
rect 22284 6196 22336 6205
rect 2780 6128 2832 6180
rect 7196 6171 7248 6180
rect 7196 6137 7205 6171
rect 7205 6137 7239 6171
rect 7239 6137 7248 6171
rect 7196 6128 7248 6137
rect 8300 6128 8352 6180
rect 9772 6171 9824 6180
rect 9772 6137 9806 6171
rect 9806 6137 9824 6171
rect 9772 6128 9824 6137
rect 14648 6128 14700 6180
rect 17316 6128 17368 6180
rect 19340 6128 19392 6180
rect 1676 6103 1728 6112
rect 1676 6069 1685 6103
rect 1685 6069 1719 6103
rect 1719 6069 1728 6103
rect 1676 6060 1728 6069
rect 3792 6060 3844 6112
rect 4252 6103 4304 6112
rect 4252 6069 4261 6103
rect 4261 6069 4295 6103
rect 4295 6069 4304 6103
rect 4252 6060 4304 6069
rect 4620 6103 4672 6112
rect 4620 6069 4629 6103
rect 4629 6069 4663 6103
rect 4663 6069 4672 6103
rect 4620 6060 4672 6069
rect 5448 6060 5500 6112
rect 6092 6060 6144 6112
rect 6460 6060 6512 6112
rect 7288 6060 7340 6112
rect 9864 6060 9916 6112
rect 12164 6103 12216 6112
rect 12164 6069 12173 6103
rect 12173 6069 12207 6103
rect 12207 6069 12216 6103
rect 12164 6060 12216 6069
rect 12440 6103 12492 6112
rect 12440 6069 12449 6103
rect 12449 6069 12483 6103
rect 12483 6069 12492 6103
rect 12900 6103 12952 6112
rect 12440 6060 12492 6069
rect 12900 6069 12909 6103
rect 12909 6069 12943 6103
rect 12943 6069 12952 6103
rect 12900 6060 12952 6069
rect 13452 6103 13504 6112
rect 13452 6069 13461 6103
rect 13461 6069 13495 6103
rect 13495 6069 13504 6103
rect 13452 6060 13504 6069
rect 15200 6060 15252 6112
rect 16304 6060 16356 6112
rect 17040 6103 17092 6112
rect 17040 6069 17049 6103
rect 17049 6069 17083 6103
rect 17083 6069 17092 6103
rect 17040 6060 17092 6069
rect 22468 6103 22520 6112
rect 22468 6069 22477 6103
rect 22477 6069 22511 6103
rect 22511 6069 22520 6103
rect 22468 6060 22520 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 3056 5856 3108 5908
rect 4804 5856 4856 5908
rect 6184 5856 6236 5908
rect 6460 5899 6512 5908
rect 6460 5865 6469 5899
rect 6469 5865 6503 5899
rect 6503 5865 6512 5899
rect 6460 5856 6512 5865
rect 7196 5856 7248 5908
rect 7932 5899 7984 5908
rect 7932 5865 7941 5899
rect 7941 5865 7975 5899
rect 7975 5865 7984 5899
rect 7932 5856 7984 5865
rect 9772 5856 9824 5908
rect 13452 5856 13504 5908
rect 14648 5856 14700 5908
rect 18144 5899 18196 5908
rect 18144 5865 18153 5899
rect 18153 5865 18187 5899
rect 18187 5865 18196 5899
rect 18144 5856 18196 5865
rect 19248 5856 19300 5908
rect 19524 5856 19576 5908
rect 20720 5856 20772 5908
rect 1768 5788 1820 5840
rect 1676 5763 1728 5772
rect 1676 5729 1710 5763
rect 1710 5729 1728 5763
rect 1676 5720 1728 5729
rect 2412 5720 2464 5772
rect 2780 5720 2832 5772
rect 4160 5720 4212 5772
rect 4344 5763 4396 5772
rect 4344 5729 4378 5763
rect 4378 5729 4396 5763
rect 4344 5720 4396 5729
rect 6920 5763 6972 5772
rect 6920 5729 6929 5763
rect 6929 5729 6963 5763
rect 6963 5729 6972 5763
rect 6920 5720 6972 5729
rect 8300 5763 8352 5772
rect 8300 5729 8309 5763
rect 8309 5729 8343 5763
rect 8343 5729 8352 5763
rect 8300 5720 8352 5729
rect 9128 5720 9180 5772
rect 10692 5720 10744 5772
rect 12348 5788 12400 5840
rect 16120 5788 16172 5840
rect 16764 5788 16816 5840
rect 19432 5788 19484 5840
rect 21456 5788 21508 5840
rect 12072 5720 12124 5772
rect 12992 5720 13044 5772
rect 15660 5763 15712 5772
rect 15660 5729 15669 5763
rect 15669 5729 15703 5763
rect 15703 5729 15712 5763
rect 15660 5720 15712 5729
rect 19984 5720 20036 5772
rect 20720 5720 20772 5772
rect 22008 5720 22060 5772
rect 22468 5720 22520 5772
rect 23296 5763 23348 5772
rect 23296 5729 23305 5763
rect 23305 5729 23339 5763
rect 23339 5729 23348 5763
rect 23296 5720 23348 5729
rect 3148 5584 3200 5636
rect 6920 5584 6972 5636
rect 7288 5652 7340 5704
rect 8576 5695 8628 5704
rect 8576 5661 8585 5695
rect 8585 5661 8619 5695
rect 8619 5661 8628 5695
rect 8576 5652 8628 5661
rect 10876 5652 10928 5704
rect 11612 5652 11664 5704
rect 16488 5652 16540 5704
rect 19340 5652 19392 5704
rect 19800 5695 19852 5704
rect 19800 5661 19809 5695
rect 19809 5661 19843 5695
rect 19843 5661 19852 5695
rect 19800 5652 19852 5661
rect 9036 5627 9088 5636
rect 9036 5593 9045 5627
rect 9045 5593 9079 5627
rect 9079 5593 9088 5627
rect 9036 5584 9088 5593
rect 13728 5584 13780 5636
rect 15844 5627 15896 5636
rect 15844 5593 15853 5627
rect 15853 5593 15887 5627
rect 15887 5593 15896 5627
rect 15844 5584 15896 5593
rect 21456 5695 21508 5704
rect 21456 5661 21465 5695
rect 21465 5661 21499 5695
rect 21499 5661 21508 5695
rect 21456 5652 21508 5661
rect 21548 5584 21600 5636
rect 3700 5559 3752 5568
rect 3700 5525 3709 5559
rect 3709 5525 3743 5559
rect 3743 5525 3752 5559
rect 3700 5516 3752 5525
rect 3792 5516 3844 5568
rect 7564 5559 7616 5568
rect 7564 5525 7573 5559
rect 7573 5525 7607 5559
rect 7607 5525 7616 5559
rect 7564 5516 7616 5525
rect 9404 5516 9456 5568
rect 9864 5516 9916 5568
rect 13268 5516 13320 5568
rect 13452 5516 13504 5568
rect 13636 5516 13688 5568
rect 15384 5516 15436 5568
rect 16672 5516 16724 5568
rect 23480 5559 23532 5568
rect 23480 5525 23489 5559
rect 23489 5525 23523 5559
rect 23523 5525 23532 5559
rect 23480 5516 23532 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 2412 5355 2464 5364
rect 2412 5321 2421 5355
rect 2421 5321 2455 5355
rect 2455 5321 2464 5355
rect 2412 5312 2464 5321
rect 2780 5244 2832 5296
rect 1584 5176 1636 5228
rect 3056 5312 3108 5364
rect 3792 5312 3844 5364
rect 4160 5312 4212 5364
rect 6092 5312 6144 5364
rect 9128 5355 9180 5364
rect 9128 5321 9137 5355
rect 9137 5321 9171 5355
rect 9171 5321 9180 5355
rect 9128 5312 9180 5321
rect 12992 5355 13044 5364
rect 12992 5321 13001 5355
rect 13001 5321 13035 5355
rect 13035 5321 13044 5355
rect 12992 5312 13044 5321
rect 14648 5312 14700 5364
rect 16488 5312 16540 5364
rect 17408 5355 17460 5364
rect 17408 5321 17417 5355
rect 17417 5321 17451 5355
rect 17451 5321 17460 5355
rect 17408 5312 17460 5321
rect 18236 5312 18288 5364
rect 20720 5312 20772 5364
rect 21456 5312 21508 5364
rect 22100 5355 22152 5364
rect 22100 5321 22109 5355
rect 22109 5321 22143 5355
rect 22143 5321 22152 5355
rect 23296 5355 23348 5364
rect 22100 5312 22152 5321
rect 23296 5321 23305 5355
rect 23305 5321 23339 5355
rect 23339 5321 23348 5355
rect 23296 5312 23348 5321
rect 3700 5176 3752 5228
rect 6184 5244 6236 5296
rect 6368 5244 6420 5296
rect 1400 5108 1452 5160
rect 4160 5108 4212 5160
rect 5448 5108 5500 5160
rect 6184 5108 6236 5160
rect 6828 5244 6880 5296
rect 12072 5244 12124 5296
rect 6828 5151 6880 5160
rect 6828 5117 6837 5151
rect 6837 5117 6871 5151
rect 6871 5117 6880 5151
rect 6828 5108 6880 5117
rect 7564 5108 7616 5160
rect 9128 5108 9180 5160
rect 9588 5151 9640 5160
rect 9588 5117 9622 5151
rect 9622 5117 9640 5151
rect 9588 5108 9640 5117
rect 6736 5040 6788 5092
rect 9956 5040 10008 5092
rect 18144 5244 18196 5296
rect 19524 5244 19576 5296
rect 22376 5287 22428 5296
rect 22376 5253 22385 5287
rect 22385 5253 22419 5287
rect 22419 5253 22428 5287
rect 22376 5244 22428 5253
rect 17776 5219 17828 5228
rect 17776 5185 17785 5219
rect 17785 5185 17819 5219
rect 17819 5185 17828 5219
rect 18604 5219 18656 5228
rect 17776 5176 17828 5185
rect 12348 5108 12400 5160
rect 12532 5151 12584 5160
rect 12532 5117 12541 5151
rect 12541 5117 12575 5151
rect 12575 5117 12584 5151
rect 12532 5108 12584 5117
rect 15660 5151 15712 5160
rect 15660 5117 15669 5151
rect 15669 5117 15703 5151
rect 15703 5117 15712 5151
rect 15660 5108 15712 5117
rect 16580 5108 16632 5160
rect 18604 5185 18613 5219
rect 18613 5185 18647 5219
rect 18647 5185 18656 5219
rect 18604 5176 18656 5185
rect 19800 5176 19852 5228
rect 20260 5176 20312 5228
rect 18512 5151 18564 5160
rect 18512 5117 18521 5151
rect 18521 5117 18555 5151
rect 18555 5117 18564 5151
rect 18512 5108 18564 5117
rect 20720 5108 20772 5160
rect 21824 5108 21876 5160
rect 22744 5151 22796 5160
rect 22744 5117 22753 5151
rect 22753 5117 22787 5151
rect 22787 5117 22796 5151
rect 22744 5108 22796 5117
rect 13636 5040 13688 5092
rect 16488 5040 16540 5092
rect 16856 5083 16908 5092
rect 16856 5049 16865 5083
rect 16865 5049 16899 5083
rect 16899 5049 16908 5083
rect 16856 5040 16908 5049
rect 3608 5015 3660 5024
rect 3608 4981 3617 5015
rect 3617 4981 3651 5015
rect 3651 4981 3660 5015
rect 3608 4972 3660 4981
rect 3884 4972 3936 5024
rect 5172 5015 5224 5024
rect 5172 4981 5181 5015
rect 5181 4981 5215 5015
rect 5215 4981 5224 5015
rect 5172 4972 5224 4981
rect 5540 5015 5592 5024
rect 5540 4981 5549 5015
rect 5549 4981 5583 5015
rect 5583 4981 5592 5015
rect 5540 4972 5592 4981
rect 5632 5015 5684 5024
rect 5632 4981 5641 5015
rect 5641 4981 5675 5015
rect 5675 4981 5684 5015
rect 6276 5015 6328 5024
rect 5632 4972 5684 4981
rect 6276 4981 6285 5015
rect 6285 4981 6319 5015
rect 6319 4981 6328 5015
rect 6276 4972 6328 4981
rect 8024 4972 8076 5024
rect 10692 5015 10744 5024
rect 10692 4981 10701 5015
rect 10701 4981 10735 5015
rect 10735 4981 10744 5015
rect 10692 4972 10744 4981
rect 11152 4972 11204 5024
rect 12716 5015 12768 5024
rect 12716 4981 12725 5015
rect 12725 4981 12759 5015
rect 12759 4981 12768 5015
rect 12716 4972 12768 4981
rect 12808 4972 12860 5024
rect 13084 4972 13136 5024
rect 16396 5015 16448 5024
rect 16396 4981 16405 5015
rect 16405 4981 16439 5015
rect 16439 4981 16448 5015
rect 16396 4972 16448 4981
rect 18972 4972 19024 5024
rect 19340 4972 19392 5024
rect 21364 5015 21416 5024
rect 21364 4981 21373 5015
rect 21373 4981 21407 5015
rect 21407 4981 21416 5015
rect 21364 4972 21416 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1768 4768 1820 4820
rect 2964 4768 3016 4820
rect 4160 4768 4212 4820
rect 4344 4811 4396 4820
rect 4344 4777 4353 4811
rect 4353 4777 4387 4811
rect 4387 4777 4396 4811
rect 4344 4768 4396 4777
rect 5172 4768 5224 4820
rect 6000 4811 6052 4820
rect 6000 4777 6009 4811
rect 6009 4777 6043 4811
rect 6043 4777 6052 4811
rect 6000 4768 6052 4777
rect 6828 4768 6880 4820
rect 7104 4811 7156 4820
rect 7104 4777 7113 4811
rect 7113 4777 7147 4811
rect 7147 4777 7156 4811
rect 7104 4768 7156 4777
rect 9128 4768 9180 4820
rect 10968 4811 11020 4820
rect 10968 4777 10977 4811
rect 10977 4777 11011 4811
rect 11011 4777 11020 4811
rect 10968 4768 11020 4777
rect 11336 4768 11388 4820
rect 11888 4768 11940 4820
rect 2780 4743 2832 4752
rect 2780 4709 2789 4743
rect 2789 4709 2823 4743
rect 2823 4709 2832 4743
rect 2780 4700 2832 4709
rect 4436 4700 4488 4752
rect 5356 4700 5408 4752
rect 6092 4700 6144 4752
rect 10508 4743 10560 4752
rect 10508 4709 10517 4743
rect 10517 4709 10551 4743
rect 10551 4709 10560 4743
rect 10508 4700 10560 4709
rect 10692 4700 10744 4752
rect 5540 4632 5592 4684
rect 6828 4632 6880 4684
rect 7196 4632 7248 4684
rect 7748 4632 7800 4684
rect 9956 4675 10008 4684
rect 9956 4641 9965 4675
rect 9965 4641 9999 4675
rect 9999 4641 10008 4675
rect 9956 4632 10008 4641
rect 10048 4632 10100 4684
rect 11704 4632 11756 4684
rect 12440 4768 12492 4820
rect 16120 4811 16172 4820
rect 16120 4777 16129 4811
rect 16129 4777 16163 4811
rect 16163 4777 16172 4811
rect 16120 4768 16172 4777
rect 16212 4768 16264 4820
rect 16948 4811 17000 4820
rect 16948 4777 16957 4811
rect 16957 4777 16991 4811
rect 16991 4777 17000 4811
rect 16948 4768 17000 4777
rect 18144 4768 18196 4820
rect 20260 4811 20312 4820
rect 20260 4777 20269 4811
rect 20269 4777 20303 4811
rect 20303 4777 20312 4811
rect 20260 4768 20312 4777
rect 21548 4811 21600 4820
rect 21548 4777 21557 4811
rect 21557 4777 21591 4811
rect 21591 4777 21600 4811
rect 21548 4768 21600 4777
rect 21824 4811 21876 4820
rect 21824 4777 21833 4811
rect 21833 4777 21867 4811
rect 21867 4777 21876 4811
rect 21824 4768 21876 4777
rect 12992 4743 13044 4752
rect 12992 4709 13001 4743
rect 13001 4709 13035 4743
rect 13035 4709 13044 4743
rect 12992 4700 13044 4709
rect 13728 4700 13780 4752
rect 19984 4700 20036 4752
rect 2964 4607 3016 4616
rect 2964 4573 2973 4607
rect 2973 4573 3007 4607
rect 3007 4573 3016 4607
rect 2964 4564 3016 4573
rect 6092 4607 6144 4616
rect 6092 4573 6101 4607
rect 6101 4573 6135 4607
rect 6135 4573 6144 4607
rect 6092 4564 6144 4573
rect 7564 4607 7616 4616
rect 7564 4573 7573 4607
rect 7573 4573 7607 4607
rect 7607 4573 7616 4607
rect 7564 4564 7616 4573
rect 2412 4539 2464 4548
rect 2412 4505 2421 4539
rect 2421 4505 2455 4539
rect 2455 4505 2464 4539
rect 2412 4496 2464 4505
rect 5632 4496 5684 4548
rect 6736 4496 6788 4548
rect 7288 4496 7340 4548
rect 10140 4564 10192 4616
rect 10692 4564 10744 4616
rect 11612 4607 11664 4616
rect 11612 4573 11621 4607
rect 11621 4573 11655 4607
rect 11655 4573 11664 4607
rect 12716 4632 12768 4684
rect 14648 4632 14700 4684
rect 15292 4675 15344 4684
rect 15292 4641 15301 4675
rect 15301 4641 15335 4675
rect 15335 4641 15344 4675
rect 15292 4632 15344 4641
rect 16856 4675 16908 4684
rect 16856 4641 16865 4675
rect 16865 4641 16899 4675
rect 16899 4641 16908 4675
rect 16856 4632 16908 4641
rect 17500 4675 17552 4684
rect 17500 4641 17509 4675
rect 17509 4641 17543 4675
rect 17543 4641 17552 4675
rect 17500 4632 17552 4641
rect 13084 4607 13136 4616
rect 11612 4564 11664 4573
rect 4620 4471 4672 4480
rect 4620 4437 4629 4471
rect 4629 4437 4663 4471
rect 4663 4437 4672 4471
rect 4620 4428 4672 4437
rect 5540 4471 5592 4480
rect 5540 4437 5549 4471
rect 5549 4437 5583 4471
rect 5583 4437 5592 4471
rect 5540 4428 5592 4437
rect 8116 4471 8168 4480
rect 8116 4437 8125 4471
rect 8125 4437 8159 4471
rect 8159 4437 8168 4471
rect 8116 4428 8168 4437
rect 8300 4428 8352 4480
rect 8852 4471 8904 4480
rect 8852 4437 8861 4471
rect 8861 4437 8895 4471
rect 8895 4437 8904 4471
rect 8852 4428 8904 4437
rect 10968 4428 11020 4480
rect 13084 4573 13093 4607
rect 13093 4573 13127 4607
rect 13127 4573 13136 4607
rect 13084 4564 13136 4573
rect 13636 4607 13688 4616
rect 13636 4573 13645 4607
rect 13645 4573 13679 4607
rect 13679 4573 13688 4607
rect 13636 4564 13688 4573
rect 13728 4564 13780 4616
rect 16580 4564 16632 4616
rect 17684 4564 17736 4616
rect 14372 4496 14424 4548
rect 15476 4539 15528 4548
rect 15476 4505 15485 4539
rect 15485 4505 15519 4539
rect 15519 4505 15528 4539
rect 15476 4496 15528 4505
rect 18052 4632 18104 4684
rect 19524 4632 19576 4684
rect 21364 4632 21416 4684
rect 18512 4607 18564 4616
rect 18512 4573 18521 4607
rect 18521 4573 18555 4607
rect 18555 4573 18564 4607
rect 18512 4564 18564 4573
rect 18604 4607 18656 4616
rect 18604 4573 18613 4607
rect 18613 4573 18647 4607
rect 18647 4573 18656 4607
rect 18604 4564 18656 4573
rect 21272 4496 21324 4548
rect 13268 4428 13320 4480
rect 17500 4428 17552 4480
rect 18328 4428 18380 4480
rect 20536 4471 20588 4480
rect 20536 4437 20545 4471
rect 20545 4437 20579 4471
rect 20579 4437 20588 4471
rect 20536 4428 20588 4437
rect 20812 4428 20864 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 3792 4267 3844 4276
rect 3792 4233 3801 4267
rect 3801 4233 3835 4267
rect 3835 4233 3844 4267
rect 3792 4224 3844 4233
rect 6000 4224 6052 4276
rect 7564 4267 7616 4276
rect 7564 4233 7573 4267
rect 7573 4233 7607 4267
rect 7607 4233 7616 4267
rect 7564 4224 7616 4233
rect 2964 4131 3016 4140
rect 2964 4097 2973 4131
rect 2973 4097 3007 4131
rect 3007 4097 3016 4131
rect 2964 4088 3016 4097
rect 7288 4156 7340 4208
rect 8116 4156 8168 4208
rect 9772 4088 9824 4140
rect 9956 4224 10008 4276
rect 11612 4224 11664 4276
rect 11704 4267 11756 4276
rect 11704 4233 11713 4267
rect 11713 4233 11747 4267
rect 11747 4233 11756 4267
rect 11704 4224 11756 4233
rect 12532 4224 12584 4276
rect 15292 4267 15344 4276
rect 15292 4233 15301 4267
rect 15301 4233 15335 4267
rect 15335 4233 15344 4267
rect 15292 4224 15344 4233
rect 16120 4224 16172 4276
rect 11152 4156 11204 4208
rect 16212 4156 16264 4208
rect 2412 3952 2464 4004
rect 3608 3952 3660 4004
rect 6000 4020 6052 4072
rect 7472 4020 7524 4072
rect 8208 4020 8260 4072
rect 8576 4020 8628 4072
rect 12164 4088 12216 4140
rect 12808 4088 12860 4140
rect 11336 4020 11388 4072
rect 13268 4088 13320 4140
rect 14004 4088 14056 4140
rect 18512 4224 18564 4276
rect 20536 4224 20588 4276
rect 21364 4224 21416 4276
rect 18788 4088 18840 4140
rect 19524 4156 19576 4208
rect 20260 4131 20312 4140
rect 20260 4097 20269 4131
rect 20269 4097 20303 4131
rect 20303 4097 20312 4131
rect 20260 4088 20312 4097
rect 13544 4020 13596 4072
rect 14372 4063 14424 4072
rect 14372 4029 14381 4063
rect 14381 4029 14415 4063
rect 14415 4029 14424 4063
rect 14372 4020 14424 4029
rect 14740 4020 14792 4072
rect 15476 4020 15528 4072
rect 4252 3952 4304 4004
rect 4896 3952 4948 4004
rect 6092 3952 6144 4004
rect 2320 3927 2372 3936
rect 2320 3893 2329 3927
rect 2329 3893 2363 3927
rect 2363 3893 2372 3927
rect 2320 3884 2372 3893
rect 2688 3927 2740 3936
rect 2688 3893 2697 3927
rect 2697 3893 2731 3927
rect 2731 3893 2740 3927
rect 2688 3884 2740 3893
rect 4344 3884 4396 3936
rect 7196 3927 7248 3936
rect 7196 3893 7205 3927
rect 7205 3893 7239 3927
rect 7239 3893 7248 3927
rect 7196 3884 7248 3893
rect 7748 3927 7800 3936
rect 7748 3893 7757 3927
rect 7757 3893 7791 3927
rect 7791 3893 7800 3927
rect 7748 3884 7800 3893
rect 7840 3884 7892 3936
rect 8852 3952 8904 4004
rect 8944 3884 8996 3936
rect 9312 3927 9364 3936
rect 9312 3893 9321 3927
rect 9321 3893 9355 3927
rect 9355 3893 9364 3927
rect 9312 3884 9364 3893
rect 9496 3884 9548 3936
rect 11244 3952 11296 4004
rect 13912 3952 13964 4004
rect 15936 3952 15988 4004
rect 16580 3952 16632 4004
rect 20168 4020 20220 4072
rect 20996 4020 21048 4072
rect 21180 4063 21232 4072
rect 21180 4029 21189 4063
rect 21189 4029 21223 4063
rect 21223 4029 21232 4063
rect 21180 4020 21232 4029
rect 22100 4063 22152 4072
rect 22100 4029 22109 4063
rect 22109 4029 22143 4063
rect 22143 4029 22152 4063
rect 22284 4063 22336 4072
rect 22100 4020 22152 4029
rect 22284 4029 22293 4063
rect 22293 4029 22327 4063
rect 22327 4029 22336 4063
rect 22284 4020 22336 4029
rect 11980 3884 12032 3936
rect 13452 3884 13504 3936
rect 16488 3884 16540 3936
rect 17408 3927 17460 3936
rect 17408 3893 17417 3927
rect 17417 3893 17451 3927
rect 17451 3893 17460 3927
rect 17408 3884 17460 3893
rect 17776 3927 17828 3936
rect 17776 3893 17785 3927
rect 17785 3893 17819 3927
rect 17819 3893 17828 3927
rect 17776 3884 17828 3893
rect 18052 3927 18104 3936
rect 18052 3893 18061 3927
rect 18061 3893 18095 3927
rect 18095 3893 18104 3927
rect 18052 3884 18104 3893
rect 19432 3927 19484 3936
rect 19432 3893 19441 3927
rect 19441 3893 19475 3927
rect 19475 3893 19484 3927
rect 22376 3952 22428 4004
rect 19432 3884 19484 3893
rect 22100 3884 22152 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1492 3680 1544 3732
rect 1860 3680 1912 3732
rect 2596 3680 2648 3732
rect 2964 3680 3016 3732
rect 3516 3680 3568 3732
rect 3608 3723 3660 3732
rect 3608 3689 3617 3723
rect 3617 3689 3651 3723
rect 3651 3689 3660 3723
rect 3608 3680 3660 3689
rect 5172 3680 5224 3732
rect 6092 3680 6144 3732
rect 7932 3680 7984 3732
rect 8760 3680 8812 3732
rect 9496 3680 9548 3732
rect 10784 3680 10836 3732
rect 11060 3680 11112 3732
rect 2228 3544 2280 3596
rect 3792 3612 3844 3664
rect 6368 3612 6420 3664
rect 7012 3612 7064 3664
rect 8208 3612 8260 3664
rect 11152 3612 11204 3664
rect 11336 3612 11388 3664
rect 12624 3680 12676 3732
rect 13084 3723 13136 3732
rect 13084 3689 13093 3723
rect 13093 3689 13127 3723
rect 13127 3689 13136 3723
rect 13084 3680 13136 3689
rect 13912 3680 13964 3732
rect 14372 3723 14424 3732
rect 14372 3689 14381 3723
rect 14381 3689 14415 3723
rect 14415 3689 14424 3723
rect 14372 3680 14424 3689
rect 14648 3723 14700 3732
rect 14648 3689 14657 3723
rect 14657 3689 14691 3723
rect 14691 3689 14700 3723
rect 14648 3680 14700 3689
rect 15936 3723 15988 3732
rect 15936 3689 15945 3723
rect 15945 3689 15979 3723
rect 15979 3689 15988 3723
rect 15936 3680 15988 3689
rect 16672 3680 16724 3732
rect 16856 3680 16908 3732
rect 17684 3680 17736 3732
rect 18696 3723 18748 3732
rect 18696 3689 18705 3723
rect 18705 3689 18739 3723
rect 18739 3689 18748 3723
rect 18696 3680 18748 3689
rect 20260 3680 20312 3732
rect 2412 3519 2464 3528
rect 2412 3485 2421 3519
rect 2421 3485 2455 3519
rect 2455 3485 2464 3519
rect 2412 3476 2464 3485
rect 1768 3383 1820 3392
rect 1768 3349 1777 3383
rect 1777 3349 1811 3383
rect 1811 3349 1820 3383
rect 1768 3340 1820 3349
rect 3424 3340 3476 3392
rect 4436 3340 4488 3392
rect 4896 3383 4948 3392
rect 4896 3349 4905 3383
rect 4905 3349 4939 3383
rect 4939 3349 4948 3383
rect 4896 3340 4948 3349
rect 7196 3544 7248 3596
rect 7932 3544 7984 3596
rect 9956 3587 10008 3596
rect 9956 3553 9965 3587
rect 9965 3553 9999 3587
rect 9999 3553 10008 3587
rect 9956 3544 10008 3553
rect 11704 3587 11756 3596
rect 6920 3476 6972 3528
rect 8484 3519 8536 3528
rect 8484 3485 8493 3519
rect 8493 3485 8527 3519
rect 8527 3485 8536 3519
rect 8484 3476 8536 3485
rect 8576 3519 8628 3528
rect 8576 3485 8585 3519
rect 8585 3485 8619 3519
rect 8619 3485 8628 3519
rect 8576 3476 8628 3485
rect 7472 3408 7524 3460
rect 7748 3340 7800 3392
rect 11704 3553 11713 3587
rect 11713 3553 11747 3587
rect 11747 3553 11756 3587
rect 13820 3612 13872 3664
rect 14556 3612 14608 3664
rect 19432 3612 19484 3664
rect 20996 3612 21048 3664
rect 11704 3544 11756 3553
rect 13452 3544 13504 3596
rect 13636 3544 13688 3596
rect 14188 3587 14240 3596
rect 14188 3553 14197 3587
rect 14197 3553 14231 3587
rect 14231 3553 14240 3587
rect 14188 3544 14240 3553
rect 11336 3476 11388 3528
rect 13728 3340 13780 3392
rect 14740 3340 14792 3392
rect 16488 3544 16540 3596
rect 18972 3544 19024 3596
rect 19524 3587 19576 3596
rect 19524 3553 19533 3587
rect 19533 3553 19567 3587
rect 19567 3553 19576 3587
rect 19524 3544 19576 3553
rect 16304 3476 16356 3528
rect 18788 3476 18840 3528
rect 16212 3408 16264 3460
rect 19156 3451 19208 3460
rect 19156 3417 19165 3451
rect 19165 3417 19199 3451
rect 19199 3417 19208 3451
rect 19156 3408 19208 3417
rect 19432 3476 19484 3528
rect 22100 3544 22152 3596
rect 22560 3544 22612 3596
rect 21456 3476 21508 3528
rect 18972 3383 19024 3392
rect 18972 3349 18981 3383
rect 18981 3349 19015 3383
rect 19015 3349 19024 3383
rect 18972 3340 19024 3349
rect 21272 3383 21324 3392
rect 21272 3349 21281 3383
rect 21281 3349 21315 3383
rect 21315 3349 21324 3383
rect 21272 3340 21324 3349
rect 21916 3340 21968 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1860 3179 1912 3188
rect 1860 3145 1869 3179
rect 1869 3145 1903 3179
rect 1903 3145 1912 3179
rect 1860 3136 1912 3145
rect 3516 3179 3568 3188
rect 3516 3145 3525 3179
rect 3525 3145 3559 3179
rect 3559 3145 3568 3179
rect 3516 3136 3568 3145
rect 4160 3136 4212 3188
rect 4528 3136 4580 3188
rect 7840 3136 7892 3188
rect 8392 3136 8444 3188
rect 9864 3136 9916 3188
rect 10784 3179 10836 3188
rect 10784 3145 10793 3179
rect 10793 3145 10827 3179
rect 10827 3145 10836 3179
rect 10784 3136 10836 3145
rect 11336 3136 11388 3188
rect 11704 3136 11756 3188
rect 14004 3179 14056 3188
rect 4436 3000 4488 3052
rect 7472 3043 7524 3052
rect 2228 2932 2280 2984
rect 2412 2975 2464 2984
rect 2412 2941 2446 2975
rect 2446 2941 2464 2975
rect 2412 2932 2464 2941
rect 4896 2932 4948 2984
rect 7472 3009 7481 3043
rect 7481 3009 7515 3043
rect 7515 3009 7524 3043
rect 7472 3000 7524 3009
rect 7748 3000 7800 3052
rect 14004 3145 14013 3179
rect 14013 3145 14047 3179
rect 14047 3145 14056 3179
rect 14004 3136 14056 3145
rect 16304 3136 16356 3188
rect 16488 3179 16540 3188
rect 16488 3145 16497 3179
rect 16497 3145 16531 3179
rect 16531 3145 16540 3179
rect 16488 3136 16540 3145
rect 17224 3136 17276 3188
rect 15108 3068 15160 3120
rect 11060 2932 11112 2984
rect 15108 2975 15160 2984
rect 15108 2941 15117 2975
rect 15117 2941 15151 2975
rect 15151 2941 15160 2975
rect 15108 2932 15160 2941
rect 4252 2864 4304 2916
rect 5264 2907 5316 2916
rect 5264 2873 5273 2907
rect 5273 2873 5307 2907
rect 5307 2873 5316 2907
rect 5264 2864 5316 2873
rect 7288 2907 7340 2916
rect 7288 2873 7297 2907
rect 7297 2873 7331 2907
rect 7331 2873 7340 2907
rect 7288 2864 7340 2873
rect 9956 2864 10008 2916
rect 13084 2864 13136 2916
rect 17592 3136 17644 3188
rect 18144 3136 18196 3188
rect 18788 3136 18840 3188
rect 19524 3136 19576 3188
rect 20628 3136 20680 3188
rect 22560 3179 22612 3188
rect 22560 3145 22569 3179
rect 22569 3145 22603 3179
rect 22603 3145 22612 3179
rect 22560 3136 22612 3145
rect 23848 3179 23900 3188
rect 23848 3145 23857 3179
rect 23857 3145 23891 3179
rect 23891 3145 23900 3179
rect 23848 3136 23900 3145
rect 18972 3000 19024 3052
rect 20168 3000 20220 3052
rect 19156 2932 19208 2984
rect 19248 2932 19300 2984
rect 21640 2975 21692 2984
rect 21640 2941 21649 2975
rect 21649 2941 21683 2975
rect 21683 2941 21692 2975
rect 21640 2932 21692 2941
rect 23664 2975 23716 2984
rect 23664 2941 23673 2975
rect 23673 2941 23707 2975
rect 23707 2941 23716 2975
rect 23664 2932 23716 2941
rect 18972 2864 19024 2916
rect 19524 2864 19576 2916
rect 6184 2839 6236 2848
rect 6184 2805 6193 2839
rect 6193 2805 6227 2839
rect 6227 2805 6236 2839
rect 6184 2796 6236 2805
rect 9588 2796 9640 2848
rect 11428 2839 11480 2848
rect 11428 2805 11437 2839
rect 11437 2805 11471 2839
rect 11471 2805 11480 2839
rect 11428 2796 11480 2805
rect 21824 2839 21876 2848
rect 21824 2805 21833 2839
rect 21833 2805 21867 2839
rect 21867 2805 21876 2839
rect 21824 2796 21876 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 3424 2592 3476 2644
rect 2872 2524 2924 2576
rect 2044 2388 2096 2440
rect 3700 2592 3752 2644
rect 3884 2635 3936 2644
rect 3884 2601 3893 2635
rect 3893 2601 3927 2635
rect 3927 2601 3936 2635
rect 3884 2592 3936 2601
rect 5448 2635 5500 2644
rect 5448 2601 5457 2635
rect 5457 2601 5491 2635
rect 5491 2601 5500 2635
rect 5448 2592 5500 2601
rect 6368 2635 6420 2644
rect 6368 2601 6377 2635
rect 6377 2601 6411 2635
rect 6411 2601 6420 2635
rect 6368 2592 6420 2601
rect 7932 2635 7984 2644
rect 7932 2601 7941 2635
rect 7941 2601 7975 2635
rect 7975 2601 7984 2635
rect 7932 2592 7984 2601
rect 8116 2635 8168 2644
rect 8116 2601 8125 2635
rect 8125 2601 8159 2635
rect 8159 2601 8168 2635
rect 8116 2592 8168 2601
rect 9588 2635 9640 2644
rect 9588 2601 9597 2635
rect 9597 2601 9631 2635
rect 9631 2601 9640 2635
rect 9588 2592 9640 2601
rect 10048 2592 10100 2644
rect 10784 2635 10836 2644
rect 10784 2601 10793 2635
rect 10793 2601 10827 2635
rect 10827 2601 10836 2635
rect 10784 2592 10836 2601
rect 4160 2524 4212 2576
rect 9772 2524 9824 2576
rect 8300 2456 8352 2508
rect 8484 2499 8536 2508
rect 8484 2465 8493 2499
rect 8493 2465 8527 2499
rect 8527 2465 8536 2499
rect 8484 2456 8536 2465
rect 9496 2456 9548 2508
rect 11980 2592 12032 2644
rect 13452 2592 13504 2644
rect 14188 2635 14240 2644
rect 14188 2601 14197 2635
rect 14197 2601 14231 2635
rect 14231 2601 14240 2635
rect 14188 2592 14240 2601
rect 14464 2592 14516 2644
rect 14740 2592 14792 2644
rect 15476 2635 15528 2644
rect 15476 2601 15485 2635
rect 15485 2601 15519 2635
rect 15519 2601 15528 2635
rect 15476 2592 15528 2601
rect 16488 2592 16540 2644
rect 17868 2592 17920 2644
rect 15292 2524 15344 2576
rect 19248 2592 19300 2644
rect 20628 2592 20680 2644
rect 21456 2635 21508 2644
rect 21456 2601 21465 2635
rect 21465 2601 21499 2635
rect 21499 2601 21508 2635
rect 21456 2592 21508 2601
rect 6920 2388 6972 2440
rect 8668 2388 8720 2440
rect 9588 2388 9640 2440
rect 10784 2388 10836 2440
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 13268 2431 13320 2440
rect 11980 2388 12032 2397
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 14740 2456 14792 2508
rect 17132 2499 17184 2508
rect 17132 2465 17141 2499
rect 17141 2465 17175 2499
rect 17175 2465 17184 2499
rect 17132 2456 17184 2465
rect 18696 2499 18748 2508
rect 18696 2465 18705 2499
rect 18705 2465 18739 2499
rect 18739 2465 18748 2499
rect 18696 2456 18748 2465
rect 19340 2456 19392 2508
rect 22192 2499 22244 2508
rect 22192 2465 22201 2499
rect 22201 2465 22235 2499
rect 22235 2465 22244 2499
rect 22192 2456 22244 2465
rect 24032 2499 24084 2508
rect 24032 2465 24041 2499
rect 24041 2465 24075 2499
rect 24075 2465 24084 2499
rect 24032 2456 24084 2465
rect 14924 2388 14976 2440
rect 15936 2388 15988 2440
rect 18880 2431 18932 2440
rect 18880 2397 18889 2431
rect 18889 2397 18923 2431
rect 18923 2397 18932 2431
rect 18880 2388 18932 2397
rect 3332 2320 3384 2372
rect 10876 2320 10928 2372
rect 11612 2363 11664 2372
rect 11612 2329 11621 2363
rect 11621 2329 11655 2363
rect 11655 2329 11664 2363
rect 11612 2320 11664 2329
rect 13728 2320 13780 2372
rect 15476 2320 15528 2372
rect 7288 2295 7340 2304
rect 7288 2261 7297 2295
rect 7297 2261 7331 2295
rect 7331 2261 7340 2295
rect 7288 2252 7340 2261
rect 15292 2295 15344 2304
rect 15292 2261 15301 2295
rect 15301 2261 15335 2295
rect 15335 2261 15344 2295
rect 15292 2252 15344 2261
rect 17316 2295 17368 2304
rect 17316 2261 17325 2295
rect 17325 2261 17359 2295
rect 17359 2261 17368 2295
rect 17316 2252 17368 2261
rect 20076 2295 20128 2304
rect 20076 2261 20085 2295
rect 20085 2261 20119 2295
rect 20119 2261 20128 2295
rect 20076 2252 20128 2261
rect 24124 2252 24176 2304
rect 24216 2295 24268 2304
rect 24216 2261 24225 2295
rect 24225 2261 24259 2295
rect 24259 2261 24268 2295
rect 24216 2252 24268 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 14648 1980 14700 2032
rect 15752 1980 15804 2032
rect 14372 1844 14424 1896
rect 18696 1844 18748 1896
<< metal2 >>
rect 294 27520 350 28000
rect 846 27520 902 28000
rect 1398 27520 1454 28000
rect 1950 27520 2006 28000
rect 2502 27520 2558 28000
rect 2778 27704 2834 27713
rect 2778 27639 2834 27648
rect 308 27418 336 27520
rect 308 27390 612 27418
rect 584 19961 612 27390
rect 860 20233 888 27520
rect 1412 24698 1440 27520
rect 1964 25514 1992 27520
rect 1964 25486 2268 25514
rect 1952 25356 2004 25362
rect 1952 25298 2004 25304
rect 1964 24721 1992 25298
rect 2136 25152 2188 25158
rect 2136 25094 2188 25100
rect 2042 24848 2098 24857
rect 2042 24783 2044 24792
rect 2096 24783 2098 24792
rect 2044 24754 2096 24760
rect 1320 24670 1440 24698
rect 1950 24712 2006 24721
rect 846 20224 902 20233
rect 846 20159 902 20168
rect 570 19952 626 19961
rect 570 19887 626 19896
rect 1320 19378 1348 24670
rect 1950 24647 2006 24656
rect 1400 24608 1452 24614
rect 1400 24550 1452 24556
rect 1412 21321 1440 24550
rect 1964 24410 1992 24647
rect 1952 24404 2004 24410
rect 1952 24346 2004 24352
rect 2044 24268 2096 24274
rect 2044 24210 2096 24216
rect 1676 24064 1728 24070
rect 1676 24006 1728 24012
rect 1584 22432 1636 22438
rect 1584 22374 1636 22380
rect 1596 21865 1624 22374
rect 1688 22098 1716 24006
rect 2056 23866 2084 24210
rect 2044 23860 2096 23866
rect 2044 23802 2096 23808
rect 2148 23304 2176 25094
rect 2056 23276 2176 23304
rect 2056 23118 2084 23276
rect 2240 23254 2268 25486
rect 2412 25356 2464 25362
rect 2412 25298 2464 25304
rect 2320 25152 2372 25158
rect 2320 25094 2372 25100
rect 2332 23866 2360 25094
rect 2424 24954 2452 25298
rect 2412 24948 2464 24954
rect 2412 24890 2464 24896
rect 2516 24834 2544 27520
rect 2424 24806 2544 24834
rect 2320 23860 2372 23866
rect 2320 23802 2372 23808
rect 2332 23322 2360 23802
rect 2320 23316 2372 23322
rect 2320 23258 2372 23264
rect 2228 23248 2280 23254
rect 2134 23216 2190 23225
rect 2228 23190 2280 23196
rect 2134 23151 2190 23160
rect 2044 23112 2096 23118
rect 1964 23072 2044 23100
rect 1860 22976 1912 22982
rect 1860 22918 1912 22924
rect 1676 22092 1728 22098
rect 1676 22034 1728 22040
rect 1582 21856 1638 21865
rect 1582 21791 1638 21800
rect 1398 21312 1454 21321
rect 1398 21247 1454 21256
rect 1398 21040 1454 21049
rect 1398 20975 1400 20984
rect 1452 20975 1454 20984
rect 1400 20946 1452 20952
rect 1688 20874 1716 22034
rect 1872 21944 1900 22918
rect 1964 22234 1992 23072
rect 2044 23054 2096 23060
rect 2148 22778 2176 23151
rect 2136 22772 2188 22778
rect 2136 22714 2188 22720
rect 2228 22636 2280 22642
rect 2228 22578 2280 22584
rect 1952 22228 2004 22234
rect 1952 22170 2004 22176
rect 2240 22166 2268 22578
rect 2318 22400 2374 22409
rect 2318 22335 2374 22344
rect 2228 22160 2280 22166
rect 2228 22102 2280 22108
rect 1872 21916 1992 21944
rect 1768 21888 1820 21894
rect 1820 21836 1900 21842
rect 1768 21830 1900 21836
rect 1780 21814 1900 21830
rect 1676 20868 1728 20874
rect 1676 20810 1728 20816
rect 1584 20800 1636 20806
rect 1584 20742 1636 20748
rect 1400 20256 1452 20262
rect 1400 20198 1452 20204
rect 1308 19372 1360 19378
rect 1308 19314 1360 19320
rect 1412 19009 1440 20198
rect 1596 19802 1624 20742
rect 1596 19774 1716 19802
rect 1584 19712 1636 19718
rect 1584 19654 1636 19660
rect 1492 19168 1544 19174
rect 1492 19110 1544 19116
rect 1398 19000 1454 19009
rect 1398 18935 1454 18944
rect 1400 18624 1452 18630
rect 1400 18566 1452 18572
rect 1412 16697 1440 18566
rect 1504 17241 1532 19110
rect 1596 18465 1624 19654
rect 1688 18834 1716 19774
rect 1676 18828 1728 18834
rect 1676 18770 1728 18776
rect 1582 18456 1638 18465
rect 1582 18391 1638 18400
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1490 17232 1546 17241
rect 1490 17167 1546 17176
rect 1492 16992 1544 16998
rect 1492 16934 1544 16940
rect 1398 16688 1454 16697
rect 1398 16623 1454 16632
rect 1400 14952 1452 14958
rect 1504 14929 1532 16934
rect 1596 16017 1624 18022
rect 1688 17882 1716 18770
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1582 16008 1638 16017
rect 1582 15943 1638 15952
rect 1584 15904 1636 15910
rect 1584 15846 1636 15852
rect 1400 14894 1452 14900
rect 1490 14920 1546 14929
rect 1412 14793 1440 14894
rect 1490 14855 1546 14864
rect 1398 14784 1454 14793
rect 1398 14719 1454 14728
rect 1398 13424 1454 13433
rect 1398 13359 1400 13368
rect 1452 13359 1454 13368
rect 1400 13330 1452 13336
rect 1596 13161 1624 15846
rect 1688 13705 1716 16730
rect 1768 16448 1820 16454
rect 1768 16390 1820 16396
rect 1780 16046 1808 16390
rect 1872 16250 1900 21814
rect 1964 21162 1992 21916
rect 2240 21554 2268 22102
rect 2332 21978 2360 22335
rect 2424 22098 2452 24806
rect 2596 24608 2648 24614
rect 2596 24550 2648 24556
rect 2504 24132 2556 24138
rect 2504 24074 2556 24080
rect 2516 23662 2544 24074
rect 2608 23662 2636 24550
rect 2792 24410 2820 27639
rect 3146 27520 3202 28000
rect 3698 27520 3754 28000
rect 4250 27520 4306 28000
rect 4802 27520 4858 28000
rect 5354 27520 5410 28000
rect 5998 27520 6054 28000
rect 6550 27520 6606 28000
rect 7102 27520 7158 28000
rect 7654 27520 7710 28000
rect 8206 27520 8262 28000
rect 8850 27520 8906 28000
rect 9402 27520 9458 28000
rect 9954 27520 10010 28000
rect 10506 27520 10562 28000
rect 11058 27520 11114 28000
rect 11702 27520 11758 28000
rect 12254 27520 12310 28000
rect 12806 27520 12862 28000
rect 13358 27520 13414 28000
rect 13910 27520 13966 28000
rect 14554 27520 14610 28000
rect 15106 27520 15162 28000
rect 15658 27520 15714 28000
rect 16210 27520 16266 28000
rect 16762 27520 16818 28000
rect 17406 27520 17462 28000
rect 17958 27520 18014 28000
rect 18510 27520 18566 28000
rect 19062 27520 19118 28000
rect 19614 27520 19670 28000
rect 20258 27520 20314 28000
rect 20810 27520 20866 28000
rect 21362 27520 21418 28000
rect 21914 27520 21970 28000
rect 22466 27520 22522 28000
rect 23110 27520 23166 28000
rect 23662 27520 23718 28000
rect 24214 27520 24270 28000
rect 24766 27520 24822 28000
rect 25318 27520 25374 28000
rect 25962 27520 26018 28000
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 3054 25392 3110 25401
rect 3054 25327 3110 25336
rect 2964 25220 3016 25226
rect 2964 25162 3016 25168
rect 2872 25152 2924 25158
rect 2872 25094 2924 25100
rect 2780 24404 2832 24410
rect 2780 24346 2832 24352
rect 2688 24064 2740 24070
rect 2688 24006 2740 24012
rect 2700 23730 2728 24006
rect 2792 23866 2820 24346
rect 2780 23860 2832 23866
rect 2780 23802 2832 23808
rect 2688 23724 2740 23730
rect 2688 23666 2740 23672
rect 2504 23656 2556 23662
rect 2504 23598 2556 23604
rect 2596 23656 2648 23662
rect 2596 23598 2648 23604
rect 2608 23474 2636 23598
rect 2608 23446 2820 23474
rect 2792 23322 2820 23446
rect 2780 23316 2832 23322
rect 2780 23258 2832 23264
rect 2596 23248 2648 23254
rect 2596 23190 2648 23196
rect 2412 22092 2464 22098
rect 2412 22034 2464 22040
rect 2332 21950 2544 21978
rect 2228 21548 2280 21554
rect 2228 21490 2280 21496
rect 2320 21412 2372 21418
rect 2320 21354 2372 21360
rect 1964 21134 2084 21162
rect 2332 21146 2360 21354
rect 1950 21040 2006 21049
rect 1950 20975 2006 20984
rect 1964 20058 1992 20975
rect 1952 20052 2004 20058
rect 1952 19994 2004 20000
rect 2056 19258 2084 21134
rect 2320 21140 2372 21146
rect 2320 21082 2372 21088
rect 2410 20496 2466 20505
rect 2410 20431 2466 20440
rect 2424 20398 2452 20431
rect 2412 20392 2464 20398
rect 2412 20334 2464 20340
rect 2424 20058 2452 20334
rect 2412 20052 2464 20058
rect 2412 19994 2464 20000
rect 2320 19916 2372 19922
rect 2320 19858 2372 19864
rect 2332 19514 2360 19858
rect 2320 19508 2372 19514
rect 2320 19450 2372 19456
rect 2320 19372 2372 19378
rect 2320 19314 2372 19320
rect 2056 19230 2176 19258
rect 2044 19168 2096 19174
rect 2044 19110 2096 19116
rect 2056 18873 2084 19110
rect 2042 18864 2098 18873
rect 2042 18799 2098 18808
rect 2044 18624 2096 18630
rect 2044 18566 2096 18572
rect 2056 18222 2084 18566
rect 2044 18216 2096 18222
rect 2044 18158 2096 18164
rect 2056 17921 2084 18158
rect 2042 17912 2098 17921
rect 2042 17847 2098 17856
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1964 17241 1992 17478
rect 1950 17232 2006 17241
rect 1950 17167 2006 17176
rect 1964 17134 1992 17167
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 1860 16244 1912 16250
rect 1860 16186 1912 16192
rect 1768 16040 1820 16046
rect 1768 15982 1820 15988
rect 1674 13696 1730 13705
rect 1674 13631 1730 13640
rect 1780 13258 1808 15982
rect 2056 15706 2084 16526
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 2042 15600 2098 15609
rect 2042 15535 2044 15544
rect 2096 15535 2098 15544
rect 2044 15506 2096 15512
rect 1952 14272 2004 14278
rect 1952 14214 2004 14220
rect 1964 13818 1992 14214
rect 2044 13864 2096 13870
rect 1964 13812 2044 13818
rect 1964 13806 2096 13812
rect 1964 13790 2084 13806
rect 1768 13252 1820 13258
rect 1768 13194 1820 13200
rect 1582 13152 1638 13161
rect 1582 13087 1638 13096
rect 1860 12640 1912 12646
rect 1582 12608 1638 12617
rect 1860 12582 1912 12588
rect 1582 12543 1638 12552
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1412 11830 1440 12174
rect 1596 11898 1624 12543
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 1400 11824 1452 11830
rect 1400 11766 1452 11772
rect 1400 11688 1452 11694
rect 1400 11630 1452 11636
rect 1412 11354 1440 11630
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1412 10033 1440 10542
rect 1688 10146 1716 12378
rect 1872 11830 1900 12582
rect 1964 12442 1992 13790
rect 2044 13728 2096 13734
rect 2044 13670 2096 13676
rect 2056 13258 2084 13670
rect 2044 13252 2096 13258
rect 2044 13194 2096 13200
rect 2044 12980 2096 12986
rect 2044 12922 2096 12928
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 1952 12300 2004 12306
rect 1952 12242 2004 12248
rect 1860 11824 1912 11830
rect 1860 11766 1912 11772
rect 1964 11354 1992 12242
rect 2056 11354 2084 12922
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 1858 10568 1914 10577
rect 1858 10503 1860 10512
rect 1912 10503 1914 10512
rect 1860 10474 1912 10480
rect 1596 10118 1716 10146
rect 1768 10124 1820 10130
rect 1398 10024 1454 10033
rect 1398 9959 1400 9968
rect 1452 9959 1454 9968
rect 1400 9930 1452 9936
rect 1492 9512 1544 9518
rect 1492 9454 1544 9460
rect 1504 9042 1532 9454
rect 1492 9036 1544 9042
rect 1492 8978 1544 8984
rect 570 7848 626 7857
rect 1596 7834 1624 10118
rect 1768 10066 1820 10072
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1688 9654 1716 9998
rect 1676 9648 1728 9654
rect 1674 9616 1676 9625
rect 1728 9616 1730 9625
rect 1674 9551 1730 9560
rect 570 7783 626 7792
rect 1504 7806 1624 7834
rect 584 7478 612 7783
rect 572 7472 624 7478
rect 572 7414 624 7420
rect 1400 7200 1452 7206
rect 1400 7142 1452 7148
rect 1412 5166 1440 7142
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 846 4312 902 4321
rect 846 4247 902 4256
rect 294 3496 350 3505
rect 294 3431 350 3440
rect 308 480 336 3431
rect 860 480 888 4247
rect 1412 4185 1440 5102
rect 1504 5001 1532 7806
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1596 5817 1624 7686
rect 1688 7410 1716 9551
rect 1780 8498 1808 10066
rect 1872 9722 1900 10474
rect 1964 10062 1992 11290
rect 2148 11218 2176 19230
rect 2228 17604 2280 17610
rect 2228 17546 2280 17552
rect 2240 17338 2268 17546
rect 2332 17490 2360 19314
rect 2332 17462 2452 17490
rect 2228 17332 2280 17338
rect 2228 17274 2280 17280
rect 2240 16810 2268 17274
rect 2240 16782 2360 16810
rect 2228 16652 2280 16658
rect 2228 16594 2280 16600
rect 2240 15706 2268 16594
rect 2332 16114 2360 16782
rect 2424 16522 2452 17462
rect 2412 16516 2464 16522
rect 2412 16458 2464 16464
rect 2320 16108 2372 16114
rect 2320 16050 2372 16056
rect 2516 15858 2544 21950
rect 2608 18714 2636 23190
rect 2688 23112 2740 23118
rect 2884 23089 2912 25094
rect 2688 23054 2740 23060
rect 2870 23080 2926 23089
rect 2700 21962 2728 23054
rect 2870 23015 2926 23024
rect 2872 22976 2924 22982
rect 2872 22918 2924 22924
rect 2884 22438 2912 22918
rect 2976 22545 3004 25162
rect 3068 25158 3096 25327
rect 3056 25152 3108 25158
rect 3056 25094 3108 25100
rect 3068 24750 3096 25094
rect 3160 24834 3188 27520
rect 3606 26616 3662 26625
rect 3606 26551 3662 26560
rect 3160 24806 3556 24834
rect 3056 24744 3108 24750
rect 3056 24686 3108 24692
rect 3332 24744 3384 24750
rect 3332 24686 3384 24692
rect 2962 22536 3018 22545
rect 2962 22471 3018 22480
rect 2872 22432 2924 22438
rect 2924 22392 3004 22420
rect 2872 22374 2924 22380
rect 2884 22309 2912 22374
rect 2688 21956 2740 21962
rect 2688 21898 2740 21904
rect 2700 21418 2728 21898
rect 2688 21412 2740 21418
rect 2688 21354 2740 21360
rect 2872 21072 2924 21078
rect 2872 21014 2924 21020
rect 2780 21004 2832 21010
rect 2780 20946 2832 20952
rect 2688 20392 2740 20398
rect 2792 20346 2820 20946
rect 2884 20369 2912 21014
rect 2976 20942 3004 22392
rect 2964 20936 3016 20942
rect 2964 20878 3016 20884
rect 2976 20602 3004 20878
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 2740 20340 2820 20346
rect 2688 20334 2820 20340
rect 2700 20318 2820 20334
rect 2870 20360 2926 20369
rect 2700 19689 2728 20318
rect 2870 20295 2872 20304
rect 2924 20295 2926 20304
rect 2872 20266 2924 20272
rect 2964 20256 3016 20262
rect 2964 20198 3016 20204
rect 2686 19680 2742 19689
rect 2686 19615 2742 19624
rect 2686 19544 2742 19553
rect 2686 19479 2742 19488
rect 2700 19174 2728 19479
rect 2976 19310 3004 20198
rect 3068 19904 3096 24686
rect 3344 24206 3372 24686
rect 3424 24608 3476 24614
rect 3424 24550 3476 24556
rect 3332 24200 3384 24206
rect 3332 24142 3384 24148
rect 3344 24070 3372 24142
rect 3332 24064 3384 24070
rect 3332 24006 3384 24012
rect 3148 23860 3200 23866
rect 3148 23802 3200 23808
rect 3240 23860 3292 23866
rect 3240 23802 3292 23808
rect 3160 19972 3188 23802
rect 3252 20262 3280 23802
rect 3344 23526 3372 24006
rect 3332 23520 3384 23526
rect 3332 23462 3384 23468
rect 3344 22982 3372 23462
rect 3332 22976 3384 22982
rect 3332 22918 3384 22924
rect 3436 21457 3464 24550
rect 3422 21448 3478 21457
rect 3422 21383 3478 21392
rect 3240 20256 3292 20262
rect 3240 20198 3292 20204
rect 3160 19944 3280 19972
rect 3068 19876 3188 19904
rect 3054 19816 3110 19825
rect 3054 19751 3056 19760
rect 3108 19751 3110 19760
rect 3056 19722 3108 19728
rect 2964 19304 3016 19310
rect 2964 19246 3016 19252
rect 2688 19168 2740 19174
rect 2688 19110 2740 19116
rect 3160 19009 3188 19876
rect 3252 19802 3280 19944
rect 3252 19774 3372 19802
rect 3240 19168 3292 19174
rect 3238 19136 3240 19145
rect 3292 19136 3294 19145
rect 3238 19071 3294 19080
rect 3146 19000 3202 19009
rect 3146 18935 3202 18944
rect 2608 18686 2820 18714
rect 2688 18624 2740 18630
rect 2688 18566 2740 18572
rect 2596 18352 2648 18358
rect 2596 18294 2648 18300
rect 2608 17678 2636 18294
rect 2700 17785 2728 18566
rect 2686 17776 2742 17785
rect 2686 17711 2742 17720
rect 2596 17672 2648 17678
rect 2596 17614 2648 17620
rect 2608 16794 2636 17614
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2596 16788 2648 16794
rect 2596 16730 2648 16736
rect 2596 16516 2648 16522
rect 2596 16458 2648 16464
rect 2332 15830 2544 15858
rect 2228 15700 2280 15706
rect 2228 15642 2280 15648
rect 2240 14618 2268 15642
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2228 14272 2280 14278
rect 2228 14214 2280 14220
rect 2240 13938 2268 14214
rect 2228 13932 2280 13938
rect 2228 13874 2280 13880
rect 2240 11529 2268 13874
rect 2332 12986 2360 15830
rect 2412 15700 2464 15706
rect 2412 15642 2464 15648
rect 2424 14482 2452 15642
rect 2608 15586 2636 16458
rect 2516 15558 2636 15586
rect 2700 15570 2728 17478
rect 2792 17218 2820 18686
rect 3160 18222 3188 18935
rect 3240 18624 3292 18630
rect 3240 18566 3292 18572
rect 3252 18290 3280 18566
rect 3344 18329 3372 19774
rect 3330 18320 3386 18329
rect 3240 18284 3292 18290
rect 3330 18255 3386 18264
rect 3240 18226 3292 18232
rect 2964 18216 3016 18222
rect 2964 18158 3016 18164
rect 3148 18216 3200 18222
rect 3148 18158 3200 18164
rect 2976 18086 3004 18158
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 2792 17190 3004 17218
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 2688 15564 2740 15570
rect 2516 15042 2544 15558
rect 2688 15506 2740 15512
rect 2596 15496 2648 15502
rect 2792 15473 2820 16390
rect 2884 15978 2912 17070
rect 2872 15972 2924 15978
rect 2872 15914 2924 15920
rect 2596 15438 2648 15444
rect 2778 15464 2834 15473
rect 2608 15162 2636 15438
rect 2778 15399 2834 15408
rect 2596 15156 2648 15162
rect 2976 15144 3004 17190
rect 3068 16998 3096 17614
rect 3252 17066 3280 18226
rect 3436 18086 3464 21383
rect 3424 18080 3476 18086
rect 3424 18022 3476 18028
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3240 17060 3292 17066
rect 3240 17002 3292 17008
rect 3056 16992 3108 16998
rect 3056 16934 3108 16940
rect 3252 16658 3280 17002
rect 3436 16794 3464 17818
rect 3424 16788 3476 16794
rect 3424 16730 3476 16736
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 3240 15428 3292 15434
rect 3240 15370 3292 15376
rect 2596 15098 2648 15104
rect 2700 15116 3004 15144
rect 2516 15014 2636 15042
rect 2412 14476 2464 14482
rect 2412 14418 2464 14424
rect 2424 13705 2452 14418
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 2410 13696 2466 13705
rect 2410 13631 2466 13640
rect 2412 13184 2464 13190
rect 2412 13126 2464 13132
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2226 11520 2282 11529
rect 2226 11455 2282 11464
rect 2136 11212 2188 11218
rect 2136 11154 2188 11160
rect 2148 11121 2176 11154
rect 2134 11112 2190 11121
rect 2134 11047 2190 11056
rect 2332 10674 2360 12378
rect 2424 11665 2452 13126
rect 2410 11656 2466 11665
rect 2410 11591 2466 11600
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2056 10266 2084 10610
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 1952 10056 2004 10062
rect 1952 9998 2004 10004
rect 1860 9716 1912 9722
rect 1860 9658 1912 9664
rect 1964 9586 1992 9998
rect 1952 9580 2004 9586
rect 1952 9522 2004 9528
rect 2044 9444 2096 9450
rect 2044 9386 2096 9392
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 2056 8090 2084 9386
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2240 8294 2268 9318
rect 2516 8634 2544 14350
rect 2608 14113 2636 15014
rect 2594 14104 2650 14113
rect 2594 14039 2650 14048
rect 2700 13394 2728 15116
rect 2870 15056 2926 15065
rect 2870 14991 2872 15000
rect 2924 14991 2926 15000
rect 2872 14962 2924 14968
rect 2870 14920 2926 14929
rect 2780 14884 2832 14890
rect 2870 14855 2926 14864
rect 2780 14826 2832 14832
rect 2688 13388 2740 13394
rect 2608 13348 2688 13376
rect 2608 12442 2636 13348
rect 2688 13330 2740 13336
rect 2792 13138 2820 14826
rect 2884 14550 2912 14855
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 2872 14544 2924 14550
rect 2872 14486 2924 14492
rect 2884 13410 2912 14486
rect 2964 14272 3016 14278
rect 2964 14214 3016 14220
rect 2976 13841 3004 14214
rect 3054 14104 3110 14113
rect 3054 14039 3110 14048
rect 3068 13870 3096 14039
rect 3056 13864 3108 13870
rect 2962 13832 3018 13841
rect 3056 13806 3108 13812
rect 2962 13767 3018 13776
rect 3068 13530 3096 13806
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 2884 13382 3096 13410
rect 2792 13110 2912 13138
rect 2688 12708 2740 12714
rect 2688 12650 2740 12656
rect 2700 12442 2728 12650
rect 2596 12436 2648 12442
rect 2596 12378 2648 12384
rect 2688 12436 2740 12442
rect 2688 12378 2740 12384
rect 2700 12322 2728 12378
rect 2608 12294 2728 12322
rect 2608 10266 2636 12294
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2792 11558 2820 11630
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2778 11248 2834 11257
rect 2778 11183 2780 11192
rect 2832 11183 2834 11192
rect 2780 11154 2832 11160
rect 2792 11098 2820 11154
rect 2700 11070 2820 11098
rect 2700 10810 2728 11070
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2792 9518 2820 9862
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2596 8356 2648 8362
rect 2596 8298 2648 8304
rect 2228 8288 2280 8294
rect 2228 8230 2280 8236
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 2056 7970 2084 8026
rect 2056 7942 2176 7970
rect 2240 7954 2268 8230
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2056 7410 2084 7822
rect 2148 7546 2176 7942
rect 2228 7948 2280 7954
rect 2228 7890 2280 7896
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 1688 6934 1716 7346
rect 1768 7268 1820 7274
rect 1768 7210 1820 7216
rect 1780 7002 1808 7210
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 1676 6928 1728 6934
rect 1676 6870 1728 6876
rect 2240 6662 2268 7890
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2516 6730 2544 7346
rect 2504 6724 2556 6730
rect 2504 6666 2556 6672
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1582 5808 1638 5817
rect 1688 5778 1716 6054
rect 1768 5840 1820 5846
rect 1768 5782 1820 5788
rect 1582 5743 1638 5752
rect 1676 5772 1728 5778
rect 1596 5234 1624 5743
rect 1676 5714 1728 5720
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1490 4992 1546 5001
rect 1490 4927 1546 4936
rect 1398 4176 1454 4185
rect 1398 4111 1454 4120
rect 1504 3738 1532 4927
rect 1780 4826 1808 5782
rect 2240 5681 2268 6598
rect 2412 5772 2464 5778
rect 2516 5760 2544 6666
rect 2464 5732 2544 5760
rect 2412 5714 2464 5720
rect 2226 5672 2282 5681
rect 2226 5607 2282 5616
rect 2424 5370 2452 5714
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 2410 4584 2466 4593
rect 2410 4519 2412 4528
rect 2464 4519 2466 4528
rect 2412 4490 2464 4496
rect 2502 4040 2558 4049
rect 2412 4004 2464 4010
rect 2502 3975 2558 3984
rect 2412 3946 2464 3952
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 1492 3732 1544 3738
rect 1492 3674 1544 3680
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 1490 3632 1546 3641
rect 1490 3567 1546 3576
rect 1504 1034 1532 3567
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 1780 1057 1808 3334
rect 1872 3194 1900 3674
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 1860 3188 1912 3194
rect 1860 3130 1912 3136
rect 2240 2990 2268 3538
rect 2228 2984 2280 2990
rect 2228 2926 2280 2932
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 2056 1873 2084 2382
rect 2042 1864 2098 1873
rect 2042 1799 2098 1808
rect 1950 1592 2006 1601
rect 1950 1527 2006 1536
rect 1412 1006 1532 1034
rect 1766 1048 1822 1057
rect 1412 480 1440 1006
rect 1766 983 1822 992
rect 1964 480 1992 1527
rect 2332 1193 2360 3878
rect 2424 3534 2452 3946
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 2424 3369 2452 3470
rect 2410 3360 2466 3369
rect 2410 3295 2466 3304
rect 2424 2990 2452 3295
rect 2412 2984 2464 2990
rect 2412 2926 2464 2932
rect 2318 1184 2374 1193
rect 2318 1119 2374 1128
rect 2516 480 2544 3975
rect 2608 3738 2636 8298
rect 2792 8294 2820 9454
rect 2884 9110 2912 13110
rect 2964 11620 3016 11626
rect 2964 11562 3016 11568
rect 2976 11150 3004 11562
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 3068 10810 3096 13382
rect 3160 12102 3188 14758
rect 3252 14482 3280 15370
rect 3528 15144 3556 24806
rect 3620 24750 3648 26551
rect 3608 24744 3660 24750
rect 3608 24686 3660 24692
rect 3608 24268 3660 24274
rect 3608 24210 3660 24216
rect 3620 24177 3648 24210
rect 3606 24168 3662 24177
rect 3606 24103 3662 24112
rect 3620 23866 3648 24103
rect 3608 23860 3660 23866
rect 3608 23802 3660 23808
rect 3608 23248 3660 23254
rect 3608 23190 3660 23196
rect 3620 22778 3648 23190
rect 3608 22772 3660 22778
rect 3608 22714 3660 22720
rect 3608 21344 3660 21350
rect 3608 21286 3660 21292
rect 3620 20942 3648 21286
rect 3608 20936 3660 20942
rect 3608 20878 3660 20884
rect 3620 20330 3648 20878
rect 3608 20324 3660 20330
rect 3608 20266 3660 20272
rect 3620 20058 3648 20266
rect 3608 20052 3660 20058
rect 3608 19994 3660 20000
rect 3608 17536 3660 17542
rect 3608 17478 3660 17484
rect 3436 15116 3556 15144
rect 3330 15056 3386 15065
rect 3330 14991 3386 15000
rect 3240 14476 3292 14482
rect 3240 14418 3292 14424
rect 3344 14074 3372 14991
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 3436 13569 3464 15116
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3528 14822 3556 14962
rect 3516 14816 3568 14822
rect 3620 14793 3648 17478
rect 3516 14758 3568 14764
rect 3606 14784 3662 14793
rect 3528 14414 3556 14758
rect 3606 14719 3662 14728
rect 3516 14408 3568 14414
rect 3516 14350 3568 14356
rect 3712 14090 3740 27520
rect 4066 25936 4122 25945
rect 4066 25871 4122 25880
rect 4080 24886 4108 25871
rect 4068 24880 4120 24886
rect 4068 24822 4120 24828
rect 3790 24576 3846 24585
rect 3790 24511 3846 24520
rect 3804 22545 3832 24511
rect 4068 24064 4120 24070
rect 4068 24006 4120 24012
rect 3974 23624 4030 23633
rect 3974 23559 3976 23568
rect 4028 23559 4030 23568
rect 3976 23530 4028 23536
rect 3976 23316 4028 23322
rect 3976 23258 4028 23264
rect 3790 22536 3846 22545
rect 3790 22471 3846 22480
rect 3792 22432 3844 22438
rect 3792 22374 3844 22380
rect 3804 22001 3832 22374
rect 3988 22098 4016 23258
rect 4080 23100 4108 24006
rect 4160 23656 4212 23662
rect 4160 23598 4212 23604
rect 4172 23254 4200 23598
rect 4160 23248 4212 23254
rect 4160 23190 4212 23196
rect 4160 23112 4212 23118
rect 4080 23072 4160 23100
rect 4160 23054 4212 23060
rect 4066 22944 4122 22953
rect 4066 22879 4122 22888
rect 3976 22092 4028 22098
rect 3976 22034 4028 22040
rect 3790 21992 3846 22001
rect 3790 21927 3846 21936
rect 3804 21078 3832 21927
rect 3792 21072 3844 21078
rect 3792 21014 3844 21020
rect 3804 20874 3832 21014
rect 3792 20868 3844 20874
rect 3792 20810 3844 20816
rect 4080 20777 4108 22879
rect 4264 22794 4292 27520
rect 4710 27160 4766 27169
rect 4710 27095 4766 27104
rect 4528 24200 4580 24206
rect 4528 24142 4580 24148
rect 4342 23760 4398 23769
rect 4342 23695 4398 23704
rect 4356 22953 4384 23695
rect 4540 23633 4568 24142
rect 4526 23624 4582 23633
rect 4526 23559 4582 23568
rect 4436 23112 4488 23118
rect 4436 23054 4488 23060
rect 4342 22944 4398 22953
rect 4342 22879 4398 22888
rect 4264 22766 4384 22794
rect 4356 22114 4384 22766
rect 4448 22166 4476 23054
rect 4347 22086 4384 22114
rect 4436 22160 4488 22166
rect 4436 22102 4488 22108
rect 4528 22092 4580 22098
rect 4347 22012 4375 22086
rect 4528 22034 4580 22040
rect 4347 21984 4384 22012
rect 4160 20800 4212 20806
rect 4066 20768 4122 20777
rect 4160 20742 4212 20748
rect 4066 20703 4122 20712
rect 4068 20392 4120 20398
rect 4068 20334 4120 20340
rect 3792 20256 3844 20262
rect 3792 20198 3844 20204
rect 3804 19718 3832 20198
rect 4080 19922 4108 20334
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 3792 19712 3844 19718
rect 3792 19654 3844 19660
rect 3804 18766 3832 19654
rect 4172 19310 4200 20742
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 3884 19168 3936 19174
rect 3884 19110 3936 19116
rect 3792 18760 3844 18766
rect 3792 18702 3844 18708
rect 3804 18426 3832 18702
rect 3792 18420 3844 18426
rect 3792 18362 3844 18368
rect 3792 15564 3844 15570
rect 3792 15506 3844 15512
rect 3804 14618 3832 15506
rect 3792 14612 3844 14618
rect 3792 14554 3844 14560
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 3528 14062 3740 14090
rect 3528 13802 3556 14062
rect 3700 13932 3752 13938
rect 3700 13874 3752 13880
rect 3608 13864 3660 13870
rect 3606 13832 3608 13841
rect 3660 13832 3662 13841
rect 3516 13796 3568 13802
rect 3606 13767 3662 13776
rect 3516 13738 3568 13744
rect 3528 13682 3556 13738
rect 3528 13654 3648 13682
rect 3422 13560 3478 13569
rect 3422 13495 3478 13504
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3240 13252 3292 13258
rect 3240 13194 3292 13200
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 3146 11792 3202 11801
rect 3146 11727 3202 11736
rect 3160 11286 3188 11727
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 3054 10160 3110 10169
rect 3054 10095 3110 10104
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 2976 9178 3004 9522
rect 3068 9217 3096 10095
rect 3148 9512 3200 9518
rect 3252 9489 3280 13194
rect 3424 12640 3476 12646
rect 3424 12582 3476 12588
rect 3436 11694 3464 12582
rect 3528 12238 3556 13466
rect 3620 13376 3648 13654
rect 3712 13530 3740 13874
rect 3700 13524 3752 13530
rect 3700 13466 3752 13472
rect 3700 13388 3752 13394
rect 3620 13348 3700 13376
rect 3700 13330 3752 13336
rect 3712 12986 3740 13330
rect 3700 12980 3752 12986
rect 3700 12922 3752 12928
rect 3516 12232 3568 12238
rect 3514 12200 3516 12209
rect 3568 12200 3570 12209
rect 3514 12135 3570 12144
rect 3528 12109 3556 12135
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3436 11558 3464 11589
rect 3424 11552 3476 11558
rect 3422 11520 3424 11529
rect 3476 11520 3478 11529
rect 3422 11455 3478 11464
rect 3436 11286 3464 11455
rect 3424 11280 3476 11286
rect 3424 11222 3476 11228
rect 3436 10674 3464 11222
rect 3514 10840 3570 10849
rect 3514 10775 3570 10784
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3422 10432 3478 10441
rect 3422 10367 3478 10376
rect 3436 10169 3464 10367
rect 3422 10160 3478 10169
rect 3422 10095 3478 10104
rect 3148 9454 3200 9460
rect 3238 9480 3294 9489
rect 3054 9208 3110 9217
rect 2964 9172 3016 9178
rect 3054 9143 3110 9152
rect 2964 9114 3016 9120
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 3160 8906 3188 9454
rect 3238 9415 3294 9424
rect 3252 9081 3280 9415
rect 3238 9072 3294 9081
rect 3238 9007 3294 9016
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3148 8900 3200 8906
rect 3148 8842 3200 8848
rect 3146 8664 3202 8673
rect 3146 8599 3202 8608
rect 3160 8498 3188 8599
rect 3252 8498 3280 8910
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 2792 7954 2820 8230
rect 3160 8090 3188 8434
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2700 5658 2728 6598
rect 2792 6186 2820 7890
rect 2962 7576 3018 7585
rect 2962 7511 2964 7520
rect 3016 7511 3018 7520
rect 2964 7482 3016 7488
rect 3436 7410 3464 10095
rect 3528 8401 3556 10775
rect 3620 10305 3648 12038
rect 3606 10296 3662 10305
rect 3662 10254 3740 10282
rect 3804 10266 3832 14350
rect 3896 13818 3924 19110
rect 4172 18902 4200 19246
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 4264 18970 4292 19110
rect 4252 18964 4304 18970
rect 4252 18906 4304 18912
rect 4160 18896 4212 18902
rect 4160 18838 4212 18844
rect 3976 18828 4028 18834
rect 3976 18770 4028 18776
rect 3988 17814 4016 18770
rect 4068 18216 4120 18222
rect 4068 18158 4120 18164
rect 3976 17808 4028 17814
rect 3976 17750 4028 17756
rect 4080 17134 4108 18158
rect 4250 17912 4306 17921
rect 4250 17847 4306 17856
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 3976 16788 4028 16794
rect 3976 16730 4028 16736
rect 3988 15638 4016 16730
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 4080 15706 4108 16390
rect 4264 15706 4292 17847
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 4252 15700 4304 15706
rect 4252 15642 4304 15648
rect 3976 15632 4028 15638
rect 3976 15574 4028 15580
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 4080 15473 4108 15506
rect 4066 15464 4122 15473
rect 4066 15399 4122 15408
rect 3974 15192 4030 15201
rect 4080 15162 4108 15399
rect 3974 15127 4030 15136
rect 4068 15156 4120 15162
rect 3988 15094 4016 15127
rect 4068 15098 4120 15104
rect 3976 15088 4028 15094
rect 3976 15030 4028 15036
rect 3988 14958 4016 15030
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 4068 14476 4120 14482
rect 4068 14418 4120 14424
rect 4080 14074 4108 14418
rect 4172 14385 4200 14758
rect 4158 14376 4214 14385
rect 4158 14311 4214 14320
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 4066 13832 4122 13841
rect 3896 13790 4016 13818
rect 3988 13530 4016 13790
rect 4066 13767 4122 13776
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 3988 13433 4016 13466
rect 3974 13424 4030 13433
rect 3974 13359 4030 13368
rect 4080 12918 4108 13767
rect 4356 13530 4384 21984
rect 4540 21146 4568 22034
rect 4620 22024 4672 22030
rect 4618 21992 4620 22001
rect 4672 21992 4674 22001
rect 4618 21927 4674 21936
rect 4724 21690 4752 27095
rect 4816 24410 4844 27520
rect 5368 25362 5396 27520
rect 5356 25356 5408 25362
rect 5356 25298 5408 25304
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6012 24562 6040 27520
rect 6184 24880 6236 24886
rect 6184 24822 6236 24828
rect 6012 24534 6132 24562
rect 4804 24404 4856 24410
rect 4804 24346 4856 24352
rect 6000 24404 6052 24410
rect 6000 24346 6052 24352
rect 5356 24132 5408 24138
rect 5356 24074 5408 24080
rect 5368 23866 5396 24074
rect 5448 24064 5500 24070
rect 5448 24006 5500 24012
rect 5356 23860 5408 23866
rect 5356 23802 5408 23808
rect 4896 23588 4948 23594
rect 4896 23530 4948 23536
rect 4908 23050 4936 23530
rect 5262 23488 5318 23497
rect 5262 23423 5318 23432
rect 5276 23322 5304 23423
rect 5264 23316 5316 23322
rect 5264 23258 5316 23264
rect 5172 23180 5224 23186
rect 5172 23122 5224 23128
rect 4896 23044 4948 23050
rect 4896 22986 4948 22992
rect 4804 22976 4856 22982
rect 4804 22918 4856 22924
rect 4712 21684 4764 21690
rect 4712 21626 4764 21632
rect 4724 21418 4752 21626
rect 4712 21412 4764 21418
rect 4712 21354 4764 21360
rect 4528 21140 4580 21146
rect 4528 21082 4580 21088
rect 4436 20256 4488 20262
rect 4436 20198 4488 20204
rect 4448 19990 4476 20198
rect 4436 19984 4488 19990
rect 4436 19926 4488 19932
rect 4436 19712 4488 19718
rect 4436 19654 4488 19660
rect 4526 19680 4582 19689
rect 4448 19378 4476 19654
rect 4526 19615 4582 19624
rect 4436 19372 4488 19378
rect 4436 19314 4488 19320
rect 4448 18902 4476 19314
rect 4436 18896 4488 18902
rect 4436 18838 4488 18844
rect 4448 18154 4476 18838
rect 4436 18148 4488 18154
rect 4436 18090 4488 18096
rect 4540 16130 4568 19615
rect 4618 18320 4674 18329
rect 4618 18255 4674 18264
rect 4632 17882 4660 18255
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 4632 17338 4660 17818
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4724 16590 4752 16934
rect 4712 16584 4764 16590
rect 4712 16526 4764 16532
rect 4724 16250 4752 16526
rect 4712 16244 4764 16250
rect 4712 16186 4764 16192
rect 4540 16102 4752 16130
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 4540 15502 4568 15846
rect 4528 15496 4580 15502
rect 4528 15438 4580 15444
rect 4540 14550 4568 15438
rect 4528 14544 4580 14550
rect 4528 14486 4580 14492
rect 4540 14074 4568 14486
rect 4528 14068 4580 14074
rect 4528 14010 4580 14016
rect 4344 13524 4396 13530
rect 4344 13466 4396 13472
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4436 13184 4488 13190
rect 4436 13126 4488 13132
rect 4068 12912 4120 12918
rect 4068 12854 4120 12860
rect 4448 12753 4476 13126
rect 4434 12744 4490 12753
rect 4434 12679 4490 12688
rect 4528 12640 4580 12646
rect 4528 12582 4580 12588
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4080 11898 4108 12242
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 4264 11937 4292 12038
rect 4250 11928 4306 11937
rect 4068 11892 4120 11898
rect 4250 11863 4306 11872
rect 4068 11834 4120 11840
rect 3974 11384 4030 11393
rect 4080 11354 4108 11834
rect 3974 11319 4030 11328
rect 4068 11348 4120 11354
rect 3988 10713 4016 11319
rect 4068 11290 4120 11296
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 3974 10704 4030 10713
rect 3884 10668 3936 10674
rect 3974 10639 4030 10648
rect 3884 10610 3936 10616
rect 3606 10231 3662 10240
rect 3514 8392 3570 8401
rect 3514 8327 3570 8336
rect 3608 8356 3660 8362
rect 3608 8298 3660 8304
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2780 6180 2832 6186
rect 2780 6122 2832 6128
rect 2792 5778 2820 6122
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2778 5672 2834 5681
rect 2700 5630 2778 5658
rect 2778 5607 2834 5616
rect 2780 5296 2832 5302
rect 2780 5238 2832 5244
rect 2792 4758 2820 5238
rect 2780 4752 2832 4758
rect 2778 4720 2780 4729
rect 2832 4720 2834 4729
rect 2778 4655 2834 4664
rect 2688 3936 2740 3942
rect 2686 3904 2688 3913
rect 2740 3904 2742 3913
rect 2686 3839 2742 3848
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 2608 2802 2636 3674
rect 2884 3618 2912 7142
rect 3422 7032 3478 7041
rect 3422 6967 3478 6976
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 3068 6254 3096 6734
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 3068 5914 3096 6190
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 2962 5672 3018 5681
rect 2962 5607 3018 5616
rect 2976 4826 3004 5607
rect 3068 5370 3096 5850
rect 3148 5636 3200 5642
rect 3148 5578 3200 5584
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 2964 4616 3016 4622
rect 3160 4604 3188 5578
rect 3016 4576 3188 4604
rect 2964 4558 3016 4564
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 2976 3738 3004 4082
rect 3436 3777 3464 6967
rect 3528 6798 3556 7686
rect 3620 7410 3648 8298
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3620 7002 3648 7346
rect 3712 7342 3740 10254
rect 3792 10260 3844 10266
rect 3792 10202 3844 10208
rect 3804 9518 3832 10202
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3896 8906 3924 10610
rect 4080 10538 4108 11018
rect 4356 10810 4384 11154
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4068 10532 4120 10538
rect 4068 10474 4120 10480
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 3884 8900 3936 8906
rect 3884 8842 3936 8848
rect 4356 7886 4384 9862
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3988 6934 4016 7686
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 3516 6792 3568 6798
rect 3988 6769 4016 6870
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 3516 6734 3568 6740
rect 3974 6760 4030 6769
rect 3974 6695 4030 6704
rect 4080 6662 4108 6802
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 3792 6112 3844 6118
rect 4080 6089 4108 6598
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 3792 6054 3844 6060
rect 4066 6080 4122 6089
rect 3804 5574 3832 6054
rect 4066 6015 4122 6024
rect 4172 5930 4200 6258
rect 4264 6118 4292 6734
rect 4342 6352 4398 6361
rect 4342 6287 4398 6296
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 4080 5902 4200 5930
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3712 5234 3740 5510
rect 3792 5364 3844 5370
rect 3792 5306 3844 5312
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 3620 4865 3648 4966
rect 3606 4856 3662 4865
rect 3606 4791 3662 4800
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 3620 3777 3648 3946
rect 3422 3768 3478 3777
rect 2964 3732 3016 3738
rect 3606 3768 3662 3777
rect 3422 3703 3478 3712
rect 3516 3732 3568 3738
rect 2964 3674 3016 3680
rect 3606 3703 3608 3712
rect 3516 3674 3568 3680
rect 3660 3703 3662 3712
rect 3608 3674 3660 3680
rect 2884 3590 3004 3618
rect 2870 2952 2926 2961
rect 2870 2887 2926 2896
rect 2608 2774 2820 2802
rect 2792 921 2820 2774
rect 2884 2582 2912 2887
rect 2872 2576 2924 2582
rect 2872 2518 2924 2524
rect 2884 1306 2912 2518
rect 2976 1465 3004 3590
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 3146 3224 3202 3233
rect 3146 3159 3202 3168
rect 3160 1986 3188 3159
rect 3436 2650 3464 3334
rect 3528 3194 3556 3674
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3712 2650 3740 5170
rect 3804 4282 3832 5306
rect 3884 5024 3936 5030
rect 3882 4992 3884 5001
rect 3936 4992 3938 5001
rect 3882 4927 3938 4936
rect 4080 4457 4108 5902
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4172 5370 4200 5714
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4160 5160 4212 5166
rect 4158 5128 4160 5137
rect 4212 5128 4214 5137
rect 4158 5063 4214 5072
rect 4172 4826 4200 5063
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4264 4706 4292 6054
rect 4356 5778 4384 6287
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4356 4826 4384 5714
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 4172 4678 4292 4706
rect 4066 4448 4122 4457
rect 4066 4383 4122 4392
rect 3792 4276 3844 4282
rect 3792 4218 3844 4224
rect 3804 3670 3832 4218
rect 4172 4049 4200 4678
rect 4158 4040 4214 4049
rect 4158 3975 4214 3984
rect 4252 4004 4304 4010
rect 4252 3946 4304 3952
rect 3792 3664 3844 3670
rect 3844 3624 3924 3652
rect 3792 3606 3844 3612
rect 3790 2816 3846 2825
rect 3790 2751 3846 2760
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3700 2644 3752 2650
rect 3700 2586 3752 2592
rect 3332 2372 3384 2378
rect 3332 2314 3384 2320
rect 3160 1958 3280 1986
rect 2962 1456 3018 1465
rect 2962 1391 3018 1400
rect 2884 1278 3188 1306
rect 2778 912 2834 921
rect 2778 847 2834 856
rect 3160 480 3188 1278
rect 3252 785 3280 1958
rect 3344 1601 3372 2314
rect 3330 1592 3386 1601
rect 3330 1527 3386 1536
rect 3804 1034 3832 2751
rect 3896 2650 3924 3624
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 4172 2582 4200 3130
rect 4264 3097 4292 3946
rect 4356 3942 4384 4762
rect 4448 4758 4476 12242
rect 4540 11801 4568 12582
rect 4632 12102 4660 13466
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4526 11792 4582 11801
rect 4526 11727 4582 11736
rect 4620 11144 4672 11150
rect 4618 11112 4620 11121
rect 4672 11112 4674 11121
rect 4618 11047 4674 11056
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4540 8430 4568 9318
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4632 8294 4660 9862
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4632 8090 4660 8230
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4540 7177 4568 7822
rect 4526 7168 4582 7177
rect 4526 7103 4582 7112
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4632 6118 4660 6802
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4436 4752 4488 4758
rect 4436 4694 4488 4700
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4344 3936 4396 3942
rect 4632 3913 4660 4422
rect 4618 3904 4674 3913
rect 4344 3878 4396 3884
rect 4540 3862 4618 3890
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4250 3088 4306 3097
rect 4448 3058 4476 3334
rect 4540 3194 4568 3862
rect 4618 3839 4674 3848
rect 4528 3188 4580 3194
rect 4724 3176 4752 16102
rect 4816 11218 4844 22918
rect 4908 22778 4936 22986
rect 4896 22772 4948 22778
rect 4896 22714 4948 22720
rect 5184 22438 5212 23122
rect 5460 22930 5488 24006
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 6012 23866 6040 24346
rect 6104 24342 6132 24534
rect 6092 24336 6144 24342
rect 6092 24278 6144 24284
rect 6104 23866 6132 24278
rect 6000 23860 6052 23866
rect 6000 23802 6052 23808
rect 6092 23860 6144 23866
rect 6092 23802 6144 23808
rect 5998 23352 6054 23361
rect 5998 23287 6054 23296
rect 5460 22902 5580 22930
rect 5552 22681 5580 22902
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5538 22672 5594 22681
rect 5538 22607 5594 22616
rect 5632 22636 5684 22642
rect 5552 22574 5580 22607
rect 5632 22578 5684 22584
rect 5540 22568 5592 22574
rect 5540 22510 5592 22516
rect 5172 22432 5224 22438
rect 5172 22374 5224 22380
rect 5184 22234 5212 22374
rect 5644 22234 5672 22578
rect 5172 22228 5224 22234
rect 5172 22170 5224 22176
rect 5632 22228 5684 22234
rect 5632 22170 5684 22176
rect 5540 22160 5592 22166
rect 5262 22128 5318 22137
rect 5540 22102 5592 22108
rect 5262 22063 5318 22072
rect 5172 21548 5224 21554
rect 5172 21490 5224 21496
rect 4988 21344 5040 21350
rect 4988 21286 5040 21292
rect 5000 21010 5028 21286
rect 4988 21004 5040 21010
rect 4988 20946 5040 20952
rect 4896 20936 4948 20942
rect 4896 20878 4948 20884
rect 4908 20262 4936 20878
rect 5184 20806 5212 21490
rect 5172 20800 5224 20806
rect 5172 20742 5224 20748
rect 4896 20256 4948 20262
rect 4896 20198 4948 20204
rect 4896 19236 4948 19242
rect 4896 19178 4948 19184
rect 4908 18222 4936 19178
rect 5080 19168 5132 19174
rect 5080 19110 5132 19116
rect 5092 18766 5120 19110
rect 5172 18964 5224 18970
rect 5172 18906 5224 18912
rect 5080 18760 5132 18766
rect 5080 18702 5132 18708
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 5080 18148 5132 18154
rect 5080 18090 5132 18096
rect 4896 17672 4948 17678
rect 4896 17614 4948 17620
rect 4908 16658 4936 17614
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 4988 16652 5040 16658
rect 4988 16594 5040 16600
rect 4896 13796 4948 13802
rect 5000 13784 5028 16594
rect 4948 13756 5028 13784
rect 4896 13738 4948 13744
rect 4894 12880 4950 12889
rect 5000 12850 5028 13756
rect 4894 12815 4950 12824
rect 4988 12844 5040 12850
rect 4908 12782 4936 12815
rect 4988 12786 5040 12792
rect 4896 12776 4948 12782
rect 4896 12718 4948 12724
rect 5092 12306 5120 18090
rect 5184 17882 5212 18906
rect 5172 17876 5224 17882
rect 5172 17818 5224 17824
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 5184 17338 5212 17682
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 5172 16720 5224 16726
rect 5172 16662 5224 16668
rect 5184 15706 5212 16662
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 5170 14784 5226 14793
rect 5170 14719 5226 14728
rect 5184 14074 5212 14719
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 5172 12844 5224 12850
rect 5172 12786 5224 12792
rect 5184 12442 5212 12786
rect 5172 12436 5224 12442
rect 5172 12378 5224 12384
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4908 11121 4936 12038
rect 4894 11112 4950 11121
rect 4894 11047 4896 11056
rect 4948 11047 4950 11056
rect 4896 11018 4948 11024
rect 4908 10987 4936 11018
rect 5276 10248 5304 22063
rect 5356 21480 5408 21486
rect 5356 21422 5408 21428
rect 5368 19310 5396 21422
rect 5552 21146 5580 22102
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 6012 21418 6040 23287
rect 6196 22778 6224 24822
rect 6564 24721 6592 27520
rect 6550 24712 6606 24721
rect 6550 24647 6606 24656
rect 6920 24608 6972 24614
rect 6748 24568 6920 24596
rect 6276 23860 6328 23866
rect 6276 23802 6328 23808
rect 6184 22772 6236 22778
rect 6184 22714 6236 22720
rect 6196 22438 6224 22714
rect 6184 22432 6236 22438
rect 6184 22374 6236 22380
rect 6000 21412 6052 21418
rect 6000 21354 6052 21360
rect 6196 21146 6224 22374
rect 5540 21140 5592 21146
rect 5540 21082 5592 21088
rect 6184 21140 6236 21146
rect 6184 21082 6236 21088
rect 6000 21072 6052 21078
rect 6000 21014 6052 21020
rect 5448 21004 5500 21010
rect 5448 20946 5500 20952
rect 5460 19310 5488 20946
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 5552 20602 5580 20742
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5540 20596 5592 20602
rect 5540 20538 5592 20544
rect 6012 20058 6040 21014
rect 6092 20868 6144 20874
rect 6092 20810 6144 20816
rect 6000 20052 6052 20058
rect 6000 19994 6052 20000
rect 6104 19786 6132 20810
rect 6196 20602 6224 21082
rect 6184 20596 6236 20602
rect 6184 20538 6236 20544
rect 6184 20256 6236 20262
rect 6184 20198 6236 20204
rect 6092 19780 6144 19786
rect 6092 19722 6144 19728
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5356 19304 5408 19310
rect 5356 19246 5408 19252
rect 5448 19304 5500 19310
rect 5448 19246 5500 19252
rect 5552 18986 5580 19654
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 6104 19514 6132 19722
rect 6092 19508 6144 19514
rect 6092 19450 6144 19456
rect 6196 19281 6224 20198
rect 6182 19272 6238 19281
rect 6182 19207 6238 19216
rect 5998 19136 6054 19145
rect 5998 19071 6054 19080
rect 5460 18958 5580 18986
rect 5460 18902 5488 18958
rect 5448 18896 5500 18902
rect 5448 18838 5500 18844
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5552 17678 5580 18022
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5632 17264 5684 17270
rect 5630 17232 5632 17241
rect 5684 17232 5686 17241
rect 5630 17167 5686 17176
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5552 16697 5580 17070
rect 5538 16688 5594 16697
rect 6012 16658 6040 19071
rect 6184 17536 6236 17542
rect 6184 17478 6236 17484
rect 5538 16623 5540 16632
rect 5592 16623 5594 16632
rect 6000 16652 6052 16658
rect 5540 16594 5592 16600
rect 6000 16594 6052 16600
rect 5356 16516 5408 16522
rect 5356 16458 5408 16464
rect 5368 16250 5396 16458
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 6012 16130 6040 16594
rect 6092 16584 6144 16590
rect 6090 16552 6092 16561
rect 6144 16552 6146 16561
rect 6090 16487 6146 16496
rect 6104 16250 6132 16487
rect 6092 16244 6144 16250
rect 6092 16186 6144 16192
rect 6012 16102 6132 16130
rect 6104 15978 6132 16102
rect 6092 15972 6144 15978
rect 6092 15914 6144 15920
rect 5724 15904 5776 15910
rect 5724 15846 5776 15852
rect 5736 15706 5764 15846
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5724 15700 5776 15706
rect 5724 15642 5776 15648
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5460 15201 5488 15302
rect 5446 15192 5502 15201
rect 5446 15127 5502 15136
rect 5552 14958 5580 15642
rect 6000 15632 6052 15638
rect 6000 15574 6052 15580
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6012 15026 6040 15574
rect 6104 15337 6132 15914
rect 6090 15328 6146 15337
rect 6090 15263 6146 15272
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 6000 15020 6052 15026
rect 6000 14962 6052 14968
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5460 13784 5488 14758
rect 6012 14618 6040 14962
rect 6000 14612 6052 14618
rect 6000 14554 6052 14560
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5552 14074 5580 14214
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 6104 13938 6132 15098
rect 6196 14929 6224 17478
rect 6182 14920 6238 14929
rect 6182 14855 6238 14864
rect 6184 14476 6236 14482
rect 6184 14418 6236 14424
rect 6196 14074 6224 14418
rect 6184 14068 6236 14074
rect 6184 14010 6236 14016
rect 6092 13932 6144 13938
rect 6092 13874 6144 13880
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 5540 13796 5592 13802
rect 5460 13756 5540 13784
rect 5356 13388 5408 13394
rect 5356 13330 5408 13336
rect 5368 10810 5396 13330
rect 5460 11354 5488 13756
rect 5540 13738 5592 13744
rect 5538 13696 5594 13705
rect 5538 13631 5594 13640
rect 5552 13530 5580 13631
rect 5920 13530 5948 13806
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5908 13524 5960 13530
rect 5908 13466 5960 13472
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 6288 13274 6316 23802
rect 6368 23656 6420 23662
rect 6368 23598 6420 23604
rect 6380 23254 6408 23598
rect 6368 23248 6420 23254
rect 6368 23190 6420 23196
rect 6380 23118 6408 23190
rect 6368 23112 6420 23118
rect 6368 23054 6420 23060
rect 6380 22778 6408 23054
rect 6368 22772 6420 22778
rect 6368 22714 6420 22720
rect 6366 22536 6422 22545
rect 6366 22471 6368 22480
rect 6420 22471 6422 22480
rect 6368 22442 6420 22448
rect 6380 20942 6408 22442
rect 6644 22092 6696 22098
rect 6644 22034 6696 22040
rect 6656 21418 6684 22034
rect 6748 21962 6776 24568
rect 6920 24550 6972 24556
rect 6920 24064 6972 24070
rect 6920 24006 6972 24012
rect 6932 23662 6960 24006
rect 6920 23656 6972 23662
rect 6920 23598 6972 23604
rect 6828 23520 6880 23526
rect 6828 23462 6880 23468
rect 6840 23254 6868 23462
rect 6828 23248 6880 23254
rect 6828 23190 6880 23196
rect 6840 22574 6868 23190
rect 7116 22794 7144 27520
rect 7668 27470 7696 27520
rect 7564 27464 7616 27470
rect 7564 27406 7616 27412
rect 7656 27464 7708 27470
rect 7656 27406 7708 27412
rect 7380 24200 7432 24206
rect 7380 24142 7432 24148
rect 7392 24070 7420 24142
rect 7380 24064 7432 24070
rect 7380 24006 7432 24012
rect 7472 24064 7524 24070
rect 7472 24006 7524 24012
rect 7392 23594 7420 24006
rect 7380 23588 7432 23594
rect 7380 23530 7432 23536
rect 7392 23186 7420 23530
rect 7484 23497 7512 24006
rect 7576 23594 7604 27406
rect 8220 24834 8248 27520
rect 7760 24806 8248 24834
rect 7564 23588 7616 23594
rect 7564 23530 7616 23536
rect 7470 23488 7526 23497
rect 7470 23423 7526 23432
rect 7380 23180 7432 23186
rect 7380 23122 7432 23128
rect 7116 22766 7328 22794
rect 6828 22568 6880 22574
rect 6828 22510 6880 22516
rect 6840 22234 6868 22510
rect 6828 22228 6880 22234
rect 6828 22170 6880 22176
rect 6828 22092 6880 22098
rect 6828 22034 6880 22040
rect 6736 21956 6788 21962
rect 6736 21898 6788 21904
rect 6840 21690 6868 22034
rect 6828 21684 6880 21690
rect 6828 21626 6880 21632
rect 6644 21412 6696 21418
rect 6644 21354 6696 21360
rect 6828 21412 6880 21418
rect 6880 21372 6960 21400
rect 6828 21354 6880 21360
rect 6368 20936 6420 20942
rect 6368 20878 6420 20884
rect 6380 20262 6408 20878
rect 6932 20777 6960 21372
rect 7012 21344 7064 21350
rect 7012 21286 7064 21292
rect 7024 21049 7052 21286
rect 7010 21040 7066 21049
rect 7010 20975 7066 20984
rect 7196 20936 7248 20942
rect 7196 20878 7248 20884
rect 6918 20768 6974 20777
rect 6918 20703 6974 20712
rect 6368 20256 6420 20262
rect 6368 20198 6420 20204
rect 6932 20058 6960 20703
rect 7208 20602 7236 20878
rect 7196 20596 7248 20602
rect 7196 20538 7248 20544
rect 7194 20360 7250 20369
rect 7300 20346 7328 22766
rect 7392 22642 7420 23122
rect 7472 22772 7524 22778
rect 7472 22714 7524 22720
rect 7380 22636 7432 22642
rect 7380 22578 7432 22584
rect 7392 21894 7420 22578
rect 7484 22438 7512 22714
rect 7472 22432 7524 22438
rect 7472 22374 7524 22380
rect 7380 21888 7432 21894
rect 7380 21830 7432 21836
rect 7392 20806 7420 21830
rect 7380 20800 7432 20806
rect 7380 20742 7432 20748
rect 7250 20318 7328 20346
rect 7380 20392 7432 20398
rect 7484 20380 7512 22374
rect 7656 21888 7708 21894
rect 7656 21830 7708 21836
rect 7564 21412 7616 21418
rect 7564 21354 7616 21360
rect 7576 21146 7604 21354
rect 7668 21350 7696 21830
rect 7656 21344 7708 21350
rect 7656 21286 7708 21292
rect 7564 21140 7616 21146
rect 7564 21082 7616 21088
rect 7432 20352 7512 20380
rect 7380 20334 7432 20340
rect 7194 20295 7250 20304
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 6644 19780 6696 19786
rect 6644 19722 6696 19728
rect 6460 18828 6512 18834
rect 6460 18770 6512 18776
rect 6368 18624 6420 18630
rect 6368 18566 6420 18572
rect 6380 15065 6408 18566
rect 6472 18154 6500 18770
rect 6656 18766 6684 19722
rect 6932 19514 6960 19994
rect 7012 19848 7064 19854
rect 7012 19790 7064 19796
rect 6920 19508 6972 19514
rect 6920 19450 6972 19456
rect 7024 19378 7052 19790
rect 7196 19508 7248 19514
rect 7196 19450 7248 19456
rect 7012 19372 7064 19378
rect 7012 19314 7064 19320
rect 7012 19236 7064 19242
rect 7012 19178 7064 19184
rect 7024 18970 7052 19178
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6644 18760 6696 18766
rect 6550 18728 6606 18737
rect 6644 18702 6696 18708
rect 6550 18663 6606 18672
rect 6460 18148 6512 18154
rect 6460 18090 6512 18096
rect 6460 17536 6512 17542
rect 6460 17478 6512 17484
rect 6472 17338 6500 17478
rect 6460 17332 6512 17338
rect 6460 17274 6512 17280
rect 6472 17134 6500 17274
rect 6460 17128 6512 17134
rect 6460 17070 6512 17076
rect 6458 15192 6514 15201
rect 6458 15127 6514 15136
rect 6366 15056 6422 15065
rect 6366 14991 6422 15000
rect 6472 14958 6500 15127
rect 6460 14952 6512 14958
rect 6460 14894 6512 14900
rect 6460 14408 6512 14414
rect 6460 14350 6512 14356
rect 6472 14074 6500 14350
rect 6460 14068 6512 14074
rect 6460 14010 6512 14016
rect 6564 13530 6592 18663
rect 6656 17814 6684 18702
rect 6748 18086 6776 18770
rect 6920 18692 6972 18698
rect 6840 18652 6920 18680
rect 6736 18080 6788 18086
rect 6736 18022 6788 18028
rect 6840 17882 6868 18652
rect 6920 18634 6972 18640
rect 7024 18290 7052 18906
rect 7012 18284 7064 18290
rect 7012 18226 7064 18232
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6644 17808 6696 17814
rect 6644 17750 6696 17756
rect 6736 17740 6788 17746
rect 6736 17682 6788 17688
rect 6748 16794 6776 17682
rect 6828 17536 6880 17542
rect 7024 17524 7052 18226
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 6880 17496 7052 17524
rect 6828 17478 6880 17484
rect 6840 17338 6868 17478
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 6656 16153 6684 16186
rect 6736 16176 6788 16182
rect 6642 16144 6698 16153
rect 6736 16118 6788 16124
rect 6642 16079 6698 16088
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 6656 15570 6684 15982
rect 6644 15564 6696 15570
rect 6644 15506 6696 15512
rect 6656 15094 6684 15506
rect 6644 15088 6696 15094
rect 6644 15030 6696 15036
rect 6656 14074 6684 15030
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6552 13524 6604 13530
rect 6552 13466 6604 13472
rect 6366 13424 6422 13433
rect 6366 13359 6368 13368
rect 6420 13359 6422 13368
rect 6368 13330 6420 13336
rect 6460 13320 6512 13326
rect 5552 12968 5580 13262
rect 6288 13246 6408 13274
rect 6460 13262 6512 13268
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5552 12940 5672 12968
rect 5644 12646 5672 12940
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5644 12481 5672 12582
rect 5630 12472 5686 12481
rect 5630 12407 5686 12416
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5552 11880 5580 12038
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5552 11852 5672 11880
rect 5540 11620 5592 11626
rect 5540 11562 5592 11568
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5356 10804 5408 10810
rect 5552 10792 5580 11562
rect 5644 11558 5672 11852
rect 6012 11626 6040 12242
rect 6000 11620 6052 11626
rect 6000 11562 6052 11568
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5644 11354 5672 11494
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 6000 11280 6052 11286
rect 6000 11222 6052 11228
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5356 10746 5408 10752
rect 5460 10764 5580 10792
rect 5184 10220 5304 10248
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 5000 9382 5028 9998
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 5000 8537 5028 9318
rect 4986 8528 5042 8537
rect 4986 8463 5042 8472
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4816 7206 4844 7822
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4816 6798 4844 7142
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 4816 5914 4844 6734
rect 5000 6458 5028 8463
rect 5184 7585 5212 10220
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 5276 9722 5304 10066
rect 5460 10062 5488 10764
rect 6012 10674 6040 11222
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 5460 9042 5488 9998
rect 5552 9926 5580 10542
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5644 10266 5672 10406
rect 5998 10296 6054 10305
rect 5632 10260 5684 10266
rect 5998 10231 6054 10240
rect 5632 10202 5684 10208
rect 5540 9920 5592 9926
rect 6012 9897 6040 10231
rect 5540 9862 5592 9868
rect 5998 9888 6054 9897
rect 5552 9178 5580 9862
rect 5622 9820 5918 9840
rect 5998 9823 6054 9832
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 5552 7750 5580 8978
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6288 8430 6316 8978
rect 6276 8424 6328 8430
rect 6276 8366 6328 8372
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 6012 7750 6040 7890
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 5170 7576 5226 7585
rect 5170 7511 5226 7520
rect 5552 7392 5580 7686
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5816 7404 5868 7410
rect 5552 7364 5764 7392
rect 5460 7274 5672 7290
rect 5460 7268 5684 7274
rect 5460 7262 5632 7268
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 5000 6254 5028 6394
rect 5184 6322 5212 6598
rect 5460 6458 5488 7262
rect 5632 7210 5684 7216
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5552 6905 5580 7142
rect 5538 6896 5594 6905
rect 5538 6831 5594 6840
rect 5736 6730 5764 7364
rect 6012 7392 6040 7686
rect 6090 7576 6146 7585
rect 6090 7511 6146 7520
rect 5868 7364 6040 7392
rect 5816 7346 5868 7352
rect 5828 6934 5856 7346
rect 6104 7274 6132 7511
rect 6092 7268 6144 7274
rect 6092 7210 6144 7216
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 5816 6928 5868 6934
rect 5816 6870 5868 6876
rect 6012 6798 6040 7142
rect 6000 6792 6052 6798
rect 6052 6752 6132 6780
rect 6000 6734 6052 6740
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 6012 6322 6040 6598
rect 6104 6390 6132 6752
rect 6092 6384 6144 6390
rect 6092 6326 6144 6332
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 6104 6118 6132 6326
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 5460 5166 5488 6054
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6104 5370 6132 6054
rect 6196 5914 6224 8230
rect 6380 7834 6408 13246
rect 6472 12918 6500 13262
rect 6564 12986 6592 13262
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6460 12912 6512 12918
rect 6460 12854 6512 12860
rect 6472 11801 6500 12854
rect 6564 11898 6592 12922
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6458 11792 6514 11801
rect 6458 11727 6514 11736
rect 6656 11694 6684 14010
rect 6748 13326 6776 16118
rect 6840 15473 6868 16934
rect 7010 16552 7066 16561
rect 7010 16487 7066 16496
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6932 15978 6960 16390
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 6826 15464 6882 15473
rect 6826 15399 6882 15408
rect 6932 15366 6960 15914
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6932 15162 6960 15302
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6840 13870 6868 14758
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6826 13560 6882 13569
rect 6826 13495 6882 13504
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6748 12442 6776 12786
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6656 11558 6684 11630
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6656 10606 6684 11494
rect 6748 11286 6776 12378
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6840 10130 6868 13495
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6932 11354 6960 11630
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6932 10198 6960 11018
rect 6920 10192 6972 10198
rect 6920 10134 6972 10140
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6552 9988 6604 9994
rect 6552 9930 6604 9936
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6288 7806 6408 7834
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5184 4826 5212 4966
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 4896 4004 4948 4010
rect 4896 3946 4948 3952
rect 4908 3398 4936 3946
rect 5184 3738 5212 4762
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 4896 3392 4948 3398
rect 4894 3360 4896 3369
rect 4948 3360 4950 3369
rect 4894 3295 4950 3304
rect 4724 3148 4844 3176
rect 4528 3130 4580 3136
rect 4250 3023 4306 3032
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4252 2916 4304 2922
rect 4252 2858 4304 2864
rect 4160 2576 4212 2582
rect 4160 2518 4212 2524
rect 4066 2000 4122 2009
rect 4066 1935 4122 1944
rect 4080 1737 4108 1935
rect 4066 1728 4122 1737
rect 4066 1663 4122 1672
rect 4172 1329 4200 2518
rect 4158 1320 4214 1329
rect 4158 1255 4214 1264
rect 3712 1006 3832 1034
rect 3238 776 3294 785
rect 3238 711 3294 720
rect 3712 480 3740 1006
rect 4264 480 4292 2858
rect 4816 480 4844 3148
rect 4908 2990 4936 3295
rect 4896 2984 4948 2990
rect 4896 2926 4948 2932
rect 5264 2916 5316 2922
rect 5264 2858 5316 2864
rect 5276 2553 5304 2858
rect 5262 2544 5318 2553
rect 5262 2479 5318 2488
rect 5368 480 5396 4694
rect 5552 4690 5580 4966
rect 5540 4684 5592 4690
rect 5460 4644 5540 4672
rect 5460 4321 5488 4644
rect 5540 4626 5592 4632
rect 5644 4554 5672 4966
rect 5998 4856 6054 4865
rect 5998 4791 6000 4800
rect 6052 4791 6054 4800
rect 6000 4762 6052 4768
rect 5632 4548 5684 4554
rect 5632 4490 5684 4496
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5446 4312 5502 4321
rect 5446 4247 5502 4256
rect 5552 3777 5580 4422
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6012 4282 6040 4762
rect 6104 4758 6132 5306
rect 6196 5302 6224 5850
rect 6184 5296 6236 5302
rect 6184 5238 6236 5244
rect 6184 5160 6236 5166
rect 6288 5137 6316 7806
rect 6368 7744 6420 7750
rect 6472 7732 6500 9318
rect 6564 9178 6592 9930
rect 6736 9716 6788 9722
rect 6840 9704 6868 10066
rect 6788 9676 6868 9704
rect 6736 9658 6788 9664
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6420 7704 6500 7732
rect 6368 7686 6420 7692
rect 6380 7206 6408 7686
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6472 6118 6500 6258
rect 6460 6112 6512 6118
rect 6460 6054 6512 6060
rect 6472 5914 6500 6054
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 6550 5536 6606 5545
rect 6550 5471 6606 5480
rect 6368 5296 6420 5302
rect 6368 5238 6420 5244
rect 6184 5102 6236 5108
rect 6274 5128 6330 5137
rect 6092 4752 6144 4758
rect 6092 4694 6144 4700
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 5538 3768 5594 3777
rect 5538 3703 5594 3712
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5446 3088 5502 3097
rect 5446 3023 5502 3032
rect 5460 2650 5488 3023
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6012 480 6040 4014
rect 6104 4010 6132 4558
rect 6092 4004 6144 4010
rect 6092 3946 6144 3952
rect 6104 3738 6132 3946
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 6196 2854 6224 5102
rect 6274 5063 6330 5072
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6184 2848 6236 2854
rect 6182 2816 6184 2825
rect 6236 2816 6238 2825
rect 6182 2751 6238 2760
rect 294 0 350 480
rect 846 0 902 480
rect 1398 0 1454 480
rect 1950 0 2006 480
rect 2502 0 2558 480
rect 3146 0 3202 480
rect 3698 0 3754 480
rect 4250 0 4306 480
rect 4802 0 4858 480
rect 5354 0 5410 480
rect 5998 0 6054 480
rect 6288 377 6316 4966
rect 6380 3670 6408 5238
rect 6368 3664 6420 3670
rect 6368 3606 6420 3612
rect 6380 2650 6408 3606
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 6564 480 6592 5471
rect 6656 4865 6684 8434
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6748 5760 6776 8366
rect 6932 8362 6960 8774
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6826 7304 6882 7313
rect 6826 7239 6882 7248
rect 6840 7206 6868 7239
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6932 7018 6960 7346
rect 6840 6990 6960 7018
rect 6840 6458 6868 6990
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6920 5772 6972 5778
rect 6748 5732 6920 5760
rect 6748 5098 6776 5732
rect 6920 5714 6972 5720
rect 6920 5636 6972 5642
rect 6920 5578 6972 5584
rect 6932 5522 6960 5578
rect 6840 5494 6960 5522
rect 6840 5302 6868 5494
rect 6828 5296 6880 5302
rect 6828 5238 6880 5244
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6736 5092 6788 5098
rect 6736 5034 6788 5040
rect 6642 4856 6698 4865
rect 6840 4826 6868 5102
rect 6642 4791 6698 4800
rect 6828 4820 6880 4826
rect 6656 3505 6684 4791
rect 6828 4762 6880 4768
rect 6828 4684 6880 4690
rect 6880 4644 6960 4672
rect 6828 4626 6880 4632
rect 6736 4548 6788 4554
rect 6736 4490 6788 4496
rect 6642 3496 6698 3505
rect 6642 3431 6698 3440
rect 6748 2825 6776 4490
rect 6932 3534 6960 4644
rect 7024 3670 7052 16487
rect 7116 13977 7144 18022
rect 7208 15201 7236 19450
rect 7300 19417 7328 20318
rect 7392 19854 7420 20334
rect 7380 19848 7432 19854
rect 7380 19790 7432 19796
rect 7286 19408 7342 19417
rect 7286 19343 7342 19352
rect 7392 18970 7420 19790
rect 7668 19514 7696 21286
rect 7656 19508 7708 19514
rect 7656 19450 7708 19456
rect 7472 19440 7524 19446
rect 7472 19382 7524 19388
rect 7380 18964 7432 18970
rect 7380 18906 7432 18912
rect 7484 18834 7512 19382
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7472 18828 7524 18834
rect 7472 18770 7524 18776
rect 7380 18148 7432 18154
rect 7380 18090 7432 18096
rect 7392 17542 7420 18090
rect 7380 17536 7432 17542
rect 7576 17513 7604 19314
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7380 17478 7432 17484
rect 7562 17504 7618 17513
rect 7392 17202 7420 17478
rect 7562 17439 7618 17448
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7472 16720 7524 16726
rect 7472 16662 7524 16668
rect 7484 16153 7512 16662
rect 7470 16144 7526 16153
rect 7470 16079 7526 16088
rect 7576 15484 7604 17439
rect 7668 17066 7696 18566
rect 7656 17060 7708 17066
rect 7656 17002 7708 17008
rect 7760 16726 7788 24806
rect 7840 24608 7892 24614
rect 7840 24550 7892 24556
rect 7852 24410 7880 24550
rect 7840 24404 7892 24410
rect 7840 24346 7892 24352
rect 8116 24200 8168 24206
rect 8116 24142 8168 24148
rect 8022 23760 8078 23769
rect 8022 23695 8078 23704
rect 7932 23588 7984 23594
rect 7932 23530 7984 23536
rect 7838 22264 7894 22273
rect 7838 22199 7894 22208
rect 7852 21146 7880 22199
rect 7840 21140 7892 21146
rect 7840 21082 7892 21088
rect 7944 19802 7972 23530
rect 8036 20097 8064 23695
rect 8128 23526 8156 24142
rect 8116 23520 8168 23526
rect 8116 23462 8168 23468
rect 8864 23361 8892 27520
rect 9416 24834 9444 27520
rect 9140 24806 9444 24834
rect 9036 24132 9088 24138
rect 9036 24074 9088 24080
rect 9048 23866 9076 24074
rect 9036 23860 9088 23866
rect 9036 23802 9088 23808
rect 8850 23352 8906 23361
rect 8850 23287 8906 23296
rect 8484 22976 8536 22982
rect 8484 22918 8536 22924
rect 8392 22704 8444 22710
rect 8390 22672 8392 22681
rect 8444 22672 8446 22681
rect 8496 22642 8524 22918
rect 8390 22607 8446 22616
rect 8484 22636 8536 22642
rect 8484 22578 8536 22584
rect 8116 22432 8168 22438
rect 8116 22374 8168 22380
rect 8484 22432 8536 22438
rect 8484 22374 8536 22380
rect 8128 21729 8156 22374
rect 8496 22234 8524 22374
rect 8484 22228 8536 22234
rect 8484 22170 8536 22176
rect 8760 22092 8812 22098
rect 8760 22034 8812 22040
rect 8772 22001 8800 22034
rect 8758 21992 8814 22001
rect 8758 21927 8814 21936
rect 8114 21720 8170 21729
rect 8114 21655 8170 21664
rect 8128 21486 8156 21655
rect 8208 21548 8260 21554
rect 8208 21490 8260 21496
rect 8116 21480 8168 21486
rect 8116 21422 8168 21428
rect 8116 20800 8168 20806
rect 8116 20742 8168 20748
rect 8022 20088 8078 20097
rect 8022 20023 8078 20032
rect 7852 19774 7972 19802
rect 7852 19446 7880 19774
rect 7932 19712 7984 19718
rect 7932 19654 7984 19660
rect 7840 19440 7892 19446
rect 7840 19382 7892 19388
rect 7944 19242 7972 19654
rect 7932 19236 7984 19242
rect 7932 19178 7984 19184
rect 7840 18760 7892 18766
rect 7840 18702 7892 18708
rect 7852 17678 7880 18702
rect 7944 18601 7972 19178
rect 8022 19000 8078 19009
rect 8022 18935 8024 18944
rect 8076 18935 8078 18944
rect 8024 18906 8076 18912
rect 7930 18592 7986 18601
rect 7930 18527 7986 18536
rect 8036 18358 8064 18906
rect 8024 18352 8076 18358
rect 8024 18294 8076 18300
rect 7840 17672 7892 17678
rect 7840 17614 7892 17620
rect 7748 16720 7800 16726
rect 7748 16662 7800 16668
rect 7840 16652 7892 16658
rect 7840 16594 7892 16600
rect 7748 16584 7800 16590
rect 7748 16526 7800 16532
rect 7760 15706 7788 16526
rect 7852 15910 7880 16594
rect 7932 16040 7984 16046
rect 7932 15982 7984 15988
rect 7840 15904 7892 15910
rect 7840 15846 7892 15852
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 7576 15456 7696 15484
rect 7194 15192 7250 15201
rect 7194 15127 7250 15136
rect 7194 15056 7250 15065
rect 7194 14991 7250 15000
rect 7208 14958 7236 14991
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7300 14278 7328 14758
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7300 14074 7328 14214
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7102 13968 7158 13977
rect 7102 13903 7158 13912
rect 7564 13932 7616 13938
rect 7564 13874 7616 13880
rect 7380 13728 7432 13734
rect 7380 13670 7432 13676
rect 7196 12640 7248 12646
rect 7196 12582 7248 12588
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7208 12345 7236 12582
rect 7300 12442 7328 12582
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7194 12336 7250 12345
rect 7194 12271 7250 12280
rect 7208 10810 7236 12271
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7116 9722 7144 10542
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7208 8498 7236 8774
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7208 6361 7236 8434
rect 7300 7410 7328 8774
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7392 7002 7420 13670
rect 7576 13530 7604 13874
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7484 11354 7512 12242
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7484 9518 7512 9862
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7484 8090 7512 9454
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7484 7410 7512 8026
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7392 6662 7420 6802
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7194 6352 7250 6361
rect 7392 6322 7420 6598
rect 7194 6287 7250 6296
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7116 4826 7144 6190
rect 7196 6180 7248 6186
rect 7196 6122 7248 6128
rect 7208 5914 7236 6122
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7300 5953 7328 6054
rect 7286 5944 7342 5953
rect 7196 5908 7248 5914
rect 7286 5879 7342 5888
rect 7196 5850 7248 5856
rect 7300 5710 7328 5879
rect 7288 5704 7340 5710
rect 7576 5658 7604 7890
rect 7288 5646 7340 5652
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7208 3942 7236 4626
rect 7300 4554 7328 5646
rect 7484 5630 7604 5658
rect 7288 4548 7340 4554
rect 7288 4490 7340 4496
rect 7300 4214 7328 4490
rect 7288 4208 7340 4214
rect 7288 4150 7340 4156
rect 7484 4078 7512 5630
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7576 5166 7604 5510
rect 7564 5160 7616 5166
rect 7564 5102 7616 5108
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 7576 4321 7604 4558
rect 7562 4312 7618 4321
rect 7562 4247 7564 4256
rect 7616 4247 7618 4256
rect 7564 4218 7616 4224
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7196 3936 7248 3942
rect 7102 3904 7158 3913
rect 7196 3878 7248 3884
rect 7102 3839 7158 3848
rect 7012 3664 7064 3670
rect 7012 3606 7064 3612
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6734 2816 6790 2825
rect 6734 2751 6790 2760
rect 6918 2544 6974 2553
rect 6918 2479 6974 2488
rect 6932 2446 6960 2479
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 7116 480 7144 3839
rect 7208 3641 7236 3878
rect 7194 3632 7250 3641
rect 7194 3567 7196 3576
rect 7248 3567 7250 3576
rect 7196 3538 7248 3544
rect 7208 3507 7236 3538
rect 7472 3460 7524 3466
rect 7472 3402 7524 3408
rect 7484 3058 7512 3402
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7286 2952 7342 2961
rect 7286 2887 7288 2896
rect 7340 2887 7342 2896
rect 7288 2858 7340 2864
rect 7288 2304 7340 2310
rect 7286 2272 7288 2281
rect 7340 2272 7342 2281
rect 7286 2207 7342 2216
rect 7668 480 7696 15456
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 7760 10742 7788 11154
rect 7748 10736 7800 10742
rect 7748 10678 7800 10684
rect 7748 8356 7800 8362
rect 7748 8298 7800 8304
rect 7760 4690 7788 8298
rect 7852 5545 7880 15846
rect 7944 15638 7972 15982
rect 7932 15632 7984 15638
rect 7932 15574 7984 15580
rect 7932 15020 7984 15026
rect 7932 14962 7984 14968
rect 7944 14618 7972 14962
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 7930 14104 7986 14113
rect 7930 14039 7986 14048
rect 7944 13870 7972 14039
rect 7932 13864 7984 13870
rect 7932 13806 7984 13812
rect 7944 13462 7972 13806
rect 7932 13456 7984 13462
rect 7932 13398 7984 13404
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 7944 12986 7972 13262
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 8036 12306 8064 13126
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 7944 9489 7972 9522
rect 7930 9480 7986 9489
rect 7930 9415 7986 9424
rect 8036 9353 8064 9862
rect 8128 9654 8156 20742
rect 8220 20618 8248 21490
rect 8392 20800 8444 20806
rect 8392 20742 8444 20748
rect 8220 20602 8340 20618
rect 8220 20596 8352 20602
rect 8220 20590 8300 20596
rect 8300 20538 8352 20544
rect 8404 20330 8432 20742
rect 8392 20324 8444 20330
rect 8392 20266 8444 20272
rect 8404 19718 8432 20266
rect 8482 19952 8538 19961
rect 8482 19887 8538 19896
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8298 19408 8354 19417
rect 8404 19378 8432 19654
rect 8298 19343 8354 19352
rect 8392 19372 8444 19378
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 8220 19009 8248 19110
rect 8206 19000 8262 19009
rect 8206 18935 8262 18944
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8220 17746 8248 18702
rect 8208 17740 8260 17746
rect 8208 17682 8260 17688
rect 8220 17202 8248 17682
rect 8208 17196 8260 17202
rect 8208 17138 8260 17144
rect 8208 17060 8260 17066
rect 8208 17002 8260 17008
rect 8220 16794 8248 17002
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 8312 14498 8340 19343
rect 8392 19314 8444 19320
rect 8404 19174 8432 19314
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8404 18426 8432 19110
rect 8392 18420 8444 18426
rect 8392 18362 8444 18368
rect 8312 14470 8432 14498
rect 8300 13728 8352 13734
rect 8300 13670 8352 13676
rect 8208 13252 8260 13258
rect 8312 13240 8340 13670
rect 8404 13530 8432 14470
rect 8496 14074 8524 19887
rect 8574 18864 8630 18873
rect 8574 18799 8630 18808
rect 8588 17338 8616 18799
rect 8576 17332 8628 17338
rect 8576 17274 8628 17280
rect 8668 17128 8720 17134
rect 8668 17070 8720 17076
rect 8680 16794 8708 17070
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8576 16040 8628 16046
rect 8576 15982 8628 15988
rect 8588 15162 8616 15982
rect 8576 15156 8628 15162
rect 8576 15098 8628 15104
rect 8588 14958 8616 15098
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8496 13802 8524 14010
rect 8484 13796 8536 13802
rect 8484 13738 8536 13744
rect 8588 13682 8616 14894
rect 8772 14006 8800 21927
rect 8850 21448 8906 21457
rect 8850 21383 8852 21392
rect 8904 21383 8906 21392
rect 8852 21354 8904 21360
rect 8944 21344 8996 21350
rect 8944 21286 8996 21292
rect 9036 21344 9088 21350
rect 9036 21286 9088 21292
rect 8850 20224 8906 20233
rect 8850 20159 8906 20168
rect 8864 18850 8892 20159
rect 8956 19310 8984 21286
rect 9048 21146 9076 21286
rect 9036 21140 9088 21146
rect 9036 21082 9088 21088
rect 9048 20058 9076 21082
rect 9036 20052 9088 20058
rect 9036 19994 9088 20000
rect 8944 19304 8996 19310
rect 8944 19246 8996 19252
rect 8956 18970 8984 19246
rect 8944 18964 8996 18970
rect 8944 18906 8996 18912
rect 8864 18822 8984 18850
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8760 14000 8812 14006
rect 8760 13942 8812 13948
rect 8864 13870 8892 14214
rect 8852 13864 8904 13870
rect 8850 13832 8852 13841
rect 8904 13832 8906 13841
rect 8850 13767 8906 13776
rect 8760 13728 8812 13734
rect 8588 13654 8708 13682
rect 8956 13682 8984 18822
rect 9036 17876 9088 17882
rect 9036 17818 9088 17824
rect 9048 16114 9076 17818
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 9140 15201 9168 24806
rect 9864 23656 9916 23662
rect 9586 23624 9642 23633
rect 9864 23598 9916 23604
rect 9586 23559 9642 23568
rect 9600 23089 9628 23559
rect 9876 23322 9904 23598
rect 9968 23474 9996 27520
rect 10520 25786 10548 27520
rect 10520 25758 10732 25786
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10704 24041 10732 25758
rect 11072 24857 11100 27520
rect 11058 24848 11114 24857
rect 11058 24783 11114 24792
rect 10782 24712 10838 24721
rect 10782 24647 10838 24656
rect 10690 24032 10746 24041
rect 10690 23967 10746 23976
rect 10796 23866 10824 24647
rect 10784 23860 10836 23866
rect 10784 23802 10836 23808
rect 10784 23656 10836 23662
rect 10784 23598 10836 23604
rect 11426 23624 11482 23633
rect 9968 23446 10180 23474
rect 9864 23316 9916 23322
rect 9864 23258 9916 23264
rect 9772 23180 9824 23186
rect 9772 23122 9824 23128
rect 9586 23080 9642 23089
rect 9586 23015 9642 23024
rect 9402 22536 9458 22545
rect 9402 22471 9458 22480
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9232 17134 9260 19110
rect 9416 18737 9444 22471
rect 9496 21888 9548 21894
rect 9496 21830 9548 21836
rect 9508 21554 9536 21830
rect 9496 21548 9548 21554
rect 9496 21490 9548 21496
rect 9508 21078 9536 21490
rect 9496 21072 9548 21078
rect 9496 21014 9548 21020
rect 9496 18896 9548 18902
rect 9496 18838 9548 18844
rect 9402 18728 9458 18737
rect 9402 18663 9458 18672
rect 9404 18624 9456 18630
rect 9404 18566 9456 18572
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 9220 17128 9272 17134
rect 9220 17070 9272 17076
rect 9324 16250 9352 18362
rect 9416 18154 9444 18566
rect 9508 18222 9536 18838
rect 9496 18216 9548 18222
rect 9496 18158 9548 18164
rect 9404 18148 9456 18154
rect 9404 18090 9456 18096
rect 9416 16522 9444 18090
rect 9508 17882 9536 18158
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9496 17672 9548 17678
rect 9494 17640 9496 17649
rect 9548 17640 9550 17649
rect 9494 17575 9550 17584
rect 9496 17196 9548 17202
rect 9496 17138 9548 17144
rect 9508 16794 9536 17138
rect 9496 16788 9548 16794
rect 9496 16730 9548 16736
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 9126 15192 9182 15201
rect 9126 15127 9182 15136
rect 9140 14113 9168 15127
rect 9324 14958 9352 16186
rect 9416 15706 9444 16458
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 9126 14104 9182 14113
rect 9126 14039 9182 14048
rect 9312 14000 9364 14006
rect 9218 13968 9274 13977
rect 9312 13942 9364 13948
rect 9218 13903 9274 13912
rect 9232 13802 9260 13903
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 8760 13670 8812 13676
rect 8574 13560 8630 13569
rect 8392 13524 8444 13530
rect 8574 13495 8630 13504
rect 8392 13466 8444 13472
rect 8392 13388 8444 13394
rect 8392 13330 8444 13336
rect 8260 13212 8340 13240
rect 8208 13194 8260 13200
rect 8220 12442 8248 13194
rect 8404 12986 8432 13330
rect 8484 13320 8536 13326
rect 8588 13297 8616 13495
rect 8484 13262 8536 13268
rect 8574 13288 8630 13297
rect 8496 13161 8524 13262
rect 8574 13223 8630 13232
rect 8482 13152 8538 13161
rect 8482 13087 8538 13096
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8680 12850 8708 13654
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 8312 11898 8340 12174
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8496 11830 8524 12174
rect 8772 11898 8800 13670
rect 8864 13654 8984 13682
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8484 11824 8536 11830
rect 8484 11766 8536 11772
rect 8496 11626 8524 11766
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8220 11354 8248 11494
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8220 10538 8248 11290
rect 8312 11218 8340 11290
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8404 10985 8432 11086
rect 8576 11008 8628 11014
rect 8390 10976 8446 10985
rect 8864 10985 8892 13654
rect 8944 13524 8996 13530
rect 8944 13466 8996 13472
rect 8956 12866 8984 13466
rect 9036 13388 9088 13394
rect 9036 13330 9088 13336
rect 9048 12986 9076 13330
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 8956 12838 9076 12866
rect 9048 12458 9076 12838
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 9039 12430 9076 12458
rect 9140 12442 9168 12786
rect 9324 12594 9352 13942
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 9416 13190 9444 13874
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9416 13025 9444 13126
rect 9402 13016 9458 13025
rect 9402 12951 9458 12960
rect 9416 12782 9444 12951
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9324 12566 9444 12594
rect 9128 12436 9180 12442
rect 9039 12356 9067 12430
rect 9128 12378 9180 12384
rect 9039 12328 9076 12356
rect 8942 11792 8998 11801
rect 8942 11727 8998 11736
rect 8956 11354 8984 11727
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 8576 10950 8628 10956
rect 8850 10976 8906 10985
rect 8390 10911 8446 10920
rect 8404 10810 8432 10911
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8208 10532 8260 10538
rect 8208 10474 8260 10480
rect 8220 10198 8248 10474
rect 8588 10198 8616 10950
rect 8850 10911 8906 10920
rect 8760 10736 8812 10742
rect 8760 10678 8812 10684
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8576 10192 8628 10198
rect 8576 10134 8628 10140
rect 8772 10130 8800 10678
rect 8760 10124 8812 10130
rect 8760 10066 8812 10072
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8116 9648 8168 9654
rect 8116 9590 8168 9596
rect 8312 9382 8340 9998
rect 8390 9480 8446 9489
rect 8390 9415 8446 9424
rect 8300 9376 8352 9382
rect 8022 9344 8078 9353
rect 8300 9318 8352 9324
rect 8022 9279 8078 9288
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 8036 9081 8064 9114
rect 8022 9072 8078 9081
rect 8022 9007 8078 9016
rect 8312 8906 8340 9318
rect 8404 9178 8432 9415
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7944 6254 7972 6598
rect 7932 6248 7984 6254
rect 7932 6190 7984 6196
rect 7930 6080 7986 6089
rect 7930 6015 7986 6024
rect 7944 5914 7972 6015
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 7838 5536 7894 5545
rect 7838 5471 7894 5480
rect 8024 5024 8076 5030
rect 8024 4966 8076 4972
rect 7748 4684 7800 4690
rect 7748 4626 7800 4632
rect 7746 4448 7802 4457
rect 7746 4383 7802 4392
rect 7760 3942 7788 4383
rect 8036 4049 8064 4966
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 8128 4214 8156 4422
rect 8116 4208 8168 4214
rect 8116 4150 8168 4156
rect 8220 4078 8248 8774
rect 8312 8634 8340 8842
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8312 8090 8340 8570
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8404 7585 8432 7686
rect 8390 7576 8446 7585
rect 8390 7511 8446 7520
rect 8496 7342 8524 7686
rect 8588 7546 8616 7822
rect 8680 7546 8708 9114
rect 8944 8832 8996 8838
rect 8944 8774 8996 8780
rect 8760 7812 8812 7818
rect 8760 7754 8812 7760
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8588 7342 8616 7482
rect 8484 7336 8536 7342
rect 8484 7278 8536 7284
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 8482 6896 8538 6905
rect 8482 6831 8484 6840
rect 8536 6831 8538 6840
rect 8484 6802 8536 6808
rect 8390 6760 8446 6769
rect 8390 6695 8446 6704
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8312 6186 8340 6598
rect 8404 6458 8432 6695
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 8298 5808 8354 5817
rect 8298 5743 8300 5752
rect 8352 5743 8354 5752
rect 8300 5714 8352 5720
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8588 5273 8616 5646
rect 8574 5264 8630 5273
rect 8574 5199 8630 5208
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8208 4072 8260 4078
rect 8022 4040 8078 4049
rect 8022 3975 8078 3984
rect 8128 4020 8208 4026
rect 8128 4014 8260 4020
rect 8128 3998 8248 4014
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7760 3058 7788 3334
rect 7852 3194 7880 3878
rect 7932 3732 7984 3738
rect 7984 3692 8064 3720
rect 7932 3674 7984 3680
rect 7932 3596 7984 3602
rect 7932 3538 7984 3544
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7944 2650 7972 3538
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 8036 1465 8064 3692
rect 8128 2650 8156 3998
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 8022 1456 8078 1465
rect 8022 1391 8078 1400
rect 7746 1320 7802 1329
rect 7746 1255 7802 1264
rect 7930 1320 7986 1329
rect 7930 1255 7986 1264
rect 7760 1057 7788 1255
rect 7746 1048 7802 1057
rect 7746 983 7802 992
rect 7944 785 7972 1255
rect 7930 776 7986 785
rect 7930 711 7986 720
rect 8220 480 8248 3606
rect 8312 3505 8340 4422
rect 8576 4072 8628 4078
rect 8574 4040 8576 4049
rect 8628 4040 8630 4049
rect 8574 3975 8630 3984
rect 8588 3534 8616 3975
rect 8484 3528 8536 3534
rect 8298 3496 8354 3505
rect 8484 3470 8536 3476
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8298 3431 8354 3440
rect 8312 2514 8340 3431
rect 8496 3369 8524 3470
rect 8482 3360 8538 3369
rect 8404 3318 8482 3346
rect 8404 3194 8432 3318
rect 8482 3295 8538 3304
rect 8680 3210 8708 6938
rect 8772 3738 8800 7754
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 8864 4185 8892 4422
rect 8850 4176 8906 4185
rect 8850 4111 8906 4120
rect 8956 4026 8984 8774
rect 9048 6798 9076 12328
rect 9416 12073 9444 12566
rect 9494 12472 9550 12481
rect 9494 12407 9550 12416
rect 9508 12374 9536 12407
rect 9496 12368 9548 12374
rect 9496 12310 9548 12316
rect 9402 12064 9458 12073
rect 9402 11999 9458 12008
rect 9416 10656 9444 11999
rect 9600 11370 9628 23015
rect 9784 22438 9812 23122
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9864 22432 9916 22438
rect 9864 22374 9916 22380
rect 9680 21956 9732 21962
rect 9680 21898 9732 21904
rect 9692 20058 9720 21898
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9692 19310 9720 19994
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9678 16688 9734 16697
rect 9678 16623 9734 16632
rect 9692 14618 9720 16623
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9692 13530 9720 14350
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9692 12345 9720 12378
rect 9678 12336 9734 12345
rect 9678 12271 9734 12280
rect 9232 10628 9444 10656
rect 9508 11342 9628 11370
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9140 9994 9168 10406
rect 9128 9988 9180 9994
rect 9128 9930 9180 9936
rect 9140 8362 9168 9930
rect 9128 8356 9180 8362
rect 9128 8298 9180 8304
rect 9140 8022 9168 8298
rect 9128 8016 9180 8022
rect 9128 7958 9180 7964
rect 9140 7478 9168 7958
rect 9232 7954 9260 10628
rect 9508 10538 9536 11342
rect 9588 11280 9640 11286
rect 9640 11228 9720 11234
rect 9588 11222 9720 11228
rect 9600 11206 9720 11222
rect 9692 10810 9720 11206
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9312 10532 9364 10538
rect 9312 10474 9364 10480
rect 9496 10532 9548 10538
rect 9496 10474 9548 10480
rect 9220 7948 9272 7954
rect 9220 7890 9272 7896
rect 9128 7472 9180 7478
rect 9128 7414 9180 7420
rect 9140 7002 9168 7414
rect 9324 7290 9352 10474
rect 9692 10062 9720 10542
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9692 9722 9720 9998
rect 9680 9716 9732 9722
rect 9508 9676 9680 9704
rect 9508 8430 9536 9676
rect 9680 9658 9732 9664
rect 9588 9580 9640 9586
rect 9640 9540 9720 9568
rect 9588 9522 9640 9528
rect 9588 9036 9640 9042
rect 9692 9024 9720 9540
rect 9784 9178 9812 22374
rect 9876 22273 9904 22374
rect 9862 22264 9918 22273
rect 9862 22199 9918 22208
rect 9864 20800 9916 20806
rect 9864 20742 9916 20748
rect 9876 20262 9904 20742
rect 9864 20256 9916 20262
rect 9864 20198 9916 20204
rect 9876 19854 9904 20198
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 9968 18902 9996 19450
rect 9956 18896 10008 18902
rect 9956 18838 10008 18844
rect 10048 18828 10100 18834
rect 10048 18770 10100 18776
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 9864 18624 9916 18630
rect 9864 18566 9916 18572
rect 9876 15586 9904 18566
rect 9968 17814 9996 18702
rect 10060 18222 10088 18770
rect 10152 18766 10180 23446
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10796 22114 10824 23598
rect 11426 23559 11482 23568
rect 11440 23526 11468 23559
rect 11428 23520 11480 23526
rect 11428 23462 11480 23468
rect 10787 22086 10824 22114
rect 10874 22128 10930 22137
rect 10787 22080 10815 22086
rect 10704 22052 10815 22080
rect 10874 22063 10876 22072
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10508 19848 10560 19854
rect 10508 19790 10560 19796
rect 10520 19514 10548 19790
rect 10508 19508 10560 19514
rect 10508 19450 10560 19456
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 10138 18592 10194 18601
rect 10138 18527 10194 18536
rect 10048 18216 10100 18222
rect 10048 18158 10100 18164
rect 9956 17808 10008 17814
rect 9954 17776 9956 17785
rect 10008 17776 10010 17785
rect 9954 17711 10010 17720
rect 10048 17128 10100 17134
rect 10046 17096 10048 17105
rect 10100 17096 10102 17105
rect 9956 17060 10008 17066
rect 10046 17031 10102 17040
rect 9956 17002 10008 17008
rect 9968 16794 9996 17002
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 10060 16250 10088 16730
rect 10152 16454 10180 18527
rect 10428 18426 10456 18702
rect 10416 18420 10468 18426
rect 10416 18362 10468 18368
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10322 17640 10378 17649
rect 10322 17575 10324 17584
rect 10376 17575 10378 17584
rect 10324 17546 10376 17552
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10704 16794 10732 22052
rect 10928 22063 10930 22072
rect 10876 22034 10928 22040
rect 10888 21690 10916 22034
rect 10968 22024 11020 22030
rect 10968 21966 11020 21972
rect 11060 22024 11112 22030
rect 11060 21966 11112 21972
rect 10876 21684 10928 21690
rect 10876 21626 10928 21632
rect 10980 21622 11008 21966
rect 11072 21894 11100 21966
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 11152 21888 11204 21894
rect 11152 21830 11204 21836
rect 10968 21616 11020 21622
rect 10966 21584 10968 21593
rect 11020 21584 11022 21593
rect 10966 21519 11022 21528
rect 10980 21493 11008 21519
rect 10968 21344 11020 21350
rect 10968 21286 11020 21292
rect 10876 20800 10928 20806
rect 10876 20742 10928 20748
rect 10888 19990 10916 20742
rect 10876 19984 10928 19990
rect 10876 19926 10928 19932
rect 10888 19378 10916 19926
rect 10876 19372 10928 19378
rect 10876 19314 10928 19320
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10796 17746 10824 19110
rect 10888 18970 10916 19314
rect 10980 19258 11008 21286
rect 11072 20602 11100 21830
rect 11164 21350 11192 21830
rect 11242 21720 11298 21729
rect 11242 21655 11298 21664
rect 11256 21486 11284 21655
rect 11428 21548 11480 21554
rect 11428 21490 11480 21496
rect 11244 21480 11296 21486
rect 11244 21422 11296 21428
rect 11152 21344 11204 21350
rect 11152 21286 11204 21292
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 11072 20058 11100 20538
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 11060 19304 11112 19310
rect 10980 19252 11060 19258
rect 10980 19246 11112 19252
rect 10980 19230 11100 19246
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 11072 18902 11100 19230
rect 11164 18970 11192 21286
rect 11440 21146 11468 21490
rect 11428 21140 11480 21146
rect 11428 21082 11480 21088
rect 11428 19372 11480 19378
rect 11428 19314 11480 19320
rect 11152 18964 11204 18970
rect 11152 18906 11204 18912
rect 11060 18896 11112 18902
rect 11060 18838 11112 18844
rect 11440 18834 11468 19314
rect 11428 18828 11480 18834
rect 11428 18770 11480 18776
rect 11060 18692 11112 18698
rect 11060 18634 11112 18640
rect 11072 18222 11100 18634
rect 11060 18216 11112 18222
rect 11060 18158 11112 18164
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 10784 17740 10836 17746
rect 10784 17682 10836 17688
rect 10796 17338 10824 17682
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 10888 17202 10916 18022
rect 10876 17196 10928 17202
rect 10876 17138 10928 17144
rect 10692 16788 10744 16794
rect 10744 16748 10916 16776
rect 10692 16730 10744 16736
rect 10232 16584 10284 16590
rect 10232 16526 10284 16532
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 10244 16130 10272 16526
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10060 16102 10272 16130
rect 9876 15558 9996 15586
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9876 14074 9904 15438
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9876 13802 9904 14010
rect 9864 13796 9916 13802
rect 9864 13738 9916 13744
rect 9968 13530 9996 15558
rect 10060 15473 10088 16102
rect 10140 15972 10192 15978
rect 10140 15914 10192 15920
rect 10152 15706 10180 15914
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10046 15464 10102 15473
rect 10046 15399 10048 15408
rect 10100 15399 10102 15408
rect 10048 15370 10100 15376
rect 10046 15328 10102 15337
rect 10046 15263 10102 15272
rect 10060 14074 10088 15263
rect 10152 15162 10180 15642
rect 10704 15484 10732 16390
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10796 15609 10824 15642
rect 10782 15600 10838 15609
rect 10782 15535 10838 15544
rect 10704 15456 10824 15484
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 10060 13870 10088 14010
rect 10152 13938 10180 15098
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10336 14074 10364 14418
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10048 13864 10100 13870
rect 10048 13806 10100 13812
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10704 13530 10732 13874
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 9968 12782 9996 13466
rect 10704 13326 10732 13466
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10704 12986 10732 13262
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10796 12866 10824 15456
rect 10704 12838 10824 12866
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10060 11898 10088 12242
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 10152 11354 10180 12378
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10336 11898 10364 12174
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 9968 10674 9996 10950
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9968 10470 9996 10610
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 10060 10282 10088 11222
rect 10322 11112 10378 11121
rect 10232 11076 10284 11082
rect 10322 11047 10378 11056
rect 10232 11018 10284 11024
rect 10244 10606 10272 11018
rect 10336 11014 10364 11047
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 10336 10606 10364 10950
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 9968 10254 10088 10282
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9692 8996 9812 9024
rect 9588 8978 9640 8984
rect 9600 8922 9628 8978
rect 9600 8894 9720 8922
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9586 7848 9642 7857
rect 9692 7818 9720 8894
rect 9784 8090 9812 8996
rect 9876 8537 9904 9862
rect 9862 8528 9918 8537
rect 9862 8463 9918 8472
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9586 7783 9642 7792
rect 9680 7812 9732 7818
rect 9494 7712 9550 7721
rect 9494 7647 9550 7656
rect 9232 7262 9352 7290
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 9036 6792 9088 6798
rect 9036 6734 9088 6740
rect 9048 6458 9076 6734
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 9128 6384 9180 6390
rect 9128 6326 9180 6332
rect 9140 5778 9168 6326
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9034 5672 9090 5681
rect 9034 5607 9036 5616
rect 9088 5607 9090 5616
rect 9036 5578 9088 5584
rect 9140 5370 9168 5714
rect 9128 5364 9180 5370
rect 9128 5306 9180 5312
rect 9140 5166 9168 5306
rect 9128 5160 9180 5166
rect 9128 5102 9180 5108
rect 9140 4826 9168 5102
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 8864 4010 8984 4026
rect 8852 4004 8984 4010
rect 8904 3998 8984 4004
rect 8852 3946 8904 3952
rect 8944 3936 8996 3942
rect 9232 3913 9260 7262
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 9416 6458 9444 6802
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9416 5574 9444 6394
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9508 5250 9536 7647
rect 9600 7274 9628 7783
rect 9680 7754 9732 7760
rect 9784 7410 9812 7890
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 9678 7168 9734 7177
rect 9678 7103 9734 7112
rect 9692 7002 9720 7103
rect 9784 7041 9812 7346
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9770 7032 9826 7041
rect 9680 6996 9732 7002
rect 9770 6967 9826 6976
rect 9680 6938 9732 6944
rect 9772 6656 9824 6662
rect 9692 6616 9772 6644
rect 9586 5536 9642 5545
rect 9586 5471 9642 5480
rect 9416 5222 9536 5250
rect 9310 4856 9366 4865
rect 9310 4791 9366 4800
rect 9324 4321 9352 4791
rect 9310 4312 9366 4321
rect 9310 4247 9366 4256
rect 9310 4040 9366 4049
rect 9310 3975 9366 3984
rect 9324 3942 9352 3975
rect 9312 3936 9364 3942
rect 8944 3878 8996 3884
rect 9218 3904 9274 3913
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8772 3641 8800 3674
rect 8758 3632 8814 3641
rect 8758 3567 8814 3576
rect 8392 3188 8444 3194
rect 8680 3182 8800 3210
rect 8392 3130 8444 3136
rect 8772 2666 8800 3182
rect 8772 2638 8892 2666
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8496 1737 8524 2450
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 8680 1737 8708 2382
rect 8482 1728 8538 1737
rect 8482 1663 8538 1672
rect 8666 1728 8722 1737
rect 8666 1663 8722 1672
rect 8864 480 8892 2638
rect 8956 1601 8984 3878
rect 9312 3878 9364 3884
rect 9218 3839 9274 3848
rect 8942 1592 8998 1601
rect 8942 1527 8998 1536
rect 9416 480 9444 5222
rect 9600 5166 9628 5471
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9508 3777 9536 3878
rect 9494 3768 9550 3777
rect 9494 3703 9496 3712
rect 9548 3703 9550 3712
rect 9496 3674 9548 3680
rect 9508 3643 9536 3674
rect 9692 2938 9720 6616
rect 9772 6598 9824 6604
rect 9876 6225 9904 7142
rect 9862 6216 9918 6225
rect 9772 6180 9824 6186
rect 9862 6151 9918 6160
rect 9772 6122 9824 6128
rect 9784 5914 9812 6122
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9876 5953 9904 6054
rect 9862 5944 9918 5953
rect 9772 5908 9824 5914
rect 9862 5879 9918 5888
rect 9772 5850 9824 5856
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 9876 4434 9904 5510
rect 9968 5409 9996 10254
rect 10230 9752 10286 9761
rect 10230 9687 10286 9696
rect 10244 9625 10272 9687
rect 10230 9616 10286 9625
rect 10230 9551 10286 9560
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 10138 9344 10194 9353
rect 10060 9217 10088 9318
rect 10138 9279 10194 9288
rect 10046 9208 10102 9217
rect 10152 9178 10180 9279
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10046 9143 10102 9152
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10046 9072 10102 9081
rect 10046 9007 10048 9016
rect 10100 9007 10102 9016
rect 10048 8978 10100 8984
rect 10152 8945 10180 9114
rect 10138 8936 10194 8945
rect 10138 8871 10194 8880
rect 10046 8528 10102 8537
rect 10046 8463 10102 8472
rect 10060 7324 10088 8463
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10152 7478 10180 7822
rect 10704 7562 10732 12838
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10796 12238 10824 12582
rect 10888 12306 10916 16748
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 10980 15162 11008 15438
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 11072 13954 11100 18158
rect 11520 18080 11572 18086
rect 11520 18022 11572 18028
rect 11428 17740 11480 17746
rect 11428 17682 11480 17688
rect 11152 17672 11204 17678
rect 11152 17614 11204 17620
rect 11164 17270 11192 17614
rect 11152 17264 11204 17270
rect 11152 17206 11204 17212
rect 11440 16998 11468 17682
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11336 15904 11388 15910
rect 11336 15846 11388 15852
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 11256 15162 11284 15642
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11348 14414 11376 15846
rect 11440 15609 11468 16934
rect 11532 15638 11560 18022
rect 11716 16794 11744 27520
rect 11796 24268 11848 24274
rect 12268 24256 12296 27520
rect 12348 24744 12400 24750
rect 12348 24686 12400 24692
rect 11796 24210 11848 24216
rect 11992 24228 12296 24256
rect 11808 23526 11836 24210
rect 11796 23520 11848 23526
rect 11796 23462 11848 23468
rect 11808 18873 11836 23462
rect 11888 20256 11940 20262
rect 11888 20198 11940 20204
rect 11900 20058 11928 20198
rect 11888 20052 11940 20058
rect 11888 19994 11940 20000
rect 11794 18864 11850 18873
rect 11794 18799 11850 18808
rect 11808 17354 11836 18799
rect 11992 18601 12020 24228
rect 12254 24168 12310 24177
rect 12254 24103 12256 24112
rect 12308 24103 12310 24112
rect 12256 24074 12308 24080
rect 12254 24032 12310 24041
rect 12254 23967 12310 23976
rect 12164 23180 12216 23186
rect 12164 23122 12216 23128
rect 12176 22574 12204 23122
rect 12164 22568 12216 22574
rect 12162 22536 12164 22545
rect 12216 22536 12218 22545
rect 12162 22471 12218 22480
rect 12164 21344 12216 21350
rect 12164 21286 12216 21292
rect 12176 19310 12204 21286
rect 12268 19961 12296 23967
rect 12360 21865 12388 24686
rect 12622 23896 12678 23905
rect 12622 23831 12624 23840
rect 12676 23831 12678 23840
rect 12624 23802 12676 23808
rect 12346 21856 12402 21865
rect 12346 21791 12402 21800
rect 12820 21593 12848 27520
rect 13372 23866 13400 27520
rect 13636 24268 13688 24274
rect 13636 24210 13688 24216
rect 13360 23860 13412 23866
rect 13360 23802 13412 23808
rect 13648 23526 13676 24210
rect 13636 23520 13688 23526
rect 13636 23462 13688 23468
rect 13648 23322 13676 23462
rect 13636 23316 13688 23322
rect 13636 23258 13688 23264
rect 13544 23112 13596 23118
rect 13544 23054 13596 23060
rect 12900 22704 12952 22710
rect 12898 22672 12900 22681
rect 12952 22672 12954 22681
rect 12898 22607 12954 22616
rect 12900 22568 12952 22574
rect 12900 22510 12952 22516
rect 12912 22137 12940 22510
rect 13556 22137 13584 23054
rect 13924 22386 13952 27520
rect 14568 27418 14596 27520
rect 14568 27390 14688 27418
rect 14278 24440 14334 24449
rect 14278 24375 14280 24384
rect 14332 24375 14334 24384
rect 14280 24346 14332 24352
rect 14004 23792 14056 23798
rect 14002 23760 14004 23769
rect 14056 23760 14058 23769
rect 14002 23695 14058 23704
rect 14556 23520 14608 23526
rect 14556 23462 14608 23468
rect 14464 22976 14516 22982
rect 14464 22918 14516 22924
rect 14476 22642 14504 22918
rect 14464 22636 14516 22642
rect 14464 22578 14516 22584
rect 14278 22536 14334 22545
rect 14278 22471 14334 22480
rect 13740 22358 13952 22386
rect 14004 22432 14056 22438
rect 14004 22374 14056 22380
rect 12898 22128 12954 22137
rect 13542 22128 13598 22137
rect 12898 22063 12954 22072
rect 13268 22092 13320 22098
rect 12806 21584 12862 21593
rect 12806 21519 12862 21528
rect 12820 20913 12848 21519
rect 12806 20904 12862 20913
rect 12806 20839 12862 20848
rect 12348 20800 12400 20806
rect 12348 20742 12400 20748
rect 12360 20505 12388 20742
rect 12346 20496 12402 20505
rect 12346 20431 12402 20440
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12544 19990 12572 20334
rect 12716 20256 12768 20262
rect 12716 20198 12768 20204
rect 12532 19984 12584 19990
rect 12254 19952 12310 19961
rect 12532 19926 12584 19932
rect 12254 19887 12310 19896
rect 12544 19786 12572 19926
rect 12622 19816 12678 19825
rect 12532 19780 12584 19786
rect 12622 19751 12678 19760
rect 12532 19722 12584 19728
rect 12636 19514 12664 19751
rect 12624 19508 12676 19514
rect 12624 19450 12676 19456
rect 12728 19446 12756 20198
rect 12716 19440 12768 19446
rect 12716 19382 12768 19388
rect 12164 19304 12216 19310
rect 12164 19246 12216 19252
rect 12254 19272 12310 19281
rect 12728 19242 12756 19382
rect 12254 19207 12310 19216
rect 12716 19236 12768 19242
rect 11978 18592 12034 18601
rect 11978 18527 12034 18536
rect 12268 18154 12296 19207
rect 12716 19178 12768 19184
rect 12728 18766 12756 19178
rect 12808 18828 12860 18834
rect 12808 18770 12860 18776
rect 12716 18760 12768 18766
rect 12716 18702 12768 18708
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12544 18222 12572 18566
rect 12728 18358 12756 18702
rect 12716 18352 12768 18358
rect 12716 18294 12768 18300
rect 12532 18216 12584 18222
rect 12360 18164 12532 18170
rect 12360 18158 12584 18164
rect 12256 18148 12308 18154
rect 12256 18090 12308 18096
rect 12360 18142 12572 18158
rect 11808 17326 12204 17354
rect 11796 17264 11848 17270
rect 11796 17206 11848 17212
rect 11704 16788 11756 16794
rect 11704 16730 11756 16736
rect 11808 16658 11836 17206
rect 12176 16708 12204 17326
rect 12360 17202 12388 18142
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12348 17196 12400 17202
rect 12348 17138 12400 17144
rect 12544 16726 12572 17478
rect 12728 17270 12756 18294
rect 12820 17338 12848 18770
rect 12912 18306 12940 22063
rect 13542 22063 13598 22072
rect 13268 22034 13320 22040
rect 13280 21894 13308 22034
rect 13636 22024 13688 22030
rect 13634 21992 13636 22001
rect 13688 21992 13690 22001
rect 13740 21962 13768 22358
rect 14016 22234 14044 22374
rect 14292 22273 14320 22471
rect 14278 22264 14334 22273
rect 13820 22228 13872 22234
rect 13820 22170 13872 22176
rect 14004 22228 14056 22234
rect 14278 22199 14334 22208
rect 14372 22228 14424 22234
rect 14004 22170 14056 22176
rect 14372 22170 14424 22176
rect 13634 21927 13690 21936
rect 13728 21956 13780 21962
rect 13268 21888 13320 21894
rect 13268 21830 13320 21836
rect 13360 21888 13412 21894
rect 13360 21830 13412 21836
rect 12992 21548 13044 21554
rect 12992 21490 13044 21496
rect 13004 21146 13032 21490
rect 13082 21448 13138 21457
rect 13082 21383 13084 21392
rect 13136 21383 13138 21392
rect 13084 21354 13136 21360
rect 13280 21146 13308 21830
rect 12992 21140 13044 21146
rect 12992 21082 13044 21088
rect 13268 21140 13320 21146
rect 13268 21082 13320 21088
rect 13004 20398 13032 21082
rect 13372 21010 13400 21830
rect 13648 21690 13676 21927
rect 13728 21898 13780 21904
rect 13636 21684 13688 21690
rect 13636 21626 13688 21632
rect 13648 21350 13676 21381
rect 13636 21344 13688 21350
rect 13740 21298 13768 21898
rect 13688 21292 13768 21298
rect 13636 21286 13768 21292
rect 13648 21270 13768 21286
rect 13360 21004 13412 21010
rect 13360 20946 13412 20952
rect 13450 20904 13506 20913
rect 13450 20839 13506 20848
rect 12992 20392 13044 20398
rect 12992 20334 13044 20340
rect 12992 20052 13044 20058
rect 12992 19994 13044 20000
rect 13004 19310 13032 19994
rect 12992 19304 13044 19310
rect 12992 19246 13044 19252
rect 13084 19168 13136 19174
rect 13084 19110 13136 19116
rect 13096 18902 13124 19110
rect 13084 18896 13136 18902
rect 13084 18838 13136 18844
rect 13096 18426 13124 18838
rect 13084 18420 13136 18426
rect 13084 18362 13136 18368
rect 13464 18306 13492 20839
rect 13648 20754 13676 21270
rect 13832 21162 13860 22170
rect 14002 22128 14058 22137
rect 14002 22063 14058 22072
rect 13740 21134 13860 21162
rect 13740 21078 13768 21134
rect 14016 21078 14044 22063
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 14108 21350 14136 21966
rect 14096 21344 14148 21350
rect 14096 21286 14148 21292
rect 13728 21072 13780 21078
rect 13728 21014 13780 21020
rect 14004 21072 14056 21078
rect 14004 21014 14056 21020
rect 14004 20936 14056 20942
rect 14004 20878 14056 20884
rect 14016 20777 14044 20878
rect 14002 20768 14058 20777
rect 13648 20726 13952 20754
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 13556 18834 13584 20198
rect 13820 19848 13872 19854
rect 13820 19790 13872 19796
rect 13832 19174 13860 19790
rect 13820 19168 13872 19174
rect 13924 19145 13952 20726
rect 14002 20703 14058 20712
rect 14016 20602 14044 20703
rect 14004 20596 14056 20602
rect 14004 20538 14056 20544
rect 14108 19310 14136 21286
rect 14186 19816 14242 19825
rect 14186 19751 14242 19760
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 13820 19110 13872 19116
rect 13910 19136 13966 19145
rect 13544 18828 13596 18834
rect 13544 18770 13596 18776
rect 13832 18329 13860 19110
rect 13910 19071 13966 19080
rect 13818 18320 13874 18329
rect 12912 18278 13032 18306
rect 13464 18278 13676 18306
rect 12808 17332 12860 17338
rect 12808 17274 12860 17280
rect 12716 17264 12768 17270
rect 12716 17206 12768 17212
rect 12084 16680 12204 16708
rect 12532 16720 12584 16726
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 11808 16250 11836 16594
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 11796 15972 11848 15978
rect 11796 15914 11848 15920
rect 11520 15632 11572 15638
rect 11426 15600 11482 15609
rect 11520 15574 11572 15580
rect 11426 15535 11482 15544
rect 11440 15502 11468 15535
rect 11428 15496 11480 15502
rect 11428 15438 11480 15444
rect 11532 15162 11560 15574
rect 11520 15156 11572 15162
rect 11520 15098 11572 15104
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11348 14074 11376 14350
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11072 13926 11376 13954
rect 11152 13796 11204 13802
rect 11152 13738 11204 13744
rect 11060 13456 11112 13462
rect 11058 13424 11060 13433
rect 11112 13424 11114 13433
rect 11058 13359 11114 13368
rect 11164 13326 11192 13738
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10796 11762 10824 12038
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10888 9761 10916 12242
rect 11164 11914 11192 13262
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 10980 11898 11192 11914
rect 10968 11892 11192 11898
rect 11020 11886 11192 11892
rect 10968 11834 11020 11840
rect 11256 11694 11284 12038
rect 11244 11688 11296 11694
rect 11150 11656 11206 11665
rect 11244 11630 11296 11636
rect 11150 11591 11152 11600
rect 11204 11591 11206 11600
rect 11152 11562 11204 11568
rect 11348 11286 11376 13926
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11440 12889 11468 13126
rect 11426 12880 11482 12889
rect 11426 12815 11482 12824
rect 11428 11688 11480 11694
rect 11428 11630 11480 11636
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 10980 10266 11008 11154
rect 11440 11014 11468 11630
rect 11428 11008 11480 11014
rect 11428 10950 11480 10956
rect 11440 10810 11468 10950
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11060 10736 11112 10742
rect 11060 10678 11112 10684
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10874 9752 10930 9761
rect 10874 9687 10930 9696
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10796 9178 10824 9318
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10888 8838 10916 9318
rect 10980 8974 11008 10202
rect 11072 9110 11100 10678
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 11060 9104 11112 9110
rect 11060 9046 11112 9052
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10888 8498 10916 8774
rect 10980 8634 11008 8910
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 11164 8378 11192 9862
rect 11336 9580 11388 9586
rect 11336 9522 11388 9528
rect 11348 9042 11376 9522
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 10980 8350 11192 8378
rect 10980 7818 11008 8350
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11164 7886 11192 8230
rect 11348 8090 11376 8978
rect 11440 8974 11468 10746
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 11440 8634 11468 8910
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 10968 7812 11020 7818
rect 10968 7754 11020 7760
rect 10704 7534 10824 7562
rect 11164 7546 11192 7822
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 10140 7472 10192 7478
rect 10140 7414 10192 7420
rect 10690 7440 10746 7449
rect 10690 7375 10746 7384
rect 10060 7296 10180 7324
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10060 6225 10088 6734
rect 10046 6216 10102 6225
rect 10046 6151 10102 6160
rect 9954 5400 10010 5409
rect 9954 5335 10010 5344
rect 9956 5092 10008 5098
rect 9956 5034 10008 5040
rect 9968 4690 9996 5034
rect 10046 4720 10102 4729
rect 9956 4684 10008 4690
rect 10046 4655 10048 4664
rect 9956 4626 10008 4632
rect 10100 4655 10102 4664
rect 10048 4626 10100 4632
rect 9968 4593 9996 4626
rect 10152 4622 10180 7296
rect 10704 7177 10732 7375
rect 10690 7168 10746 7177
rect 10289 7100 10585 7120
rect 10690 7103 10746 7112
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10796 7002 10824 7534
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 10966 7440 11022 7449
rect 10966 7375 10968 7384
rect 11020 7375 11022 7384
rect 10968 7346 11020 7352
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 10784 6996 10836 7002
rect 10784 6938 10836 6944
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10244 6458 10272 6734
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10244 6361 10272 6394
rect 10230 6352 10286 6361
rect 10230 6287 10286 6296
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10704 5030 10732 5714
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10704 4758 10732 4966
rect 10508 4752 10560 4758
rect 10506 4720 10508 4729
rect 10692 4752 10744 4758
rect 10560 4720 10562 4729
rect 10692 4694 10744 4700
rect 10506 4655 10562 4664
rect 10140 4616 10192 4622
rect 9954 4584 10010 4593
rect 10140 4558 10192 4564
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 9954 4519 10010 4528
rect 9876 4406 10180 4434
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 9772 4140 9824 4146
rect 9824 4100 9904 4128
rect 9772 4082 9824 4088
rect 9770 3632 9826 3641
rect 9770 3567 9826 3576
rect 9508 2910 9720 2938
rect 9508 2514 9536 2910
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9600 2650 9628 2790
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9600 2446 9628 2586
rect 9784 2582 9812 3567
rect 9876 3194 9904 4100
rect 9968 3602 9996 4218
rect 10046 4040 10102 4049
rect 10046 3975 10102 3984
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9968 2922 9996 3538
rect 9956 2916 10008 2922
rect 9956 2858 10008 2864
rect 9954 2816 10010 2825
rect 9954 2751 10010 2760
rect 9772 2576 9824 2582
rect 9772 2518 9824 2524
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 9968 480 9996 2751
rect 10060 2650 10088 3975
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 10152 2145 10180 4406
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10704 2632 10732 4558
rect 10796 3738 10824 6734
rect 10888 6662 10916 7278
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 11072 6882 11100 7210
rect 10980 6854 11100 6882
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10980 6089 11008 6854
rect 11256 6746 11284 7686
rect 11348 7410 11376 8026
rect 11428 7744 11480 7750
rect 11428 7686 11480 7692
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11072 6718 11284 6746
rect 10966 6080 11022 6089
rect 10966 6015 11022 6024
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 10796 2650 10824 3130
rect 10520 2604 10732 2632
rect 10784 2644 10836 2650
rect 10138 2136 10194 2145
rect 10138 2071 10194 2080
rect 10520 480 10548 2604
rect 10784 2586 10836 2592
rect 10796 2446 10824 2586
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 10888 2378 10916 5646
rect 10980 4826 11008 6015
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 10980 3720 11008 4422
rect 11072 4049 11100 6718
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11256 5681 11284 6598
rect 11242 5672 11298 5681
rect 11242 5607 11298 5616
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 11164 4214 11192 4966
rect 11348 4826 11376 7142
rect 11440 6798 11468 7686
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11152 4208 11204 4214
rect 11152 4150 11204 4156
rect 11058 4040 11114 4049
rect 11058 3975 11114 3984
rect 11060 3732 11112 3738
rect 10980 3692 11060 3720
rect 11060 3674 11112 3680
rect 11072 2990 11100 3674
rect 11164 3670 11192 4150
rect 11348 4078 11376 4762
rect 11336 4072 11388 4078
rect 11242 4040 11298 4049
rect 11336 4014 11388 4020
rect 11242 3975 11244 3984
rect 11296 3975 11298 3984
rect 11244 3946 11296 3952
rect 11242 3904 11298 3913
rect 11242 3839 11298 3848
rect 11152 3664 11204 3670
rect 11152 3606 11204 3612
rect 11256 3097 11284 3839
rect 11336 3664 11388 3670
rect 11336 3606 11388 3612
rect 11348 3534 11376 3606
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11348 3194 11376 3470
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 11242 3088 11298 3097
rect 11242 3023 11298 3032
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 11428 2848 11480 2854
rect 11426 2816 11428 2825
rect 11480 2816 11482 2825
rect 11426 2751 11482 2760
rect 10876 2372 10928 2378
rect 10876 2314 10928 2320
rect 11532 1442 11560 13330
rect 11702 12336 11758 12345
rect 11612 12300 11664 12306
rect 11702 12271 11704 12280
rect 11612 12242 11664 12248
rect 11756 12271 11758 12280
rect 11704 12242 11756 12248
rect 11624 12073 11652 12242
rect 11610 12064 11666 12073
rect 11610 11999 11666 12008
rect 11624 11898 11652 11999
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11716 11830 11744 12242
rect 11704 11824 11756 11830
rect 11704 11766 11756 11772
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 11624 10266 11652 10406
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11808 9994 11836 15914
rect 11992 15910 12020 16594
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 12084 13138 12112 16680
rect 12532 16662 12584 16668
rect 12806 15736 12862 15745
rect 12440 15700 12492 15706
rect 12806 15671 12808 15680
rect 12440 15642 12492 15648
rect 12860 15671 12862 15680
rect 12808 15642 12860 15648
rect 12452 15314 12480 15642
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12360 15286 12480 15314
rect 12360 15162 12388 15286
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 12728 14890 12756 15506
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12716 14884 12768 14890
rect 12716 14826 12768 14832
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 12164 14272 12216 14278
rect 12164 14214 12216 14220
rect 12176 13462 12204 14214
rect 12268 14074 12296 14418
rect 12716 14408 12768 14414
rect 12820 14396 12848 14894
rect 12768 14368 12848 14396
rect 12716 14350 12768 14356
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12164 13456 12216 13462
rect 12164 13398 12216 13404
rect 12176 13258 12204 13398
rect 12164 13252 12216 13258
rect 12164 13194 12216 13200
rect 12084 13110 12204 13138
rect 11886 13016 11942 13025
rect 11886 12951 11942 12960
rect 11900 12617 11928 12951
rect 11886 12608 11942 12617
rect 11886 12543 11942 12552
rect 11900 12238 11928 12543
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11794 9752 11850 9761
rect 11794 9687 11850 9696
rect 11612 9444 11664 9450
rect 11612 9386 11664 9392
rect 11624 7018 11652 9386
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11716 8090 11744 9318
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11624 6990 11744 7018
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11624 5710 11652 6802
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11716 4690 11744 6990
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11624 4282 11652 4558
rect 11716 4282 11744 4626
rect 11612 4276 11664 4282
rect 11612 4218 11664 4224
rect 11704 4276 11756 4282
rect 11704 4218 11756 4224
rect 11704 3596 11756 3602
rect 11704 3538 11756 3544
rect 11716 3194 11744 3538
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11808 2496 11836 9687
rect 11992 9489 12020 9862
rect 11978 9480 12034 9489
rect 11978 9415 12034 9424
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11900 8634 11928 8978
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11900 8537 11928 8570
rect 11886 8528 11942 8537
rect 11886 8463 11942 8472
rect 12084 8090 12112 9114
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12176 7970 12204 13110
rect 12452 12850 12480 14282
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12544 13802 12572 14214
rect 12728 14074 12756 14350
rect 12716 14068 12768 14074
rect 12636 14028 12716 14056
rect 12532 13796 12584 13802
rect 12532 13738 12584 13744
rect 12544 12986 12572 13738
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12452 11354 12480 12786
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12544 10962 12572 11834
rect 12636 11694 12664 14028
rect 12716 14010 12768 14016
rect 12714 13832 12770 13841
rect 12714 13767 12770 13776
rect 12728 11778 12756 13767
rect 12808 13456 12860 13462
rect 12808 13398 12860 13404
rect 12820 13297 12848 13398
rect 12806 13288 12862 13297
rect 12806 13223 12862 13232
rect 12820 11898 12848 13223
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 12912 12782 12940 13126
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 12912 12442 12940 12718
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12728 11750 12940 11778
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12716 11620 12768 11626
rect 12716 11562 12768 11568
rect 12728 11082 12756 11562
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12544 10934 12664 10962
rect 12636 10606 12664 10934
rect 12806 10840 12862 10849
rect 12806 10775 12862 10784
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12636 10266 12664 10542
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12452 9466 12480 10066
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12636 9722 12664 9998
rect 12728 9722 12756 10406
rect 12820 9761 12848 10775
rect 12806 9752 12862 9761
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12716 9716 12768 9722
rect 12806 9687 12862 9696
rect 12716 9658 12768 9664
rect 12360 9438 12480 9466
rect 12360 9382 12388 9438
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12438 8256 12494 8265
rect 12438 8191 12494 8200
rect 12176 7942 12388 7970
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 12268 7546 12296 7822
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12360 7478 12388 7942
rect 12348 7472 12400 7478
rect 12268 7420 12348 7426
rect 12268 7414 12400 7420
rect 12268 7398 12388 7414
rect 12452 7410 12480 8191
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 11900 6458 11928 6734
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11900 4826 11928 6394
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12072 5772 12124 5778
rect 12072 5714 12124 5720
rect 12084 5302 12112 5714
rect 12072 5296 12124 5302
rect 12072 5238 12124 5244
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 12176 4146 12204 6054
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 11992 2650 12020 3878
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 11716 2468 11836 2496
rect 11978 2544 12034 2553
rect 11978 2479 12034 2488
rect 12162 2544 12218 2553
rect 12162 2479 12218 2488
rect 11610 2408 11666 2417
rect 11610 2343 11612 2352
rect 11664 2343 11666 2352
rect 11612 2314 11664 2320
rect 11072 1414 11560 1442
rect 11072 480 11100 1414
rect 11716 480 11744 2468
rect 11992 2446 12020 2479
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 12176 1737 12204 2479
rect 12162 1728 12218 1737
rect 12162 1663 12218 1672
rect 12268 480 12296 7398
rect 12360 7349 12388 7398
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12820 6848 12848 9687
rect 12728 6820 12848 6848
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12544 6322 12572 6598
rect 12532 6316 12584 6322
rect 12584 6276 12664 6304
rect 12532 6258 12584 6264
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12348 5840 12400 5846
rect 12348 5782 12400 5788
rect 12360 5166 12388 5782
rect 12348 5160 12400 5166
rect 12348 5102 12400 5108
rect 12452 4826 12480 6054
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12544 4282 12572 5102
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12636 3738 12664 6276
rect 12728 5114 12756 6820
rect 12806 6760 12862 6769
rect 12806 6695 12808 6704
rect 12860 6695 12862 6704
rect 12808 6666 12860 6672
rect 12912 6474 12940 11750
rect 13004 10849 13032 18278
rect 13176 17536 13228 17542
rect 13176 17478 13228 17484
rect 13188 17066 13216 17478
rect 13358 17232 13414 17241
rect 13358 17167 13414 17176
rect 13176 17060 13228 17066
rect 13176 17002 13228 17008
rect 13188 16946 13216 17002
rect 13096 16918 13216 16946
rect 13096 16794 13124 16918
rect 13084 16788 13136 16794
rect 13084 16730 13136 16736
rect 13096 16697 13124 16730
rect 13082 16688 13138 16697
rect 13082 16623 13138 16632
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 13096 15162 13124 15438
rect 13084 15156 13136 15162
rect 13084 15098 13136 15104
rect 13268 14884 13320 14890
rect 13268 14826 13320 14832
rect 13084 12368 13136 12374
rect 13084 12310 13136 12316
rect 13096 11694 13124 12310
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 13280 11540 13308 14826
rect 13372 12481 13400 17167
rect 13452 14884 13504 14890
rect 13452 14826 13504 14832
rect 13464 13326 13492 14826
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13556 13326 13584 14418
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13464 12850 13492 13262
rect 13556 12986 13584 13262
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 13556 12730 13584 12922
rect 13464 12702 13584 12730
rect 13358 12472 13414 12481
rect 13358 12407 13414 12416
rect 13464 12238 13492 12702
rect 13648 12594 13676 18278
rect 13728 18284 13780 18290
rect 14200 18306 14228 19751
rect 14200 18278 14320 18306
rect 13818 18255 13874 18264
rect 13728 18226 13780 18232
rect 13740 17354 13768 18226
rect 14188 18148 14240 18154
rect 14188 18090 14240 18096
rect 14004 18080 14056 18086
rect 14004 18022 14056 18028
rect 13740 17338 13952 17354
rect 13740 17332 13964 17338
rect 13740 17326 13912 17332
rect 13912 17274 13964 17280
rect 13924 15978 13952 17274
rect 13912 15972 13964 15978
rect 13912 15914 13964 15920
rect 13924 15706 13952 15914
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 13832 14074 13860 15506
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 13924 14074 13952 14350
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13912 14068 13964 14074
rect 13912 14010 13964 14016
rect 13924 13954 13952 14010
rect 13832 13926 13952 13954
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13740 13530 13768 13670
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13740 12753 13768 13330
rect 13726 12744 13782 12753
rect 13726 12679 13782 12688
rect 13832 12594 13860 13926
rect 14016 13818 14044 18022
rect 14200 17542 14228 18090
rect 14188 17536 14240 17542
rect 14188 17478 14240 17484
rect 14096 14884 14148 14890
rect 14096 14826 14148 14832
rect 14108 14618 14136 14826
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 14094 14512 14150 14521
rect 14094 14447 14150 14456
rect 13556 12566 13676 12594
rect 13740 12566 13860 12594
rect 13924 13790 14044 13818
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13452 11552 13504 11558
rect 13280 11512 13400 11540
rect 13266 11384 13322 11393
rect 13266 11319 13268 11328
rect 13320 11319 13322 11328
rect 13268 11290 13320 11296
rect 13084 11008 13136 11014
rect 13084 10950 13136 10956
rect 12990 10840 13046 10849
rect 12990 10775 13046 10784
rect 12990 10704 13046 10713
rect 13096 10674 13124 10950
rect 13174 10704 13230 10713
rect 12990 10639 13046 10648
rect 13084 10668 13136 10674
rect 13004 10305 13032 10639
rect 13174 10639 13230 10648
rect 13084 10610 13136 10616
rect 12990 10296 13046 10305
rect 12990 10231 13046 10240
rect 13096 8922 13124 10610
rect 13188 10606 13216 10639
rect 13176 10600 13228 10606
rect 13176 10542 13228 10548
rect 13268 10056 13320 10062
rect 13004 8894 13124 8922
rect 13188 10016 13268 10044
rect 13004 8537 13032 8894
rect 13084 8832 13136 8838
rect 13084 8774 13136 8780
rect 12990 8528 13046 8537
rect 12990 8463 13046 8472
rect 13096 8362 13124 8774
rect 13084 8356 13136 8362
rect 13084 8298 13136 8304
rect 13096 7886 13124 8298
rect 13188 8090 13216 10016
rect 13268 9998 13320 10004
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 13280 7954 13308 9658
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 13174 7712 13230 7721
rect 13174 7647 13230 7656
rect 13188 7410 13216 7647
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 12912 6446 13124 6474
rect 12990 6352 13046 6361
rect 12990 6287 13046 6296
rect 12900 6112 12952 6118
rect 12898 6080 12900 6089
rect 12952 6080 12954 6089
rect 12898 6015 12954 6024
rect 13004 5778 13032 6287
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 13004 5370 13032 5714
rect 12992 5364 13044 5370
rect 12992 5306 13044 5312
rect 12728 5086 12940 5114
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12808 5024 12860 5030
rect 12808 4966 12860 4972
rect 12728 4690 12756 4966
rect 12716 4684 12768 4690
rect 12716 4626 12768 4632
rect 12820 4146 12848 4966
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 12912 4026 12940 5086
rect 13096 5030 13124 6446
rect 13280 5574 13308 6734
rect 13268 5568 13320 5574
rect 13268 5510 13320 5516
rect 13084 5024 13136 5030
rect 13084 4966 13136 4972
rect 13174 4856 13230 4865
rect 13174 4791 13230 4800
rect 12992 4752 13044 4758
rect 12992 4694 13044 4700
rect 13004 4457 13032 4694
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 12990 4448 13046 4457
rect 12990 4383 13046 4392
rect 12820 3998 12940 4026
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12820 480 12848 3998
rect 13096 3738 13124 4558
rect 13188 4185 13216 4791
rect 13268 4480 13320 4486
rect 13268 4422 13320 4428
rect 13174 4176 13230 4185
rect 13280 4146 13308 4422
rect 13174 4111 13230 4120
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 13096 2922 13124 3674
rect 13084 2916 13136 2922
rect 13084 2858 13136 2864
rect 13280 2446 13308 4082
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 13372 480 13400 11512
rect 13452 11494 13504 11500
rect 13464 11150 13492 11494
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13464 10810 13492 11086
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13464 9450 13492 9998
rect 13452 9444 13504 9450
rect 13452 9386 13504 9392
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13464 6118 13492 6734
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13464 5914 13492 6054
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 13450 5808 13506 5817
rect 13450 5743 13506 5752
rect 13464 5574 13492 5743
rect 13452 5568 13504 5574
rect 13452 5510 13504 5516
rect 13556 4162 13584 12566
rect 13634 12472 13690 12481
rect 13634 12407 13690 12416
rect 13648 9994 13676 12407
rect 13740 12374 13768 12566
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13740 11354 13768 12106
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13832 11558 13860 12038
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13924 11370 13952 13790
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 14016 12986 14044 13466
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14108 12866 14136 14447
rect 14016 12838 14136 12866
rect 14016 11506 14044 12838
rect 14096 12640 14148 12646
rect 14096 12582 14148 12588
rect 14108 12306 14136 12582
rect 14096 12300 14148 12306
rect 14096 12242 14148 12248
rect 14108 11898 14136 12242
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14200 11812 14228 17478
rect 14292 15065 14320 18278
rect 14278 15056 14334 15065
rect 14278 14991 14334 15000
rect 14292 14521 14320 14991
rect 14278 14512 14334 14521
rect 14278 14447 14334 14456
rect 14384 11914 14412 22170
rect 14476 22098 14504 22578
rect 14568 22506 14596 23462
rect 14556 22500 14608 22506
rect 14556 22442 14608 22448
rect 14464 22092 14516 22098
rect 14464 22034 14516 22040
rect 14476 20942 14504 22034
rect 14556 21888 14608 21894
rect 14556 21830 14608 21836
rect 14568 21418 14596 21830
rect 14556 21412 14608 21418
rect 14556 21354 14608 21360
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14464 19780 14516 19786
rect 14464 19722 14516 19728
rect 14476 19310 14504 19722
rect 14568 19514 14596 21354
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14554 19408 14610 19417
rect 14554 19343 14610 19352
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 14476 18970 14504 19246
rect 14464 18964 14516 18970
rect 14464 18906 14516 18912
rect 14476 18290 14504 18906
rect 14464 18284 14516 18290
rect 14464 18226 14516 18232
rect 14476 17882 14504 18226
rect 14464 17876 14516 17882
rect 14464 17818 14516 17824
rect 14568 15706 14596 19343
rect 14660 18154 14688 27390
rect 15120 25242 15148 27520
rect 14844 25214 15148 25242
rect 14844 23322 14872 25214
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15476 24404 15528 24410
rect 15476 24346 15528 24352
rect 15488 24313 15516 24346
rect 15474 24304 15530 24313
rect 15292 24268 15344 24274
rect 15474 24239 15530 24248
rect 15292 24210 15344 24216
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15108 23792 15160 23798
rect 15106 23760 15108 23769
rect 15160 23760 15162 23769
rect 15106 23695 15162 23704
rect 15304 23526 15332 24210
rect 15672 23866 15700 27520
rect 16118 24848 16174 24857
rect 16118 24783 16174 24792
rect 16132 24614 16160 24783
rect 16120 24608 16172 24614
rect 16120 24550 16172 24556
rect 16224 24449 16252 27520
rect 16776 24721 16804 27520
rect 16762 24712 16818 24721
rect 16762 24647 16818 24656
rect 17420 24449 17448 27520
rect 17972 24857 18000 27520
rect 17958 24848 18014 24857
rect 17958 24783 18014 24792
rect 18142 24848 18198 24857
rect 18142 24783 18198 24792
rect 16210 24440 16266 24449
rect 16210 24375 16266 24384
rect 16394 24440 16450 24449
rect 16394 24375 16450 24384
rect 17406 24440 17462 24449
rect 17406 24375 17462 24384
rect 17774 24440 17830 24449
rect 17774 24375 17830 24384
rect 15660 23860 15712 23866
rect 15660 23802 15712 23808
rect 15292 23520 15344 23526
rect 15292 23462 15344 23468
rect 14832 23316 14884 23322
rect 14832 23258 14884 23264
rect 14844 22658 14872 23258
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14752 22630 14872 22658
rect 14752 22438 14780 22630
rect 14832 22500 14884 22506
rect 14832 22442 14884 22448
rect 14740 22432 14792 22438
rect 14740 22374 14792 22380
rect 14752 22234 14780 22374
rect 14740 22228 14792 22234
rect 14740 22170 14792 22176
rect 14844 22114 14872 22442
rect 14752 22086 14872 22114
rect 14752 22012 14780 22086
rect 14752 21984 14872 22012
rect 14740 21004 14792 21010
rect 14740 20946 14792 20952
rect 14752 20602 14780 20946
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14740 19984 14792 19990
rect 14740 19926 14792 19932
rect 14648 18148 14700 18154
rect 14648 18090 14700 18096
rect 14752 18086 14780 19926
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14464 15360 14516 15366
rect 14464 15302 14516 15308
rect 14476 12442 14504 15302
rect 14738 13968 14794 13977
rect 14738 13903 14794 13912
rect 14556 13388 14608 13394
rect 14556 13330 14608 13336
rect 14568 13161 14596 13330
rect 14752 13326 14780 13903
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 14554 13152 14610 13161
rect 14554 13087 14610 13096
rect 14568 12986 14596 13087
rect 14752 12986 14780 13262
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 14740 12980 14792 12986
rect 14740 12922 14792 12928
rect 14646 12880 14702 12889
rect 14646 12815 14702 12824
rect 14464 12436 14516 12442
rect 14464 12378 14516 12384
rect 14384 11886 14596 11914
rect 14660 11898 14688 12815
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14752 11937 14780 12038
rect 14738 11928 14794 11937
rect 14200 11784 14504 11812
rect 14278 11656 14334 11665
rect 14278 11591 14334 11600
rect 14016 11478 14136 11506
rect 13728 11348 13780 11354
rect 13924 11342 14044 11370
rect 13728 11290 13780 11296
rect 13912 11280 13964 11286
rect 13910 11248 13912 11257
rect 13964 11248 13966 11257
rect 13910 11183 13966 11192
rect 13820 10600 13872 10606
rect 13818 10568 13820 10577
rect 13872 10568 13874 10577
rect 13818 10503 13874 10512
rect 13912 10464 13964 10470
rect 13818 10432 13874 10441
rect 13912 10406 13964 10412
rect 13818 10367 13874 10376
rect 13832 10266 13860 10367
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13924 10033 13952 10406
rect 13910 10024 13966 10033
rect 13636 9988 13688 9994
rect 13910 9959 13966 9968
rect 13636 9930 13688 9936
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13648 9382 13676 9454
rect 13912 9444 13964 9450
rect 13912 9386 13964 9392
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13648 8634 13676 9318
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 13728 8084 13780 8090
rect 13832 8072 13860 8910
rect 13924 8838 13952 9386
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 13924 8634 13952 8774
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 13780 8044 13860 8072
rect 13728 8026 13780 8032
rect 13740 7546 13768 8026
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13924 7546 13952 7822
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 14016 7274 14044 11342
rect 14108 7410 14136 11478
rect 14292 11354 14320 11591
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 14370 10432 14426 10441
rect 14370 10367 14426 10376
rect 14188 10192 14240 10198
rect 14186 10160 14188 10169
rect 14240 10160 14242 10169
rect 14186 10095 14242 10104
rect 14278 8528 14334 8537
rect 14278 8463 14334 8472
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 14004 7268 14056 7274
rect 14004 7210 14056 7216
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13634 5944 13690 5953
rect 13634 5879 13690 5888
rect 13648 5574 13676 5879
rect 13728 5636 13780 5642
rect 13728 5578 13780 5584
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13648 5098 13676 5510
rect 13636 5092 13688 5098
rect 13636 5034 13688 5040
rect 13648 4622 13676 5034
rect 13740 4758 13768 5578
rect 13728 4752 13780 4758
rect 13728 4694 13780 4700
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13464 4134 13584 4162
rect 13634 4176 13690 4185
rect 13464 3942 13492 4134
rect 13634 4111 13690 4120
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13452 3596 13504 3602
rect 13452 3538 13504 3544
rect 13464 2650 13492 3538
rect 13556 2689 13584 4014
rect 13648 3602 13676 4111
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 13740 3398 13768 4558
rect 13832 3670 13860 6258
rect 13910 5672 13966 5681
rect 13910 5607 13966 5616
rect 13924 4010 13952 5607
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 13912 4004 13964 4010
rect 13912 3946 13964 3952
rect 13924 3738 13952 3946
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 13820 3664 13872 3670
rect 13820 3606 13872 3612
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13542 2680 13598 2689
rect 13452 2644 13504 2650
rect 13542 2615 13598 2624
rect 13452 2586 13504 2592
rect 13740 2378 13768 3334
rect 14016 3194 14044 4082
rect 14004 3188 14056 3194
rect 14004 3130 14056 3136
rect 14108 2802 14136 7142
rect 14200 5001 14228 7686
rect 14292 7410 14320 8463
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14292 7002 14320 7346
rect 14384 7206 14412 10367
rect 14476 7410 14504 11784
rect 14568 10010 14596 11886
rect 14648 11892 14700 11898
rect 14738 11863 14794 11872
rect 14648 11834 14700 11840
rect 14752 11762 14780 11863
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14844 11558 14872 21984
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15304 19990 15332 23462
rect 15384 23180 15436 23186
rect 15384 23122 15436 23128
rect 15396 22438 15424 23122
rect 15476 22976 15528 22982
rect 15474 22944 15476 22953
rect 15528 22944 15530 22953
rect 15474 22879 15530 22888
rect 16408 22778 16436 24375
rect 16856 24268 16908 24274
rect 16856 24210 16908 24216
rect 17408 24268 17460 24274
rect 17408 24210 17460 24216
rect 16868 23526 16896 24210
rect 17038 24032 17094 24041
rect 17038 23967 17094 23976
rect 17052 23866 17080 23967
rect 17040 23860 17092 23866
rect 17040 23802 17092 23808
rect 17420 23662 17448 24210
rect 17788 24138 17816 24375
rect 18156 24177 18184 24783
rect 18524 24410 18552 27520
rect 18878 24712 18934 24721
rect 18878 24647 18934 24656
rect 18892 24410 18920 24647
rect 18512 24404 18564 24410
rect 18512 24346 18564 24352
rect 18880 24404 18932 24410
rect 18880 24346 18932 24352
rect 18972 24268 19024 24274
rect 18972 24210 19024 24216
rect 18142 24168 18198 24177
rect 17776 24132 17828 24138
rect 18142 24103 18198 24112
rect 17776 24074 17828 24080
rect 18234 23896 18290 23905
rect 18234 23831 18236 23840
rect 18288 23831 18290 23840
rect 18236 23802 18288 23808
rect 17408 23656 17460 23662
rect 17408 23598 17460 23604
rect 16856 23520 16908 23526
rect 16856 23462 16908 23468
rect 17222 23488 17278 23497
rect 16868 22778 16896 23462
rect 17222 23423 17278 23432
rect 17236 23322 17264 23423
rect 17224 23316 17276 23322
rect 17224 23258 17276 23264
rect 17040 23180 17092 23186
rect 17040 23122 17092 23128
rect 17052 23089 17080 23122
rect 17038 23080 17094 23089
rect 17038 23015 17094 23024
rect 17052 22778 17080 23015
rect 16396 22772 16448 22778
rect 16396 22714 16448 22720
rect 16856 22772 16908 22778
rect 16856 22714 16908 22720
rect 17040 22772 17092 22778
rect 17040 22714 17092 22720
rect 15476 22568 15528 22574
rect 15476 22510 15528 22516
rect 15384 22432 15436 22438
rect 15384 22374 15436 22380
rect 15292 19984 15344 19990
rect 15292 19926 15344 19932
rect 15108 19916 15160 19922
rect 15108 19858 15160 19864
rect 15120 19802 15148 19858
rect 15120 19774 15332 19802
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15304 18970 15332 19774
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 15396 18630 15424 22374
rect 15488 19417 15516 22510
rect 15568 22092 15620 22098
rect 15568 22034 15620 22040
rect 15580 21690 15608 22034
rect 16670 21992 16726 22001
rect 16670 21927 16672 21936
rect 16724 21927 16726 21936
rect 16672 21898 16724 21904
rect 15568 21684 15620 21690
rect 15568 21626 15620 21632
rect 15580 21146 15608 21626
rect 15568 21140 15620 21146
rect 15568 21082 15620 21088
rect 15580 20602 15608 21082
rect 15568 20596 15620 20602
rect 15568 20538 15620 20544
rect 15750 19952 15806 19961
rect 15750 19887 15806 19896
rect 15474 19408 15530 19417
rect 15474 19343 15530 19352
rect 15384 18624 15436 18630
rect 15384 18566 15436 18572
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15658 17368 15714 17377
rect 15658 17303 15714 17312
rect 15672 16658 15700 17303
rect 15764 16794 15792 19887
rect 17314 18728 17370 18737
rect 17314 18663 17370 18672
rect 16210 17776 16266 17785
rect 16210 17711 16266 17720
rect 16026 17096 16082 17105
rect 16026 17031 16082 17040
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 15660 16652 15712 16658
rect 15660 16594 15712 16600
rect 15292 16448 15344 16454
rect 15292 16390 15344 16396
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 15120 15609 15148 15846
rect 15304 15745 15332 16390
rect 15672 16046 15700 16594
rect 15764 16182 15792 16730
rect 15934 16688 15990 16697
rect 15934 16623 15990 16632
rect 15948 16590 15976 16623
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 15948 16250 15976 16526
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 15752 16176 15804 16182
rect 15752 16118 15804 16124
rect 15660 16040 15712 16046
rect 15660 15982 15712 15988
rect 15290 15736 15346 15745
rect 15290 15671 15346 15680
rect 15752 15632 15804 15638
rect 15106 15600 15162 15609
rect 15752 15574 15804 15580
rect 15106 15535 15162 15544
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15764 14822 15792 15574
rect 15936 15564 15988 15570
rect 15936 15506 15988 15512
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 14936 14618 14964 14758
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15396 13870 15424 14758
rect 15568 14544 15620 14550
rect 15568 14486 15620 14492
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15488 13530 15516 14214
rect 15580 13870 15608 14486
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15568 13864 15620 13870
rect 15568 13806 15620 13812
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15580 13394 15608 13806
rect 15672 13530 15700 14418
rect 15660 13524 15712 13530
rect 15660 13466 15712 13472
rect 15764 13394 15792 14758
rect 15856 14550 15884 15438
rect 15948 14822 15976 15506
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15844 14544 15896 14550
rect 15844 14486 15896 14492
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15568 13252 15620 13258
rect 15568 13194 15620 13200
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15212 12730 15240 12786
rect 15120 12702 15240 12730
rect 15120 12442 15148 12702
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14832 11552 14884 11558
rect 14646 11520 14702 11529
rect 14832 11494 14884 11500
rect 14646 11455 14702 11464
rect 14660 11014 14688 11455
rect 14738 11248 14794 11257
rect 14738 11183 14794 11192
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14660 10810 14688 10950
rect 14752 10810 14780 11183
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 14740 10804 14792 10810
rect 14740 10746 14792 10752
rect 14568 9982 14688 10010
rect 14556 9920 14608 9926
rect 14554 9888 14556 9897
rect 14608 9888 14610 9897
rect 14554 9823 14610 9832
rect 14556 8968 14608 8974
rect 14554 8936 14556 8945
rect 14608 8936 14610 8945
rect 14554 8871 14610 8880
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14464 7268 14516 7274
rect 14464 7210 14516 7216
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 14292 6662 14320 6802
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14292 6089 14320 6598
rect 14278 6080 14334 6089
rect 14278 6015 14334 6024
rect 14186 4992 14242 5001
rect 14186 4927 14242 4936
rect 14200 3602 14228 4927
rect 14372 4548 14424 4554
rect 14372 4490 14424 4496
rect 14384 4078 14412 4490
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14384 3641 14412 3674
rect 14370 3632 14426 3641
rect 14188 3596 14240 3602
rect 14370 3567 14426 3576
rect 14188 3538 14240 3544
rect 14186 3224 14242 3233
rect 14186 3159 14242 3168
rect 14016 2774 14136 2802
rect 14016 2666 14044 2774
rect 13924 2638 14044 2666
rect 14200 2650 14228 3159
rect 14476 3108 14504 7210
rect 14660 7154 14688 9982
rect 14568 7126 14688 7154
rect 14568 3670 14596 7126
rect 14646 7032 14702 7041
rect 14646 6967 14702 6976
rect 14660 6186 14688 6967
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14648 6180 14700 6186
rect 14648 6122 14700 6128
rect 14660 5914 14688 6122
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14660 5370 14688 5850
rect 14648 5364 14700 5370
rect 14648 5306 14700 5312
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 14660 3738 14688 4626
rect 14752 4078 14780 6598
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14556 3664 14608 3670
rect 14556 3606 14608 3612
rect 14568 3233 14596 3606
rect 14740 3392 14792 3398
rect 14740 3334 14792 3340
rect 14554 3224 14610 3233
rect 14554 3159 14610 3168
rect 14476 3080 14596 3108
rect 14568 2802 14596 3080
rect 14559 2774 14596 2802
rect 14559 2666 14587 2774
rect 14188 2644 14240 2650
rect 13728 2372 13780 2378
rect 13728 2314 13780 2320
rect 13924 480 13952 2638
rect 14188 2586 14240 2592
rect 14464 2644 14516 2650
rect 14559 2638 14596 2666
rect 14752 2650 14780 3334
rect 14844 3108 14872 11494
rect 14922 11384 14978 11393
rect 14922 11319 14924 11328
rect 14976 11319 14978 11328
rect 14924 11290 14976 11296
rect 15304 11150 15332 12038
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15304 10792 15332 11086
rect 15120 10764 15332 10792
rect 15120 10266 15148 10764
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15396 9654 15424 11698
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15488 11218 15516 11494
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 14924 9104 14976 9110
rect 14922 9072 14924 9081
rect 14976 9072 14978 9081
rect 14922 9007 14978 9016
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15290 7848 15346 7857
rect 15290 7783 15346 7792
rect 15474 7848 15530 7857
rect 15474 7783 15530 7792
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15304 7478 15332 7783
rect 15488 7546 15516 7783
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15292 7472 15344 7478
rect 15292 7414 15344 7420
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 15120 6746 15148 7346
rect 15488 7342 15516 7482
rect 15476 7336 15528 7342
rect 15476 7278 15528 7284
rect 15120 6718 15332 6746
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15212 5681 15240 6054
rect 15198 5672 15254 5681
rect 15198 5607 15254 5616
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15304 4690 15332 6718
rect 15384 5568 15436 5574
rect 15382 5536 15384 5545
rect 15436 5536 15438 5545
rect 15382 5471 15438 5480
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15304 4282 15332 4626
rect 15474 4584 15530 4593
rect 15474 4519 15476 4528
rect 15528 4519 15530 4528
rect 15476 4490 15528 4496
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 15476 4072 15528 4078
rect 15476 4014 15528 4020
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15108 3120 15160 3126
rect 14844 3080 14964 3108
rect 14464 2586 14516 2592
rect 14476 2281 14504 2586
rect 14462 2272 14518 2281
rect 14462 2207 14518 2216
rect 14372 1896 14424 1902
rect 14370 1864 14372 1873
rect 14424 1864 14426 1873
rect 14370 1799 14426 1808
rect 14568 480 14596 2638
rect 14740 2644 14792 2650
rect 14936 2632 14964 3080
rect 15108 3062 15160 3068
rect 15120 2990 15148 3062
rect 15108 2984 15160 2990
rect 15108 2926 15160 2932
rect 15488 2650 15516 4014
rect 14740 2586 14792 2592
rect 14844 2604 14964 2632
rect 15476 2644 15528 2650
rect 14738 2544 14794 2553
rect 14738 2479 14740 2488
rect 14792 2479 14794 2488
rect 14740 2450 14792 2456
rect 14648 2032 14700 2038
rect 14646 2000 14648 2009
rect 14844 2020 14872 2604
rect 15476 2586 15528 2592
rect 15292 2576 15344 2582
rect 14922 2544 14978 2553
rect 15292 2518 15344 2524
rect 14922 2479 14978 2488
rect 14936 2446 14964 2479
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 15304 2310 15332 2518
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14700 2000 14702 2009
rect 14844 1992 15148 2020
rect 14646 1935 14702 1944
rect 15120 480 15148 1992
rect 15304 1601 15332 2246
rect 15488 2145 15516 2314
rect 15474 2136 15530 2145
rect 15474 2071 15530 2080
rect 15290 1592 15346 1601
rect 15290 1527 15346 1536
rect 15580 626 15608 13194
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15856 12442 15884 13126
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 15750 12336 15806 12345
rect 15750 12271 15752 12280
rect 15804 12271 15806 12280
rect 15752 12242 15804 12248
rect 15764 11830 15792 12242
rect 15856 11898 15884 12378
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 15752 11824 15804 11830
rect 15752 11766 15804 11772
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15658 11112 15714 11121
rect 15658 11047 15660 11056
rect 15712 11047 15714 11056
rect 15660 11018 15712 11024
rect 15764 10538 15792 11154
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 15752 10532 15804 10538
rect 15752 10474 15804 10480
rect 15764 10266 15792 10474
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15856 10062 15884 10746
rect 15948 10713 15976 14758
rect 16040 13258 16068 17031
rect 16120 16176 16172 16182
rect 16120 16118 16172 16124
rect 16028 13252 16080 13258
rect 16028 13194 16080 13200
rect 16132 13138 16160 16118
rect 16224 15201 16252 17711
rect 17130 16552 17186 16561
rect 17130 16487 17186 16496
rect 16210 15192 16266 15201
rect 16210 15127 16266 15136
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16684 14414 16712 14758
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16224 13326 16252 13670
rect 16684 13530 16712 14350
rect 16672 13524 16724 13530
rect 16672 13466 16724 13472
rect 16684 13326 16712 13466
rect 16212 13320 16264 13326
rect 16212 13262 16264 13268
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16040 13110 16160 13138
rect 16040 12322 16068 13110
rect 16224 12782 16252 13262
rect 16764 13184 16816 13190
rect 16764 13126 16816 13132
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 16488 12708 16540 12714
rect 16488 12650 16540 12656
rect 16040 12294 16160 12322
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 16040 11218 16068 12174
rect 16028 11212 16080 11218
rect 16028 11154 16080 11160
rect 15934 10704 15990 10713
rect 15934 10639 15990 10648
rect 15936 10124 15988 10130
rect 15936 10066 15988 10072
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15948 9926 15976 10066
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 15936 9920 15988 9926
rect 15936 9862 15988 9868
rect 15948 9110 15976 9862
rect 16040 9518 16068 9998
rect 16028 9512 16080 9518
rect 16028 9454 16080 9460
rect 15936 9104 15988 9110
rect 15936 9046 15988 9052
rect 16040 9042 16068 9454
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15856 8294 15884 8434
rect 15936 8424 15988 8430
rect 15934 8392 15936 8401
rect 15988 8392 15990 8401
rect 15934 8327 15990 8336
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 15672 7546 15700 7822
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 15764 7206 15792 7686
rect 15856 7410 15884 8230
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15672 5166 15700 5714
rect 15660 5160 15712 5166
rect 15658 5128 15660 5137
rect 15712 5128 15714 5137
rect 15658 5063 15714 5072
rect 15764 2038 15792 7142
rect 16040 6798 16068 8978
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 16040 6458 16068 6734
rect 16028 6452 16080 6458
rect 16028 6394 16080 6400
rect 16132 5930 16160 12294
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16408 11354 16436 12038
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16304 11144 16356 11150
rect 16304 11086 16356 11092
rect 16316 10130 16344 11086
rect 16500 10810 16528 12650
rect 16776 11529 16804 13126
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16868 12238 16896 12582
rect 17038 12336 17094 12345
rect 17038 12271 17040 12280
rect 17092 12271 17094 12280
rect 17040 12242 17092 12248
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 17040 12164 17092 12170
rect 17040 12106 17092 12112
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 16762 11520 16818 11529
rect 16762 11455 16818 11464
rect 16960 11257 16988 12038
rect 17052 11558 17080 12106
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 16946 11248 17002 11257
rect 16946 11183 17002 11192
rect 16488 10804 16540 10810
rect 16488 10746 16540 10752
rect 16764 10464 16816 10470
rect 16764 10406 16816 10412
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 16304 9648 16356 9654
rect 16302 9616 16304 9625
rect 16356 9616 16358 9625
rect 16776 9586 16804 10406
rect 17052 10033 17080 11494
rect 17144 11286 17172 16487
rect 17222 16144 17278 16153
rect 17222 16079 17278 16088
rect 17132 11280 17184 11286
rect 17132 11222 17184 11228
rect 17038 10024 17094 10033
rect 17038 9959 17094 9968
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 16302 9551 16358 9560
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16776 9110 16804 9522
rect 16764 9104 16816 9110
rect 16764 9046 16816 9052
rect 16960 9042 16988 9862
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16396 8560 16448 8566
rect 16396 8502 16448 8508
rect 16408 8090 16436 8502
rect 16500 8362 16528 8910
rect 16684 8634 16712 8978
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 16396 7812 16448 7818
rect 16396 7754 16448 7760
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 16316 6934 16344 7346
rect 16304 6928 16356 6934
rect 16304 6870 16356 6876
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 16040 5902 16160 5930
rect 15842 5672 15898 5681
rect 15842 5607 15844 5616
rect 15896 5607 15898 5616
rect 15844 5578 15896 5584
rect 16040 4865 16068 5902
rect 16120 5840 16172 5846
rect 16120 5782 16172 5788
rect 16026 4856 16082 4865
rect 16132 4826 16160 5782
rect 16224 4826 16252 6598
rect 16304 6112 16356 6118
rect 16408 6100 16436 7754
rect 16500 6866 16528 8298
rect 16960 8090 16988 8978
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 16488 6452 16540 6458
rect 16488 6394 16540 6400
rect 16356 6072 16436 6100
rect 16304 6054 16356 6060
rect 16500 5710 16528 6394
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16500 5370 16528 5646
rect 16488 5364 16540 5370
rect 16316 5324 16488 5352
rect 16026 4791 16082 4800
rect 16120 4820 16172 4826
rect 16120 4762 16172 4768
rect 16212 4820 16264 4826
rect 16212 4762 16264 4768
rect 16132 4282 16160 4762
rect 16120 4276 16172 4282
rect 16120 4218 16172 4224
rect 16224 4214 16252 4762
rect 16212 4208 16264 4214
rect 16212 4150 16264 4156
rect 15936 4004 15988 4010
rect 15936 3946 15988 3952
rect 15948 3738 15976 3946
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 15948 2446 15976 3674
rect 16316 3534 16344 5324
rect 16488 5306 16540 5312
rect 16592 5166 16620 7686
rect 16776 7206 16804 7822
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16776 7002 16804 7142
rect 16764 6996 16816 7002
rect 16764 6938 16816 6944
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16684 5574 16712 6802
rect 16776 5846 16804 6938
rect 16856 6248 16908 6254
rect 16854 6216 16856 6225
rect 16908 6216 16910 6225
rect 16854 6151 16910 6160
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 16764 5840 16816 5846
rect 16764 5782 16816 5788
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16946 5536 17002 5545
rect 16580 5160 16632 5166
rect 16580 5102 16632 5108
rect 16488 5092 16540 5098
rect 16488 5034 16540 5040
rect 16396 5024 16448 5030
rect 16394 4992 16396 5001
rect 16448 4992 16450 5001
rect 16394 4927 16450 4936
rect 16500 3942 16528 5034
rect 16684 4978 16712 5510
rect 16946 5471 17002 5480
rect 16854 5128 16910 5137
rect 16854 5063 16856 5072
rect 16908 5063 16910 5072
rect 16856 5034 16908 5040
rect 16592 4950 16712 4978
rect 16592 4622 16620 4950
rect 16960 4826 16988 5471
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 16856 4684 16908 4690
rect 16856 4626 16908 4632
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16592 4010 16620 4558
rect 16580 4004 16632 4010
rect 16580 3946 16632 3952
rect 16488 3936 16540 3942
rect 16488 3878 16540 3884
rect 16868 3738 16896 4626
rect 17052 4457 17080 6054
rect 17038 4448 17094 4457
rect 17038 4383 17094 4392
rect 16672 3732 16724 3738
rect 16672 3674 16724 3680
rect 16856 3732 16908 3738
rect 16856 3674 16908 3680
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 16212 3460 16264 3466
rect 16212 3402 16264 3408
rect 15936 2440 15988 2446
rect 15936 2382 15988 2388
rect 15752 2032 15804 2038
rect 15752 1974 15804 1980
rect 15580 598 15700 626
rect 15672 480 15700 598
rect 16224 480 16252 3402
rect 16316 3194 16344 3470
rect 16500 3194 16528 3538
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16500 2650 16528 3130
rect 16488 2644 16540 2650
rect 16488 2586 16540 2592
rect 16684 2553 16712 3674
rect 17236 3194 17264 16079
rect 17328 13530 17356 18663
rect 17420 17649 17448 23598
rect 18984 23526 19012 24210
rect 17592 23520 17644 23526
rect 17592 23462 17644 23468
rect 18604 23520 18656 23526
rect 18604 23462 18656 23468
rect 18972 23520 19024 23526
rect 19076 23497 19104 27520
rect 19628 25786 19656 27520
rect 19444 25758 19656 25786
rect 19444 24449 19472 25758
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19430 24440 19486 24449
rect 19622 24432 19918 24452
rect 19430 24375 19486 24384
rect 19706 24032 19762 24041
rect 19706 23967 19762 23976
rect 19720 23866 19748 23967
rect 20272 23905 20300 27520
rect 20824 24721 20852 27520
rect 20810 24712 20866 24721
rect 20810 24647 20866 24656
rect 20812 24268 20864 24274
rect 20812 24210 20864 24216
rect 20258 23896 20314 23905
rect 19708 23860 19760 23866
rect 20258 23831 20314 23840
rect 19708 23802 19760 23808
rect 19432 23656 19484 23662
rect 19432 23598 19484 23604
rect 18972 23462 19024 23468
rect 19062 23488 19118 23497
rect 17604 21457 17632 23462
rect 18236 23180 18288 23186
rect 18236 23122 18288 23128
rect 18248 22438 18276 23122
rect 18512 22500 18564 22506
rect 18512 22442 18564 22448
rect 18236 22432 18288 22438
rect 18236 22374 18288 22380
rect 17590 21448 17646 21457
rect 17590 21383 17646 21392
rect 17498 19136 17554 19145
rect 17498 19071 17554 19080
rect 17406 17640 17462 17649
rect 17406 17575 17462 17584
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 17328 12345 17356 13466
rect 17420 13462 17448 17575
rect 17408 13456 17460 13462
rect 17408 13398 17460 13404
rect 17420 12986 17448 13398
rect 17408 12980 17460 12986
rect 17408 12922 17460 12928
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 17314 12336 17370 12345
rect 17314 12271 17370 12280
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17328 11694 17356 12174
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 17328 6186 17356 11630
rect 17420 11218 17448 12378
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17420 10470 17448 11154
rect 17408 10464 17460 10470
rect 17406 10432 17408 10441
rect 17460 10432 17462 10441
rect 17406 10367 17462 10376
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17420 9178 17448 9318
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17316 6180 17368 6186
rect 17316 6122 17368 6128
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 16762 2816 16818 2825
rect 16762 2751 16818 2760
rect 16670 2544 16726 2553
rect 16670 2479 16726 2488
rect 16684 2009 16712 2479
rect 16670 2000 16726 2009
rect 16670 1935 16726 1944
rect 16776 480 16804 2751
rect 17130 2680 17186 2689
rect 17130 2615 17186 2624
rect 17144 2514 17172 2615
rect 17132 2508 17184 2514
rect 17132 2450 17184 2456
rect 17328 2394 17356 6122
rect 17406 5400 17462 5409
rect 17406 5335 17408 5344
rect 17460 5335 17462 5344
rect 17408 5306 17460 5312
rect 17512 4842 17540 19071
rect 17604 12442 17632 21383
rect 18248 17241 18276 22374
rect 18234 17232 18290 17241
rect 18234 17167 18290 17176
rect 18326 13424 18382 13433
rect 18326 13359 18382 13368
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17696 12322 17724 13262
rect 18340 12782 18368 13359
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 18064 12442 18092 12718
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 17604 12294 17724 12322
rect 17604 12238 17632 12294
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 17604 11558 17632 12174
rect 17592 11552 17644 11558
rect 17592 11494 17644 11500
rect 18050 11384 18106 11393
rect 18050 11319 18106 11328
rect 17868 11144 17920 11150
rect 17920 11092 18000 11098
rect 17868 11086 18000 11092
rect 17880 11070 18000 11086
rect 17972 9586 18000 11070
rect 18064 10810 18092 11319
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 18236 10532 18288 10538
rect 18236 10474 18288 10480
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 18064 10305 18092 10406
rect 18050 10296 18106 10305
rect 18050 10231 18052 10240
rect 18104 10231 18106 10240
rect 18052 10202 18104 10208
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 17592 9512 17644 9518
rect 17592 9454 17644 9460
rect 17604 8090 17632 9454
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17788 8430 17816 9318
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 17972 8537 18000 8774
rect 18064 8634 18092 10202
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 17958 8528 18014 8537
rect 17958 8463 18014 8472
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17776 8016 17828 8022
rect 17776 7958 17828 7964
rect 17788 5352 17816 7958
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17880 7274 17908 7822
rect 17972 7342 18000 7890
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 17868 7268 17920 7274
rect 17868 7210 17920 7216
rect 18064 6497 18092 8230
rect 18248 7154 18276 10474
rect 18524 10266 18552 22442
rect 18616 16561 18644 23462
rect 18984 23322 19012 23462
rect 19062 23423 19118 23432
rect 18972 23316 19024 23322
rect 18972 23258 19024 23264
rect 19340 22568 19392 22574
rect 19338 22536 19340 22545
rect 19392 22536 19394 22545
rect 19338 22471 19394 22480
rect 19444 19825 19472 23598
rect 20824 23526 20852 24210
rect 21376 24041 21404 27520
rect 21362 24032 21418 24041
rect 21362 23967 21418 23976
rect 21362 23896 21418 23905
rect 21362 23831 21364 23840
rect 21416 23831 21418 23840
rect 21364 23802 21416 23808
rect 21088 23656 21140 23662
rect 21088 23598 21140 23604
rect 20812 23520 20864 23526
rect 20812 23462 20864 23468
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19430 19816 19486 19825
rect 19430 19751 19486 19760
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 20824 17377 20852 23462
rect 21100 23322 21128 23598
rect 21088 23316 21140 23322
rect 21088 23258 21140 23264
rect 20902 23216 20958 23225
rect 20902 23151 20904 23160
rect 20956 23151 20958 23160
rect 20904 23122 20956 23128
rect 20916 22778 20944 23122
rect 21928 22953 21956 27520
rect 22480 24410 22508 27520
rect 22468 24404 22520 24410
rect 22468 24346 22520 24352
rect 23124 23905 23152 27520
rect 23110 23896 23166 23905
rect 23110 23831 23166 23840
rect 23480 23656 23532 23662
rect 23676 23633 23704 27520
rect 24228 24857 24256 27520
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24214 24848 24270 24857
rect 24214 24783 24270 24792
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 23480 23598 23532 23604
rect 23662 23624 23718 23633
rect 23492 23322 23520 23598
rect 23662 23559 23718 23568
rect 23570 23352 23626 23361
rect 23480 23316 23532 23322
rect 23570 23287 23626 23296
rect 23480 23258 23532 23264
rect 22192 23180 22244 23186
rect 22192 23122 22244 23128
rect 21914 22944 21970 22953
rect 21914 22879 21970 22888
rect 20904 22772 20956 22778
rect 20904 22714 20956 22720
rect 22204 22574 22232 23122
rect 22192 22568 22244 22574
rect 22192 22510 22244 22516
rect 23584 22001 23612 23287
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24780 22681 24808 27520
rect 25332 23866 25360 27520
rect 25976 24177 26004 27520
rect 26528 24313 26556 27520
rect 26514 24304 26570 24313
rect 26514 24239 26570 24248
rect 25962 24168 26018 24177
rect 25962 24103 26018 24112
rect 25320 23860 25372 23866
rect 25320 23802 25372 23808
rect 27080 23769 27108 27520
rect 27066 23760 27122 23769
rect 27066 23695 27122 23704
rect 24766 22672 24822 22681
rect 24766 22607 24822 22616
rect 23570 21992 23626 22001
rect 23570 21927 23626 21936
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 27632 18737 27660 27520
rect 27618 18728 27674 18737
rect 27618 18663 27674 18672
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 20810 17368 20866 17377
rect 24289 17360 24585 17380
rect 20810 17303 20866 17312
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 18602 16552 18658 16561
rect 18602 16487 18658 16496
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 19338 15192 19394 15201
rect 24289 15184 24585 15204
rect 19338 15127 19394 15136
rect 18604 11552 18656 11558
rect 18604 11494 18656 11500
rect 18616 11014 18644 11494
rect 18970 11112 19026 11121
rect 18970 11047 19026 11056
rect 18604 11008 18656 11014
rect 18604 10950 18656 10956
rect 18616 10674 18644 10950
rect 18604 10668 18656 10674
rect 18604 10610 18656 10616
rect 18984 10266 19012 11047
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 18972 10260 19024 10266
rect 18972 10202 19024 10208
rect 18880 10124 18932 10130
rect 18880 10066 18932 10072
rect 18892 9625 18920 10066
rect 19064 10056 19116 10062
rect 19064 9998 19116 10004
rect 19076 9722 19104 9998
rect 19352 9722 19380 15127
rect 19522 15056 19578 15065
rect 19522 14991 19578 15000
rect 19432 12640 19484 12646
rect 19430 12608 19432 12617
rect 19484 12608 19486 12617
rect 19430 12543 19486 12552
rect 19432 10260 19484 10266
rect 19432 10202 19484 10208
rect 19064 9716 19116 9722
rect 19064 9658 19116 9664
rect 19340 9716 19392 9722
rect 19340 9658 19392 9664
rect 19444 9654 19472 10202
rect 18972 9648 19024 9654
rect 18878 9616 18934 9625
rect 18604 9580 18656 9586
rect 19432 9648 19484 9654
rect 18972 9590 19024 9596
rect 19338 9616 19394 9625
rect 18878 9551 18934 9560
rect 18604 9522 18656 9528
rect 18616 8838 18644 9522
rect 18984 9178 19012 9590
rect 19432 9590 19484 9596
rect 19338 9551 19394 9560
rect 19352 9178 19380 9551
rect 18972 9172 19024 9178
rect 18972 9114 19024 9120
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 18420 8356 18472 8362
rect 18420 8298 18472 8304
rect 18432 8265 18460 8298
rect 18418 8256 18474 8265
rect 18418 8191 18474 8200
rect 18616 7886 18644 8774
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18328 7812 18380 7818
rect 18328 7754 18380 7760
rect 18340 7478 18368 7754
rect 18604 7744 18656 7750
rect 18708 7698 18736 8434
rect 18656 7692 18736 7698
rect 18604 7686 18736 7692
rect 18616 7670 18736 7686
rect 18328 7472 18380 7478
rect 18328 7414 18380 7420
rect 18510 7440 18566 7449
rect 18510 7375 18512 7384
rect 18564 7375 18566 7384
rect 18512 7346 18564 7352
rect 18420 7336 18472 7342
rect 18420 7278 18472 7284
rect 18326 7168 18382 7177
rect 18248 7126 18326 7154
rect 18326 7103 18382 7112
rect 18432 7002 18460 7278
rect 18512 7268 18564 7274
rect 18512 7210 18564 7216
rect 18420 6996 18472 7002
rect 18420 6938 18472 6944
rect 18050 6488 18106 6497
rect 18050 6423 18106 6432
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 18156 5914 18184 6190
rect 18234 6080 18290 6089
rect 18234 6015 18290 6024
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 17958 5672 18014 5681
rect 17958 5607 18014 5616
rect 17788 5324 17908 5352
rect 17774 5264 17830 5273
rect 17774 5199 17776 5208
rect 17828 5199 17830 5208
rect 17776 5170 17828 5176
rect 17512 4814 17632 4842
rect 17498 4720 17554 4729
rect 17498 4655 17500 4664
rect 17552 4655 17554 4664
rect 17500 4626 17552 4632
rect 17500 4480 17552 4486
rect 17500 4422 17552 4428
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17420 2961 17448 3878
rect 17406 2952 17462 2961
rect 17406 2887 17462 2896
rect 17236 2366 17356 2394
rect 17236 1329 17264 2366
rect 17316 2304 17368 2310
rect 17512 2258 17540 4422
rect 17604 3194 17632 4814
rect 17684 4616 17736 4622
rect 17684 4558 17736 4564
rect 17696 3738 17724 4558
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17684 3732 17736 3738
rect 17684 3674 17736 3680
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17788 3097 17816 3878
rect 17774 3088 17830 3097
rect 17774 3023 17830 3032
rect 17880 2650 17908 5324
rect 17868 2644 17920 2650
rect 17868 2586 17920 2592
rect 17316 2246 17368 2252
rect 17328 1465 17356 2246
rect 17420 2230 17540 2258
rect 17314 1456 17370 1465
rect 17314 1391 17370 1400
rect 17222 1320 17278 1329
rect 17222 1255 17278 1264
rect 17420 480 17448 2230
rect 17972 480 18000 5607
rect 18156 5302 18184 5850
rect 18248 5370 18276 6015
rect 18326 5808 18382 5817
rect 18326 5743 18382 5752
rect 18236 5364 18288 5370
rect 18236 5306 18288 5312
rect 18144 5296 18196 5302
rect 18144 5238 18196 5244
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 18052 4684 18104 4690
rect 18052 4626 18104 4632
rect 18064 4049 18092 4626
rect 18050 4040 18106 4049
rect 18050 3975 18106 3984
rect 18064 3942 18092 3975
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 18156 3194 18184 4762
rect 18340 4486 18368 5743
rect 18524 5273 18552 7210
rect 18616 6361 18644 7670
rect 18788 7404 18840 7410
rect 18788 7346 18840 7352
rect 19340 7404 19392 7410
rect 19340 7346 19392 7352
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18602 6352 18658 6361
rect 18602 6287 18658 6296
rect 18708 6254 18736 6598
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 18510 5264 18566 5273
rect 18510 5199 18566 5208
rect 18604 5228 18656 5234
rect 18524 5166 18552 5199
rect 18604 5170 18656 5176
rect 18512 5160 18564 5166
rect 18512 5102 18564 5108
rect 18616 4622 18644 5170
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18524 4282 18552 4558
rect 18512 4276 18564 4282
rect 18512 4218 18564 4224
rect 18800 4146 18828 7346
rect 19246 7168 19302 7177
rect 19246 7103 19302 7112
rect 19260 7002 19288 7103
rect 19352 7041 19380 7346
rect 19338 7032 19394 7041
rect 19248 6996 19300 7002
rect 19338 6967 19394 6976
rect 19248 6938 19300 6944
rect 19260 5914 19288 6938
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19352 6186 19380 6734
rect 19444 6390 19472 6734
rect 19432 6384 19484 6390
rect 19430 6352 19432 6361
rect 19484 6352 19486 6361
rect 19430 6287 19486 6296
rect 19340 6180 19392 6186
rect 19340 6122 19392 6128
rect 19444 6066 19472 6287
rect 19352 6038 19472 6066
rect 19248 5908 19300 5914
rect 19248 5850 19300 5856
rect 19352 5710 19380 6038
rect 19430 5944 19486 5953
rect 19536 5914 19564 14991
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 20076 7744 20128 7750
rect 20076 7686 20128 7692
rect 20088 7206 20116 7686
rect 19984 7200 20036 7206
rect 19984 7142 20036 7148
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19996 6662 20024 7142
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19996 6458 20024 6598
rect 19984 6452 20036 6458
rect 19984 6394 20036 6400
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19430 5879 19486 5888
rect 19524 5908 19576 5914
rect 19444 5846 19472 5879
rect 19524 5850 19576 5856
rect 19432 5840 19484 5846
rect 19432 5782 19484 5788
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19536 5302 19564 5850
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 19800 5704 19852 5710
rect 19800 5646 19852 5652
rect 19524 5296 19576 5302
rect 19524 5238 19576 5244
rect 18972 5024 19024 5030
rect 18972 4966 19024 4972
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 18984 4185 19012 4966
rect 19062 4448 19118 4457
rect 19062 4383 19118 4392
rect 18970 4176 19026 4185
rect 18788 4140 18840 4146
rect 18708 4100 18788 4128
rect 18708 3738 18736 4100
rect 18970 4111 19026 4120
rect 18788 4082 18840 4088
rect 18786 3904 18842 3913
rect 18786 3839 18842 3848
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 18800 3534 18828 3839
rect 18972 3596 19024 3602
rect 18972 3538 19024 3544
rect 18788 3528 18840 3534
rect 18788 3470 18840 3476
rect 18510 3224 18566 3233
rect 18144 3188 18196 3194
rect 18800 3194 18828 3470
rect 18984 3398 19012 3538
rect 18972 3392 19024 3398
rect 18972 3334 19024 3340
rect 18510 3159 18566 3168
rect 18788 3188 18840 3194
rect 18144 3130 18196 3136
rect 18524 480 18552 3159
rect 18788 3130 18840 3136
rect 18984 3058 19012 3334
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 18972 2916 19024 2922
rect 18972 2858 19024 2864
rect 18984 2553 19012 2858
rect 18970 2544 19026 2553
rect 18696 2508 18748 2514
rect 18970 2479 19026 2488
rect 18696 2450 18748 2456
rect 18708 1902 18736 2450
rect 18880 2440 18932 2446
rect 18880 2382 18932 2388
rect 18696 1896 18748 1902
rect 18696 1838 18748 1844
rect 18892 1601 18920 2382
rect 18970 2000 19026 2009
rect 18970 1935 19026 1944
rect 18984 1737 19012 1935
rect 18970 1728 19026 1737
rect 18970 1663 19026 1672
rect 18878 1592 18934 1601
rect 18878 1527 18934 1536
rect 19076 480 19104 4383
rect 19352 4321 19380 4966
rect 19536 4690 19564 5238
rect 19812 5234 19840 5646
rect 19800 5228 19852 5234
rect 19800 5170 19852 5176
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19996 4758 20024 5714
rect 19984 4752 20036 4758
rect 19984 4694 20036 4700
rect 19524 4684 19576 4690
rect 19524 4626 19576 4632
rect 19338 4312 19394 4321
rect 19338 4247 19394 4256
rect 19536 4214 19564 4626
rect 19524 4208 19576 4214
rect 19524 4150 19576 4156
rect 20180 4078 20208 9658
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 20536 7472 20588 7478
rect 20536 7414 20588 7420
rect 20260 5228 20312 5234
rect 20260 5170 20312 5176
rect 20272 4826 20300 5170
rect 20548 5148 20576 7414
rect 22282 7304 22338 7313
rect 22282 7239 22338 7248
rect 20628 7200 20680 7206
rect 20680 7160 20760 7188
rect 20628 7142 20680 7148
rect 20732 5914 20760 7160
rect 22190 6760 22246 6769
rect 20996 6724 21048 6730
rect 22190 6695 22246 6704
rect 20996 6666 21048 6672
rect 20902 6488 20958 6497
rect 20902 6423 20958 6432
rect 20916 6254 20944 6423
rect 21008 6322 21036 6666
rect 20996 6316 21048 6322
rect 20996 6258 21048 6264
rect 21456 6316 21508 6322
rect 21456 6258 21508 6264
rect 20904 6248 20956 6254
rect 20904 6190 20956 6196
rect 20720 5908 20772 5914
rect 20720 5850 20772 5856
rect 21468 5846 21496 6258
rect 21456 5840 21508 5846
rect 21456 5782 21508 5788
rect 20720 5772 20772 5778
rect 20720 5714 20772 5720
rect 20732 5370 20760 5714
rect 21468 5710 21496 5782
rect 22008 5772 22060 5778
rect 22008 5714 22060 5720
rect 21456 5704 21508 5710
rect 21456 5646 21508 5652
rect 21468 5370 21496 5646
rect 21548 5636 21600 5642
rect 21548 5578 21600 5584
rect 20720 5364 20772 5370
rect 20720 5306 20772 5312
rect 21456 5364 21508 5370
rect 21456 5306 21508 5312
rect 20720 5160 20772 5166
rect 20548 5120 20720 5148
rect 20720 5102 20772 5108
rect 21364 5024 21416 5030
rect 21364 4966 21416 4972
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 21178 4720 21234 4729
rect 21376 4690 21404 4966
rect 21560 4826 21588 5578
rect 21638 5400 21694 5409
rect 22020 5386 22048 5714
rect 22020 5370 22140 5386
rect 22020 5364 22152 5370
rect 22020 5358 22100 5364
rect 21638 5335 21694 5344
rect 21548 4820 21600 4826
rect 21548 4762 21600 4768
rect 21652 4729 21680 5335
rect 22100 5306 22152 5312
rect 21824 5160 21876 5166
rect 21824 5102 21876 5108
rect 21836 4826 21864 5102
rect 22204 4842 22232 6695
rect 22296 6254 22324 7239
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 22468 6112 22520 6118
rect 22468 6054 22520 6060
rect 22480 5778 22508 6054
rect 22468 5772 22520 5778
rect 22468 5714 22520 5720
rect 23296 5772 23348 5778
rect 23296 5714 23348 5720
rect 23308 5370 23336 5714
rect 23480 5568 23532 5574
rect 23480 5510 23532 5516
rect 23296 5364 23348 5370
rect 23296 5306 23348 5312
rect 22376 5296 22428 5302
rect 22374 5264 22376 5273
rect 22428 5264 22430 5273
rect 22374 5199 22430 5208
rect 22744 5160 22796 5166
rect 22742 5128 22744 5137
rect 22796 5128 22798 5137
rect 22742 5063 22798 5072
rect 21824 4820 21876 4826
rect 22204 4814 22324 4842
rect 21824 4762 21876 4768
rect 21638 4720 21694 4729
rect 21178 4655 21234 4664
rect 21364 4684 21416 4690
rect 20536 4480 20588 4486
rect 20536 4422 20588 4428
rect 20812 4480 20864 4486
rect 20812 4422 20864 4428
rect 20548 4282 20576 4422
rect 20536 4276 20588 4282
rect 20536 4218 20588 4224
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 20168 4072 20220 4078
rect 20168 4014 20220 4020
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 19444 3670 19472 3878
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 20272 3738 20300 4082
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 19432 3528 19484 3534
rect 19154 3496 19210 3505
rect 19432 3470 19484 3476
rect 19154 3431 19156 3440
rect 19208 3431 19210 3440
rect 19156 3402 19208 3408
rect 19156 2984 19208 2990
rect 19156 2926 19208 2932
rect 19248 2984 19300 2990
rect 19248 2926 19300 2932
rect 19168 2496 19196 2926
rect 19260 2650 19288 2926
rect 19248 2644 19300 2650
rect 19248 2586 19300 2592
rect 19340 2508 19392 2514
rect 19168 2468 19340 2496
rect 19340 2450 19392 2456
rect 19444 1193 19472 3470
rect 19536 3194 19564 3538
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 20628 3188 20680 3194
rect 20628 3130 20680 3136
rect 20168 3052 20220 3058
rect 20168 2994 20220 3000
rect 19524 2916 19576 2922
rect 19524 2858 19576 2864
rect 19430 1184 19486 1193
rect 19430 1119 19486 1128
rect 19536 921 19564 2858
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 20076 2304 20128 2310
rect 20076 2246 20128 2252
rect 20088 1601 20116 2246
rect 20074 1592 20130 1601
rect 20074 1527 20130 1536
rect 19614 1456 19670 1465
rect 19614 1391 19670 1400
rect 19522 912 19578 921
rect 19522 847 19578 856
rect 19628 480 19656 1391
rect 20180 1057 20208 2994
rect 20640 2650 20668 3130
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 20258 1456 20314 1465
rect 20258 1391 20314 1400
rect 20166 1048 20222 1057
rect 20166 983 20222 992
rect 20272 480 20300 1391
rect 20824 480 20852 4422
rect 21192 4078 21220 4655
rect 21638 4655 21694 4664
rect 21364 4626 21416 4632
rect 21272 4548 21324 4554
rect 21272 4490 21324 4496
rect 20996 4072 21048 4078
rect 20996 4014 21048 4020
rect 21180 4072 21232 4078
rect 21180 4014 21232 4020
rect 21008 3670 21036 4014
rect 20996 3664 21048 3670
rect 20996 3606 21048 3612
rect 21284 3618 21312 4490
rect 21376 4282 21404 4626
rect 21364 4276 21416 4282
rect 21364 4218 21416 4224
rect 22296 4078 22324 4814
rect 22100 4072 22152 4078
rect 22098 4040 22100 4049
rect 22284 4072 22336 4078
rect 22152 4040 22154 4049
rect 23492 4049 23520 5510
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24214 4584 24270 4593
rect 24214 4519 24270 4528
rect 22284 4014 22336 4020
rect 23478 4040 23534 4049
rect 22098 3975 22154 3984
rect 22376 4004 22428 4010
rect 23478 3975 23534 3984
rect 22376 3946 22428 3952
rect 22100 3936 22152 3942
rect 22100 3878 22152 3884
rect 21284 3590 21404 3618
rect 22112 3602 22140 3878
rect 21272 3392 21324 3398
rect 21272 3334 21324 3340
rect 21284 2961 21312 3334
rect 21270 2952 21326 2961
rect 21270 2887 21326 2896
rect 21376 480 21404 3590
rect 22100 3596 22152 3602
rect 22100 3538 22152 3544
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 21468 2650 21496 3470
rect 21916 3392 21968 3398
rect 21916 3334 21968 3340
rect 21638 3088 21694 3097
rect 21638 3023 21694 3032
rect 21652 2990 21680 3023
rect 21640 2984 21692 2990
rect 21640 2926 21692 2932
rect 21824 2848 21876 2854
rect 21822 2816 21824 2825
rect 21876 2816 21878 2825
rect 21822 2751 21878 2760
rect 21456 2644 21508 2650
rect 21456 2586 21508 2592
rect 21928 480 21956 3334
rect 22192 2508 22244 2514
rect 22192 2450 22244 2456
rect 22204 2281 22232 2450
rect 22190 2272 22246 2281
rect 22190 2207 22246 2216
rect 22388 1442 22416 3946
rect 24228 3641 24256 4519
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 25318 4040 25374 4049
rect 25318 3975 25374 3984
rect 23662 3632 23718 3641
rect 22560 3596 22612 3602
rect 23662 3567 23718 3576
rect 24214 3632 24270 3641
rect 24214 3567 24270 3576
rect 22560 3538 22612 3544
rect 22572 3194 22600 3538
rect 22560 3188 22612 3194
rect 22560 3130 22612 3136
rect 23676 2990 23704 3567
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 23846 3224 23902 3233
rect 24289 3216 24585 3236
rect 23846 3159 23848 3168
rect 23900 3159 23902 3168
rect 23848 3130 23900 3136
rect 23664 2984 23716 2990
rect 23110 2952 23166 2961
rect 23664 2926 23716 2932
rect 23110 2887 23166 2896
rect 22388 1414 22508 1442
rect 22480 480 22508 1414
rect 23124 480 23152 2887
rect 23662 2816 23718 2825
rect 23662 2751 23718 2760
rect 23676 480 23704 2751
rect 24030 2544 24086 2553
rect 24030 2479 24032 2488
rect 24084 2479 24086 2488
rect 24032 2450 24084 2456
rect 24766 2408 24822 2417
rect 24766 2343 24822 2352
rect 24124 2304 24176 2310
rect 24124 2246 24176 2252
rect 24216 2304 24268 2310
rect 24216 2246 24268 2252
rect 24136 1170 24164 2246
rect 24228 1465 24256 2246
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24214 1456 24270 1465
rect 24214 1391 24270 1400
rect 24136 1142 24256 1170
rect 24228 480 24256 1142
rect 24780 480 24808 2343
rect 25332 480 25360 3975
rect 26514 3632 26570 3641
rect 26514 3567 26570 3576
rect 25962 1592 26018 1601
rect 25962 1527 26018 1536
rect 25976 480 26004 1527
rect 26528 480 26556 3567
rect 27066 2000 27122 2009
rect 27066 1935 27122 1944
rect 27080 480 27108 1935
rect 27618 1728 27674 1737
rect 27618 1663 27674 1672
rect 27632 480 27660 1663
rect 6274 368 6330 377
rect 6274 303 6330 312
rect 6550 0 6606 480
rect 7102 0 7158 480
rect 7654 0 7710 480
rect 8206 0 8262 480
rect 8850 0 8906 480
rect 9402 0 9458 480
rect 9954 0 10010 480
rect 10506 0 10562 480
rect 11058 0 11114 480
rect 11702 0 11758 480
rect 12254 0 12310 480
rect 12806 0 12862 480
rect 13358 0 13414 480
rect 13910 0 13966 480
rect 14554 0 14610 480
rect 15106 0 15162 480
rect 15658 0 15714 480
rect 16210 0 16266 480
rect 16762 0 16818 480
rect 17406 0 17462 480
rect 17958 0 18014 480
rect 18510 0 18566 480
rect 19062 0 19118 480
rect 19614 0 19670 480
rect 20258 0 20314 480
rect 20810 0 20866 480
rect 21362 0 21418 480
rect 21914 0 21970 480
rect 22466 0 22522 480
rect 23110 0 23166 480
rect 23662 0 23718 480
rect 24214 0 24270 480
rect 24766 0 24822 480
rect 25318 0 25374 480
rect 25962 0 26018 480
rect 26514 0 26570 480
rect 27066 0 27122 480
rect 27618 0 27674 480
<< via2 >>
rect 2778 27648 2834 27704
rect 2042 24812 2098 24848
rect 2042 24792 2044 24812
rect 2044 24792 2096 24812
rect 2096 24792 2098 24812
rect 846 20168 902 20224
rect 570 19896 626 19952
rect 1950 24656 2006 24712
rect 2134 23160 2190 23216
rect 1582 21800 1638 21856
rect 1398 21256 1454 21312
rect 1398 21004 1454 21040
rect 1398 20984 1400 21004
rect 1400 20984 1452 21004
rect 1452 20984 1454 21004
rect 2318 22344 2374 22400
rect 1398 18944 1454 19000
rect 1582 18400 1638 18456
rect 1490 17176 1546 17232
rect 1398 16632 1454 16688
rect 1582 15952 1638 16008
rect 1490 14864 1546 14920
rect 1398 14728 1454 14784
rect 1398 13388 1454 13424
rect 1398 13368 1400 13388
rect 1400 13368 1452 13388
rect 1452 13368 1454 13388
rect 3054 25336 3110 25392
rect 1950 20984 2006 21040
rect 2410 20440 2466 20496
rect 2042 18808 2098 18864
rect 2042 17856 2098 17912
rect 1950 17176 2006 17232
rect 1674 13640 1730 13696
rect 2042 15564 2098 15600
rect 2042 15544 2044 15564
rect 2044 15544 2096 15564
rect 2096 15544 2098 15564
rect 1582 13096 1638 13152
rect 1582 12552 1638 12608
rect 1858 10532 1914 10568
rect 1858 10512 1860 10532
rect 1860 10512 1912 10532
rect 1912 10512 1914 10532
rect 1398 9988 1454 10024
rect 1398 9968 1400 9988
rect 1400 9968 1452 9988
rect 1452 9968 1454 9988
rect 570 7792 626 7848
rect 1674 9596 1676 9616
rect 1676 9596 1728 9616
rect 1728 9596 1730 9616
rect 1674 9560 1730 9596
rect 846 4256 902 4312
rect 294 3440 350 3496
rect 2870 23024 2926 23080
rect 3606 26560 3662 26616
rect 2962 22480 3018 22536
rect 2870 20324 2926 20360
rect 2870 20304 2872 20324
rect 2872 20304 2924 20324
rect 2924 20304 2926 20324
rect 2686 19624 2742 19680
rect 2686 19488 2742 19544
rect 3422 21392 3478 21448
rect 3054 19780 3110 19816
rect 3054 19760 3056 19780
rect 3056 19760 3108 19780
rect 3108 19760 3110 19780
rect 3238 19116 3240 19136
rect 3240 19116 3292 19136
rect 3292 19116 3294 19136
rect 3238 19080 3294 19116
rect 3146 18944 3202 19000
rect 2686 17720 2742 17776
rect 3330 18264 3386 18320
rect 2778 15408 2834 15464
rect 2410 13640 2466 13696
rect 2226 11464 2282 11520
rect 2134 11056 2190 11112
rect 2410 11600 2466 11656
rect 2594 14048 2650 14104
rect 2870 15020 2926 15056
rect 2870 15000 2872 15020
rect 2872 15000 2924 15020
rect 2924 15000 2926 15020
rect 2870 14864 2926 14920
rect 3054 14048 3110 14104
rect 2962 13776 3018 13832
rect 2778 11212 2834 11248
rect 2778 11192 2780 11212
rect 2780 11192 2832 11212
rect 2832 11192 2834 11212
rect 1582 5752 1638 5808
rect 1490 4936 1546 4992
rect 1398 4120 1454 4176
rect 2226 5616 2282 5672
rect 2410 4548 2466 4584
rect 2410 4528 2412 4548
rect 2412 4528 2464 4548
rect 2464 4528 2466 4548
rect 2502 3984 2558 4040
rect 1490 3576 1546 3632
rect 2042 1808 2098 1864
rect 1950 1536 2006 1592
rect 1766 992 1822 1048
rect 2410 3304 2466 3360
rect 2318 1128 2374 1184
rect 3606 24112 3662 24168
rect 3330 15000 3386 15056
rect 3606 14728 3662 14784
rect 4066 25880 4122 25936
rect 3790 24520 3846 24576
rect 3974 23588 4030 23624
rect 3974 23568 3976 23588
rect 3976 23568 4028 23588
rect 4028 23568 4030 23588
rect 3790 22480 3846 22536
rect 4066 22888 4122 22944
rect 3790 21936 3846 21992
rect 4710 27104 4766 27160
rect 4342 23704 4398 23760
rect 4526 23568 4582 23624
rect 4342 22888 4398 22944
rect 4066 20712 4122 20768
rect 3606 13812 3608 13832
rect 3608 13812 3660 13832
rect 3660 13812 3662 13832
rect 3606 13776 3662 13812
rect 3422 13504 3478 13560
rect 3146 11736 3202 11792
rect 3054 10104 3110 10160
rect 3514 12180 3516 12200
rect 3516 12180 3568 12200
rect 3568 12180 3570 12200
rect 3514 12144 3570 12180
rect 3422 11500 3424 11520
rect 3424 11500 3476 11520
rect 3476 11500 3478 11520
rect 3422 11464 3478 11500
rect 3514 10784 3570 10840
rect 3422 10376 3478 10432
rect 3422 10104 3478 10160
rect 3054 9152 3110 9208
rect 3238 9424 3294 9480
rect 3238 9016 3294 9072
rect 3146 8608 3202 8664
rect 2962 7540 3018 7576
rect 2962 7520 2964 7540
rect 2964 7520 3016 7540
rect 3016 7520 3018 7540
rect 3606 10240 3662 10296
rect 4250 17856 4306 17912
rect 4066 15408 4122 15464
rect 3974 15136 4030 15192
rect 4158 14320 4214 14376
rect 4066 13776 4122 13832
rect 3974 13368 4030 13424
rect 4618 21972 4620 21992
rect 4620 21972 4672 21992
rect 4672 21972 4674 21992
rect 4618 21936 4674 21972
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5262 23432 5318 23488
rect 4526 19624 4582 19680
rect 4618 18264 4674 18320
rect 4434 12688 4490 12744
rect 4250 11872 4306 11928
rect 3974 11328 4030 11384
rect 3974 10648 4030 10704
rect 3514 8336 3570 8392
rect 2778 5616 2834 5672
rect 2778 4700 2780 4720
rect 2780 4700 2832 4720
rect 2832 4700 2834 4720
rect 2778 4664 2834 4700
rect 2686 3884 2688 3904
rect 2688 3884 2740 3904
rect 2740 3884 2742 3904
rect 2686 3848 2742 3884
rect 3422 6976 3478 7032
rect 2962 5616 3018 5672
rect 3974 6704 4030 6760
rect 4066 6024 4122 6080
rect 4342 6296 4398 6352
rect 3606 4800 3662 4856
rect 3422 3712 3478 3768
rect 3606 3732 3662 3768
rect 3606 3712 3608 3732
rect 3608 3712 3660 3732
rect 3660 3712 3662 3732
rect 2870 2896 2926 2952
rect 3146 3168 3202 3224
rect 3882 4972 3884 4992
rect 3884 4972 3936 4992
rect 3936 4972 3938 4992
rect 3882 4936 3938 4972
rect 4158 5108 4160 5128
rect 4160 5108 4212 5128
rect 4212 5108 4214 5128
rect 4158 5072 4214 5108
rect 4066 4392 4122 4448
rect 4158 3984 4214 4040
rect 3790 2760 3846 2816
rect 2962 1400 3018 1456
rect 2778 856 2834 912
rect 3330 1536 3386 1592
rect 4526 11736 4582 11792
rect 4618 11092 4620 11112
rect 4620 11092 4672 11112
rect 4672 11092 4674 11112
rect 4618 11056 4674 11092
rect 4526 7112 4582 7168
rect 4250 3032 4306 3088
rect 4618 3848 4674 3904
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5998 23296 6054 23352
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5538 22616 5594 22672
rect 5262 22072 5318 22128
rect 4894 12824 4950 12880
rect 5170 14728 5226 14784
rect 4894 11076 4950 11112
rect 4894 11056 4896 11076
rect 4896 11056 4948 11076
rect 4948 11056 4950 11076
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 6550 24656 6606 24712
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 6182 19216 6238 19272
rect 5998 19080 6054 19136
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5630 17212 5632 17232
rect 5632 17212 5684 17232
rect 5684 17212 5686 17232
rect 5630 17176 5686 17212
rect 5538 16652 5594 16688
rect 5538 16632 5540 16652
rect 5540 16632 5592 16652
rect 5592 16632 5594 16652
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 6090 16532 6092 16552
rect 6092 16532 6144 16552
rect 6144 16532 6146 16552
rect 6090 16496 6146 16532
rect 5446 15136 5502 15192
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 6090 15272 6146 15328
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 6182 14864 6238 14920
rect 5538 13640 5594 13696
rect 6366 22500 6422 22536
rect 6366 22480 6368 22500
rect 6368 22480 6420 22500
rect 6420 22480 6422 22500
rect 7470 23432 7526 23488
rect 7010 20984 7066 21040
rect 6918 20712 6974 20768
rect 7194 20304 7250 20360
rect 6550 18672 6606 18728
rect 6458 15136 6514 15192
rect 6366 15000 6422 15056
rect 6642 16088 6698 16144
rect 6366 13388 6422 13424
rect 6366 13368 6368 13388
rect 6368 13368 6420 13388
rect 6420 13368 6422 13388
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5630 12416 5686 12472
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 4986 8472 5042 8528
rect 5998 10240 6054 10296
rect 5998 9832 6054 9888
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5170 7520 5226 7576
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5538 6840 5594 6896
rect 6090 7520 6146 7576
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 6458 11736 6514 11792
rect 7010 16496 7066 16552
rect 6826 15408 6882 15464
rect 6826 13504 6882 13560
rect 4894 3340 4896 3360
rect 4896 3340 4948 3360
rect 4948 3340 4950 3360
rect 4894 3304 4950 3340
rect 4066 1944 4122 2000
rect 4066 1672 4122 1728
rect 4158 1264 4214 1320
rect 3238 720 3294 776
rect 5262 2488 5318 2544
rect 5998 4820 6054 4856
rect 5998 4800 6000 4820
rect 6000 4800 6052 4820
rect 6052 4800 6054 4820
rect 5446 4256 5502 4312
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 6550 5480 6606 5536
rect 5538 3712 5594 3768
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5446 3032 5502 3088
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6274 5072 6330 5128
rect 6182 2796 6184 2816
rect 6184 2796 6236 2816
rect 6236 2796 6238 2816
rect 6182 2760 6238 2796
rect 6826 7248 6882 7304
rect 6642 4800 6698 4856
rect 6642 3440 6698 3496
rect 7286 19352 7342 19408
rect 7562 17448 7618 17504
rect 7470 16088 7526 16144
rect 8022 23704 8078 23760
rect 7838 22208 7894 22264
rect 8850 23296 8906 23352
rect 8390 22652 8392 22672
rect 8392 22652 8444 22672
rect 8444 22652 8446 22672
rect 8390 22616 8446 22652
rect 8758 21936 8814 21992
rect 8114 21664 8170 21720
rect 8022 20032 8078 20088
rect 8022 18964 8078 19000
rect 8022 18944 8024 18964
rect 8024 18944 8076 18964
rect 8076 18944 8078 18964
rect 7930 18536 7986 18592
rect 7194 15136 7250 15192
rect 7194 15000 7250 15056
rect 7102 13912 7158 13968
rect 7194 12280 7250 12336
rect 7194 6296 7250 6352
rect 7286 5888 7342 5944
rect 7562 4276 7618 4312
rect 7562 4256 7564 4276
rect 7564 4256 7616 4276
rect 7616 4256 7618 4276
rect 7102 3848 7158 3904
rect 6734 2760 6790 2816
rect 6918 2488 6974 2544
rect 7194 3596 7250 3632
rect 7194 3576 7196 3596
rect 7196 3576 7248 3596
rect 7248 3576 7250 3596
rect 7286 2916 7342 2952
rect 7286 2896 7288 2916
rect 7288 2896 7340 2916
rect 7340 2896 7342 2916
rect 7286 2252 7288 2272
rect 7288 2252 7340 2272
rect 7340 2252 7342 2272
rect 7286 2216 7342 2252
rect 7930 14048 7986 14104
rect 7930 9424 7986 9480
rect 8482 19896 8538 19952
rect 8298 19352 8354 19408
rect 8206 18944 8262 19000
rect 8574 18808 8630 18864
rect 8850 21412 8906 21448
rect 8850 21392 8852 21412
rect 8852 21392 8904 21412
rect 8904 21392 8906 21412
rect 8850 20168 8906 20224
rect 8850 13812 8852 13832
rect 8852 13812 8904 13832
rect 8904 13812 8906 13832
rect 8850 13776 8906 13812
rect 9586 23568 9642 23624
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 11058 24792 11114 24848
rect 10782 24656 10838 24712
rect 10690 23976 10746 24032
rect 9586 23024 9642 23080
rect 9402 22480 9458 22536
rect 9402 18672 9458 18728
rect 9494 17620 9496 17640
rect 9496 17620 9548 17640
rect 9548 17620 9550 17640
rect 9494 17584 9550 17620
rect 9126 15136 9182 15192
rect 9126 14048 9182 14104
rect 9218 13912 9274 13968
rect 8574 13504 8630 13560
rect 8574 13232 8630 13288
rect 8482 13096 8538 13152
rect 8390 10920 8446 10976
rect 9402 12960 9458 13016
rect 8942 11736 8998 11792
rect 8850 10920 8906 10976
rect 8390 9424 8446 9480
rect 8022 9288 8078 9344
rect 8022 9016 8078 9072
rect 7930 6024 7986 6080
rect 7838 5480 7894 5536
rect 7746 4392 7802 4448
rect 8390 7520 8446 7576
rect 8482 6860 8538 6896
rect 8482 6840 8484 6860
rect 8484 6840 8536 6860
rect 8536 6840 8538 6860
rect 8390 6704 8446 6760
rect 8298 5772 8354 5808
rect 8298 5752 8300 5772
rect 8300 5752 8352 5772
rect 8352 5752 8354 5772
rect 8574 5208 8630 5264
rect 8022 3984 8078 4040
rect 8022 1400 8078 1456
rect 7746 1264 7802 1320
rect 7930 1264 7986 1320
rect 7746 992 7802 1048
rect 7930 720 7986 776
rect 8574 4020 8576 4040
rect 8576 4020 8628 4040
rect 8628 4020 8630 4040
rect 8574 3984 8630 4020
rect 8298 3440 8354 3496
rect 8482 3304 8538 3360
rect 8850 4120 8906 4176
rect 9494 12416 9550 12472
rect 9402 12008 9458 12064
rect 9678 16632 9734 16688
rect 9678 12280 9734 12336
rect 9862 22208 9918 22264
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 11426 23568 11482 23624
rect 10874 22092 10930 22128
rect 10874 22072 10876 22092
rect 10876 22072 10928 22092
rect 10928 22072 10930 22092
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10138 18536 10194 18592
rect 9954 17756 9956 17776
rect 9956 17756 10008 17776
rect 10008 17756 10010 17776
rect 9954 17720 10010 17756
rect 10046 17076 10048 17096
rect 10048 17076 10100 17096
rect 10100 17076 10102 17096
rect 10046 17040 10102 17076
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10322 17604 10378 17640
rect 10322 17584 10324 17604
rect 10324 17584 10376 17604
rect 10376 17584 10378 17604
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10966 21564 10968 21584
rect 10968 21564 11020 21584
rect 11020 21564 11022 21584
rect 10966 21528 11022 21564
rect 11242 21664 11298 21720
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10046 15428 10102 15464
rect 10046 15408 10048 15428
rect 10048 15408 10100 15428
rect 10100 15408 10102 15428
rect 10046 15272 10102 15328
rect 10782 15544 10838 15600
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10322 11056 10378 11112
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 9586 7792 9642 7848
rect 9862 8472 9918 8528
rect 9494 7656 9550 7712
rect 9034 5636 9090 5672
rect 9034 5616 9036 5636
rect 9036 5616 9088 5636
rect 9088 5616 9090 5636
rect 9678 7112 9734 7168
rect 9770 6976 9826 7032
rect 9586 5480 9642 5536
rect 9310 4800 9366 4856
rect 9310 4256 9366 4312
rect 9310 3984 9366 4040
rect 8758 3576 8814 3632
rect 8482 1672 8538 1728
rect 8666 1672 8722 1728
rect 9218 3848 9274 3904
rect 8942 1536 8998 1592
rect 9494 3732 9550 3768
rect 9494 3712 9496 3732
rect 9496 3712 9548 3732
rect 9548 3712 9550 3732
rect 9862 6160 9918 6216
rect 9862 5888 9918 5944
rect 10230 9696 10286 9752
rect 10230 9560 10286 9616
rect 10138 9288 10194 9344
rect 10046 9152 10102 9208
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10046 9036 10102 9072
rect 10046 9016 10048 9036
rect 10048 9016 10100 9036
rect 10100 9016 10102 9036
rect 10138 8880 10194 8936
rect 10046 8472 10102 8528
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 11794 18808 11850 18864
rect 12254 24132 12310 24168
rect 12254 24112 12256 24132
rect 12256 24112 12308 24132
rect 12308 24112 12310 24132
rect 12254 23976 12310 24032
rect 12162 22516 12164 22536
rect 12164 22516 12216 22536
rect 12216 22516 12218 22536
rect 12162 22480 12218 22516
rect 12622 23860 12678 23896
rect 12622 23840 12624 23860
rect 12624 23840 12676 23860
rect 12676 23840 12678 23860
rect 12346 21800 12402 21856
rect 12898 22652 12900 22672
rect 12900 22652 12952 22672
rect 12952 22652 12954 22672
rect 12898 22616 12954 22652
rect 14278 24404 14334 24440
rect 14278 24384 14280 24404
rect 14280 24384 14332 24404
rect 14332 24384 14334 24404
rect 14002 23740 14004 23760
rect 14004 23740 14056 23760
rect 14056 23740 14058 23760
rect 14002 23704 14058 23740
rect 14278 22480 14334 22536
rect 12898 22072 12954 22128
rect 12806 21528 12862 21584
rect 12806 20848 12862 20904
rect 12346 20440 12402 20496
rect 12254 19896 12310 19952
rect 12622 19760 12678 19816
rect 12254 19216 12310 19272
rect 11978 18536 12034 18592
rect 13542 22072 13598 22128
rect 13634 21972 13636 21992
rect 13636 21972 13688 21992
rect 13688 21972 13690 21992
rect 13634 21936 13690 21972
rect 14278 22208 14334 22264
rect 13082 21412 13138 21448
rect 13082 21392 13084 21412
rect 13084 21392 13136 21412
rect 13136 21392 13138 21412
rect 13450 20848 13506 20904
rect 14002 22072 14058 22128
rect 14002 20712 14058 20768
rect 14186 19760 14242 19816
rect 13910 19080 13966 19136
rect 11426 15544 11482 15600
rect 11058 13404 11060 13424
rect 11060 13404 11112 13424
rect 11112 13404 11114 13424
rect 11058 13368 11114 13404
rect 11150 11620 11206 11656
rect 11150 11600 11152 11620
rect 11152 11600 11204 11620
rect 11204 11600 11206 11620
rect 11426 12824 11482 12880
rect 10874 9696 10930 9752
rect 10690 7384 10746 7440
rect 10046 6160 10102 6216
rect 9954 5344 10010 5400
rect 10046 4684 10102 4720
rect 10046 4664 10048 4684
rect 10048 4664 10100 4684
rect 10100 4664 10102 4684
rect 10690 7112 10746 7168
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10966 7404 11022 7440
rect 10966 7384 10968 7404
rect 10968 7384 11020 7404
rect 11020 7384 11022 7404
rect 10230 6296 10286 6352
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10506 4700 10508 4720
rect 10508 4700 10560 4720
rect 10560 4700 10562 4720
rect 10506 4664 10562 4700
rect 9954 4528 10010 4584
rect 9770 3576 9826 3632
rect 10046 3984 10102 4040
rect 9954 2760 10010 2816
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10966 6024 11022 6080
rect 10138 2080 10194 2136
rect 11242 5616 11298 5672
rect 11058 3984 11114 4040
rect 11242 4004 11298 4040
rect 11242 3984 11244 4004
rect 11244 3984 11296 4004
rect 11296 3984 11298 4004
rect 11242 3848 11298 3904
rect 11242 3032 11298 3088
rect 11426 2796 11428 2816
rect 11428 2796 11480 2816
rect 11480 2796 11482 2816
rect 11426 2760 11482 2796
rect 11702 12300 11758 12336
rect 11702 12280 11704 12300
rect 11704 12280 11756 12300
rect 11756 12280 11758 12300
rect 11610 12008 11666 12064
rect 12806 15700 12862 15736
rect 12806 15680 12808 15700
rect 12808 15680 12860 15700
rect 12860 15680 12862 15700
rect 11886 12960 11942 13016
rect 11886 12552 11942 12608
rect 11794 9696 11850 9752
rect 11978 9424 12034 9480
rect 11886 8472 11942 8528
rect 12714 13776 12770 13832
rect 12806 13232 12862 13288
rect 12806 10784 12862 10840
rect 12806 9696 12862 9752
rect 12438 8200 12494 8256
rect 11978 2488 12034 2544
rect 12162 2488 12218 2544
rect 11610 2372 11666 2408
rect 11610 2352 11612 2372
rect 11612 2352 11664 2372
rect 11664 2352 11666 2372
rect 12162 1672 12218 1728
rect 12806 6724 12862 6760
rect 12806 6704 12808 6724
rect 12808 6704 12860 6724
rect 12860 6704 12862 6724
rect 13358 17176 13414 17232
rect 13082 16632 13138 16688
rect 13358 12416 13414 12472
rect 13818 18264 13874 18320
rect 13726 12688 13782 12744
rect 14094 14456 14150 14512
rect 13266 11348 13322 11384
rect 13266 11328 13268 11348
rect 13268 11328 13320 11348
rect 13320 11328 13322 11348
rect 12990 10784 13046 10840
rect 12990 10648 13046 10704
rect 13174 10648 13230 10704
rect 12990 10240 13046 10296
rect 12990 8472 13046 8528
rect 13174 7656 13230 7712
rect 12990 6296 13046 6352
rect 12898 6060 12900 6080
rect 12900 6060 12952 6080
rect 12952 6060 12954 6080
rect 12898 6024 12954 6060
rect 13174 4800 13230 4856
rect 12990 4392 13046 4448
rect 13174 4120 13230 4176
rect 13450 5752 13506 5808
rect 13634 12416 13690 12472
rect 14278 15000 14334 15056
rect 14278 14456 14334 14512
rect 14554 19352 14610 19408
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 15474 24248 15530 24304
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 15106 23740 15108 23760
rect 15108 23740 15160 23760
rect 15160 23740 15162 23760
rect 15106 23704 15162 23740
rect 16118 24792 16174 24848
rect 16762 24656 16818 24712
rect 17958 24792 18014 24848
rect 18142 24792 18198 24848
rect 16210 24384 16266 24440
rect 16394 24384 16450 24440
rect 17406 24384 17462 24440
rect 17774 24384 17830 24440
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14738 13912 14794 13968
rect 14554 13096 14610 13152
rect 14646 12824 14702 12880
rect 14278 11600 14334 11656
rect 13910 11228 13912 11248
rect 13912 11228 13964 11248
rect 13964 11228 13966 11248
rect 13910 11192 13966 11228
rect 13818 10548 13820 10568
rect 13820 10548 13872 10568
rect 13872 10548 13874 10568
rect 13818 10512 13874 10548
rect 13818 10376 13874 10432
rect 13910 9968 13966 10024
rect 14370 10376 14426 10432
rect 14186 10140 14188 10160
rect 14188 10140 14240 10160
rect 14240 10140 14242 10160
rect 14186 10104 14242 10140
rect 14278 8472 14334 8528
rect 13634 5888 13690 5944
rect 13634 4120 13690 4176
rect 13910 5616 13966 5672
rect 13542 2624 13598 2680
rect 14738 11872 14794 11928
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 15474 22924 15476 22944
rect 15476 22924 15528 22944
rect 15528 22924 15530 22944
rect 15474 22888 15530 22924
rect 17038 23976 17094 24032
rect 18878 24656 18934 24712
rect 18142 24112 18198 24168
rect 18234 23860 18290 23896
rect 18234 23840 18236 23860
rect 18236 23840 18288 23860
rect 18288 23840 18290 23860
rect 17222 23432 17278 23488
rect 17038 23024 17094 23080
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 16670 21956 16726 21992
rect 16670 21936 16672 21956
rect 16672 21936 16724 21956
rect 16724 21936 16726 21956
rect 15750 19896 15806 19952
rect 15474 19352 15530 19408
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 15658 17312 15714 17368
rect 17314 18672 17370 18728
rect 16210 17720 16266 17776
rect 16026 17040 16082 17096
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 15934 16632 15990 16688
rect 15290 15680 15346 15736
rect 15106 15544 15162 15600
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14646 11464 14702 11520
rect 14738 11192 14794 11248
rect 14554 9868 14556 9888
rect 14556 9868 14608 9888
rect 14608 9868 14610 9888
rect 14554 9832 14610 9868
rect 14554 8916 14556 8936
rect 14556 8916 14608 8936
rect 14608 8916 14610 8936
rect 14554 8880 14610 8916
rect 14278 6024 14334 6080
rect 14186 4936 14242 4992
rect 14370 3576 14426 3632
rect 14186 3168 14242 3224
rect 14646 6976 14702 7032
rect 14554 3168 14610 3224
rect 14922 11348 14978 11384
rect 14922 11328 14924 11348
rect 14924 11328 14976 11348
rect 14976 11328 14978 11348
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14922 9052 14924 9072
rect 14924 9052 14976 9072
rect 14976 9052 14978 9072
rect 14922 9016 14978 9052
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 15290 7792 15346 7848
rect 15474 7792 15530 7848
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 15198 5616 15254 5672
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15382 5516 15384 5536
rect 15384 5516 15436 5536
rect 15436 5516 15438 5536
rect 15382 5480 15438 5516
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15474 4548 15530 4584
rect 15474 4528 15476 4548
rect 15476 4528 15528 4548
rect 15528 4528 15530 4548
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14462 2216 14518 2272
rect 14370 1844 14372 1864
rect 14372 1844 14424 1864
rect 14424 1844 14426 1864
rect 14370 1808 14426 1844
rect 14738 2508 14794 2544
rect 14738 2488 14740 2508
rect 14740 2488 14792 2508
rect 14792 2488 14794 2508
rect 14922 2488 14978 2544
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 14646 1980 14648 2000
rect 14648 1980 14700 2000
rect 14700 1980 14702 2000
rect 14646 1944 14702 1980
rect 15474 2080 15530 2136
rect 15290 1536 15346 1592
rect 15750 12300 15806 12336
rect 15750 12280 15752 12300
rect 15752 12280 15804 12300
rect 15804 12280 15806 12300
rect 15658 11076 15714 11112
rect 15658 11056 15660 11076
rect 15660 11056 15712 11076
rect 15712 11056 15714 11076
rect 17130 16496 17186 16552
rect 16210 15136 16266 15192
rect 15934 10648 15990 10704
rect 15934 8372 15936 8392
rect 15936 8372 15988 8392
rect 15988 8372 15990 8392
rect 15934 8336 15990 8372
rect 15658 5108 15660 5128
rect 15660 5108 15712 5128
rect 15712 5108 15714 5128
rect 15658 5072 15714 5108
rect 17038 12300 17094 12336
rect 17038 12280 17040 12300
rect 17040 12280 17092 12300
rect 17092 12280 17094 12300
rect 16762 11464 16818 11520
rect 16946 11192 17002 11248
rect 16302 9596 16304 9616
rect 16304 9596 16356 9616
rect 16356 9596 16358 9616
rect 16302 9560 16358 9596
rect 17222 16088 17278 16144
rect 17038 9968 17094 10024
rect 15842 5636 15898 5672
rect 15842 5616 15844 5636
rect 15844 5616 15896 5636
rect 15896 5616 15898 5636
rect 16026 4800 16082 4856
rect 16854 6196 16856 6216
rect 16856 6196 16908 6216
rect 16908 6196 16910 6216
rect 16854 6160 16910 6196
rect 16394 4972 16396 4992
rect 16396 4972 16448 4992
rect 16448 4972 16450 4992
rect 16394 4936 16450 4972
rect 16946 5480 17002 5536
rect 16854 5092 16910 5128
rect 16854 5072 16856 5092
rect 16856 5072 16908 5092
rect 16908 5072 16910 5092
rect 17038 4392 17094 4448
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19430 24384 19486 24440
rect 19706 23976 19762 24032
rect 20810 24656 20866 24712
rect 20258 23840 20314 23896
rect 17590 21392 17646 21448
rect 17498 19080 17554 19136
rect 17406 17584 17462 17640
rect 17314 12280 17370 12336
rect 17406 10412 17408 10432
rect 17408 10412 17460 10432
rect 17460 10412 17462 10432
rect 17406 10376 17462 10412
rect 16762 2760 16818 2816
rect 16670 2488 16726 2544
rect 16670 1944 16726 2000
rect 17130 2624 17186 2680
rect 17406 5364 17462 5400
rect 17406 5344 17408 5364
rect 17408 5344 17460 5364
rect 17460 5344 17462 5364
rect 18234 17176 18290 17232
rect 18326 13368 18382 13424
rect 18050 11328 18106 11384
rect 18050 10260 18106 10296
rect 18050 10240 18052 10260
rect 18052 10240 18104 10260
rect 18104 10240 18106 10260
rect 17958 8472 18014 8528
rect 19062 23432 19118 23488
rect 19338 22516 19340 22536
rect 19340 22516 19392 22536
rect 19392 22516 19394 22536
rect 19338 22480 19394 22516
rect 21362 23976 21418 24032
rect 21362 23860 21418 23896
rect 21362 23840 21364 23860
rect 21364 23840 21416 23860
rect 21416 23840 21418 23860
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19430 19760 19486 19816
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 20902 23180 20958 23216
rect 20902 23160 20904 23180
rect 20904 23160 20956 23180
rect 20956 23160 20958 23180
rect 23110 23840 23166 23896
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24214 24792 24270 24848
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 23662 23568 23718 23624
rect 23570 23296 23626 23352
rect 21914 22888 21970 22944
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 26514 24248 26570 24304
rect 25962 24112 26018 24168
rect 27066 23704 27122 23760
rect 24766 22616 24822 22672
rect 23570 21936 23626 21992
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 27618 18672 27674 18728
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 20810 17312 20866 17368
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 18602 16496 18658 16552
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 19338 15136 19394 15192
rect 18970 11056 19026 11112
rect 19522 15000 19578 15056
rect 19430 12588 19432 12608
rect 19432 12588 19484 12608
rect 19484 12588 19486 12608
rect 19430 12552 19486 12588
rect 18878 9560 18934 9616
rect 19338 9560 19394 9616
rect 18418 8200 18474 8256
rect 18510 7404 18566 7440
rect 18510 7384 18512 7404
rect 18512 7384 18564 7404
rect 18564 7384 18566 7404
rect 18326 7112 18382 7168
rect 18050 6432 18106 6488
rect 18234 6024 18290 6080
rect 17958 5616 18014 5672
rect 17774 5228 17830 5264
rect 17774 5208 17776 5228
rect 17776 5208 17828 5228
rect 17828 5208 17830 5228
rect 17498 4684 17554 4720
rect 17498 4664 17500 4684
rect 17500 4664 17552 4684
rect 17552 4664 17554 4684
rect 17406 2896 17462 2952
rect 17774 3032 17830 3088
rect 17314 1400 17370 1456
rect 17222 1264 17278 1320
rect 18326 5752 18382 5808
rect 18050 3984 18106 4040
rect 18602 6296 18658 6352
rect 18510 5208 18566 5264
rect 19246 7112 19302 7168
rect 19338 6976 19394 7032
rect 19430 6332 19432 6352
rect 19432 6332 19484 6352
rect 19484 6332 19486 6352
rect 19430 6296 19486 6332
rect 19430 5888 19486 5944
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19062 4392 19118 4448
rect 18970 4120 19026 4176
rect 18786 3848 18842 3904
rect 18510 3168 18566 3224
rect 18970 2488 19026 2544
rect 18970 1944 19026 2000
rect 18970 1672 19026 1728
rect 18878 1536 18934 1592
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19338 4256 19394 4312
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 22282 7248 22338 7304
rect 22190 6704 22246 6760
rect 20902 6432 20958 6488
rect 21178 4664 21234 4720
rect 21638 5344 21694 5400
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 22374 5244 22376 5264
rect 22376 5244 22428 5264
rect 22428 5244 22430 5264
rect 22374 5208 22430 5244
rect 22742 5108 22744 5128
rect 22744 5108 22796 5128
rect 22796 5108 22798 5128
rect 22742 5072 22798 5108
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19154 3460 19210 3496
rect 19154 3440 19156 3460
rect 19156 3440 19208 3460
rect 19208 3440 19210 3460
rect 19430 1128 19486 1184
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20074 1536 20130 1592
rect 19614 1400 19670 1456
rect 19522 856 19578 912
rect 20258 1400 20314 1456
rect 20166 992 20222 1048
rect 21638 4664 21694 4720
rect 22098 4020 22100 4040
rect 22100 4020 22152 4040
rect 22152 4020 22154 4040
rect 22098 3984 22154 4020
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24214 4528 24270 4584
rect 23478 3984 23534 4040
rect 21270 2896 21326 2952
rect 21638 3032 21694 3088
rect 21822 2796 21824 2816
rect 21824 2796 21876 2816
rect 21876 2796 21878 2816
rect 21822 2760 21878 2796
rect 22190 2216 22246 2272
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 25318 3984 25374 4040
rect 23662 3576 23718 3632
rect 24214 3576 24270 3632
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 23846 3188 23902 3224
rect 23846 3168 23848 3188
rect 23848 3168 23900 3188
rect 23900 3168 23902 3188
rect 23110 2896 23166 2952
rect 23662 2760 23718 2816
rect 24030 2508 24086 2544
rect 24030 2488 24032 2508
rect 24032 2488 24084 2508
rect 24084 2488 24086 2508
rect 24766 2352 24822 2408
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 24214 1400 24270 1456
rect 26514 3576 26570 3632
rect 25962 1536 26018 1592
rect 27066 1944 27122 2000
rect 27618 1672 27674 1728
rect 6274 312 6330 368
<< metal3 >>
rect 0 27706 480 27736
rect 2773 27706 2839 27709
rect 0 27704 2839 27706
rect 0 27648 2778 27704
rect 2834 27648 2839 27704
rect 0 27646 2839 27648
rect 0 27616 480 27646
rect 2773 27643 2839 27646
rect 0 27162 480 27192
rect 4705 27162 4771 27165
rect 0 27160 4771 27162
rect 0 27104 4710 27160
rect 4766 27104 4771 27160
rect 0 27102 4771 27104
rect 0 27072 480 27102
rect 4705 27099 4771 27102
rect 0 26618 480 26648
rect 3601 26618 3667 26621
rect 0 26616 3667 26618
rect 0 26560 3606 26616
rect 3662 26560 3667 26616
rect 0 26558 3667 26560
rect 0 26528 480 26558
rect 3601 26555 3667 26558
rect 0 25938 480 25968
rect 4061 25938 4127 25941
rect 0 25936 4127 25938
rect 0 25880 4066 25936
rect 4122 25880 4127 25936
rect 0 25878 4127 25880
rect 0 25848 480 25878
rect 4061 25875 4127 25878
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25394 480 25424
rect 3049 25394 3115 25397
rect 0 25392 3115 25394
rect 0 25336 3054 25392
rect 3110 25336 3115 25392
rect 0 25334 3115 25336
rect 0 25304 480 25334
rect 3049 25331 3115 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 0 24850 480 24880
rect 2037 24850 2103 24853
rect 11053 24850 11119 24853
rect 0 24790 1226 24850
rect 0 24760 480 24790
rect 1166 24578 1226 24790
rect 2037 24848 11119 24850
rect 2037 24792 2042 24848
rect 2098 24792 11058 24848
rect 11114 24792 11119 24848
rect 2037 24790 11119 24792
rect 2037 24787 2103 24790
rect 11053 24787 11119 24790
rect 16113 24850 16179 24853
rect 17953 24850 18019 24853
rect 16113 24848 18019 24850
rect 16113 24792 16118 24848
rect 16174 24792 17958 24848
rect 18014 24792 18019 24848
rect 16113 24790 18019 24792
rect 16113 24787 16179 24790
rect 17953 24787 18019 24790
rect 18137 24850 18203 24853
rect 24209 24850 24275 24853
rect 18137 24848 24275 24850
rect 18137 24792 18142 24848
rect 18198 24792 24214 24848
rect 24270 24792 24275 24848
rect 18137 24790 24275 24792
rect 18137 24787 18203 24790
rect 24209 24787 24275 24790
rect 1945 24714 2011 24717
rect 6545 24714 6611 24717
rect 1945 24712 6611 24714
rect 1945 24656 1950 24712
rect 2006 24656 6550 24712
rect 6606 24656 6611 24712
rect 1945 24654 6611 24656
rect 1945 24651 2011 24654
rect 6545 24651 6611 24654
rect 10777 24714 10843 24717
rect 16757 24714 16823 24717
rect 10777 24712 16823 24714
rect 10777 24656 10782 24712
rect 10838 24656 16762 24712
rect 16818 24656 16823 24712
rect 10777 24654 16823 24656
rect 10777 24651 10843 24654
rect 16757 24651 16823 24654
rect 18873 24714 18939 24717
rect 20805 24714 20871 24717
rect 18873 24712 20871 24714
rect 18873 24656 18878 24712
rect 18934 24656 20810 24712
rect 20866 24656 20871 24712
rect 18873 24654 20871 24656
rect 18873 24651 18939 24654
rect 20805 24651 20871 24654
rect 3785 24578 3851 24581
rect 1166 24576 3851 24578
rect 1166 24520 3790 24576
rect 3846 24520 3851 24576
rect 1166 24518 3851 24520
rect 3785 24515 3851 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 14273 24442 14339 24445
rect 16205 24442 16271 24445
rect 14273 24440 16271 24442
rect 14273 24384 14278 24440
rect 14334 24384 16210 24440
rect 16266 24384 16271 24440
rect 14273 24382 16271 24384
rect 14273 24379 14339 24382
rect 16205 24379 16271 24382
rect 16389 24442 16455 24445
rect 17401 24442 17467 24445
rect 16389 24440 17467 24442
rect 16389 24384 16394 24440
rect 16450 24384 17406 24440
rect 17462 24384 17467 24440
rect 16389 24382 17467 24384
rect 16389 24379 16455 24382
rect 17401 24379 17467 24382
rect 17769 24442 17835 24445
rect 19425 24442 19491 24445
rect 17769 24440 19491 24442
rect 17769 24384 17774 24440
rect 17830 24384 19430 24440
rect 19486 24384 19491 24440
rect 17769 24382 19491 24384
rect 17769 24379 17835 24382
rect 19425 24379 19491 24382
rect 15469 24306 15535 24309
rect 26509 24306 26575 24309
rect 15469 24304 26575 24306
rect 15469 24248 15474 24304
rect 15530 24248 26514 24304
rect 26570 24248 26575 24304
rect 15469 24246 26575 24248
rect 15469 24243 15535 24246
rect 26509 24243 26575 24246
rect 0 24170 480 24200
rect 3601 24170 3667 24173
rect 0 24168 3667 24170
rect 0 24112 3606 24168
rect 3662 24112 3667 24168
rect 0 24110 3667 24112
rect 0 24080 480 24110
rect 3601 24107 3667 24110
rect 12249 24170 12315 24173
rect 18137 24170 18203 24173
rect 25957 24170 26023 24173
rect 12249 24168 18203 24170
rect 12249 24112 12254 24168
rect 12310 24112 18142 24168
rect 18198 24112 18203 24168
rect 12249 24110 18203 24112
rect 12249 24107 12315 24110
rect 18137 24107 18203 24110
rect 19566 24168 26023 24170
rect 19566 24112 25962 24168
rect 26018 24112 26023 24168
rect 19566 24110 26023 24112
rect 10685 24034 10751 24037
rect 12249 24034 12315 24037
rect 10685 24032 12315 24034
rect 10685 23976 10690 24032
rect 10746 23976 12254 24032
rect 12310 23976 12315 24032
rect 10685 23974 12315 23976
rect 10685 23971 10751 23974
rect 12249 23971 12315 23974
rect 17033 24034 17099 24037
rect 19566 24034 19626 24110
rect 25957 24107 26023 24110
rect 17033 24032 19626 24034
rect 17033 23976 17038 24032
rect 17094 23976 19626 24032
rect 17033 23974 19626 23976
rect 19701 24034 19767 24037
rect 21357 24034 21423 24037
rect 19701 24032 21423 24034
rect 19701 23976 19706 24032
rect 19762 23976 21362 24032
rect 21418 23976 21423 24032
rect 19701 23974 21423 23976
rect 17033 23971 17099 23974
rect 19701 23971 19767 23974
rect 21357 23971 21423 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 12617 23898 12683 23901
rect 6134 23896 12683 23898
rect 6134 23840 12622 23896
rect 12678 23840 12683 23896
rect 6134 23838 12683 23840
rect 4337 23762 4403 23765
rect 6134 23762 6194 23838
rect 12617 23835 12683 23838
rect 18229 23898 18295 23901
rect 20253 23898 20319 23901
rect 18229 23896 20319 23898
rect 18229 23840 18234 23896
rect 18290 23840 20258 23896
rect 20314 23840 20319 23896
rect 18229 23838 20319 23840
rect 18229 23835 18295 23838
rect 20253 23835 20319 23838
rect 21357 23898 21423 23901
rect 23105 23898 23171 23901
rect 21357 23896 23171 23898
rect 21357 23840 21362 23896
rect 21418 23840 23110 23896
rect 23166 23840 23171 23896
rect 21357 23838 23171 23840
rect 21357 23835 21423 23838
rect 23105 23835 23171 23838
rect 4337 23760 6194 23762
rect 4337 23704 4342 23760
rect 4398 23704 6194 23760
rect 4337 23702 6194 23704
rect 8017 23762 8083 23765
rect 13997 23762 14063 23765
rect 8017 23760 14063 23762
rect 8017 23704 8022 23760
rect 8078 23704 14002 23760
rect 14058 23704 14063 23760
rect 8017 23702 14063 23704
rect 4337 23699 4403 23702
rect 8017 23699 8083 23702
rect 13997 23699 14063 23702
rect 15101 23762 15167 23765
rect 27061 23762 27127 23765
rect 15101 23760 27127 23762
rect 15101 23704 15106 23760
rect 15162 23704 27066 23760
rect 27122 23704 27127 23760
rect 15101 23702 27127 23704
rect 15101 23699 15167 23702
rect 27061 23699 27127 23702
rect 0 23626 480 23656
rect 3969 23626 4035 23629
rect 4521 23626 4587 23629
rect 9581 23626 9647 23629
rect 0 23566 3848 23626
rect 0 23536 480 23566
rect 3788 23354 3848 23566
rect 3969 23624 9647 23626
rect 3969 23568 3974 23624
rect 4030 23568 4526 23624
rect 4582 23568 9586 23624
rect 9642 23568 9647 23624
rect 3969 23566 9647 23568
rect 3969 23563 4035 23566
rect 4521 23563 4587 23566
rect 9581 23563 9647 23566
rect 11421 23626 11487 23629
rect 23657 23626 23723 23629
rect 11421 23624 23723 23626
rect 11421 23568 11426 23624
rect 11482 23568 23662 23624
rect 23718 23568 23723 23624
rect 11421 23566 23723 23568
rect 11421 23563 11487 23566
rect 23657 23563 23723 23566
rect 5257 23490 5323 23493
rect 7465 23490 7531 23493
rect 5257 23488 7531 23490
rect 5257 23432 5262 23488
rect 5318 23432 7470 23488
rect 7526 23432 7531 23488
rect 5257 23430 7531 23432
rect 5257 23427 5323 23430
rect 7465 23427 7531 23430
rect 17217 23490 17283 23493
rect 19057 23490 19123 23493
rect 17217 23488 19123 23490
rect 17217 23432 17222 23488
rect 17278 23432 19062 23488
rect 19118 23432 19123 23488
rect 17217 23430 19123 23432
rect 17217 23427 17283 23430
rect 19057 23427 19123 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 5993 23354 6059 23357
rect 8845 23354 8911 23357
rect 3788 23352 6059 23354
rect 3788 23296 5998 23352
rect 6054 23296 6059 23352
rect 3788 23294 6059 23296
rect 5993 23291 6059 23294
rect 6134 23352 8911 23354
rect 6134 23296 8850 23352
rect 8906 23296 8911 23352
rect 6134 23294 8911 23296
rect 2129 23218 2195 23221
rect 6134 23218 6194 23294
rect 8845 23291 8911 23294
rect 23565 23354 23631 23357
rect 27520 23354 28000 23384
rect 23565 23352 28000 23354
rect 23565 23296 23570 23352
rect 23626 23296 28000 23352
rect 23565 23294 28000 23296
rect 23565 23291 23631 23294
rect 27520 23264 28000 23294
rect 20897 23218 20963 23221
rect 2129 23216 6194 23218
rect 2129 23160 2134 23216
rect 2190 23160 6194 23216
rect 2129 23158 6194 23160
rect 8526 23216 20963 23218
rect 8526 23160 20902 23216
rect 20958 23160 20963 23216
rect 8526 23158 20963 23160
rect 2129 23155 2195 23158
rect 0 23082 480 23112
rect 2865 23082 2931 23085
rect 0 23080 2931 23082
rect 0 23024 2870 23080
rect 2926 23024 2931 23080
rect 0 23022 2931 23024
rect 0 22992 480 23022
rect 2865 23019 2931 23022
rect 4061 22946 4127 22949
rect 4337 22946 4403 22949
rect 4061 22944 4403 22946
rect 4061 22888 4066 22944
rect 4122 22888 4342 22944
rect 4398 22888 4403 22944
rect 4061 22886 4403 22888
rect 4061 22883 4127 22886
rect 4337 22883 4403 22886
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 5533 22674 5599 22677
rect 8385 22674 8451 22677
rect 5533 22672 8451 22674
rect 5533 22616 5538 22672
rect 5594 22616 8390 22672
rect 8446 22616 8451 22672
rect 5533 22614 8451 22616
rect 5533 22611 5599 22614
rect 8385 22611 8451 22614
rect 0 22538 480 22568
rect 2957 22538 3023 22541
rect 0 22536 3023 22538
rect 0 22480 2962 22536
rect 3018 22480 3023 22536
rect 0 22478 3023 22480
rect 0 22448 480 22478
rect 2957 22475 3023 22478
rect 3785 22538 3851 22541
rect 6361 22538 6427 22541
rect 3785 22536 6427 22538
rect 3785 22480 3790 22536
rect 3846 22480 6366 22536
rect 6422 22480 6427 22536
rect 3785 22478 6427 22480
rect 3785 22475 3851 22478
rect 6361 22475 6427 22478
rect 2313 22402 2379 22405
rect 8526 22402 8586 23158
rect 20897 23155 20963 23158
rect 9581 23082 9647 23085
rect 17033 23082 17099 23085
rect 9581 23080 17099 23082
rect 9581 23024 9586 23080
rect 9642 23024 17038 23080
rect 17094 23024 17099 23080
rect 9581 23022 17099 23024
rect 9581 23019 9647 23022
rect 17033 23019 17099 23022
rect 15469 22946 15535 22949
rect 21909 22946 21975 22949
rect 15469 22944 21975 22946
rect 15469 22888 15474 22944
rect 15530 22888 21914 22944
rect 21970 22888 21975 22944
rect 15469 22886 21975 22888
rect 15469 22883 15535 22886
rect 21909 22883 21975 22886
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 19382 22716 19626 22776
rect 12893 22674 12959 22677
rect 19382 22674 19442 22716
rect 12893 22672 19442 22674
rect 12893 22616 12898 22672
rect 12954 22616 19442 22672
rect 12893 22614 19442 22616
rect 19566 22674 19626 22716
rect 24761 22674 24827 22677
rect 19566 22672 24827 22674
rect 19566 22616 24766 22672
rect 24822 22616 24827 22672
rect 19566 22614 24827 22616
rect 12893 22611 12959 22614
rect 24761 22611 24827 22614
rect 9397 22538 9463 22541
rect 12157 22538 12223 22541
rect 9397 22536 12223 22538
rect 9397 22480 9402 22536
rect 9458 22480 12162 22536
rect 12218 22480 12223 22536
rect 9397 22478 12223 22480
rect 9397 22475 9463 22478
rect 12157 22475 12223 22478
rect 14273 22538 14339 22541
rect 19333 22538 19399 22541
rect 14273 22536 19399 22538
rect 14273 22480 14278 22536
rect 14334 22480 19338 22536
rect 19394 22480 19399 22536
rect 14273 22478 19399 22480
rect 14273 22475 14339 22478
rect 19333 22475 19399 22478
rect 2313 22400 8586 22402
rect 2313 22344 2318 22400
rect 2374 22344 8586 22400
rect 2313 22342 8586 22344
rect 2313 22339 2379 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 7833 22266 7899 22269
rect 9857 22266 9923 22269
rect 14273 22266 14339 22269
rect 7833 22264 9923 22266
rect 7833 22208 7838 22264
rect 7894 22208 9862 22264
rect 9918 22208 9923 22264
rect 7833 22206 9923 22208
rect 7833 22203 7899 22206
rect 9857 22203 9923 22206
rect 10734 22264 14339 22266
rect 10734 22208 14278 22264
rect 14334 22208 14339 22264
rect 10734 22206 14339 22208
rect 5257 22130 5323 22133
rect 10734 22130 10794 22206
rect 14273 22203 14339 22206
rect 5257 22128 10794 22130
rect 5257 22072 5262 22128
rect 5318 22072 10794 22128
rect 5257 22070 10794 22072
rect 10869 22130 10935 22133
rect 12893 22130 12959 22133
rect 10869 22128 12959 22130
rect 10869 22072 10874 22128
rect 10930 22072 12898 22128
rect 12954 22072 12959 22128
rect 10869 22070 12959 22072
rect 5257 22067 5323 22070
rect 10869 22067 10935 22070
rect 12893 22067 12959 22070
rect 13537 22130 13603 22133
rect 13997 22130 14063 22133
rect 13537 22128 14063 22130
rect 13537 22072 13542 22128
rect 13598 22072 14002 22128
rect 14058 22072 14063 22128
rect 13537 22070 14063 22072
rect 13537 22067 13603 22070
rect 13997 22067 14063 22070
rect 3785 21994 3851 21997
rect 4613 21994 4679 21997
rect 3785 21992 4679 21994
rect 3785 21936 3790 21992
rect 3846 21936 4618 21992
rect 4674 21936 4679 21992
rect 3785 21934 4679 21936
rect 3785 21931 3851 21934
rect 4613 21931 4679 21934
rect 8753 21994 8819 21997
rect 13629 21994 13695 21997
rect 16665 21994 16731 21997
rect 23565 21994 23631 21997
rect 8753 21992 9460 21994
rect 8753 21936 8758 21992
rect 8814 21960 9460 21992
rect 13629 21992 23631 21994
rect 8814 21936 9644 21960
rect 8753 21934 9644 21936
rect 8753 21931 8819 21934
rect 9400 21900 9644 21934
rect 13629 21936 13634 21992
rect 13690 21936 16670 21992
rect 16726 21936 23570 21992
rect 23626 21936 23631 21992
rect 13629 21934 23631 21936
rect 13629 21931 13695 21934
rect 16665 21931 16731 21934
rect 23565 21931 23631 21934
rect 0 21858 480 21888
rect 1577 21858 1643 21861
rect 0 21856 1643 21858
rect 0 21800 1582 21856
rect 1638 21800 1643 21856
rect 0 21798 1643 21800
rect 9584 21858 9644 21900
rect 12341 21858 12407 21861
rect 9584 21856 12407 21858
rect 9584 21800 12346 21856
rect 12402 21800 12407 21856
rect 9584 21798 12407 21800
rect 0 21768 480 21798
rect 1577 21795 1643 21798
rect 12341 21795 12407 21798
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 8109 21722 8175 21725
rect 11237 21722 11303 21725
rect 8109 21720 11303 21722
rect 8109 21664 8114 21720
rect 8170 21664 11242 21720
rect 11298 21664 11303 21720
rect 8109 21662 11303 21664
rect 8109 21659 8175 21662
rect 11237 21659 11303 21662
rect 10961 21586 11027 21589
rect 12801 21586 12867 21589
rect 10961 21584 12867 21586
rect 10961 21528 10966 21584
rect 11022 21528 12806 21584
rect 12862 21528 12867 21584
rect 10961 21526 12867 21528
rect 10961 21523 11027 21526
rect 12801 21523 12867 21526
rect 3417 21450 3483 21453
rect 8845 21450 8911 21453
rect 3417 21448 8911 21450
rect 3417 21392 3422 21448
rect 3478 21392 8850 21448
rect 8906 21392 8911 21448
rect 3417 21390 8911 21392
rect 3417 21387 3483 21390
rect 8845 21387 8911 21390
rect 13077 21450 13143 21453
rect 17585 21450 17651 21453
rect 13077 21448 17651 21450
rect 13077 21392 13082 21448
rect 13138 21392 17590 21448
rect 17646 21392 17651 21448
rect 13077 21390 17651 21392
rect 13077 21387 13143 21390
rect 17585 21387 17651 21390
rect 0 21314 480 21344
rect 1393 21314 1459 21317
rect 0 21312 1459 21314
rect 0 21256 1398 21312
rect 1454 21256 1459 21312
rect 0 21254 1459 21256
rect 0 21224 480 21254
rect 1393 21251 1459 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 1393 21042 1459 21045
rect 1945 21042 2011 21045
rect 7005 21042 7071 21045
rect 1393 21040 7071 21042
rect 1393 20984 1398 21040
rect 1454 20984 1950 21040
rect 2006 20984 7010 21040
rect 7066 20984 7071 21040
rect 1393 20982 7071 20984
rect 1393 20979 1459 20982
rect 1945 20979 2011 20982
rect 7005 20979 7071 20982
rect 12801 20906 12867 20909
rect 13445 20906 13511 20909
rect 12801 20904 13511 20906
rect 12801 20848 12806 20904
rect 12862 20848 13450 20904
rect 13506 20848 13511 20904
rect 12801 20846 13511 20848
rect 12801 20843 12867 20846
rect 13445 20843 13511 20846
rect 0 20770 480 20800
rect 4061 20770 4127 20773
rect 0 20768 4127 20770
rect 0 20712 4066 20768
rect 4122 20712 4127 20768
rect 0 20710 4127 20712
rect 0 20680 480 20710
rect 4061 20707 4127 20710
rect 6913 20770 6979 20773
rect 13997 20770 14063 20773
rect 6913 20768 14063 20770
rect 6913 20712 6918 20768
rect 6974 20712 14002 20768
rect 14058 20712 14063 20768
rect 6913 20710 14063 20712
rect 6913 20707 6979 20710
rect 13997 20707 14063 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 2405 20498 2471 20501
rect 12341 20498 12407 20501
rect 2405 20496 12407 20498
rect 2405 20440 2410 20496
rect 2466 20440 12346 20496
rect 12402 20440 12407 20496
rect 2405 20438 12407 20440
rect 2405 20435 2471 20438
rect 12341 20435 12407 20438
rect 2865 20362 2931 20365
rect 7189 20362 7255 20365
rect 2865 20360 7255 20362
rect 2865 20304 2870 20360
rect 2926 20304 7194 20360
rect 7250 20304 7255 20360
rect 2865 20302 7255 20304
rect 2865 20299 2931 20302
rect 7189 20299 7255 20302
rect 841 20226 907 20229
rect 8845 20226 8911 20229
rect 841 20224 8911 20226
rect 841 20168 846 20224
rect 902 20168 8850 20224
rect 8906 20168 8911 20224
rect 841 20166 8911 20168
rect 841 20163 907 20166
rect 8845 20163 8911 20166
rect 10277 20160 10597 20161
rect 0 20090 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 8017 20090 8083 20093
rect 0 20088 8083 20090
rect 0 20032 8022 20088
rect 8078 20032 8083 20088
rect 0 20030 8083 20032
rect 0 20000 480 20030
rect 8017 20027 8083 20030
rect 565 19954 631 19957
rect 8477 19954 8543 19957
rect 565 19952 8543 19954
rect 565 19896 570 19952
rect 626 19896 8482 19952
rect 8538 19896 8543 19952
rect 565 19894 8543 19896
rect 565 19891 631 19894
rect 8477 19891 8543 19894
rect 12249 19954 12315 19957
rect 15745 19954 15811 19957
rect 12249 19952 15811 19954
rect 12249 19896 12254 19952
rect 12310 19896 15750 19952
rect 15806 19896 15811 19952
rect 12249 19894 15811 19896
rect 12249 19891 12315 19894
rect 15745 19891 15811 19894
rect 3049 19818 3115 19821
rect 12617 19818 12683 19821
rect 3049 19816 12683 19818
rect 3049 19760 3054 19816
rect 3110 19760 12622 19816
rect 12678 19760 12683 19816
rect 3049 19758 12683 19760
rect 3049 19755 3115 19758
rect 12617 19755 12683 19758
rect 14181 19818 14247 19821
rect 19425 19818 19491 19821
rect 14181 19816 19491 19818
rect 14181 19760 14186 19816
rect 14242 19760 19430 19816
rect 19486 19760 19491 19816
rect 14181 19758 19491 19760
rect 14181 19755 14247 19758
rect 19425 19755 19491 19758
rect 2681 19682 2747 19685
rect 4521 19682 4587 19685
rect 2681 19680 4587 19682
rect 2681 19624 2686 19680
rect 2742 19624 4526 19680
rect 4582 19624 4587 19680
rect 2681 19622 4587 19624
rect 2681 19619 2747 19622
rect 4521 19619 4587 19622
rect 5610 19616 5930 19617
rect 0 19546 480 19576
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 2681 19546 2747 19549
rect 0 19544 2747 19546
rect 0 19488 2686 19544
rect 2742 19488 2747 19544
rect 0 19486 2747 19488
rect 0 19456 480 19486
rect 2681 19483 2747 19486
rect 7281 19410 7347 19413
rect 8293 19410 8359 19413
rect 7281 19408 8359 19410
rect 7281 19352 7286 19408
rect 7342 19352 8298 19408
rect 8354 19352 8359 19408
rect 7281 19350 8359 19352
rect 7281 19347 7347 19350
rect 8293 19347 8359 19350
rect 14549 19410 14615 19413
rect 15469 19410 15535 19413
rect 14549 19408 15535 19410
rect 14549 19352 14554 19408
rect 14610 19352 15474 19408
rect 15530 19352 15535 19408
rect 14549 19350 15535 19352
rect 14549 19347 14615 19350
rect 15469 19347 15535 19350
rect 6177 19274 6243 19277
rect 12249 19274 12315 19277
rect 6177 19272 12315 19274
rect 6177 19216 6182 19272
rect 6238 19216 12254 19272
rect 12310 19216 12315 19272
rect 6177 19214 12315 19216
rect 6177 19211 6243 19214
rect 12249 19211 12315 19214
rect 3233 19138 3299 19141
rect 5993 19138 6059 19141
rect 3233 19136 6059 19138
rect 3233 19080 3238 19136
rect 3294 19080 5998 19136
rect 6054 19080 6059 19136
rect 3233 19078 6059 19080
rect 3233 19075 3299 19078
rect 5993 19075 6059 19078
rect 13905 19138 13971 19141
rect 17493 19138 17559 19141
rect 13905 19136 17559 19138
rect 13905 19080 13910 19136
rect 13966 19080 17498 19136
rect 17554 19080 17559 19136
rect 13905 19078 17559 19080
rect 13905 19075 13971 19078
rect 17493 19075 17559 19078
rect 10277 19072 10597 19073
rect 0 19002 480 19032
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 1393 19002 1459 19005
rect 0 19000 1459 19002
rect 0 18944 1398 19000
rect 1454 18944 1459 19000
rect 0 18942 1459 18944
rect 0 18912 480 18942
rect 1393 18939 1459 18942
rect 3141 19002 3207 19005
rect 8017 19002 8083 19005
rect 3141 19000 8083 19002
rect 3141 18944 3146 19000
rect 3202 18944 8022 19000
rect 8078 18944 8083 19000
rect 3141 18942 8083 18944
rect 3141 18939 3207 18942
rect 8017 18939 8083 18942
rect 8201 19002 8267 19005
rect 8201 19000 8770 19002
rect 8201 18944 8206 19000
rect 8262 18944 8770 19000
rect 8201 18942 8770 18944
rect 8201 18939 8267 18942
rect 2037 18866 2103 18869
rect 8569 18866 8635 18869
rect 2037 18864 8635 18866
rect 2037 18808 2042 18864
rect 2098 18808 8574 18864
rect 8630 18808 8635 18864
rect 2037 18806 8635 18808
rect 8710 18866 8770 18942
rect 11789 18866 11855 18869
rect 8710 18864 11855 18866
rect 8710 18808 11794 18864
rect 11850 18808 11855 18864
rect 8710 18806 11855 18808
rect 2037 18803 2103 18806
rect 8569 18803 8635 18806
rect 11789 18803 11855 18806
rect 6545 18730 6611 18733
rect 9397 18730 9463 18733
rect 6545 18728 9463 18730
rect 6545 18672 6550 18728
rect 6606 18672 9402 18728
rect 9458 18672 9463 18728
rect 6545 18670 9463 18672
rect 6545 18667 6611 18670
rect 9397 18667 9463 18670
rect 17309 18730 17375 18733
rect 27613 18730 27679 18733
rect 17309 18728 27679 18730
rect 17309 18672 17314 18728
rect 17370 18672 27618 18728
rect 27674 18672 27679 18728
rect 17309 18670 27679 18672
rect 17309 18667 17375 18670
rect 27613 18667 27679 18670
rect 7925 18594 7991 18597
rect 10133 18594 10199 18597
rect 11973 18594 12039 18597
rect 7925 18592 12039 18594
rect 7925 18536 7930 18592
rect 7986 18536 10138 18592
rect 10194 18536 11978 18592
rect 12034 18536 12039 18592
rect 7925 18534 12039 18536
rect 7925 18531 7991 18534
rect 10133 18531 10199 18534
rect 11973 18531 12039 18534
rect 5610 18528 5930 18529
rect 0 18458 480 18488
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 1577 18458 1643 18461
rect 0 18456 1643 18458
rect 0 18400 1582 18456
rect 1638 18400 1643 18456
rect 0 18398 1643 18400
rect 0 18368 480 18398
rect 1577 18395 1643 18398
rect 3325 18322 3391 18325
rect 4613 18322 4679 18325
rect 13813 18322 13879 18325
rect 3325 18320 13879 18322
rect 3325 18264 3330 18320
rect 3386 18264 4618 18320
rect 4674 18264 13818 18320
rect 13874 18264 13879 18320
rect 3325 18262 13879 18264
rect 3325 18259 3391 18262
rect 4613 18259 4679 18262
rect 13813 18259 13879 18262
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 2037 17914 2103 17917
rect 4245 17914 4311 17917
rect 2037 17912 4311 17914
rect 2037 17856 2042 17912
rect 2098 17856 4250 17912
rect 4306 17856 4311 17912
rect 2037 17854 4311 17856
rect 2037 17851 2103 17854
rect 4245 17851 4311 17854
rect 0 17778 480 17808
rect 2681 17778 2747 17781
rect 0 17776 2747 17778
rect 0 17720 2686 17776
rect 2742 17720 2747 17776
rect 0 17718 2747 17720
rect 0 17688 480 17718
rect 2681 17715 2747 17718
rect 9949 17778 10015 17781
rect 16205 17778 16271 17781
rect 9949 17776 16271 17778
rect 9949 17720 9954 17776
rect 10010 17720 16210 17776
rect 16266 17720 16271 17776
rect 9949 17718 16271 17720
rect 9949 17715 10015 17718
rect 16205 17715 16271 17718
rect 9489 17642 9555 17645
rect 10317 17642 10383 17645
rect 17401 17642 17467 17645
rect 9489 17640 10383 17642
rect 9489 17584 9494 17640
rect 9550 17584 10322 17640
rect 10378 17584 10383 17640
rect 9489 17582 10383 17584
rect 9489 17579 9555 17582
rect 10317 17579 10383 17582
rect 14782 17640 17467 17642
rect 14782 17584 17406 17640
rect 17462 17584 17467 17640
rect 14782 17582 17467 17584
rect 7557 17506 7623 17509
rect 14782 17506 14842 17582
rect 17401 17579 17467 17582
rect 7557 17504 14842 17506
rect 7557 17448 7562 17504
rect 7618 17448 14842 17504
rect 7557 17446 14842 17448
rect 7557 17443 7623 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 15653 17370 15719 17373
rect 20805 17370 20871 17373
rect 15653 17368 20871 17370
rect 15653 17312 15658 17368
rect 15714 17312 20810 17368
rect 20866 17312 20871 17368
rect 15653 17310 20871 17312
rect 15653 17307 15719 17310
rect 20805 17307 20871 17310
rect 0 17234 480 17264
rect 1485 17234 1551 17237
rect 0 17232 1551 17234
rect 0 17176 1490 17232
rect 1546 17176 1551 17232
rect 0 17174 1551 17176
rect 0 17144 480 17174
rect 1485 17171 1551 17174
rect 1945 17234 2011 17237
rect 5625 17234 5691 17237
rect 1945 17232 5691 17234
rect 1945 17176 1950 17232
rect 2006 17176 5630 17232
rect 5686 17176 5691 17232
rect 1945 17174 5691 17176
rect 1945 17171 2011 17174
rect 5625 17171 5691 17174
rect 13353 17234 13419 17237
rect 18229 17234 18295 17237
rect 13353 17232 18295 17234
rect 13353 17176 13358 17232
rect 13414 17176 18234 17232
rect 18290 17176 18295 17232
rect 13353 17174 18295 17176
rect 13353 17171 13419 17174
rect 18229 17171 18295 17174
rect 10041 17098 10107 17101
rect 16021 17098 16087 17101
rect 10041 17096 16087 17098
rect 10041 17040 10046 17096
rect 10102 17040 16026 17096
rect 16082 17040 16087 17096
rect 10041 17038 16087 17040
rect 10041 17035 10107 17038
rect 16021 17035 16087 17038
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 0 16690 480 16720
rect 1393 16690 1459 16693
rect 0 16688 1459 16690
rect 0 16632 1398 16688
rect 1454 16632 1459 16688
rect 0 16630 1459 16632
rect 0 16600 480 16630
rect 1393 16627 1459 16630
rect 5533 16690 5599 16693
rect 9673 16690 9739 16693
rect 5533 16688 9739 16690
rect 5533 16632 5538 16688
rect 5594 16632 9678 16688
rect 9734 16632 9739 16688
rect 5533 16630 9739 16632
rect 5533 16627 5599 16630
rect 9673 16627 9739 16630
rect 13077 16690 13143 16693
rect 15929 16690 15995 16693
rect 13077 16688 15995 16690
rect 13077 16632 13082 16688
rect 13138 16632 15934 16688
rect 15990 16632 15995 16688
rect 13077 16630 15995 16632
rect 13077 16627 13143 16630
rect 15929 16627 15995 16630
rect 6085 16554 6151 16557
rect 7005 16554 7071 16557
rect 17125 16554 17191 16557
rect 18597 16554 18663 16557
rect 6085 16552 18663 16554
rect 6085 16496 6090 16552
rect 6146 16496 7010 16552
rect 7066 16496 17130 16552
rect 17186 16496 18602 16552
rect 18658 16496 18663 16552
rect 6085 16494 18663 16496
rect 6085 16491 6151 16494
rect 7005 16491 7071 16494
rect 17125 16491 17191 16494
rect 18597 16491 18663 16494
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 6637 16146 6703 16149
rect 7465 16146 7531 16149
rect 17217 16146 17283 16149
rect 6637 16144 17283 16146
rect 6637 16088 6642 16144
rect 6698 16088 7470 16144
rect 7526 16088 17222 16144
rect 17278 16088 17283 16144
rect 6637 16086 17283 16088
rect 6637 16083 6703 16086
rect 7465 16083 7531 16086
rect 17217 16083 17283 16086
rect 0 16010 480 16040
rect 1577 16010 1643 16013
rect 0 16008 1643 16010
rect 0 15952 1582 16008
rect 1638 15952 1643 16008
rect 0 15950 1643 15952
rect 0 15920 480 15950
rect 1577 15947 1643 15950
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 12801 15738 12867 15741
rect 15285 15738 15351 15741
rect 12801 15736 15351 15738
rect 12801 15680 12806 15736
rect 12862 15680 15290 15736
rect 15346 15680 15351 15736
rect 12801 15678 15351 15680
rect 12801 15675 12867 15678
rect 15285 15675 15351 15678
rect 2037 15602 2103 15605
rect 10777 15602 10843 15605
rect 2037 15600 10843 15602
rect 2037 15544 2042 15600
rect 2098 15544 10782 15600
rect 10838 15544 10843 15600
rect 2037 15542 10843 15544
rect 2037 15539 2103 15542
rect 10777 15539 10843 15542
rect 11421 15602 11487 15605
rect 15101 15602 15167 15605
rect 11421 15600 15167 15602
rect 11421 15544 11426 15600
rect 11482 15544 15106 15600
rect 15162 15544 15167 15600
rect 11421 15542 15167 15544
rect 11421 15539 11487 15542
rect 15101 15539 15167 15542
rect 0 15466 480 15496
rect 2773 15466 2839 15469
rect 0 15464 2839 15466
rect 0 15408 2778 15464
rect 2834 15408 2839 15464
rect 0 15406 2839 15408
rect 0 15376 480 15406
rect 2773 15403 2839 15406
rect 4061 15466 4127 15469
rect 6821 15466 6887 15469
rect 10041 15468 10107 15469
rect 4061 15464 6887 15466
rect 4061 15408 4066 15464
rect 4122 15408 6826 15464
rect 6882 15408 6887 15464
rect 4061 15406 6887 15408
rect 4061 15403 4127 15406
rect 6821 15403 6887 15406
rect 9990 15404 9996 15468
rect 10060 15466 10107 15468
rect 10060 15464 10152 15466
rect 10102 15408 10152 15464
rect 10060 15406 10152 15408
rect 10060 15404 10107 15406
rect 10041 15403 10107 15404
rect 6085 15330 6151 15333
rect 10041 15330 10107 15333
rect 6085 15328 10107 15330
rect 6085 15272 6090 15328
rect 6146 15272 10046 15328
rect 10102 15272 10107 15328
rect 6085 15270 10107 15272
rect 6085 15267 6151 15270
rect 10041 15267 10107 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 3969 15194 4035 15197
rect 5441 15194 5507 15197
rect 3969 15192 5507 15194
rect 3969 15136 3974 15192
rect 4030 15136 5446 15192
rect 5502 15136 5507 15192
rect 3969 15134 5507 15136
rect 3969 15131 4035 15134
rect 5441 15131 5507 15134
rect 6453 15194 6519 15197
rect 7189 15194 7255 15197
rect 6453 15192 7255 15194
rect 6453 15136 6458 15192
rect 6514 15136 7194 15192
rect 7250 15136 7255 15192
rect 6453 15134 7255 15136
rect 6453 15131 6519 15134
rect 7189 15131 7255 15134
rect 9121 15194 9187 15197
rect 16205 15194 16271 15197
rect 19333 15194 19399 15197
rect 9121 15192 14842 15194
rect 9121 15136 9126 15192
rect 9182 15136 14842 15192
rect 9121 15134 14842 15136
rect 9121 15131 9187 15134
rect 2865 15058 2931 15061
rect 3325 15058 3391 15061
rect 6361 15058 6427 15061
rect 2865 15056 6427 15058
rect 2865 15000 2870 15056
rect 2926 15000 3330 15056
rect 3386 15000 6366 15056
rect 6422 15000 6427 15056
rect 2865 14998 6427 15000
rect 2865 14995 2931 14998
rect 3325 14995 3391 14998
rect 6361 14995 6427 14998
rect 7189 15058 7255 15061
rect 14273 15058 14339 15061
rect 7189 15056 14339 15058
rect 7189 15000 7194 15056
rect 7250 15000 14278 15056
rect 14334 15000 14339 15056
rect 7189 14998 14339 15000
rect 14782 15058 14842 15134
rect 16205 15192 19399 15194
rect 16205 15136 16210 15192
rect 16266 15136 19338 15192
rect 19394 15136 19399 15192
rect 16205 15134 19399 15136
rect 16205 15131 16271 15134
rect 19333 15131 19399 15134
rect 19517 15058 19583 15061
rect 14782 15056 19583 15058
rect 14782 15000 19522 15056
rect 19578 15000 19583 15056
rect 14782 14998 19583 15000
rect 7189 14995 7255 14998
rect 14273 14995 14339 14998
rect 19517 14995 19583 14998
rect 0 14922 480 14952
rect 1485 14922 1551 14925
rect 0 14920 1551 14922
rect 0 14864 1490 14920
rect 1546 14864 1551 14920
rect 0 14862 1551 14864
rect 0 14832 480 14862
rect 1485 14859 1551 14862
rect 2865 14922 2931 14925
rect 6177 14922 6243 14925
rect 2865 14920 6243 14922
rect 2865 14864 2870 14920
rect 2926 14864 6182 14920
rect 6238 14864 6243 14920
rect 2865 14862 6243 14864
rect 2865 14859 2931 14862
rect 6177 14859 6243 14862
rect 1393 14786 1459 14789
rect 3601 14786 3667 14789
rect 5165 14786 5231 14789
rect 1393 14784 5231 14786
rect 1393 14728 1398 14784
rect 1454 14728 3606 14784
rect 3662 14728 5170 14784
rect 5226 14728 5231 14784
rect 1393 14726 5231 14728
rect 1393 14723 1459 14726
rect 3601 14723 3667 14726
rect 5165 14723 5231 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 14089 14514 14155 14517
rect 14273 14514 14339 14517
rect 14089 14512 14339 14514
rect 14089 14456 14094 14512
rect 14150 14456 14278 14512
rect 14334 14456 14339 14512
rect 14089 14454 14339 14456
rect 14089 14451 14155 14454
rect 14273 14451 14339 14454
rect 0 14378 480 14408
rect 4153 14378 4219 14381
rect 0 14376 4219 14378
rect 0 14320 4158 14376
rect 4214 14320 4219 14376
rect 0 14318 4219 14320
rect 0 14288 480 14318
rect 4153 14315 4219 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 2589 14106 2655 14109
rect 3049 14106 3115 14109
rect 2589 14104 3115 14106
rect 2589 14048 2594 14104
rect 2650 14048 3054 14104
rect 3110 14048 3115 14104
rect 2589 14046 3115 14048
rect 2589 14043 2655 14046
rect 3049 14043 3115 14046
rect 7925 14106 7991 14109
rect 9121 14106 9187 14109
rect 7925 14104 9187 14106
rect 7925 14048 7930 14104
rect 7986 14048 9126 14104
rect 9182 14048 9187 14104
rect 7925 14046 9187 14048
rect 7925 14043 7991 14046
rect 9121 14043 9187 14046
rect 7097 13970 7163 13973
rect 9213 13970 9279 13973
rect 14733 13970 14799 13973
rect 27520 13970 28000 14000
rect 7097 13968 9138 13970
rect 7097 13912 7102 13968
rect 7158 13912 9138 13968
rect 7097 13910 9138 13912
rect 7097 13907 7163 13910
rect 2957 13834 3023 13837
rect 3366 13834 3372 13836
rect 2957 13832 3372 13834
rect 2957 13776 2962 13832
rect 3018 13776 3372 13832
rect 2957 13774 3372 13776
rect 2957 13771 3023 13774
rect 3366 13772 3372 13774
rect 3436 13772 3442 13836
rect 3601 13834 3667 13837
rect 4061 13834 4127 13837
rect 8845 13834 8911 13837
rect 3601 13832 8911 13834
rect 3601 13776 3606 13832
rect 3662 13776 4066 13832
rect 4122 13776 8850 13832
rect 8906 13776 8911 13832
rect 3601 13774 8911 13776
rect 9078 13834 9138 13910
rect 9213 13968 14799 13970
rect 9213 13912 9218 13968
rect 9274 13912 14738 13968
rect 14794 13912 14799 13968
rect 9213 13910 14799 13912
rect 9213 13907 9279 13910
rect 14733 13907 14799 13910
rect 23614 13910 28000 13970
rect 12709 13834 12775 13837
rect 9078 13832 12775 13834
rect 9078 13776 12714 13832
rect 12770 13776 12775 13832
rect 9078 13774 12775 13776
rect 3601 13771 3667 13774
rect 4061 13771 4127 13774
rect 8845 13771 8911 13774
rect 12709 13771 12775 13774
rect 0 13698 480 13728
rect 1669 13698 1735 13701
rect 0 13696 1735 13698
rect 0 13640 1674 13696
rect 1730 13640 1735 13696
rect 0 13638 1735 13640
rect 0 13608 480 13638
rect 1669 13635 1735 13638
rect 2405 13698 2471 13701
rect 5533 13698 5599 13701
rect 2405 13696 5599 13698
rect 2405 13640 2410 13696
rect 2466 13640 5538 13696
rect 5594 13640 5599 13696
rect 2405 13638 5599 13640
rect 2405 13635 2471 13638
rect 5533 13635 5599 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 3417 13562 3483 13565
rect 6821 13562 6887 13565
rect 8569 13562 8635 13565
rect 3417 13560 8635 13562
rect 3417 13504 3422 13560
rect 3478 13504 6826 13560
rect 6882 13504 8574 13560
rect 8630 13504 8635 13560
rect 3417 13502 8635 13504
rect 3417 13499 3483 13502
rect 6821 13499 6887 13502
rect 8569 13499 8635 13502
rect 1393 13426 1459 13429
rect 3969 13426 4035 13429
rect 1393 13424 4035 13426
rect 1393 13368 1398 13424
rect 1454 13368 3974 13424
rect 4030 13368 4035 13424
rect 1393 13366 4035 13368
rect 1393 13363 1459 13366
rect 3969 13363 4035 13366
rect 6361 13426 6427 13429
rect 11053 13426 11119 13429
rect 6361 13424 11119 13426
rect 6361 13368 6366 13424
rect 6422 13368 11058 13424
rect 11114 13368 11119 13424
rect 6361 13366 11119 13368
rect 6361 13363 6427 13366
rect 11053 13363 11119 13366
rect 18321 13426 18387 13429
rect 23614 13426 23674 13910
rect 27520 13880 28000 13910
rect 18321 13424 23674 13426
rect 18321 13368 18326 13424
rect 18382 13368 23674 13424
rect 18321 13366 23674 13368
rect 18321 13363 18387 13366
rect 8569 13290 8635 13293
rect 12801 13290 12867 13293
rect 8569 13288 12867 13290
rect 8569 13232 8574 13288
rect 8630 13232 12806 13288
rect 12862 13232 12867 13288
rect 8569 13230 12867 13232
rect 8569 13227 8635 13230
rect 12801 13227 12867 13230
rect 0 13154 480 13184
rect 1577 13154 1643 13157
rect 0 13152 1643 13154
rect 0 13096 1582 13152
rect 1638 13096 1643 13152
rect 0 13094 1643 13096
rect 0 13064 480 13094
rect 1577 13091 1643 13094
rect 8477 13154 8543 13157
rect 14549 13154 14615 13157
rect 8477 13152 14615 13154
rect 8477 13096 8482 13152
rect 8538 13096 14554 13152
rect 14610 13096 14615 13152
rect 8477 13094 14615 13096
rect 8477 13091 8543 13094
rect 14549 13091 14615 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 9397 13018 9463 13021
rect 11881 13018 11947 13021
rect 9397 13016 11947 13018
rect 9397 12960 9402 13016
rect 9458 12960 11886 13016
rect 11942 12960 11947 13016
rect 9397 12958 11947 12960
rect 9397 12955 9463 12958
rect 11881 12955 11947 12958
rect 4889 12882 4955 12885
rect 11421 12882 11487 12885
rect 14641 12882 14707 12885
rect 4889 12880 14707 12882
rect 4889 12824 4894 12880
rect 4950 12824 11426 12880
rect 11482 12824 14646 12880
rect 14702 12824 14707 12880
rect 4889 12822 14707 12824
rect 4889 12819 4955 12822
rect 11421 12819 11487 12822
rect 14641 12819 14707 12822
rect 4429 12746 4495 12749
rect 13721 12746 13787 12749
rect 4429 12744 13787 12746
rect 4429 12688 4434 12744
rect 4490 12688 13726 12744
rect 13782 12688 13787 12744
rect 4429 12686 13787 12688
rect 4429 12683 4495 12686
rect 13721 12683 13787 12686
rect 0 12610 480 12640
rect 1577 12610 1643 12613
rect 0 12608 1643 12610
rect 0 12552 1582 12608
rect 1638 12552 1643 12608
rect 0 12550 1643 12552
rect 0 12520 480 12550
rect 1577 12547 1643 12550
rect 11881 12610 11947 12613
rect 19425 12610 19491 12613
rect 11881 12608 19491 12610
rect 11881 12552 11886 12608
rect 11942 12552 19430 12608
rect 19486 12552 19491 12608
rect 11881 12550 19491 12552
rect 11881 12547 11947 12550
rect 19425 12547 19491 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 5625 12474 5691 12477
rect 9489 12474 9555 12477
rect 5625 12472 9555 12474
rect 5625 12416 5630 12472
rect 5686 12416 9494 12472
rect 9550 12416 9555 12472
rect 5625 12414 9555 12416
rect 5625 12411 5691 12414
rect 9489 12411 9555 12414
rect 13353 12474 13419 12477
rect 13629 12474 13695 12477
rect 13353 12472 13695 12474
rect 13353 12416 13358 12472
rect 13414 12416 13634 12472
rect 13690 12416 13695 12472
rect 13353 12414 13695 12416
rect 13353 12411 13419 12414
rect 13629 12411 13695 12414
rect 7189 12338 7255 12341
rect 9673 12338 9739 12341
rect 7189 12336 9739 12338
rect 7189 12280 7194 12336
rect 7250 12280 9678 12336
rect 9734 12280 9739 12336
rect 7189 12278 9739 12280
rect 7189 12275 7255 12278
rect 9673 12275 9739 12278
rect 11697 12338 11763 12341
rect 15745 12338 15811 12341
rect 11697 12336 15811 12338
rect 11697 12280 11702 12336
rect 11758 12280 15750 12336
rect 15806 12280 15811 12336
rect 11697 12278 15811 12280
rect 11697 12275 11763 12278
rect 15745 12275 15811 12278
rect 17033 12338 17099 12341
rect 17309 12338 17375 12341
rect 17033 12336 17375 12338
rect 17033 12280 17038 12336
rect 17094 12280 17314 12336
rect 17370 12280 17375 12336
rect 17033 12278 17375 12280
rect 17033 12275 17099 12278
rect 17309 12275 17375 12278
rect 3509 12202 3575 12205
rect 3509 12200 11944 12202
rect 3509 12144 3514 12200
rect 3570 12144 11944 12200
rect 3509 12142 11944 12144
rect 3509 12139 3575 12142
rect 9397 12066 9463 12069
rect 11605 12066 11671 12069
rect 9397 12064 11671 12066
rect 9397 12008 9402 12064
rect 9458 12008 11610 12064
rect 11666 12008 11671 12064
rect 9397 12006 11671 12008
rect 9397 12003 9463 12006
rect 11605 12003 11671 12006
rect 5610 12000 5930 12001
rect 0 11930 480 11960
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 4245 11930 4311 11933
rect 11094 11930 11100 11932
rect 0 11928 4311 11930
rect 0 11872 4250 11928
rect 4306 11872 4311 11928
rect 0 11870 4311 11872
rect 0 11840 480 11870
rect 4245 11867 4311 11870
rect 6134 11870 11100 11930
rect 3141 11794 3207 11797
rect 4521 11794 4587 11797
rect 6134 11794 6194 11870
rect 11094 11868 11100 11870
rect 11164 11868 11170 11932
rect 11884 11930 11944 12142
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 14733 11930 14799 11933
rect 11884 11928 14799 11930
rect 11884 11872 14738 11928
rect 14794 11872 14799 11928
rect 11884 11870 14799 11872
rect 14733 11867 14799 11870
rect 3141 11792 6194 11794
rect 3141 11736 3146 11792
rect 3202 11736 4526 11792
rect 4582 11736 6194 11792
rect 3141 11734 6194 11736
rect 6453 11794 6519 11797
rect 8937 11794 9003 11797
rect 6453 11792 9003 11794
rect 6453 11736 6458 11792
rect 6514 11736 8942 11792
rect 8998 11736 9003 11792
rect 6453 11734 9003 11736
rect 3141 11731 3207 11734
rect 4521 11731 4587 11734
rect 6453 11731 6519 11734
rect 8937 11731 9003 11734
rect 2405 11658 2471 11661
rect 11145 11658 11211 11661
rect 14273 11658 14339 11661
rect 2405 11656 14339 11658
rect 2405 11600 2410 11656
rect 2466 11600 11150 11656
rect 11206 11600 14278 11656
rect 14334 11600 14339 11656
rect 2405 11598 14339 11600
rect 2405 11595 2471 11598
rect 11145 11595 11211 11598
rect 14273 11595 14339 11598
rect 2221 11522 2287 11525
rect 3417 11522 3483 11525
rect 2221 11520 3483 11522
rect 2221 11464 2226 11520
rect 2282 11464 3422 11520
rect 3478 11464 3483 11520
rect 2221 11462 3483 11464
rect 2221 11459 2287 11462
rect 3417 11459 3483 11462
rect 14641 11522 14707 11525
rect 16757 11522 16823 11525
rect 14641 11520 16823 11522
rect 14641 11464 14646 11520
rect 14702 11464 16762 11520
rect 16818 11464 16823 11520
rect 14641 11462 16823 11464
rect 14641 11459 14707 11462
rect 16757 11459 16823 11462
rect 10277 11456 10597 11457
rect 0 11386 480 11416
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 3969 11386 4035 11389
rect 0 11384 4035 11386
rect 0 11328 3974 11384
rect 4030 11328 4035 11384
rect 0 11326 4035 11328
rect 0 11296 480 11326
rect 3969 11323 4035 11326
rect 13261 11386 13327 11389
rect 14917 11386 14983 11389
rect 18045 11386 18111 11389
rect 13261 11384 14796 11386
rect 13261 11328 13266 11384
rect 13322 11328 14796 11384
rect 13261 11326 14796 11328
rect 13261 11323 13327 11326
rect 14736 11253 14796 11326
rect 14917 11384 18111 11386
rect 14917 11328 14922 11384
rect 14978 11328 18050 11384
rect 18106 11328 18111 11384
rect 14917 11326 18111 11328
rect 14917 11323 14983 11326
rect 18045 11323 18111 11326
rect 2773 11250 2839 11253
rect 13905 11250 13971 11253
rect 2773 11248 13971 11250
rect 2773 11192 2778 11248
rect 2834 11192 13910 11248
rect 13966 11192 13971 11248
rect 2773 11190 13971 11192
rect 2773 11187 2839 11190
rect 13905 11187 13971 11190
rect 14733 11250 14799 11253
rect 16941 11250 17007 11253
rect 14733 11248 17007 11250
rect 14733 11192 14738 11248
rect 14794 11192 16946 11248
rect 17002 11192 17007 11248
rect 14733 11190 17007 11192
rect 14733 11187 14799 11190
rect 16941 11187 17007 11190
rect 2129 11114 2195 11117
rect 4613 11114 4679 11117
rect 2129 11112 4679 11114
rect 2129 11056 2134 11112
rect 2190 11056 4618 11112
rect 4674 11056 4679 11112
rect 2129 11054 4679 11056
rect 2129 11051 2195 11054
rect 4613 11051 4679 11054
rect 4889 11114 4955 11117
rect 10317 11114 10383 11117
rect 4889 11112 10383 11114
rect 4889 11056 4894 11112
rect 4950 11056 10322 11112
rect 10378 11056 10383 11112
rect 4889 11054 10383 11056
rect 4889 11051 4955 11054
rect 10317 11051 10383 11054
rect 15653 11114 15719 11117
rect 18965 11114 19031 11117
rect 15653 11112 19031 11114
rect 15653 11056 15658 11112
rect 15714 11056 18970 11112
rect 19026 11056 19031 11112
rect 15653 11054 19031 11056
rect 15653 11051 15719 11054
rect 18965 11051 19031 11054
rect 8385 10978 8451 10981
rect 8845 10978 8911 10981
rect 8385 10976 13186 10978
rect 8385 10920 8390 10976
rect 8446 10920 8850 10976
rect 8906 10920 13186 10976
rect 8385 10918 13186 10920
rect 8385 10915 8451 10918
rect 8845 10915 8911 10918
rect 5610 10912 5930 10913
rect 0 10842 480 10872
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 3509 10842 3575 10845
rect 0 10840 3575 10842
rect 0 10784 3514 10840
rect 3570 10784 3575 10840
rect 0 10782 3575 10784
rect 0 10752 480 10782
rect 3509 10779 3575 10782
rect 12801 10842 12867 10845
rect 12985 10842 13051 10845
rect 12801 10840 13051 10842
rect 12801 10784 12806 10840
rect 12862 10784 12990 10840
rect 13046 10784 13051 10840
rect 12801 10782 13051 10784
rect 12801 10779 12867 10782
rect 12985 10779 13051 10782
rect 13126 10709 13186 10918
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 3969 10706 4035 10709
rect 12985 10706 13051 10709
rect 3969 10704 13051 10706
rect 3969 10648 3974 10704
rect 4030 10648 12990 10704
rect 13046 10648 13051 10704
rect 3969 10646 13051 10648
rect 13126 10706 13235 10709
rect 15929 10706 15995 10709
rect 13126 10704 15995 10706
rect 13126 10648 13174 10704
rect 13230 10648 15934 10704
rect 15990 10648 15995 10704
rect 13126 10646 15995 10648
rect 3969 10643 4035 10646
rect 12985 10643 13051 10646
rect 13169 10643 13235 10646
rect 15929 10643 15995 10646
rect 1853 10570 1919 10573
rect 13813 10570 13879 10573
rect 1853 10568 13879 10570
rect 1853 10512 1858 10568
rect 1914 10512 13818 10568
rect 13874 10512 13879 10568
rect 1853 10510 13879 10512
rect 1853 10507 1919 10510
rect 13813 10507 13879 10510
rect 3417 10436 3483 10437
rect 3366 10372 3372 10436
rect 3436 10434 3483 10436
rect 3436 10432 3528 10434
rect 3478 10376 3528 10432
rect 3436 10374 3528 10376
rect 3436 10372 3483 10374
rect 11094 10372 11100 10436
rect 11164 10434 11170 10436
rect 13813 10434 13879 10437
rect 11164 10432 13879 10434
rect 11164 10376 13818 10432
rect 13874 10376 13879 10432
rect 11164 10374 13879 10376
rect 11164 10372 11170 10374
rect 3417 10371 3483 10372
rect 13813 10371 13879 10374
rect 14365 10434 14431 10437
rect 17401 10434 17467 10437
rect 14365 10432 17467 10434
rect 14365 10376 14370 10432
rect 14426 10376 17406 10432
rect 17462 10376 17467 10432
rect 14365 10374 17467 10376
rect 14365 10371 14431 10374
rect 17401 10371 17467 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 3601 10298 3667 10301
rect 5993 10298 6059 10301
rect 3601 10296 6059 10298
rect 3601 10240 3606 10296
rect 3662 10240 5998 10296
rect 6054 10240 6059 10296
rect 3601 10238 6059 10240
rect 3601 10235 3667 10238
rect 5993 10235 6059 10238
rect 12985 10298 13051 10301
rect 18045 10298 18111 10301
rect 12985 10296 18111 10298
rect 12985 10240 12990 10296
rect 13046 10240 18050 10296
rect 18106 10240 18111 10296
rect 12985 10238 18111 10240
rect 12985 10235 13051 10238
rect 18045 10235 18111 10238
rect 0 10162 480 10192
rect 3049 10162 3115 10165
rect 0 10160 3115 10162
rect 0 10104 3054 10160
rect 3110 10104 3115 10160
rect 0 10102 3115 10104
rect 0 10072 480 10102
rect 3049 10099 3115 10102
rect 3417 10162 3483 10165
rect 14181 10162 14247 10165
rect 3417 10160 14247 10162
rect 3417 10104 3422 10160
rect 3478 10104 14186 10160
rect 14242 10104 14247 10160
rect 3417 10102 14247 10104
rect 3417 10099 3483 10102
rect 14181 10099 14247 10102
rect 1393 10026 1459 10029
rect 13905 10026 13971 10029
rect 17033 10026 17099 10029
rect 1393 10024 13971 10026
rect 1393 9968 1398 10024
rect 1454 9968 13910 10024
rect 13966 9968 13971 10024
rect 1393 9966 13971 9968
rect 1393 9963 1459 9966
rect 13905 9963 13971 9966
rect 14782 10024 17099 10026
rect 14782 9968 17038 10024
rect 17094 9968 17099 10024
rect 14782 9966 17099 9968
rect 5993 9890 6059 9893
rect 14549 9890 14615 9893
rect 5993 9888 14615 9890
rect 5993 9832 5998 9888
rect 6054 9832 14554 9888
rect 14610 9832 14615 9888
rect 5993 9830 14615 9832
rect 5993 9827 6059 9830
rect 14549 9827 14615 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 9990 9692 9996 9756
rect 10060 9754 10066 9756
rect 10225 9754 10291 9757
rect 10060 9752 10291 9754
rect 10060 9696 10230 9752
rect 10286 9696 10291 9752
rect 10060 9694 10291 9696
rect 10060 9692 10066 9694
rect 10225 9691 10291 9694
rect 10869 9754 10935 9757
rect 11789 9754 11855 9757
rect 10869 9752 11855 9754
rect 10869 9696 10874 9752
rect 10930 9696 11794 9752
rect 11850 9696 11855 9752
rect 10869 9694 11855 9696
rect 10869 9691 10935 9694
rect 11789 9691 11855 9694
rect 12801 9754 12867 9757
rect 14782 9754 14842 9966
rect 17033 9963 17099 9966
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 12801 9752 14842 9754
rect 12801 9696 12806 9752
rect 12862 9696 14842 9752
rect 12801 9694 14842 9696
rect 12801 9691 12867 9694
rect 0 9618 480 9648
rect 1669 9618 1735 9621
rect 0 9616 1735 9618
rect 0 9560 1674 9616
rect 1730 9560 1735 9616
rect 0 9558 1735 9560
rect 0 9528 480 9558
rect 1669 9555 1735 9558
rect 9622 9556 9628 9620
rect 9692 9618 9698 9620
rect 10225 9618 10291 9621
rect 9692 9616 10291 9618
rect 9692 9560 10230 9616
rect 10286 9560 10291 9616
rect 9692 9558 10291 9560
rect 9692 9556 9698 9558
rect 10225 9555 10291 9558
rect 16297 9618 16363 9621
rect 18873 9618 18939 9621
rect 19333 9618 19399 9621
rect 16297 9616 19399 9618
rect 16297 9560 16302 9616
rect 16358 9560 18878 9616
rect 18934 9560 19338 9616
rect 19394 9560 19399 9616
rect 16297 9558 19399 9560
rect 16297 9555 16363 9558
rect 18873 9555 18939 9558
rect 19333 9555 19399 9558
rect 3233 9482 3299 9485
rect 7925 9482 7991 9485
rect 3233 9480 7991 9482
rect 3233 9424 3238 9480
rect 3294 9424 7930 9480
rect 7986 9424 7991 9480
rect 3233 9422 7991 9424
rect 3233 9419 3299 9422
rect 7925 9419 7991 9422
rect 8385 9482 8451 9485
rect 11973 9482 12039 9485
rect 8385 9480 12039 9482
rect 8385 9424 8390 9480
rect 8446 9424 11978 9480
rect 12034 9424 12039 9480
rect 8385 9422 12039 9424
rect 8385 9419 8451 9422
rect 11973 9419 12039 9422
rect 8017 9346 8083 9349
rect 10133 9346 10199 9349
rect 8017 9344 10199 9346
rect 8017 9288 8022 9344
rect 8078 9288 10138 9344
rect 10194 9288 10199 9344
rect 8017 9286 10199 9288
rect 8017 9283 8083 9286
rect 10133 9283 10199 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 3049 9210 3115 9213
rect 10041 9210 10107 9213
rect 3049 9208 10107 9210
rect 3049 9152 3054 9208
rect 3110 9152 10046 9208
rect 10102 9152 10107 9208
rect 3049 9150 10107 9152
rect 3049 9147 3115 9150
rect 10041 9147 10107 9150
rect 0 9074 480 9104
rect 3233 9074 3299 9077
rect 0 9072 3299 9074
rect 0 9016 3238 9072
rect 3294 9016 3299 9072
rect 0 9014 3299 9016
rect 0 8984 480 9014
rect 3233 9011 3299 9014
rect 8017 9074 8083 9077
rect 10041 9074 10107 9077
rect 14917 9074 14983 9077
rect 8017 9072 14983 9074
rect 8017 9016 8022 9072
rect 8078 9016 10046 9072
rect 10102 9016 14922 9072
rect 14978 9016 14983 9072
rect 8017 9014 14983 9016
rect 8017 9011 8083 9014
rect 10041 9011 10107 9014
rect 14917 9011 14983 9014
rect 10133 8938 10199 8941
rect 14549 8938 14615 8941
rect 10133 8936 14615 8938
rect 10133 8880 10138 8936
rect 10194 8880 14554 8936
rect 14610 8880 14615 8936
rect 10133 8878 14615 8880
rect 10133 8875 10199 8878
rect 14549 8875 14615 8878
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 3141 8666 3207 8669
rect 3141 8664 5274 8666
rect 3141 8608 3146 8664
rect 3202 8608 5274 8664
rect 3141 8606 5274 8608
rect 3141 8603 3207 8606
rect 0 8530 480 8560
rect 4981 8530 5047 8533
rect 0 8528 5047 8530
rect 0 8472 4986 8528
rect 5042 8472 5047 8528
rect 0 8470 5047 8472
rect 5214 8530 5274 8606
rect 9857 8530 9923 8533
rect 10041 8530 10107 8533
rect 5214 8528 10107 8530
rect 5214 8472 9862 8528
rect 9918 8472 10046 8528
rect 10102 8472 10107 8528
rect 5214 8470 10107 8472
rect 0 8440 480 8470
rect 4981 8467 5047 8470
rect 9857 8467 9923 8470
rect 10041 8467 10107 8470
rect 11881 8530 11947 8533
rect 12985 8530 13051 8533
rect 14273 8530 14339 8533
rect 17953 8530 18019 8533
rect 11881 8528 18019 8530
rect 11881 8472 11886 8528
rect 11942 8472 12990 8528
rect 13046 8472 14278 8528
rect 14334 8472 17958 8528
rect 18014 8472 18019 8528
rect 11881 8470 18019 8472
rect 11881 8467 11947 8470
rect 12985 8467 13051 8470
rect 14273 8467 14339 8470
rect 17953 8467 18019 8470
rect 3509 8394 3575 8397
rect 15929 8394 15995 8397
rect 3509 8392 15995 8394
rect 3509 8336 3514 8392
rect 3570 8336 15934 8392
rect 15990 8336 15995 8392
rect 3509 8334 15995 8336
rect 3509 8331 3575 8334
rect 15929 8331 15995 8334
rect 12433 8258 12499 8261
rect 18413 8258 18479 8261
rect 12433 8256 18479 8258
rect 12433 8200 12438 8256
rect 12494 8200 18418 8256
rect 18474 8200 18479 8256
rect 12433 8198 18479 8200
rect 12433 8195 12499 8198
rect 18413 8195 18479 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 0 7850 480 7880
rect 565 7850 631 7853
rect 0 7848 631 7850
rect 0 7792 570 7848
rect 626 7792 631 7848
rect 0 7790 631 7792
rect 0 7760 480 7790
rect 565 7787 631 7790
rect 9581 7850 9647 7853
rect 15285 7850 15351 7853
rect 15469 7852 15535 7853
rect 15469 7850 15516 7852
rect 9581 7848 15351 7850
rect 9581 7792 9586 7848
rect 9642 7792 15290 7848
rect 15346 7792 15351 7848
rect 9581 7790 15351 7792
rect 15424 7848 15516 7850
rect 15424 7792 15474 7848
rect 15424 7790 15516 7792
rect 9581 7787 9647 7790
rect 15285 7787 15351 7790
rect 15469 7788 15516 7790
rect 15580 7788 15586 7852
rect 15469 7787 15535 7788
rect 9489 7714 9555 7717
rect 13169 7714 13235 7717
rect 9489 7712 13235 7714
rect 9489 7656 9494 7712
rect 9550 7656 13174 7712
rect 13230 7656 13235 7712
rect 9489 7654 13235 7656
rect 9489 7651 9555 7654
rect 13169 7651 13235 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 2957 7578 3023 7581
rect 5165 7578 5231 7581
rect 2957 7576 5231 7578
rect 2957 7520 2962 7576
rect 3018 7520 5170 7576
rect 5226 7520 5231 7576
rect 2957 7518 5231 7520
rect 2957 7515 3023 7518
rect 5165 7515 5231 7518
rect 6085 7578 6151 7581
rect 8385 7578 8451 7581
rect 6085 7576 8451 7578
rect 6085 7520 6090 7576
rect 6146 7520 8390 7576
rect 8446 7520 8451 7576
rect 6085 7518 8451 7520
rect 6085 7515 6151 7518
rect 8385 7515 8451 7518
rect 10685 7442 10751 7445
rect 4846 7440 10751 7442
rect 4846 7384 10690 7440
rect 10746 7384 10751 7440
rect 4846 7382 10751 7384
rect 0 7306 480 7336
rect 4846 7306 4906 7382
rect 10685 7379 10751 7382
rect 10961 7442 11027 7445
rect 18505 7442 18571 7445
rect 10961 7440 18571 7442
rect 10961 7384 10966 7440
rect 11022 7384 18510 7440
rect 18566 7384 18571 7440
rect 10961 7382 18571 7384
rect 10961 7379 11027 7382
rect 18505 7379 18571 7382
rect 0 7246 4906 7306
rect 6821 7306 6887 7309
rect 22277 7306 22343 7309
rect 6821 7304 22343 7306
rect 6821 7248 6826 7304
rect 6882 7248 22282 7304
rect 22338 7248 22343 7304
rect 6821 7246 22343 7248
rect 0 7216 480 7246
rect 6821 7243 6887 7246
rect 22277 7243 22343 7246
rect 4521 7170 4587 7173
rect 9673 7170 9739 7173
rect 4521 7168 9739 7170
rect 4521 7112 4526 7168
rect 4582 7112 9678 7168
rect 9734 7112 9739 7168
rect 4521 7110 9739 7112
rect 4521 7107 4587 7110
rect 9673 7107 9739 7110
rect 10685 7170 10751 7173
rect 18321 7170 18387 7173
rect 19241 7170 19307 7173
rect 10685 7168 19307 7170
rect 10685 7112 10690 7168
rect 10746 7112 18326 7168
rect 18382 7112 19246 7168
rect 19302 7112 19307 7168
rect 10685 7110 19307 7112
rect 10685 7107 10751 7110
rect 18321 7107 18387 7110
rect 19241 7107 19307 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 3417 7034 3483 7037
rect 9765 7034 9831 7037
rect 3417 7032 9831 7034
rect 3417 6976 3422 7032
rect 3478 6976 9770 7032
rect 9826 6976 9831 7032
rect 3417 6974 9831 6976
rect 3417 6971 3483 6974
rect 9765 6971 9831 6974
rect 14641 7034 14707 7037
rect 19333 7034 19399 7037
rect 14641 7032 19399 7034
rect 14641 6976 14646 7032
rect 14702 6976 19338 7032
rect 19394 6976 19399 7032
rect 14641 6974 19399 6976
rect 14641 6971 14707 6974
rect 19333 6971 19399 6974
rect 5533 6898 5599 6901
rect 8477 6898 8543 6901
rect 5533 6896 8543 6898
rect 5533 6840 5538 6896
rect 5594 6840 8482 6896
rect 8538 6840 8543 6896
rect 5533 6838 8543 6840
rect 5533 6835 5599 6838
rect 8477 6835 8543 6838
rect 0 6762 480 6792
rect 3734 6762 3740 6764
rect 0 6702 3740 6762
rect 0 6672 480 6702
rect 3734 6700 3740 6702
rect 3804 6700 3810 6764
rect 3969 6762 4035 6765
rect 8385 6762 8451 6765
rect 3969 6760 8451 6762
rect 3969 6704 3974 6760
rect 4030 6704 8390 6760
rect 8446 6704 8451 6760
rect 3969 6702 8451 6704
rect 3969 6699 4035 6702
rect 8385 6699 8451 6702
rect 12801 6762 12867 6765
rect 22185 6762 22251 6765
rect 12801 6760 22251 6762
rect 12801 6704 12806 6760
rect 12862 6704 22190 6760
rect 22246 6704 22251 6760
rect 12801 6702 22251 6704
rect 12801 6699 12867 6702
rect 22185 6699 22251 6702
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 18045 6490 18111 6493
rect 20897 6490 20963 6493
rect 18045 6488 20963 6490
rect 18045 6432 18050 6488
rect 18106 6432 20902 6488
rect 20958 6432 20963 6488
rect 18045 6430 20963 6432
rect 18045 6427 18111 6430
rect 20897 6427 20963 6430
rect 4337 6354 4403 6357
rect 7189 6354 7255 6357
rect 10225 6354 10291 6357
rect 4337 6352 10291 6354
rect 4337 6296 4342 6352
rect 4398 6296 7194 6352
rect 7250 6296 10230 6352
rect 10286 6296 10291 6352
rect 4337 6294 10291 6296
rect 4337 6291 4403 6294
rect 7189 6291 7255 6294
rect 10225 6291 10291 6294
rect 12985 6354 13051 6357
rect 18597 6354 18663 6357
rect 19425 6354 19491 6357
rect 12985 6352 19491 6354
rect 12985 6296 12990 6352
rect 13046 6296 18602 6352
rect 18658 6296 19430 6352
rect 19486 6296 19491 6352
rect 12985 6294 19491 6296
rect 12985 6291 13051 6294
rect 18597 6291 18663 6294
rect 19425 6291 19491 6294
rect 9857 6218 9923 6221
rect 2776 6216 9923 6218
rect 2776 6160 9862 6216
rect 9918 6160 9923 6216
rect 2776 6158 9923 6160
rect 2776 6116 2836 6158
rect 9857 6155 9923 6158
rect 10041 6218 10107 6221
rect 16849 6218 16915 6221
rect 10041 6216 16915 6218
rect 10041 6160 10046 6216
rect 10102 6160 16854 6216
rect 16910 6160 16915 6216
rect 10041 6158 16915 6160
rect 10041 6155 10107 6158
rect 16849 6155 16915 6158
rect 0 6082 480 6112
rect 2684 6082 2836 6116
rect 0 6056 2836 6082
rect 4061 6082 4127 6085
rect 7925 6082 7991 6085
rect 4061 6080 7991 6082
rect 0 6022 2744 6056
rect 4061 6024 4066 6080
rect 4122 6024 7930 6080
rect 7986 6024 7991 6080
rect 4061 6022 7991 6024
rect 0 5992 480 6022
rect 4061 6019 4127 6022
rect 7925 6019 7991 6022
rect 10961 6082 11027 6085
rect 12893 6082 12959 6085
rect 10961 6080 12959 6082
rect 10961 6024 10966 6080
rect 11022 6024 12898 6080
rect 12954 6024 12959 6080
rect 10961 6022 12959 6024
rect 10961 6019 11027 6022
rect 12893 6019 12959 6022
rect 14273 6082 14339 6085
rect 18229 6082 18295 6085
rect 14273 6080 18295 6082
rect 14273 6024 14278 6080
rect 14334 6024 18234 6080
rect 18290 6024 18295 6080
rect 14273 6022 18295 6024
rect 14273 6019 14339 6022
rect 18229 6019 18295 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 7281 5946 7347 5949
rect 9857 5946 9923 5949
rect 7281 5944 9923 5946
rect 7281 5888 7286 5944
rect 7342 5888 9862 5944
rect 9918 5888 9923 5944
rect 7281 5886 9923 5888
rect 7281 5883 7347 5886
rect 9857 5883 9923 5886
rect 13629 5946 13695 5949
rect 19425 5946 19491 5949
rect 13629 5944 19491 5946
rect 13629 5888 13634 5944
rect 13690 5888 19430 5944
rect 19486 5888 19491 5944
rect 13629 5886 19491 5888
rect 13629 5883 13695 5886
rect 19425 5883 19491 5886
rect 1577 5810 1643 5813
rect 8293 5810 8359 5813
rect 1577 5808 8359 5810
rect 1577 5752 1582 5808
rect 1638 5752 8298 5808
rect 8354 5752 8359 5808
rect 1577 5750 8359 5752
rect 1577 5747 1643 5750
rect 8293 5747 8359 5750
rect 13445 5810 13511 5813
rect 18321 5810 18387 5813
rect 13445 5808 18387 5810
rect 13445 5752 13450 5808
rect 13506 5752 18326 5808
rect 18382 5752 18387 5808
rect 13445 5750 18387 5752
rect 13445 5747 13511 5750
rect 18321 5747 18387 5750
rect 2221 5674 2287 5677
rect 2086 5672 2287 5674
rect 2086 5616 2226 5672
rect 2282 5616 2287 5672
rect 2086 5614 2287 5616
rect 0 5538 480 5568
rect 2086 5538 2146 5614
rect 2221 5611 2287 5614
rect 2773 5674 2839 5677
rect 2957 5674 3023 5677
rect 9029 5674 9095 5677
rect 2773 5672 9095 5674
rect 2773 5616 2778 5672
rect 2834 5616 2962 5672
rect 3018 5616 9034 5672
rect 9090 5616 9095 5672
rect 2773 5614 9095 5616
rect 2773 5611 2839 5614
rect 2957 5611 3023 5614
rect 9029 5611 9095 5614
rect 11237 5674 11303 5677
rect 13905 5674 13971 5677
rect 15193 5674 15259 5677
rect 11237 5672 13971 5674
rect 11237 5616 11242 5672
rect 11298 5616 13910 5672
rect 13966 5616 13971 5672
rect 11237 5614 13971 5616
rect 11237 5611 11303 5614
rect 13905 5611 13971 5614
rect 14782 5672 15259 5674
rect 14782 5616 15198 5672
rect 15254 5616 15259 5672
rect 14782 5614 15259 5616
rect 0 5478 2146 5538
rect 6545 5538 6611 5541
rect 7833 5538 7899 5541
rect 6545 5536 7899 5538
rect 6545 5480 6550 5536
rect 6606 5480 7838 5536
rect 7894 5480 7899 5536
rect 6545 5478 7899 5480
rect 0 5448 480 5478
rect 6545 5475 6611 5478
rect 7833 5475 7899 5478
rect 9581 5538 9647 5541
rect 14782 5538 14842 5614
rect 15193 5611 15259 5614
rect 15837 5674 15903 5677
rect 17953 5674 18019 5677
rect 15837 5672 18019 5674
rect 15837 5616 15842 5672
rect 15898 5616 17958 5672
rect 18014 5616 18019 5672
rect 15837 5614 18019 5616
rect 15837 5611 15903 5614
rect 17953 5611 18019 5614
rect 9581 5536 14842 5538
rect 9581 5480 9586 5536
rect 9642 5480 14842 5536
rect 9581 5478 14842 5480
rect 15377 5538 15443 5541
rect 16941 5538 17007 5541
rect 15377 5536 17007 5538
rect 15377 5480 15382 5536
rect 15438 5480 16946 5536
rect 17002 5480 17007 5536
rect 15377 5478 17007 5480
rect 9581 5475 9647 5478
rect 15377 5475 15443 5478
rect 16941 5475 17007 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 9949 5404 10015 5405
rect 9949 5400 9996 5404
rect 10060 5402 10066 5404
rect 17401 5402 17467 5405
rect 21633 5402 21699 5405
rect 9949 5344 9954 5400
rect 9949 5340 9996 5344
rect 10060 5342 10106 5402
rect 17401 5400 21699 5402
rect 17401 5344 17406 5400
rect 17462 5344 21638 5400
rect 21694 5344 21699 5400
rect 17401 5342 21699 5344
rect 10060 5340 10066 5342
rect 9949 5339 10015 5340
rect 17401 5339 17467 5342
rect 21633 5339 21699 5342
rect 8569 5266 8635 5269
rect 17769 5266 17835 5269
rect 8569 5264 17835 5266
rect 8569 5208 8574 5264
rect 8630 5208 17774 5264
rect 17830 5208 17835 5264
rect 8569 5206 17835 5208
rect 8569 5203 8635 5206
rect 17769 5203 17835 5206
rect 18505 5266 18571 5269
rect 22369 5266 22435 5269
rect 18505 5264 22435 5266
rect 18505 5208 18510 5264
rect 18566 5208 22374 5264
rect 22430 5208 22435 5264
rect 18505 5206 22435 5208
rect 18505 5203 18571 5206
rect 22369 5203 22435 5206
rect 4153 5130 4219 5133
rect 6269 5130 6335 5133
rect 15653 5130 15719 5133
rect 4153 5128 15719 5130
rect 4153 5072 4158 5128
rect 4214 5072 6274 5128
rect 6330 5072 15658 5128
rect 15714 5072 15719 5128
rect 4153 5070 15719 5072
rect 4153 5067 4219 5070
rect 6269 5067 6335 5070
rect 15653 5067 15719 5070
rect 16849 5130 16915 5133
rect 22737 5130 22803 5133
rect 16849 5128 22803 5130
rect 16849 5072 16854 5128
rect 16910 5072 22742 5128
rect 22798 5072 22803 5128
rect 16849 5070 22803 5072
rect 16849 5067 16915 5070
rect 22737 5067 22803 5070
rect 0 4994 480 5024
rect 1485 4994 1551 4997
rect 0 4992 1551 4994
rect 0 4936 1490 4992
rect 1546 4936 1551 4992
rect 0 4934 1551 4936
rect 0 4904 480 4934
rect 1485 4931 1551 4934
rect 3877 4994 3943 4997
rect 9622 4994 9628 4996
rect 3877 4992 9628 4994
rect 3877 4936 3882 4992
rect 3938 4936 9628 4992
rect 3877 4934 9628 4936
rect 3877 4931 3943 4934
rect 9622 4932 9628 4934
rect 9692 4932 9698 4996
rect 14181 4994 14247 4997
rect 16389 4994 16455 4997
rect 14181 4992 16455 4994
rect 14181 4936 14186 4992
rect 14242 4936 16394 4992
rect 16450 4936 16455 4992
rect 14181 4934 16455 4936
rect 14181 4931 14247 4934
rect 16389 4931 16455 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 3601 4858 3667 4861
rect 5993 4858 6059 4861
rect 3601 4856 6059 4858
rect 3601 4800 3606 4856
rect 3662 4800 5998 4856
rect 6054 4800 6059 4856
rect 3601 4798 6059 4800
rect 3601 4795 3667 4798
rect 5993 4795 6059 4798
rect 6637 4858 6703 4861
rect 9305 4858 9371 4861
rect 6637 4856 9371 4858
rect 6637 4800 6642 4856
rect 6698 4800 9310 4856
rect 9366 4800 9371 4856
rect 6637 4798 9371 4800
rect 6637 4795 6703 4798
rect 9305 4795 9371 4798
rect 13169 4858 13235 4861
rect 16021 4858 16087 4861
rect 13169 4856 19488 4858
rect 13169 4800 13174 4856
rect 13230 4800 16026 4856
rect 16082 4800 19488 4856
rect 13169 4798 19488 4800
rect 13169 4795 13235 4798
rect 16021 4795 16087 4798
rect 2773 4722 2839 4725
rect 10041 4722 10107 4725
rect 2773 4720 10107 4722
rect 2773 4664 2778 4720
rect 2834 4664 10046 4720
rect 10102 4664 10107 4720
rect 2773 4662 10107 4664
rect 2773 4659 2839 4662
rect 10041 4659 10107 4662
rect 10501 4722 10567 4725
rect 17493 4722 17559 4725
rect 10501 4720 17559 4722
rect 10501 4664 10506 4720
rect 10562 4664 17498 4720
rect 17554 4664 17559 4720
rect 10501 4662 17559 4664
rect 19428 4722 19488 4798
rect 21173 4722 21239 4725
rect 19428 4720 21239 4722
rect 19428 4664 21178 4720
rect 21234 4664 21239 4720
rect 19428 4662 21239 4664
rect 10501 4659 10567 4662
rect 17493 4659 17559 4662
rect 21173 4659 21239 4662
rect 21633 4722 21699 4725
rect 27520 4722 28000 4752
rect 21633 4720 28000 4722
rect 21633 4664 21638 4720
rect 21694 4664 28000 4720
rect 21633 4662 28000 4664
rect 21633 4659 21699 4662
rect 27520 4632 28000 4662
rect 2405 4586 2471 4589
rect 9949 4586 10015 4589
rect 2405 4584 10015 4586
rect 2405 4528 2410 4584
rect 2466 4528 9954 4584
rect 10010 4528 10015 4584
rect 2405 4526 10015 4528
rect 2405 4523 2471 4526
rect 9949 4523 10015 4526
rect 15469 4586 15535 4589
rect 24209 4586 24275 4589
rect 15469 4584 24275 4586
rect 15469 4528 15474 4584
rect 15530 4528 24214 4584
rect 24270 4528 24275 4584
rect 15469 4526 24275 4528
rect 15469 4523 15535 4526
rect 24209 4523 24275 4526
rect 0 4450 480 4480
rect 4061 4450 4127 4453
rect 0 4448 4127 4450
rect 0 4392 4066 4448
rect 4122 4392 4127 4448
rect 0 4390 4127 4392
rect 0 4360 480 4390
rect 4061 4387 4127 4390
rect 7741 4450 7807 4453
rect 12985 4450 13051 4453
rect 7741 4448 13051 4450
rect 7741 4392 7746 4448
rect 7802 4392 12990 4448
rect 13046 4392 13051 4448
rect 7741 4390 13051 4392
rect 7741 4387 7807 4390
rect 12985 4387 13051 4390
rect 17033 4450 17099 4453
rect 19057 4450 19123 4453
rect 17033 4448 19123 4450
rect 17033 4392 17038 4448
rect 17094 4392 19062 4448
rect 19118 4392 19123 4448
rect 17033 4390 19123 4392
rect 17033 4387 17099 4390
rect 19057 4387 19123 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 841 4314 907 4317
rect 5441 4314 5507 4317
rect 841 4312 5507 4314
rect 841 4256 846 4312
rect 902 4256 5446 4312
rect 5502 4256 5507 4312
rect 841 4254 5507 4256
rect 841 4251 907 4254
rect 5441 4251 5507 4254
rect 7557 4314 7623 4317
rect 9305 4314 9371 4317
rect 19333 4314 19399 4317
rect 7557 4312 9138 4314
rect 7557 4256 7562 4312
rect 7618 4256 9138 4312
rect 7557 4254 9138 4256
rect 7557 4251 7623 4254
rect 1393 4178 1459 4181
rect 8845 4178 8911 4181
rect 1393 4176 8911 4178
rect 1393 4120 1398 4176
rect 1454 4120 8850 4176
rect 8906 4120 8911 4176
rect 1393 4118 8911 4120
rect 9078 4178 9138 4254
rect 9305 4312 13692 4314
rect 9305 4256 9310 4312
rect 9366 4256 13692 4312
rect 9305 4254 13692 4256
rect 9305 4251 9371 4254
rect 13632 4181 13692 4254
rect 15334 4312 19399 4314
rect 15334 4256 19338 4312
rect 19394 4256 19399 4312
rect 15334 4254 19399 4256
rect 13169 4178 13235 4181
rect 9078 4176 13235 4178
rect 9078 4120 13174 4176
rect 13230 4120 13235 4176
rect 9078 4118 13235 4120
rect 1393 4115 1459 4118
rect 8845 4115 8911 4118
rect 13169 4115 13235 4118
rect 13629 4178 13695 4181
rect 15334 4178 15394 4254
rect 19333 4251 19399 4254
rect 18965 4178 19031 4181
rect 13629 4176 15394 4178
rect 13629 4120 13634 4176
rect 13690 4120 15394 4176
rect 13629 4118 15394 4120
rect 17910 4176 19031 4178
rect 17910 4120 18970 4176
rect 19026 4120 19031 4176
rect 17910 4118 19031 4120
rect 13629 4115 13695 4118
rect 2497 4042 2563 4045
rect 4153 4042 4219 4045
rect 8017 4042 8083 4045
rect 8569 4042 8635 4045
rect 2497 4040 6976 4042
rect 2497 3984 2502 4040
rect 2558 3984 4158 4040
rect 4214 3984 6976 4040
rect 2497 3982 6976 3984
rect 2497 3979 2563 3982
rect 4153 3979 4219 3982
rect 2681 3906 2747 3909
rect 4613 3906 4679 3909
rect 2681 3904 4679 3906
rect 2681 3848 2686 3904
rect 2742 3848 4618 3904
rect 4674 3848 4679 3904
rect 2681 3846 4679 3848
rect 2681 3843 2747 3846
rect 4613 3843 4679 3846
rect 0 3770 480 3800
rect 3417 3770 3483 3773
rect 0 3768 3483 3770
rect 0 3712 3422 3768
rect 3478 3712 3483 3768
rect 0 3710 3483 3712
rect 0 3680 480 3710
rect 3417 3707 3483 3710
rect 3601 3770 3667 3773
rect 5533 3770 5599 3773
rect 3601 3768 5599 3770
rect 3601 3712 3606 3768
rect 3662 3712 5538 3768
rect 5594 3712 5599 3768
rect 3601 3710 5599 3712
rect 6916 3770 6976 3982
rect 8017 4040 8635 4042
rect 8017 3984 8022 4040
rect 8078 3984 8574 4040
rect 8630 3984 8635 4040
rect 8017 3982 8635 3984
rect 8017 3979 8083 3982
rect 8569 3979 8635 3982
rect 9305 4042 9371 4045
rect 10041 4042 10107 4045
rect 11053 4042 11119 4045
rect 9305 4040 11119 4042
rect 9305 3984 9310 4040
rect 9366 3984 10046 4040
rect 10102 3984 11058 4040
rect 11114 3984 11119 4040
rect 9305 3982 11119 3984
rect 9305 3979 9371 3982
rect 10041 3979 10107 3982
rect 11053 3979 11119 3982
rect 11237 4042 11303 4045
rect 17910 4042 17970 4118
rect 18965 4115 19031 4118
rect 11237 4040 17970 4042
rect 11237 3984 11242 4040
rect 11298 3984 17970 4040
rect 11237 3982 17970 3984
rect 18045 4042 18111 4045
rect 22093 4042 22159 4045
rect 18045 4040 22159 4042
rect 18045 3984 18050 4040
rect 18106 3984 22098 4040
rect 22154 3984 22159 4040
rect 18045 3982 22159 3984
rect 11237 3979 11303 3982
rect 18045 3979 18111 3982
rect 22093 3979 22159 3982
rect 23473 4042 23539 4045
rect 25313 4042 25379 4045
rect 23473 4040 25379 4042
rect 23473 3984 23478 4040
rect 23534 3984 25318 4040
rect 25374 3984 25379 4040
rect 23473 3982 25379 3984
rect 23473 3979 23539 3982
rect 25313 3979 25379 3982
rect 7097 3906 7163 3909
rect 9213 3906 9279 3909
rect 7097 3904 9279 3906
rect 7097 3848 7102 3904
rect 7158 3848 9218 3904
rect 9274 3848 9279 3904
rect 7097 3846 9279 3848
rect 7097 3843 7163 3846
rect 9213 3843 9279 3846
rect 11237 3906 11303 3909
rect 18781 3906 18847 3909
rect 11237 3904 18847 3906
rect 11237 3848 11242 3904
rect 11298 3848 18786 3904
rect 18842 3848 18847 3904
rect 11237 3846 18847 3848
rect 11237 3843 11303 3846
rect 18781 3843 18847 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 9489 3770 9555 3773
rect 6916 3768 9555 3770
rect 6916 3712 9494 3768
rect 9550 3712 9555 3768
rect 6916 3710 9555 3712
rect 3601 3707 3667 3710
rect 5533 3707 5599 3710
rect 9489 3707 9555 3710
rect 1485 3634 1551 3637
rect 7189 3634 7255 3637
rect 1485 3632 7255 3634
rect 1485 3576 1490 3632
rect 1546 3576 7194 3632
rect 7250 3576 7255 3632
rect 1485 3574 7255 3576
rect 1485 3571 1551 3574
rect 7189 3571 7255 3574
rect 8753 3634 8819 3637
rect 9765 3634 9831 3637
rect 8753 3632 9831 3634
rect 8753 3576 8758 3632
rect 8814 3576 9770 3632
rect 9826 3576 9831 3632
rect 8753 3574 9831 3576
rect 8753 3571 8819 3574
rect 9765 3571 9831 3574
rect 14365 3634 14431 3637
rect 23657 3634 23723 3637
rect 14365 3632 23723 3634
rect 14365 3576 14370 3632
rect 14426 3576 23662 3632
rect 23718 3576 23723 3632
rect 14365 3574 23723 3576
rect 14365 3571 14431 3574
rect 23657 3571 23723 3574
rect 24209 3634 24275 3637
rect 26509 3634 26575 3637
rect 24209 3632 26575 3634
rect 24209 3576 24214 3632
rect 24270 3576 26514 3632
rect 26570 3576 26575 3632
rect 24209 3574 26575 3576
rect 24209 3571 24275 3574
rect 26509 3571 26575 3574
rect 289 3498 355 3501
rect 6637 3498 6703 3501
rect 289 3496 6703 3498
rect 289 3440 294 3496
rect 350 3440 6642 3496
rect 6698 3440 6703 3496
rect 289 3438 6703 3440
rect 289 3435 355 3438
rect 6637 3435 6703 3438
rect 8293 3498 8359 3501
rect 19149 3498 19215 3501
rect 8293 3496 19215 3498
rect 8293 3440 8298 3496
rect 8354 3440 19154 3496
rect 19210 3440 19215 3496
rect 8293 3438 19215 3440
rect 8293 3435 8359 3438
rect 19149 3435 19215 3438
rect 2405 3362 2471 3365
rect 4889 3362 4955 3365
rect 2405 3360 4955 3362
rect 2405 3304 2410 3360
rect 2466 3304 4894 3360
rect 4950 3304 4955 3360
rect 2405 3302 4955 3304
rect 2405 3299 2471 3302
rect 4889 3299 4955 3302
rect 8477 3362 8543 3365
rect 8477 3360 14842 3362
rect 8477 3304 8482 3360
rect 8538 3304 14842 3360
rect 8477 3302 14842 3304
rect 8477 3299 8543 3302
rect 5610 3296 5930 3297
rect 0 3226 480 3256
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 3141 3226 3207 3229
rect 0 3224 3207 3226
rect 0 3168 3146 3224
rect 3202 3168 3207 3224
rect 0 3166 3207 3168
rect 0 3136 480 3166
rect 3141 3163 3207 3166
rect 14181 3226 14247 3229
rect 14549 3226 14615 3229
rect 14181 3224 14615 3226
rect 14181 3168 14186 3224
rect 14242 3168 14554 3224
rect 14610 3168 14615 3224
rect 14181 3166 14615 3168
rect 14181 3163 14247 3166
rect 14549 3163 14615 3166
rect 4245 3090 4311 3093
rect 5441 3090 5507 3093
rect 11237 3090 11303 3093
rect 4245 3088 11303 3090
rect 4245 3032 4250 3088
rect 4306 3032 5446 3088
rect 5502 3032 11242 3088
rect 11298 3032 11303 3088
rect 4245 3030 11303 3032
rect 14782 3090 14842 3302
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 18505 3226 18571 3229
rect 23841 3226 23907 3229
rect 18505 3224 23907 3226
rect 18505 3168 18510 3224
rect 18566 3168 23846 3224
rect 23902 3168 23907 3224
rect 18505 3166 23907 3168
rect 18505 3163 18571 3166
rect 23841 3163 23907 3166
rect 17769 3090 17835 3093
rect 21633 3092 21699 3093
rect 14782 3088 17835 3090
rect 14782 3032 17774 3088
rect 17830 3032 17835 3088
rect 14782 3030 17835 3032
rect 4245 3027 4311 3030
rect 5441 3027 5507 3030
rect 11237 3027 11303 3030
rect 17769 3027 17835 3030
rect 21582 3028 21588 3092
rect 21652 3090 21699 3092
rect 21652 3088 21744 3090
rect 21694 3032 21744 3088
rect 21652 3030 21744 3032
rect 21652 3028 21699 3030
rect 21633 3027 21699 3028
rect 2865 2954 2931 2957
rect 7281 2954 7347 2957
rect 17401 2954 17467 2957
rect 2865 2952 17467 2954
rect 2865 2896 2870 2952
rect 2926 2896 7286 2952
rect 7342 2896 17406 2952
rect 17462 2896 17467 2952
rect 2865 2894 17467 2896
rect 2865 2891 2931 2894
rect 7281 2891 7347 2894
rect 17401 2891 17467 2894
rect 21265 2954 21331 2957
rect 23105 2954 23171 2957
rect 21265 2952 23171 2954
rect 21265 2896 21270 2952
rect 21326 2896 23110 2952
rect 23166 2896 23171 2952
rect 21265 2894 23171 2896
rect 21265 2891 21331 2894
rect 23105 2891 23171 2894
rect 3785 2818 3851 2821
rect 6177 2818 6243 2821
rect 3785 2816 6243 2818
rect 3785 2760 3790 2816
rect 3846 2760 6182 2816
rect 6238 2760 6243 2816
rect 3785 2758 6243 2760
rect 3785 2755 3851 2758
rect 6177 2755 6243 2758
rect 6729 2818 6795 2821
rect 9949 2820 10015 2821
rect 9949 2818 9996 2820
rect 6729 2816 7850 2818
rect 6729 2760 6734 2816
rect 6790 2760 7850 2816
rect 6729 2758 7850 2760
rect 9904 2816 9996 2818
rect 9904 2760 9954 2816
rect 9904 2758 9996 2760
rect 6729 2755 6795 2758
rect 0 2682 480 2712
rect 0 2622 1226 2682
rect 0 2592 480 2622
rect 1166 2410 1226 2622
rect 5257 2546 5323 2549
rect 6913 2546 6979 2549
rect 5257 2544 6979 2546
rect 5257 2488 5262 2544
rect 5318 2488 6918 2544
rect 6974 2488 6979 2544
rect 5257 2486 6979 2488
rect 7790 2546 7850 2758
rect 9949 2756 9996 2758
rect 10060 2756 10066 2820
rect 11421 2818 11487 2821
rect 16757 2818 16823 2821
rect 11421 2816 16823 2818
rect 11421 2760 11426 2816
rect 11482 2760 16762 2816
rect 16818 2760 16823 2816
rect 11421 2758 16823 2760
rect 9949 2755 10015 2756
rect 11421 2755 11487 2758
rect 16757 2755 16823 2758
rect 21817 2818 21883 2821
rect 23657 2818 23723 2821
rect 21817 2816 23723 2818
rect 21817 2760 21822 2816
rect 21878 2760 23662 2816
rect 23718 2760 23723 2816
rect 21817 2758 23723 2760
rect 21817 2755 21883 2758
rect 23657 2755 23723 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 13537 2682 13603 2685
rect 17125 2682 17191 2685
rect 13537 2680 17191 2682
rect 13537 2624 13542 2680
rect 13598 2624 17130 2680
rect 17186 2624 17191 2680
rect 13537 2622 17191 2624
rect 13537 2619 13603 2622
rect 17125 2619 17191 2622
rect 11973 2546 12039 2549
rect 7790 2544 12039 2546
rect 7790 2488 11978 2544
rect 12034 2488 12039 2544
rect 7790 2486 12039 2488
rect 5257 2483 5323 2486
rect 6913 2483 6979 2486
rect 11973 2483 12039 2486
rect 12157 2546 12223 2549
rect 14733 2546 14799 2549
rect 12157 2544 14799 2546
rect 12157 2488 12162 2544
rect 12218 2488 14738 2544
rect 14794 2488 14799 2544
rect 12157 2486 14799 2488
rect 12157 2483 12223 2486
rect 14733 2483 14799 2486
rect 14917 2546 14983 2549
rect 16665 2546 16731 2549
rect 14917 2544 16731 2546
rect 14917 2488 14922 2544
rect 14978 2488 16670 2544
rect 16726 2488 16731 2544
rect 14917 2486 16731 2488
rect 14917 2483 14983 2486
rect 16665 2483 16731 2486
rect 18965 2546 19031 2549
rect 24025 2546 24091 2549
rect 18965 2544 24091 2546
rect 18965 2488 18970 2544
rect 19026 2488 24030 2544
rect 24086 2488 24091 2544
rect 18965 2486 24091 2488
rect 18965 2483 19031 2486
rect 24025 2483 24091 2486
rect 11605 2410 11671 2413
rect 24761 2410 24827 2413
rect 1166 2350 7114 2410
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 0 2002 480 2032
rect 4061 2002 4127 2005
rect 0 2000 4127 2002
rect 0 1944 4066 2000
rect 4122 1944 4127 2000
rect 0 1942 4127 1944
rect 7054 2002 7114 2350
rect 11605 2408 24827 2410
rect 11605 2352 11610 2408
rect 11666 2352 24766 2408
rect 24822 2352 24827 2408
rect 11605 2350 24827 2352
rect 11605 2347 11671 2350
rect 24761 2347 24827 2350
rect 7281 2274 7347 2277
rect 14457 2274 14523 2277
rect 22185 2274 22251 2277
rect 7281 2272 14523 2274
rect 7281 2216 7286 2272
rect 7342 2216 14462 2272
rect 14518 2216 14523 2272
rect 7281 2214 14523 2216
rect 7281 2211 7347 2214
rect 14457 2211 14523 2214
rect 15334 2272 22251 2274
rect 15334 2216 22190 2272
rect 22246 2216 22251 2272
rect 15334 2214 22251 2216
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 10133 2138 10199 2141
rect 10133 2136 14842 2138
rect 10133 2080 10138 2136
rect 10194 2080 14842 2136
rect 10133 2078 14842 2080
rect 10133 2075 10199 2078
rect 14641 2002 14707 2005
rect 7054 2000 14707 2002
rect 7054 1944 14646 2000
rect 14702 1944 14707 2000
rect 7054 1942 14707 1944
rect 14782 2002 14842 2078
rect 15334 2002 15394 2214
rect 22185 2211 22251 2214
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 15469 2138 15535 2141
rect 15469 2136 24042 2138
rect 15469 2080 15474 2136
rect 15530 2080 24042 2136
rect 15469 2078 24042 2080
rect 15469 2075 15535 2078
rect 14782 1942 15394 2002
rect 16665 2002 16731 2005
rect 18965 2002 19031 2005
rect 16665 2000 19031 2002
rect 16665 1944 16670 2000
rect 16726 1944 18970 2000
rect 19026 1944 19031 2000
rect 16665 1942 19031 1944
rect 23982 2002 24042 2078
rect 27061 2002 27127 2005
rect 23982 2000 27127 2002
rect 23982 1944 27066 2000
rect 27122 1944 27127 2000
rect 23982 1942 27127 1944
rect 0 1912 480 1942
rect 4061 1939 4127 1942
rect 14641 1939 14707 1942
rect 16665 1939 16731 1942
rect 18965 1939 19031 1942
rect 27061 1939 27127 1942
rect 2037 1866 2103 1869
rect 14365 1866 14431 1869
rect 2037 1864 14431 1866
rect 2037 1808 2042 1864
rect 2098 1808 14370 1864
rect 14426 1808 14431 1864
rect 2037 1806 14431 1808
rect 2037 1803 2103 1806
rect 14365 1803 14431 1806
rect 4061 1730 4127 1733
rect 8477 1730 8543 1733
rect 4061 1728 8543 1730
rect 4061 1672 4066 1728
rect 4122 1672 8482 1728
rect 8538 1672 8543 1728
rect 4061 1670 8543 1672
rect 4061 1667 4127 1670
rect 8477 1667 8543 1670
rect 8661 1730 8727 1733
rect 12157 1730 12223 1733
rect 8661 1728 12223 1730
rect 8661 1672 8666 1728
rect 8722 1672 12162 1728
rect 12218 1672 12223 1728
rect 8661 1670 12223 1672
rect 8661 1667 8727 1670
rect 12157 1667 12223 1670
rect 18965 1730 19031 1733
rect 27613 1730 27679 1733
rect 18965 1728 27679 1730
rect 18965 1672 18970 1728
rect 19026 1672 27618 1728
rect 27674 1672 27679 1728
rect 18965 1670 27679 1672
rect 18965 1667 19031 1670
rect 27613 1667 27679 1670
rect 1945 1594 2011 1597
rect 3325 1594 3391 1597
rect 8937 1594 9003 1597
rect 15285 1594 15351 1597
rect 18873 1594 18939 1597
rect 1945 1592 15351 1594
rect 1945 1536 1950 1592
rect 2006 1536 3330 1592
rect 3386 1536 8942 1592
rect 8998 1536 15290 1592
rect 15346 1536 15351 1592
rect 1945 1534 15351 1536
rect 1945 1531 2011 1534
rect 3325 1531 3391 1534
rect 8937 1531 9003 1534
rect 15285 1531 15351 1534
rect 17174 1592 18939 1594
rect 17174 1536 18878 1592
rect 18934 1536 18939 1592
rect 17174 1534 18939 1536
rect 0 1458 480 1488
rect 2957 1458 3023 1461
rect 0 1456 3023 1458
rect 0 1400 2962 1456
rect 3018 1400 3023 1456
rect 0 1398 3023 1400
rect 0 1368 480 1398
rect 2957 1395 3023 1398
rect 8017 1458 8083 1461
rect 17174 1458 17234 1534
rect 18873 1531 18939 1534
rect 20069 1594 20135 1597
rect 25957 1594 26023 1597
rect 20069 1592 26023 1594
rect 20069 1536 20074 1592
rect 20130 1536 25962 1592
rect 26018 1536 26023 1592
rect 20069 1534 26023 1536
rect 20069 1531 20135 1534
rect 25957 1531 26023 1534
rect 8017 1456 17234 1458
rect 8017 1400 8022 1456
rect 8078 1400 17234 1456
rect 8017 1398 17234 1400
rect 17309 1458 17375 1461
rect 19609 1458 19675 1461
rect 17309 1456 19675 1458
rect 17309 1400 17314 1456
rect 17370 1400 19614 1456
rect 19670 1400 19675 1456
rect 17309 1398 19675 1400
rect 8017 1395 8083 1398
rect 17309 1395 17375 1398
rect 19609 1395 19675 1398
rect 20253 1458 20319 1461
rect 24209 1458 24275 1461
rect 20253 1456 24275 1458
rect 20253 1400 20258 1456
rect 20314 1400 24214 1456
rect 24270 1400 24275 1456
rect 20253 1398 24275 1400
rect 20253 1395 20319 1398
rect 24209 1395 24275 1398
rect 4153 1322 4219 1325
rect 7741 1322 7807 1325
rect 4153 1320 7807 1322
rect 4153 1264 4158 1320
rect 4214 1264 7746 1320
rect 7802 1264 7807 1320
rect 4153 1262 7807 1264
rect 4153 1259 4219 1262
rect 7741 1259 7807 1262
rect 7925 1322 7991 1325
rect 17217 1322 17283 1325
rect 7925 1320 17283 1322
rect 7925 1264 7930 1320
rect 7986 1264 17222 1320
rect 17278 1264 17283 1320
rect 7925 1262 17283 1264
rect 7925 1259 7991 1262
rect 17217 1259 17283 1262
rect 2313 1186 2379 1189
rect 19425 1186 19491 1189
rect 2313 1184 19491 1186
rect 2313 1128 2318 1184
rect 2374 1128 19430 1184
rect 19486 1128 19491 1184
rect 2313 1126 19491 1128
rect 2313 1123 2379 1126
rect 19425 1123 19491 1126
rect 1761 1050 1827 1053
rect 7741 1050 7807 1053
rect 20161 1050 20227 1053
rect 1761 1048 7666 1050
rect 1761 992 1766 1048
rect 1822 992 7666 1048
rect 1761 990 7666 992
rect 1761 987 1827 990
rect 0 914 480 944
rect 2773 914 2839 917
rect 0 912 2839 914
rect 0 856 2778 912
rect 2834 856 2839 912
rect 0 854 2839 856
rect 7606 914 7666 990
rect 7741 1048 20227 1050
rect 7741 992 7746 1048
rect 7802 992 20166 1048
rect 20222 992 20227 1048
rect 7741 990 20227 992
rect 7741 987 7807 990
rect 20161 987 20227 990
rect 19517 914 19583 917
rect 7606 912 19583 914
rect 7606 856 19522 912
rect 19578 856 19583 912
rect 7606 854 19583 856
rect 0 824 480 854
rect 2773 851 2839 854
rect 19517 851 19583 854
rect 3233 778 3299 781
rect 7925 778 7991 781
rect 3233 776 7991 778
rect 3233 720 3238 776
rect 3294 720 7930 776
rect 7986 720 7991 776
rect 3233 718 7991 720
rect 3233 715 3299 718
rect 7925 715 7991 718
rect 0 370 480 400
rect 6269 370 6335 373
rect 0 368 6335 370
rect 0 312 6274 368
rect 6330 312 6335 368
rect 0 310 6335 312
rect 0 280 480 310
rect 6269 307 6335 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 9996 15464 10060 15468
rect 9996 15408 10046 15464
rect 10046 15408 10060 15464
rect 9996 15404 10060 15408
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 3372 13772 3436 13836
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 11100 11868 11164 11932
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 3372 10432 3436 10436
rect 3372 10376 3422 10432
rect 3422 10376 3436 10432
rect 3372 10372 3436 10376
rect 11100 10372 11164 10436
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 9996 9692 10060 9756
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 9628 9556 9692 9620
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 15516 7848 15580 7852
rect 15516 7792 15530 7848
rect 15530 7792 15580 7848
rect 15516 7788 15580 7792
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 3740 6700 3804 6764
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 9996 5400 10060 5404
rect 9996 5344 10010 5400
rect 10010 5344 10060 5400
rect 9996 5340 10060 5344
rect 9628 4932 9692 4996
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 21588 3088 21652 3092
rect 21588 3032 21638 3088
rect 21638 3032 21652 3088
rect 21588 3028 21652 3032
rect 9996 2816 10060 2820
rect 9996 2760 10010 2816
rect 10010 2760 10060 2816
rect 9996 2756 10060 2760
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 9995 15468 10061 15469
rect 9995 15404 9996 15468
rect 10060 15404 10061 15468
rect 9995 15403 10061 15404
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 3371 13836 3437 13837
rect 3371 13772 3372 13836
rect 3436 13772 3437 13836
rect 3371 13771 3437 13772
rect 3374 10437 3434 13771
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 3371 10436 3437 10437
rect 3371 10372 3372 10436
rect 3436 10372 3437 10436
rect 3371 10371 3437 10372
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 9998 9757 10058 15403
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 11099 11932 11165 11933
rect 11099 11868 11100 11932
rect 11164 11868 11165 11932
rect 11099 11867 11165 11868
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 11102 10437 11162 11867
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 11099 10436 11165 10437
rect 11099 10372 11100 10436
rect 11164 10372 11165 10436
rect 11099 10371 11165 10372
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 9995 9756 10061 9757
rect 9995 9692 9996 9756
rect 10060 9692 10061 9756
rect 9995 9691 10061 9692
rect 9627 9620 9693 9621
rect 9627 9556 9628 9620
rect 9692 9556 9693 9620
rect 9627 9555 9693 9556
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 3742 6765 3802 7702
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 3739 6764 3805 6765
rect 3739 6700 3740 6764
rect 3804 6700 3805 6764
rect 3739 6699 3805 6700
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 9630 4997 9690 9555
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 9995 5404 10061 5405
rect 9995 5340 9996 5404
rect 10060 5340 10061 5404
rect 9995 5339 10061 5340
rect 9627 4996 9693 4997
rect 9627 4932 9628 4996
rect 9692 4932 9693 4996
rect 9627 4931 9693 4932
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 9630 3178 9690 4931
rect 9998 2821 10058 5339
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 9995 2820 10061 2821
rect 9995 2756 9996 2820
rect 10060 2756 10061 2820
rect 9995 2755 10061 2756
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 3654 7702 3890 7938
rect 9542 2942 9778 3178
rect 15430 7852 15666 7938
rect 15430 7788 15516 7852
rect 15516 7788 15580 7852
rect 15580 7788 15666 7852
rect 15430 7702 15666 7788
rect 21502 3092 21738 3178
rect 21502 3028 21588 3092
rect 21588 3028 21652 3092
rect 21652 3028 21738 3092
rect 21502 2942 21738 3028
<< metal5 >>
rect 3612 7938 15708 7980
rect 3612 7702 3654 7938
rect 3890 7702 15430 7938
rect 15666 7702 15708 7938
rect 3612 7660 15708 7702
rect 9500 3178 21780 3220
rect 9500 2942 9542 3178
rect 9778 2942 21502 3178
rect 21738 2942 21780 3178
rect 9500 2900 21780 2942
use scs8hd_fill_2  FILLER_1_9 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_6
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_conb_1  _041_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l1_in_2_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_2_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_38 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_34
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_30
timestamp 1586364061
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4876 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 5980 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_51
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_50
timestamp 1586364061
transform 1 0 5704 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_54
timestamp 1586364061
transform 1 0 6072 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6348 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_55
timestamp 1586364061
transform 1 0 6164 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_59
timestamp 1586364061
transform 1 0 6532 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_68
timestamp 1586364061
transform 1 0 7360 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l1_in_4_
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use scs8hd_buf_1  mux_bottom_track_1.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7084 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_77
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_71
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l1_in_5_
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_102
timestamp 1586364061
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_106
timestamp 1586364061
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_107
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _092_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _078_
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_decap_3  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 12604 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_1_148
timestamp 1586364061
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_144
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _074_
timestamp 1586364061
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15088 0 1 2720
box -38 -48 1786 592
use scs8hd_buf_2  _087_
timestamp 1586364061
transform 1 0 17112 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_165
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_0_171
timestamp 1586364061
transform 1 0 16836 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_decap_3  FILLER_1_198
timestamp 1586364061
transform 1 0 19320 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _076_
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 20424 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_210
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 20608 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_212
timestamp 1586364061
transform 1 0 20608 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 20976 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 20792 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_216
timestamp 1586364061
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_214
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_218
timestamp 1586364061
transform 1 0 21160 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_227
timestamp 1586364061
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_222
timestamp 1586364061
transform 1 0 21528 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_222 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21528 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 21344 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _080_
timestamp 1586364061
transform 1 0 21620 0 1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_235 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 22724 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_231
timestamp 1586364061
transform 1 0 22356 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_233
timestamp 1586364061
transform 1 0 22540 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_228
timestamp 1586364061
transform 1 0 22080 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 22540 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 22724 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _079_
timestamp 1586364061
transform 1 0 22172 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_0_237
timestamp 1586364061
transform 1 0 22908 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_1_243
timestamp 1586364061
transform 1 0 23460 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_245
timestamp 1586364061
transform 1 0 23644 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_buf_2  _089_
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_249
timestamp 1586364061
transform 1 0 24012 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_253
timestamp 1586364061
transform 1 0 24380 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _086_
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_253 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_257
timestamp 1586364061
transform 1 0 24748 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_0_269
timestamp 1586364061
transform 1 0 25852 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_265
timestamp 1586364061
transform 1 0 25484 0 1 2720
box -38 -48 1142 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 2760 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_16
timestamp 1586364061
transform 1 0 2576 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_24
timestamp 1586364061
transform 1 0 3312 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_20
timestamp 1586364061
transform 1 0 2944 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 3128 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_28
timestamp 1586364061
transform 1 0 3680 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3496 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_39
timestamp 1586364061
transform 1 0 4692 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_36
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 4508 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5520 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 5336 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_43
timestamp 1586364061
transform 1 0 5060 0 -1 3808
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_67
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_71
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10120 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 9292 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9844 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_91
timestamp 1586364061
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_97
timestamp 1586364061
transform 1 0 10028 0 -1 3808
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 11684 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_107
timestamp 1586364061
transform 1 0 10948 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_112
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_134
timestamp 1586364061
transform 1 0 13432 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_138
timestamp 1586364061
transform 1 0 13800 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _093_
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_1  mux_bottom_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_158
timestamp 1586364061
transform 1 0 15640 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 15824 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_162
timestamp 1586364061
transform 1 0 16008 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1586364061
transform 1 0 19136 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18952 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_188
timestamp 1586364061
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_192
timestamp 1586364061
transform 1 0 18768 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _081_
timestamp 1586364061
transform 1 0 21068 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 20148 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 20516 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_205
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_209
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_213
timestamp 1586364061
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _083_
timestamp 1586364061
transform 1 0 22172 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_221
timestamp 1586364061
transform 1 0 21436 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_2_233
timestamp 1586364061
transform 1 0 22540 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_245
timestamp 1586364061
transform 1 0 23644 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_257
timestamp 1586364061
transform 1 0 24748 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_2_269
timestamp 1586364061
transform 1 0 25852 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2300 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 2116 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_9
timestamp 1586364061
transform 1 0 1932 0 1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 3864 0 1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3680 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3312 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_22
timestamp 1586364061
transform 1 0 3128 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_26
timestamp 1586364061
transform 1 0 3496 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_49
timestamp 1586364061
transform 1 0 5612 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1586364061
transform 1 0 7728 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7084 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7452 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_67
timestamp 1586364061
transform 1 0 7268 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_71
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 8740 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_81
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_85
timestamp 1586364061
transform 1 0 8924 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 406 592
use scs8hd_conb_1  _046_
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 11684 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_102
timestamp 1586364061
transform 1 0 10488 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_105
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_109
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_113
timestamp 1586364061
transform 1 0 11500 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_117
timestamp 1586364061
transform 1 0 11868 0 1 3808
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_136
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_149
timestamp 1586364061
transform 1 0 14812 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_153
timestamp 1586364061
transform 1 0 15180 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1586364061
transform 1 0 16100 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15916 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_160
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_172
timestamp 1586364061
transform 1 0 16928 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_176
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_197
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _082_
timestamp 1586364061
transform 1 0 21160 0 1 3808
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 20976 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_210
timestamp 1586364061
transform 1 0 20424 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_214
timestamp 1586364061
transform 1 0 20792 0 1 3808
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22264 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 22080 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22724 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_222
timestamp 1586364061
transform 1 0 21528 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_226
timestamp 1586364061
transform 1 0 21896 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_233
timestamp 1586364061
transform 1 0 22540 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_237
timestamp 1586364061
transform 1 0 22908 0 1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_243
timestamp 1586364061
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_11
timestamp 1586364061
transform 1 0 2116 0 -1 4896
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 4600 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_29
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_36
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5520 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_40
timestamp 1586364061
transform 1 0 4784 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_46
timestamp 1586364061
transform 1 0 5336 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_57
timestamp 1586364061
transform 1 0 6348 0 -1 4896
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7084 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 8096 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_61
timestamp 1586364061
transform 1 0 6716 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_64
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_74
timestamp 1586364061
transform 1 0 7912 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_78
timestamp 1586364061
transform 1 0 8280 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_82
timestamp 1586364061
transform 1 0 8648 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_86
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9292 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_91
timestamp 1586364061
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_buf_1  mux_bottom_track_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 9936 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_99
timestamp 1586364061
transform 1 0 10212 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l1_in_6_
timestamp 1586364061
transform 1 0 10948 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 10396 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_103
timestamp 1586364061
transform 1 0 10580 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_116
timestamp 1586364061
transform 1 0 11776 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1586364061
transform 1 0 12512 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 13524 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12328 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_120
timestamp 1586364061
transform 1 0 12144 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_133
timestamp 1586364061
transform 1 0 13340 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_137
timestamp 1586364061
transform 1 0 13708 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_2  _075_
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use scs8hd_buf_2  _091_
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 13892 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_158
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16468 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_162
timestamp 1586364061
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_165
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_176
timestamp 1586364061
transform 1 0 17296 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_180
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_193
timestamp 1586364061
transform 1 0 18860 0 -1 4896
box -38 -48 406 592
use scs8hd_buf_2  _084_
timestamp 1586364061
transform 1 0 19596 0 -1 4896
box -38 -48 406 592
use scs8hd_buf_2  _085_
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 20148 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20516 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_199
timestamp 1586364061
transform 1 0 19412 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_205
timestamp 1586364061
transform 1 0 19964 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_209
timestamp 1586364061
transform 1 0 20332 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_213
timestamp 1586364061
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 21436 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21804 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_219
timestamp 1586364061
transform 1 0 21252 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_223
timestamp 1586364061
transform 1 0 21620 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_12
timestamp 1586364061
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_16
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_20
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_24
timestamp 1586364061
transform 1 0 3312 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_36
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_40
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9292 0 1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_81
timestamp 1586364061
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_85
timestamp 1586364061
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_108
timestamp 1586364061
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_112
timestamp 1586364061
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_116
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1786 592
use scs8hd_buf_1  mux_bottom_track_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12512 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_131
timestamp 1586364061
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_154
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_160
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_175
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_197
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 866 592
use scs8hd_buf_1  mux_bottom_track_17.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 21160 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_210
timestamp 1586364061
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_214
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21620 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21988 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 22724 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_221
timestamp 1586364061
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_225
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_229
timestamp 1586364061
transform 1 0 22172 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_233
timestamp 1586364061
transform 1 0 22540 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_237
timestamp 1586364061
transform 1 0 22908 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 23276 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_243
timestamp 1586364061
transform 1 0 23460 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 1786 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_29
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_26
timestamp 1586364061
transform 1 0 3496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_22
timestamp 1586364061
transform 1 0 3128 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_35
timestamp 1586364061
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_31
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 4508 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_55
timestamp 1586364061
transform 1 0 6164 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_51
timestamp 1586364061
transform 1 0 5796 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6348 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 5980 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1586364061
transform 1 0 6532 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 7544 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_72
timestamp 1586364061
transform 1 0 7728 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 7912 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_76
timestamp 1586364061
transform 1 0 8096 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 8280 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_79
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _043_
timestamp 1586364061
transform 1 0 8556 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_83
timestamp 1586364061
transform 1 0 8740 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_87
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11960 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_112
timestamp 1586364061
transform 1 0 11408 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_116
timestamp 1586364061
transform 1 0 11776 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12144 0 -1 5984
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_136
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_140
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_139
timestamp 1586364061
transform 1 0 13892 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14260 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14076 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 15456 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_buf_2  _090_
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 1786 592
use scs8hd_decap_3  FILLER_7_168
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_162
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_168
timestamp 1586364061
transform 1 0 16560 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_162
timestamp 1586364061
transform 1 0 16008 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _088_
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 16744 0 -1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 18860 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_189
timestamp 1586364061
transform 1 0 18492 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_195
timestamp 1586364061
transform 1 0 19044 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_207
timestamp 1586364061
transform 1 0 20148 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_203
timestamp 1586364061
transform 1 0 19780 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 19964 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_213
timestamp 1586364061
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_210
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 20332 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1586364061
transform 1 0 20516 0 1 5984
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use scs8hd_buf_1  mux_bottom_track_33.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22264 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 21528 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22724 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_224
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_6_236
timestamp 1586364061
transform 1 0 22816 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_224
timestamp 1586364061
transform 1 0 21712 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_233
timestamp 1586364061
transform 1 0 22540 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_237
timestamp 1586364061
transform 1 0 22908 0 1 5984
box -38 -48 590 592
use scs8hd_buf_2  _077_
timestamp 1586364061
transform 1 0 23276 0 -1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_240
timestamp 1586364061
transform 1 0 23184 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_245
timestamp 1586364061
transform 1 0 23644 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_257
timestamp 1586364061
transform 1 0 24748 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_243
timestamp 1586364061
transform 1 0 23460 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_269
timestamp 1586364061
transform 1 0 25852 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_conb_1  _044_
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5980 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_46
timestamp 1586364061
transform 1 0 5336 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_50
timestamp 1586364061
transform 1 0 5704 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 7912 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8280 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_72
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_76
timestamp 1586364061
transform 1 0 8096 0 -1 7072
box -38 -48 222 592
use scs8hd_conb_1  _045_
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 8924 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_83
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_87
timestamp 1586364061
transform 1 0 9108 0 -1 7072
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_107
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_8_119
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_125
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_136
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_140
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_148
timestamp 1586364061
transform 1 0 14720 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_144
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14536 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_158
timestamp 1586364061
transform 1 0 15640 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 130 592
use scs8hd_conb_1  _047_
timestamp 1586364061
transform 1 0 15364 0 -1 7072
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_162
timestamp 1586364061
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_165
timestamp 1586364061
transform 1 0 16284 0 -1 7072
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 18308 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_185
timestamp 1586364061
transform 1 0 18124 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_189
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 20516 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 19872 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_206
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_210
timestamp 1586364061
transform 1 0 20424 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_12
timestamp 1586364061
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_16
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_29
timestamp 1586364061
transform 1 0 3772 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_33
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_37
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_41
timestamp 1586364061
transform 1 0 4876 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_78
timestamp 1586364061
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1586364061
transform 1 0 8648 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 8464 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_91
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_95
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_99
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _042_
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_126
timestamp 1586364061
transform 1 0 12696 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_132
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1586364061
transform 1 0 15640 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_145
timestamp 1586364061
transform 1 0 14444 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_149
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_154
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_167
timestamp 1586364061
transform 1 0 16468 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_177
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_181
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_197
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_210
timestamp 1586364061
transform 1 0 20424 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_222
timestamp 1586364061
transform 1 0 21528 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_234
timestamp 1586364061
transform 1 0 22632 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_242
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 2668 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_12
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_16
timestamp 1586364061
transform 1 0 2576 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_19
timestamp 1586364061
transform 1 0 2852 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3036 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6072 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 5796 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_45
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_49
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_53
timestamp 1586364061
transform 1 0 5980 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_73
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_77
timestamp 1586364061
transform 1 0 8188 0 -1 8160
box -38 -48 222 592
use scs8hd_conb_1  _036_
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1586364061
transform 1 0 11684 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11500 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_107
timestamp 1586364061
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_111
timestamp 1586364061
transform 1 0 11316 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_124
timestamp 1586364061
transform 1 0 12512 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_128
timestamp 1586364061
transform 1 0 12880 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_131
timestamp 1586364061
transform 1 0 13156 0 -1 8160
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 15640 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14260 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1586364061
transform 1 0 16008 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 17388 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17020 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_160
timestamp 1586364061
transform 1 0 15824 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_171
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_175
timestamp 1586364061
transform 1 0 17204 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1586364061
transform 1 0 17572 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 18952 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_188
timestamp 1586364061
transform 1 0 18400 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_192
timestamp 1586364061
transform 1 0 18768 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_196
timestamp 1586364061
transform 1 0 19136 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 19596 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_200
timestamp 1586364061
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_203
timestamp 1586364061
transform 1 0 19780 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_211
timestamp 1586364061
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_conb_1  _037_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 1840 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_6
timestamp 1586364061
transform 1 0 1656 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_10
timestamp 1586364061
transform 1 0 2024 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_14
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_26
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_30
timestamp 1586364061
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_75
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_78
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 8648 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use scs8hd_conb_1  _035_
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_101
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_105
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12972 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12788 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 15180 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_148
timestamp 1586364061
transform 1 0 14720 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_152
timestamp 1586364061
transform 1 0 15088 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_155
timestamp 1586364061
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1586364061
transform 1 0 16100 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_172
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_176
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l1_in_3_
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_180
timestamp 1586364061
transform 1 0 17664 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_197
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_209
timestamp 1586364061
transform 1 0 20332 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_221
timestamp 1586364061
transform 1 0 21436 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_233
timestamp 1586364061
transform 1 0 22540 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_11_241
timestamp 1586364061
transform 1 0 23276 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 1472 0 -1 9248
box -38 -48 1786 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 130 592
use scs8hd_conb_1  _038_
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4508 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_35
timestamp 1586364061
transform 1 0 4324 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_39
timestamp 1586364061
transform 1 0 4692 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 5428 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_43
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 7544 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_60
timestamp 1586364061
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_64
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_72
timestamp 1586364061
transform 1 0 7728 0 -1 9248
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11776 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 11592 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11132 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_107
timestamp 1586364061
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_111
timestamp 1586364061
transform 1 0 11316 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_135
timestamp 1586364061
transform 1 0 13524 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_140
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_144
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 14536 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_148
timestamp 1586364061
transform 1 0 14720 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 14904 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_152
timestamp 1586364061
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 15456 0 -1 9248
box -38 -48 222 592
use scs8hd_conb_1  _040_
timestamp 1586364061
transform 1 0 15640 0 -1 9248
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16652 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 16468 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_161
timestamp 1586364061
transform 1 0 15916 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_165
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 18952 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 19320 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_188
timestamp 1586364061
transform 1 0 18400 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_192
timestamp 1586364061
transform 1 0 18768 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_196
timestamp 1586364061
transform 1 0 19136 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_200
timestamp 1586364061
transform 1 0 19504 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_12_212
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_24.mux_l1_in_3_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 866 592
use scs8hd_mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 866 592
use scs8hd_decap_4  FILLER_14_16
timestamp 1586364061
transform 1 0 2576 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_12
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_16
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_12
timestamp 1586364061
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_20
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_20
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 3036 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_36
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 4600 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 3036 0 1 9248
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_14_40
timestamp 1586364061
transform 1 0 4784 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_44
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_40
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 866 592
use scs8hd_conb_1  _034_
timestamp 1586364061
transform 1 0 5520 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_54
timestamp 1586364061
transform 1 0 6072 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_50
timestamp 1586364061
transform 1 0 5704 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6440 0 -1 10336
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1786 592
use scs8hd_mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_67
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_71
timestamp 1586364061
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_85
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_81
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_91
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_13_101
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_16.mux_l1_in_3_
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_116
timestamp 1586364061
transform 1 0 11776 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_112
timestamp 1586364061
transform 1 0 11408 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 11592 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_120
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 12788 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_136
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_134
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_129
timestamp 1586364061
transform 1 0 12972 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_14_140
timestamp 1586364061
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14168 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_148
timestamp 1586364061
transform 1 0 14720 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_144
timestamp 1586364061
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14536 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_158
timestamp 1586364061
transform 1 0 15640 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_157
timestamp 1586364061
transform 1 0 15548 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 15456 0 -1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 16008 0 -1 10336
box -38 -48 1786 592
use scs8hd_mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1586364061
transform 1 0 16284 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 15824 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_161
timestamp 1586364061
transform 1 0 15916 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_164
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_174
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_186
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_181
timestamp 1586364061
transform 1 0 17756 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1586364061
transform 1 0 18492 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_12  FILLER_14_198
timestamp 1586364061
transform 1 0 19320 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 19780 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_201
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_205
timestamp 1586364061
transform 1 0 19964 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_210
timestamp 1586364061
transform 1 0 20424 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_229
timestamp 1586364061
transform 1 0 22172 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_241
timestamp 1586364061
transform 1 0 23276 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2668 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_12
timestamp 1586364061
transform 1 0 2208 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_16
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_19
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1586364061
transform 1 0 3220 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_32
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_36
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_40
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7728 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7544 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_68
timestamp 1586364061
transform 1 0 7360 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_91
timestamp 1586364061
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_95
timestamp 1586364061
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_108
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_112
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_116
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_136
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 14536 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 14904 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_140
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_144
timestamp 1586364061
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_148
timestamp 1586364061
transform 1 0 14720 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_152
timestamp 1586364061
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_4.mux_l1_in_6_
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_205
timestamp 1586364061
transform 1 0 19964 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_217
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_229
timestamp 1586364061
transform 1 0 22172 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_241
timestamp 1586364061
transform 1 0 23276 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_buf_1  mux_left_track_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_10
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_1  mux_left_track_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 4140 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 4600 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_36
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_40
timestamp 1586364061
transform 1 0 4784 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_46
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7912 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_66
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_70
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 8924 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_83
timestamp 1586364061
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_87
timestamp 1586364061
transform 1 0 9108 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_97
timestamp 1586364061
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10396 0 -1 11424
box -38 -48 1786 592
use scs8hd_mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_120
timestamp 1586364061
transform 1 0 12144 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_137
timestamp 1586364061
transform 1 0 13708 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14260 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 13892 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_149
timestamp 1586364061
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15640 0 -1 11424
box -38 -48 866 592
use scs8hd_mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 17204 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 17020 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 16652 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_167
timestamp 1586364061
transform 1 0 16468 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_171
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_184
timestamp 1586364061
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_188
timestamp 1586364061
transform 1 0 18400 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_200
timestamp 1586364061
transform 1 0 19504 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_16_212
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_buf_2  _072_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 2852 0 1 11424
box -38 -48 1786 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 2668 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_11
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_38
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 5336 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_42
timestamp 1586364061
transform 1 0 4968 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_48
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_52
timestamp 1586364061
transform 1 0 5888 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_81
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_85
timestamp 1586364061
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_89
timestamp 1586364061
transform 1 0 9292 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_95
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_99
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12512 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1586364061
transform 1 0 14996 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_143
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_160
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_164
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_168
timestamp 1586364061
transform 1 0 16560 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_174
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_178
timestamp 1586364061
transform 1 0 17480 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 17664 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_182
timestamp 1586364061
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1786 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_buf_2  _073_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3312 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3680 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_22
timestamp 1586364061
transform 1 0 3128 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_26
timestamp 1586364061
transform 1 0 3496 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_30
timestamp 1586364061
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_36
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 4968 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_40
timestamp 1586364061
transform 1 0 4784 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7820 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 7636 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 7268 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_65
timestamp 1586364061
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_69
timestamp 1586364061
transform 1 0 7452 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_82
timestamp 1586364061
transform 1 0 8648 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_86
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_89
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_106
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_119
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12512 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 13800 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_123
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_126
timestamp 1586364061
transform 1 0 12696 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_136
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15364 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_140
timestamp 1586364061
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_144
timestamp 1586364061
transform 1 0 14352 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_4.mux_l1_in_5_
timestamp 1586364061
transform 1 0 16928 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 16744 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_164
timestamp 1586364061
transform 1 0 16192 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_168
timestamp 1586364061
transform 1 0 16560 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18032 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_181
timestamp 1586364061
transform 1 0 17756 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_186
timestamp 1586364061
transform 1 0 18216 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_198
timestamp 1586364061
transform 1 0 19320 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_210
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_6
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 1840 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_buf_1  mux_left_track_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_10
timestamp 1586364061
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 2024 0 1 12512
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_29
timestamp 1586364061
transform 1 0 3772 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_33
timestamp 1586364061
transform 1 0 4140 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 4232 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1586364061
transform 1 0 4416 0 -1 13600
box -38 -48 866 592
use scs8hd_mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4508 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_49
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_45
timestamp 1586364061
transform 1 0 5244 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_46
timestamp 1586364061
transform 1 0 5336 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 5428 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_55
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 406 592
use scs8hd_decap_3  FILLER_19_50
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_62
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_20_72
timestamp 1586364061
transform 1 0 7728 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_77
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7544 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9108 0 1 12512
box -38 -48 1786 592
use scs8hd_mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_81
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 406 592
use scs8hd_decap_3  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_89
timestamp 1586364061
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_106
timestamp 1586364061
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11040 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_114
timestamp 1586364061
transform 1 0 11592 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_110
timestamp 1586364061
transform 1 0 11224 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 11408 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 11776 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 12788 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1586364061
transform 1 0 12512 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_137
timestamp 1586364061
transform 1 0 13708 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_133
timestamp 1586364061
transform 1 0 13340 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 13156 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 13340 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_146
timestamp 1586364061
transform 1 0 14536 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_142
timestamp 1586364061
transform 1 0 14168 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_148
timestamp 1586364061
transform 1 0 14720 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_144
timestamp 1586364061
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 13892 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 14536 0 1 12512
box -38 -48 222 592
use scs8hd_conb_1  _039_
timestamp 1586364061
transform 1 0 14076 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_150
timestamp 1586364061
transform 1 0 14904 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_152
timestamp 1586364061
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 1786 592
use scs8hd_mux2_1  mux_top_track_4.mux_l1_in_4_
timestamp 1586364061
transform 1 0 16836 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 16652 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_163
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_167
timestamp 1586364061
transform 1 0 16468 0 -1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_192
timestamp 1586364061
transform 1 0 18768 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_203
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_215
timestamp 1586364061
transform 1 0 20884 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_204
timestamp 1586364061
transform 1 0 19872 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_212
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_227
timestamp 1586364061
transform 1 0 21988 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_239
timestamp 1586364061
transform 1 0 23092 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_243
timestamp 1586364061
transform 1 0 23460 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_263
timestamp 1586364061
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1586364061
transform 1 0 1564 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_14
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_18
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 3128 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4140 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4508 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_31
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_35
timestamp 1586364061
transform 1 0 4324 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7176 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6992 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_75
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_79
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 9752 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_92
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_96
timestamp 1586364061
transform 1 0 9936 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_11.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10304 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 11316 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_109
timestamp 1586364061
transform 1 0 11132 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_113
timestamp 1586364061
transform 1 0 11500 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12696 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 13064 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_128
timestamp 1586364061
transform 1 0 12880 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14812 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 14260 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_141
timestamp 1586364061
transform 1 0 14076 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_145
timestamp 1586364061
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_168
timestamp 1586364061
transform 1 0 16560 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_172
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_21_180
timestamp 1586364061
transform 1 0 17664 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_buf_1  mux_left_track_7.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_6
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_10
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6532 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5980 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6348 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_51
timestamp 1586364061
transform 1 0 5796 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_55
timestamp 1586364061
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_78
timestamp 1586364061
transform 1 0 8280 0 -1 14688
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_11.mux_l3_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_82
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_85
timestamp 1586364061
transform 1 0 8924 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_89
timestamp 1586364061
transform 1 0 9292 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11776 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_102
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_106
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_114
timestamp 1586364061
transform 1 0 11592 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_118
timestamp 1586364061
transform 1 0 11960 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12696 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 12512 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 12144 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_122
timestamp 1586364061
transform 1 0 12328 0 -1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_151
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_175
timestamp 1586364061
transform 1 0 17204 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_187
timestamp 1586364061
transform 1 0 18308 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_199
timestamp 1586364061
transform 1 0 19412 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_22_211
timestamp 1586364061
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_263
timestamp 1586364061
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_buf_1  mux_left_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2208 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_6
timestamp 1586364061
transform 1 0 1656 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_10
timestamp 1586364061
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use scs8hd_buf_2  _069_
timestamp 1586364061
transform 1 0 3956 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_23
timestamp 1586364061
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_35
timestamp 1586364061
transform 1 0 4324 0 1 14688
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_40
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_71
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_75
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_79
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_11.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_102
timestamp 1586364061
transform 1 0 10488 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_107
timestamp 1586364061
transform 1 0 10948 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_111
timestamp 1586364061
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_115
timestamp 1586364061
transform 1 0 11684 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_119
timestamp 1586364061
transform 1 0 12052 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_127
timestamp 1586364061
transform 1 0 12788 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12604 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12972 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_131
timestamp 1586364061
transform 1 0 13156 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 13708 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 13892 0 1 14688
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_23_158
timestamp 1586364061
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16560 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_162
timestamp 1586364061
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_166
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_170
timestamp 1586364061
transform 1 0 16744 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_23_182
timestamp 1586364061
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_232
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_buf_1  mux_left_track_13.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_6
timestamp 1586364061
transform 1 0 1656 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_10
timestamp 1586364061
transform 1 0 2024 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_1  mux_left_track_15.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 4508 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_35
timestamp 1586364061
transform 1 0 4324 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_39
timestamp 1586364061
transform 1 0 4692 0 -1 15776
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 5796 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 5520 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_43
timestamp 1586364061
transform 1 0 5060 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_46
timestamp 1586364061
transform 1 0 5336 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_50
timestamp 1586364061
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 7728 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8096 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_70
timestamp 1586364061
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_74
timestamp 1586364061
transform 1 0 7912 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_78
timestamp 1586364061
transform 1 0 8280 0 -1 15776
box -38 -48 314 592
use scs8hd_conb_1  _049_
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9936 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_98
timestamp 1586364061
transform 1 0 10120 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_13.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 10304 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_114
timestamp 1586364061
transform 1 0 11592 0 -1 15776
box -38 -48 774 592
use scs8hd_mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12328 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 13708 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_131
timestamp 1586364061
transform 1 0 13156 0 -1 15776
box -38 -48 590 592
use scs8hd_mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use scs8hd_buf_1  mux_top_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 14168 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_139
timestamp 1586364061
transform 1 0 13892 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_149
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_175
timestamp 1586364061
transform 1 0 17204 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_187
timestamp 1586364061
transform 1 0 18308 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_199
timestamp 1586364061
transform 1 0 19412 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_24_211
timestamp 1586364061
transform 1 0 20516 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_buf_2  _071_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_7.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 1786 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 2208 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_11
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_14
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_37
timestamp 1586364061
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _033_
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_41
timestamp 1586364061
transform 1 0 4876 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_46
timestamp 1586364061
transform 1 0 5336 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_11.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 7176 0 1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6992 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_11.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 9292 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_85
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_91
timestamp 1586364061
transform 1 0 9476 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_13.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 13708 0 1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_156
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_160
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_164
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_168
timestamp 1586364061
transform 1 0 16560 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_25_180
timestamp 1586364061
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_220
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_2  _070_
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use scs8hd_buf_2  _068_
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_7
timestamp 1586364061
transform 1 0 1748 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 1932 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_12
timestamp 1586364061
transform 1 0 2208 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_11
timestamp 1586364061
transform 1 0 2116 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 2300 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 2024 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_16
timestamp 1586364061
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_19
timestamp 1586364061
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use scs8hd_buf_2  _067_
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_7.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 2944 0 1 16864
box -38 -48 1786 592
use scs8hd_mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_43
timestamp 1586364061
transform 1 0 5060 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_45
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 5428 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 5244 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 4876 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1586364061
transform 1 0 5612 0 -1 16864
box -38 -48 866 592
use scs8hd_buf_1  mux_left_track_11.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 5428 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_54
timestamp 1586364061
transform 1 0 6072 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_50
timestamp 1586364061
transform 1 0 5704 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_58
timestamp 1586364061
transform 1 0 6440 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_62
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6624 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 866 592
use scs8hd_mux2_1  mux_left_track_15.mux_l3_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_75
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_71
timestamp 1586364061
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_79
timestamp 1586364061
transform 1 0 8372 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_75
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 8188 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  mux_left_track_19.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_82
timestamp 1586364061
transform 1 0 8648 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_89
timestamp 1586364061
transform 1 0 9292 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_26_83
timestamp 1586364061
transform 1 0 8740 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 8556 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8832 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_99
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9384 0 1 16864
box -38 -48 866 592
use scs8hd_mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9936 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_6  FILLER_27_103
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 590 592
use scs8hd_decap_8  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11132 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_113
timestamp 1586364061
transform 1 0 11500 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_conb_1  _050_
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_13.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 11684 0 -1 16864
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_left_track_13.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13064 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_23.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12696 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_134
timestamp 1586364061
transform 1 0 13432 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_128
timestamp 1586364061
transform 1 0 12880 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_26_146
timestamp 1586364061
transform 1 0 14536 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_26_152
timestamp 1586364061
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_151
timestamp 1586364061
transform 1 0 14996 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_175
timestamp 1586364061
transform 1 0 17204 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_163
timestamp 1586364061
transform 1 0 16100 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_175
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_187
timestamp 1586364061
transform 1 0 18308 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_199
timestamp 1586364061
transform 1 0 19412 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_26_211
timestamp 1586364061
transform 1 0 20516 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_conb_1  _032_
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 1840 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_6
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_10
timestamp 1586364061
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_7.mux_l1_in_3_
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use scs8hd_conb_1  _051_
timestamp 1586364061
transform 1 0 5612 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6440 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6072 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 5060 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 5428 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_41
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_45
timestamp 1586364061
transform 1 0 5244 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_52
timestamp 1586364061
transform 1 0 5888 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_15.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6624 0 -1 17952
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_28_79
timestamp 1586364061
transform 1 0 8372 0 -1 17952
box -38 -48 774 592
use scs8hd_buf_1  mux_left_track_21.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 10120 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9844 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_87
timestamp 1586364061
transform 1 0 9108 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_97
timestamp 1586364061
transform 1 0 10028 0 -1 17952
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_15.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 11132 0 -1 17952
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_28_101
timestamp 1586364061
transform 1 0 10396 0 -1 17952
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 13248 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_128
timestamp 1586364061
transform 1 0 12880 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_6  FILLER_28_134
timestamp 1586364061
transform 1 0 13432 0 -1 17952
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13984 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_142
timestamp 1586364061
transform 1 0 14168 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_146
timestamp 1586364061
transform 1 0 14536 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_152
timestamp 1586364061
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_buf_2  _066_
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_7.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2668 0 1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_13
timestamp 1586364061
transform 1 0 2300 0 1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_7.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3680 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_26
timestamp 1586364061
transform 1 0 3496 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_30
timestamp 1586364061
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6992 0 1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_15.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9476 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9292 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_83
timestamp 1586364061
transform 1 0 8740 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_87
timestamp 1586364061
transform 1 0 9108 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_13.mux_l2_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_23.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 866 592
use scs8hd_decap_12  FILLER_29_149
timestamp 1586364061
transform 1 0 14812 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_161
timestamp 1586364061
transform 1 0 15916 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_173
timestamp 1586364061
transform 1 0 17020 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_181
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_buf_2  _063_
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 406 592
use scs8hd_buf_2  _065_
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 1932 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 2300 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_11
timestamp 1586364061
transform 1 0 2116 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_19
timestamp 1586364061
transform 1 0 2852 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 3036 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_36
timestamp 1586364061
transform 1 0 4416 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4232 0 -1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4508 0 -1 19040
box -38 -48 866 592
use scs8hd_mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 6072 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 5520 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_46
timestamp 1586364061
transform 1 0 5336 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_50
timestamp 1586364061
transform 1 0 5704 0 -1 19040
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_15.mux_l2_in_1_
timestamp 1586364061
transform 1 0 7636 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 7084 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_63
timestamp 1586364061
transform 1 0 6900 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_67
timestamp 1586364061
transform 1 0 7268 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_2  FILLER_30_88
timestamp 1586364061
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use scs8hd_conb_1  _027_
timestamp 1586364061
transform 1 0 11224 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_21.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11040 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 11684 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12052 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_106
timestamp 1586364061
transform 1 0 10856 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_113
timestamp 1586364061
transform 1 0 11500 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_23.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12696 0 -1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_121
timestamp 1586364061
transform 1 0 12236 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_125
timestamp 1586364061
transform 1 0 12604 0 -1 19040
box -38 -48 130 592
use scs8hd_conb_1  _028_
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_12  FILLER_30_157
timestamp 1586364061
transform 1 0 15548 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_169
timestamp 1586364061
transform 1 0 16652 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_181
timestamp 1586364061
transform 1 0 17756 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_193
timestamp 1586364061
transform 1 0 18860 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_205
timestamp 1586364061
transform 1 0 19964 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_213
timestamp 1586364061
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_buf_2  _060_
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 406 592
use scs8hd_buf_2  _064_
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 2300 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_11
timestamp 1586364061
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_19
timestamp 1586364061
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 3036 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_23
timestamp 1586364061
transform 1 0 3220 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_38
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_42
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 222 592
use scs8hd_conb_1  _031_
timestamp 1586364061
transform 1 0 5336 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_49
timestamp 1586364061
transform 1 0 5612 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7452 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6992 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_66
timestamp 1586364061
transform 1 0 7176 0 1 19040
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9200 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8648 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_80
timestamp 1586364061
transform 1 0 8464 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_84
timestamp 1586364061
transform 1 0 8832 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_97
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_21.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10488 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_101
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_104
timestamp 1586364061
transform 1 0 10672 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12604 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_134
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_138
timestamp 1586364061
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_23.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14168 0 1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_23.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_161
timestamp 1586364061
transform 1 0 15916 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_173
timestamp 1586364061
transform 1 0 17020 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_181
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_buf_2  _062_
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use scs8hd_buf_1  mux_left_track_23.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1932 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 2300 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_7
timestamp 1586364061
transform 1 0 1748 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_11
timestamp 1586364061
transform 1 0 2116 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_18
timestamp 1586364061
transform 1 0 2760 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2944 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_22
timestamp 1586364061
transform 1 0 3128 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 6532 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 5980 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_51
timestamp 1586364061
transform 1 0 5796 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_55
timestamp 1586364061
transform 1 0 6164 0 -1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7636 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8004 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8372 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_73
timestamp 1586364061
transform 1 0 7820 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_77
timestamp 1586364061
transform 1 0 8188 0 -1 20128
box -38 -48 222 592
use scs8hd_conb_1  _053_
timestamp 1586364061
transform 1 0 8556 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_19.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9844 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_19.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10212 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_90
timestamp 1586364061
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_97
timestamp 1586364061
transform 1 0 10028 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_21.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10488 0 -1 20128
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_32_101
timestamp 1586364061
transform 1 0 10396 0 -1 20128
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_23.mux_l1_in_1_
timestamp 1586364061
transform 1 0 13524 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 13340 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_21.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_121
timestamp 1586364061
transform 1 0 12236 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_125
timestamp 1586364061
transform 1 0 12604 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_131
timestamp 1586364061
transform 1 0 13156 0 -1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_23.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14536 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_144
timestamp 1586364061
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_148
timestamp 1586364061
transform 1 0 14720 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_152
timestamp 1586364061
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_6
timestamp 1586364061
transform 1 0 1656 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 1840 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_buf_1  mux_left_track_17.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use scs8hd_buf_2  _061_
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_10
timestamp 1586364061
transform 1 0 2024 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_16
timestamp 1586364061
transform 1 0 2576 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_12
timestamp 1586364061
transform 1 0 2208 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 2024 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 2208 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2760 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2392 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_23
timestamp 1586364061
transform 1 0 3220 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_20
timestamp 1586364061
transform 1 0 2944 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3404 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3220 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4324 0 -1 21216
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 3404 0 1 20128
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_34_48
timestamp 1586364061
transform 1 0 5520 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_44
timestamp 1586364061
transform 1 0 5152 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 5520 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 5336 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_58
timestamp 1586364061
transform 1 0 6440 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_54
timestamp 1586364061
transform 1 0 6072 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_50
timestamp 1586364061
transform 1 0 5704 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 5704 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 6256 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 5888 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 5888 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_65
timestamp 1586364061
transform 1 0 7084 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_61
timestamp 1586364061
transform 1 0 6716 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6900 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 7268 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 7176 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7452 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_78
timestamp 1586364061
transform 1 0 8280 0 -1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7360 0 1 20128
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_34_87
timestamp 1586364061
transform 1 0 9108 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_3  FILLER_34_82
timestamp 1586364061
transform 1 0 8648 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_87
timestamp 1586364061
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_19.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9292 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 8924 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_91
timestamp 1586364061
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_91
timestamp 1586364061
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_19.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_19.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_left_track_19.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9844 0 1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 11592 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_114
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_112
timestamp 1586364061
transform 1 0 11408 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_116
timestamp 1586364061
transform 1 0 11776 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_127
timestamp 1586364061
transform 1 0 12788 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_123
timestamp 1586364061
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12604 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_21.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_buf_1  mux_left_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12144 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_131
timestamp 1586364061
transform 1 0 13156 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13340 0 -1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1586364061
transform 1 0 13524 0 -1 21216
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_21.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_34_144
timestamp 1586364061
transform 1 0 14352 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_146
timestamp 1586364061
transform 1 0 14536 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_142
timestamp 1586364061
transform 1 0 14168 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 14352 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_152
timestamp 1586364061
transform 1 0 15088 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_150
timestamp 1586364061
transform 1 0 14904 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 15456 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 15088 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_158
timestamp 1586364061
transform 1 0 15640 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_154
timestamp 1586364061
transform 1 0 15272 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_166
timestamp 1586364061
transform 1 0 16376 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_33_178
timestamp 1586364061
transform 1 0 17480 0 1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_170
timestamp 1586364061
transform 1 0 16744 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_182
timestamp 1586364061
transform 1 0 17848 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_182
timestamp 1586364061
transform 1 0 17848 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_194
timestamp 1586364061
transform 1 0 18952 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_206
timestamp 1586364061
transform 1 0 20056 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 2208 0 1 21216
box -38 -48 1786 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 2024 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 1564 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_7
timestamp 1586364061
transform 1 0 1748 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 4324 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_31
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_37
timestamp 1586364061
transform 1 0 4508 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1586364061
transform 1 0 4876 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_50
timestamp 1586364061
transform 1 0 5704 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_55
timestamp 1586364061
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6992 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8372 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_73
timestamp 1586364061
transform 1 0 7820 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_77
timestamp 1586364061
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_19.mux_l1_in_1_
timestamp 1586364061
transform 1 0 8924 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 8740 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_81
timestamp 1586364061
transform 1 0 8556 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_94
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_21.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10488 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_100
timestamp 1586364061
transform 1 0 10304 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_104
timestamp 1586364061
transform 1 0 10672 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_114
timestamp 1586364061
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_132
timestamp 1586364061
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_136
timestamp 1586364061
transform 1 0 13616 0 1 21216
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14168 0 1 21216
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13984 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 16100 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_161
timestamp 1586364061
transform 1 0 15916 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_165
timestamp 1586364061
transform 1 0 16284 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_177
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1786 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_22
timestamp 1586364061
transform 1 0 3128 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 6348 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6164 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 5520 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_41
timestamp 1586364061
transform 1 0 4876 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_46
timestamp 1586364061
transform 1 0 5336 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_50
timestamp 1586364061
transform 1 0 5704 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_54
timestamp 1586364061
transform 1 0 6072 0 -1 22304
box -38 -48 130 592
use scs8hd_conb_1  _048_
timestamp 1586364061
transform 1 0 7912 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 8372 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 7728 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_66
timestamp 1586364061
transform 1 0 7176 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_70
timestamp 1586364061
transform 1 0 7544 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_77
timestamp 1586364061
transform 1 0 8188 0 -1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8924 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_81
timestamp 1586364061
transform 1 0 8556 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_4  FILLER_36_87
timestamp 1586364061
transform 1 0 9108 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_91
timestamp 1586364061
transform 1 0 9476 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_99
timestamp 1586364061
transform 1 0 10212 0 -1 22304
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10488 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 11500 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10304 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_111
timestamp 1586364061
transform 1 0 11316 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_115
timestamp 1586364061
transform 1 0 11684 0 -1 22304
box -38 -48 774 592
use scs8hd_mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13340 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12420 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 13156 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14352 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_142
timestamp 1586364061
transform 1 0 14168 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_146
timestamp 1586364061
transform 1 0 14536 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_152
timestamp 1586364061
transform 1 0 15088 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_173
timestamp 1586364061
transform 1 0 17020 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_185
timestamp 1586364061
transform 1 0 18124 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_197
timestamp 1586364061
transform 1 0 19228 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_209
timestamp 1586364061
transform 1 0 20332 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_213
timestamp 1586364061
transform 1 0 20700 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_buf_2  _056_
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 2668 0 1 22304
box -38 -48 1786 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__056__A
timestamp 1586364061
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_11
timestamp 1586364061
transform 1 0 2116 0 1 22304
box -38 -48 406 592
use scs8hd_decap_4  FILLER_37_36
timestamp 1586364061
transform 1 0 4416 0 1 22304
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4784 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_42
timestamp 1586364061
transform 1 0 4968 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_53
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_57
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use scs8hd_mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1586364061
transform 1 0 8372 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_71
timestamp 1586364061
transform 1 0 7636 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_75
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use scs8hd_conb_1  _052_
timestamp 1586364061
transform 1 0 9936 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 9660 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_88
timestamp 1586364061
transform 1 0 9200 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_92
timestamp 1586364061
transform 1 0 9568 0 1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_37_95
timestamp 1586364061
transform 1 0 9844 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_99
timestamp 1586364061
transform 1 0 10212 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_111
timestamp 1586364061
transform 1 0 11316 0 1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_37_119
timestamp 1586364061
transform 1 0 12052 0 1 22304
box -38 -48 130 592
use scs8hd_buf_2  _098_
timestamp 1586364061
transform 1 0 12696 0 1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 13248 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13800 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_130
timestamp 1586364061
transform 1 0 13064 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_134
timestamp 1586364061
transform 1 0 13432 0 1 22304
box -38 -48 406 592
use scs8hd_buf_2  _111_
timestamp 1586364061
transform 1 0 15548 0 1 22304
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13984 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 15272 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_149
timestamp 1586364061
transform 1 0 14812 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_153
timestamp 1586364061
transform 1 0 15180 0 1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_37_156
timestamp 1586364061
transform 1 0 15456 0 1 22304
box -38 -48 130 592
use scs8hd_buf_1  mux_top_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16652 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 17112 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 16100 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17480 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_161
timestamp 1586364061
transform 1 0 15916 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_165
timestamp 1586364061
transform 1 0 16284 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_172
timestamp 1586364061
transform 1 0 16928 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_176
timestamp 1586364061
transform 1 0 17296 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18216 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_180
timestamp 1586364061
transform 1 0 17664 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_188
timestamp 1586364061
transform 1 0 18400 0 1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20884 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_200
timestamp 1586364061
transform 1 0 19504 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_37_212
timestamp 1586364061
transform 1 0 20608 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_217
timestamp 1586364061
transform 1 0 21068 0 1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22172 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_231
timestamp 1586364061
transform 1 0 22356 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_37_243
timestamp 1586364061
transform 1 0 23460 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 1748 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 1564 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 2760 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_16
timestamp 1586364061
transform 1 0 2576 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_24
timestamp 1586364061
transform 1 0 3312 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_20
timestamp 1586364061
transform 1 0 2944 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 3128 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_28
timestamp 1586364061
transform 1 0 3680 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4232 0 -1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_36
timestamp 1586364061
transform 1 0 4416 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4600 0 -1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6348 0 -1 23392
box -38 -48 1786 592
use scs8hd_mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 4784 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5888 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_49
timestamp 1586364061
transform 1 0 5612 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_38_54
timestamp 1586364061
transform 1 0 6072 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 8372 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_76
timestamp 1586364061
transform 1 0 8096 0 -1 23392
box -38 -48 314 592
use scs8hd_buf_1  mux_top_track_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_81
timestamp 1586364061
transform 1 0 8556 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_38_89
timestamp 1586364061
transform 1 0 9292 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_96
timestamp 1586364061
transform 1 0 9936 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_108
timestamp 1586364061
transform 1 0 11040 0 -1 23392
box -38 -48 1142 592
use scs8hd_conb_1  _029_
timestamp 1586364061
transform 1 0 13524 0 -1 23392
box -38 -48 314 592
use scs8hd_buf_1  mux_top_track_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12512 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_38_120
timestamp 1586364061
transform 1 0 12144 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_38_127
timestamp 1586364061
transform 1 0 12788 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_38_138
timestamp 1586364061
transform 1 0 13800 0 -1 23392
box -38 -48 222 592
use scs8hd_buf_2  _103_
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13984 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14352 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_142
timestamp 1586364061
transform 1 0 14168 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_146
timestamp 1586364061
transform 1 0 14536 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_38_152
timestamp 1586364061
transform 1 0 15088 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_158
timestamp 1586364061
transform 1 0 15640 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_2  _108_
timestamp 1586364061
transform 1 0 17020 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  FILLER_38_170
timestamp 1586364061
transform 1 0 16744 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_177
timestamp 1586364061
transform 1 0 17388 0 -1 23392
box -38 -48 774 592
use scs8hd_buf_1  mux_top_track_16.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18124 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_188
timestamp 1586364061
transform 1 0 18400 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_1  mux_top_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_200
timestamp 1586364061
transform 1 0 19504 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_38_212
timestamp 1586364061
transform 1 0 20608 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_218
timestamp 1586364061
transform 1 0 21160 0 -1 23392
box -38 -48 774 592
use scs8hd_buf_1  mux_top_track_32.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22172 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_38_226
timestamp 1586364061
transform 1 0 21896 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_232
timestamp 1586364061
transform 1 0 22448 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_244
timestamp 1586364061
transform 1 0 23552 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_256
timestamp 1586364061
transform 1 0 24656 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_38_268
timestamp 1586364061
transform 1 0 25760 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_38_274
timestamp 1586364061
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_6
timestamp 1586364061
transform 1 0 1656 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_7
timestamp 1586364061
transform 1 0 1748 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 1564 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__A
timestamp 1586364061
transform 1 0 1840 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_conb_1  _030_
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_10
timestamp 1586364061
transform 1 0 2024 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 2208 0 -1 24480
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2116 0 1 23392
box -38 -48 866 592
use scs8hd_mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1586364061
transform 1 0 2392 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_23
timestamp 1586364061
transform 1 0 3220 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_28
timestamp 1586364061
transform 1 0 3680 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_24
timestamp 1586364061
transform 1 0 3312 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_20
timestamp 1586364061
transform 1 0 2944 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 3772 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 3404 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 3128 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 3496 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 3864 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4048 0 1 23392
box -38 -48 1786 592
use scs8hd_mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5888 0 -1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_55
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_41
timestamp 1586364061
transform 1 0 4876 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_6  FILLER_40_46
timestamp 1586364061
transform 1 0 5336 0 -1 24480
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1786 592
use scs8hd_mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7452 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6900 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7268 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_61
timestamp 1586364061
transform 1 0 6716 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_65
timestamp 1586364061
transform 1 0 7084 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_78
timestamp 1586364061
transform 1 0 8280 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_89
timestamp 1586364061
transform 1 0 9292 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_85
timestamp 1586364061
transform 1 0 8924 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_81
timestamp 1586364061
transform 1 0 8556 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9108 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 8740 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_90
timestamp 1586364061
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_97
timestamp 1586364061
transform 1 0 10028 0 1 23392
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_buf_2  _112_
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_39_106
timestamp 1586364061
transform 1 0 10856 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_102
timestamp 1586364061
transform 1 0 10488 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 10672 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_118
timestamp 1586364061
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_114
timestamp 1586364061
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _100_
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _099_
timestamp 1586364061
transform 1 0 12052 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_39_127
timestamp 1586364061
transform 1 0 12788 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_buf_2  _058_
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 406 592
use scs8hd_decap_6  FILLER_40_135
timestamp 1586364061
transform 1 0 13524 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_131
timestamp 1586364061
transform 1 0 13156 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 13616 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 12972 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _059_
timestamp 1586364061
transform 1 0 13800 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_123
timestamp 1586364061
transform 1 0 12420 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_145
timestamp 1586364061
transform 1 0 14444 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_146
timestamp 1586364061
transform 1 0 14536 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_142
timestamp 1586364061
transform 1 0 14168 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 14352 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _113_
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_154
timestamp 1586364061
transform 1 0 15272 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 14720 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 15456 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_buf_2  _095_
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _094_
timestamp 1586364061
transform 1 0 14904 0 1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_40_158
timestamp 1586364061
transform 1 0 15640 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_8  FILLER_39_158
timestamp 1586364061
transform 1 0 15640 0 1 23392
box -38 -48 774 592
use scs8hd_buf_2  _096_
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _109_
timestamp 1586364061
transform 1 0 16468 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 16468 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_166
timestamp 1586364061
transform 1 0 16376 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_169
timestamp 1586364061
transform 1 0 16652 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_175
timestamp 1586364061
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_40_171
timestamp 1586364061
transform 1 0 16836 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_8  FILLER_40_183
timestamp 1586364061
transform 1 0 17940 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_188
timestamp 1586364061
transform 1 0 18400 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_179
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_buf_2  _107_
timestamp 1586364061
transform 1 0 17572 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _106_
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use scs8hd_decap_3  FILLER_39_196
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_192
timestamp 1586364061
transform 1 0 18768 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 18952 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 18584 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _105_
timestamp 1586364061
transform 1 0 18676 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_195
timestamp 1586364061
transform 1 0 19044 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_40_207
timestamp 1586364061
transform 1 0 20148 0 -1 24480
box -38 -48 590 592
use scs8hd_decap_8  FILLER_39_207
timestamp 1586364061
transform 1 0 20148 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_203
timestamp 1586364061
transform 1 0 19780 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 19964 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _104_
timestamp 1586364061
transform 1 0 19412 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_213
timestamp 1586364061
transform 1 0 20700 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 20884 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_buf_2  _102_
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_217
timestamp 1586364061
transform 1 0 21068 0 1 23392
box -38 -48 130 592
use scs8hd_buf_2  _101_
timestamp 1586364061
transform 1 0 21160 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 21712 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_222
timestamp 1586364061
transform 1 0 21528 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_226
timestamp 1586364061
transform 1 0 21896 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_39_238
timestamp 1586364061
transform 1 0 23000 0 1 23392
box -38 -48 590 592
use scs8hd_decap_12  FILLER_40_219
timestamp 1586364061
transform 1 0 21252 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_231
timestamp 1586364061
transform 1 0 22356 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _097_
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 24196 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_249
timestamp 1586364061
transform 1 0 24012 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_253
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_243
timestamp 1586364061
transform 1 0 23460 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_255
timestamp 1586364061
transform 1 0 24564 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_265
timestamp 1586364061
transform 1 0 25484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_267
timestamp 1586364061
transform 1 0 25668 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_buf_2  _057_
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2576 0 1 24480
box -38 -48 866 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 1932 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__A
timestamp 1586364061
transform 1 0 2392 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_7
timestamp 1586364061
transform 1 0 1748 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_11
timestamp 1586364061
transform 1 0 2116 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_25
timestamp 1586364061
transform 1 0 3404 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_29
timestamp 1586364061
transform 1 0 3772 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_41
timestamp 1586364061
transform 1 0 4876 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_53
timestamp 1586364061
transform 1 0 5980 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 7452 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_41_68
timestamp 1586364061
transform 1 0 7360 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_71
timestamp 1586364061
transform 1 0 7636 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_83
timestamp 1586364061
transform 1 0 8740 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_95
timestamp 1586364061
transform 1 0 9844 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_107
timestamp 1586364061
transform 1 0 10948 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_41_119
timestamp 1586364061
transform 1 0 12052 0 1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _110_
timestamp 1586364061
transform 1 0 15916 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 16468 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_165
timestamp 1586364061
transform 1 0 16284 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_169
timestamp 1586364061
transform 1 0 16652 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_181
timestamp 1586364061
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_buf_2  _054_
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 406 592
use scs8hd_buf_2  _055_
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 1932 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 2300 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_7
timestamp 1586364061
transform 1 0 1748 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_11
timestamp 1586364061
transform 1 0 2116 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_19
timestamp 1586364061
transform 1 0 2852 0 -1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 3036 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_23
timestamp 1586364061
transform 1 0 3220 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_34_
port 0 nsew default input
rlabel metal2 s 846 0 902 480 6 bottom_left_grid_pin_35_
port 1 nsew default input
rlabel metal2 s 1398 0 1454 480 6 bottom_left_grid_pin_36_
port 2 nsew default input
rlabel metal2 s 1950 0 2006 480 6 bottom_left_grid_pin_37_
port 3 nsew default input
rlabel metal2 s 2502 0 2558 480 6 bottom_left_grid_pin_38_
port 4 nsew default input
rlabel metal2 s 3146 0 3202 480 6 bottom_left_grid_pin_39_
port 5 nsew default input
rlabel metal2 s 3698 0 3754 480 6 bottom_left_grid_pin_40_
port 6 nsew default input
rlabel metal2 s 4250 0 4306 480 6 bottom_left_grid_pin_41_
port 7 nsew default input
rlabel metal2 s 27618 0 27674 480 6 bottom_right_grid_pin_1_
port 8 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 ccff_head
port 9 nsew default input
rlabel metal3 s 27520 23264 28000 23384 6 ccff_tail
port 10 nsew default tristate
rlabel metal3 s 0 280 480 400 6 chanx_left_in[0]
port 11 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[10]
port 12 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[11]
port 13 nsew default input
rlabel metal3 s 0 7216 480 7336 6 chanx_left_in[12]
port 14 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[13]
port 15 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[14]
port 16 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[15]
port 17 nsew default input
rlabel metal3 s 0 9528 480 9648 6 chanx_left_in[16]
port 18 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[17]
port 19 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[18]
port 20 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[19]
port 21 nsew default input
rlabel metal3 s 0 824 480 944 6 chanx_left_in[1]
port 22 nsew default input
rlabel metal3 s 0 1368 480 1488 6 chanx_left_in[2]
port 23 nsew default input
rlabel metal3 s 0 1912 480 2032 6 chanx_left_in[3]
port 24 nsew default input
rlabel metal3 s 0 2592 480 2712 6 chanx_left_in[4]
port 25 nsew default input
rlabel metal3 s 0 3136 480 3256 6 chanx_left_in[5]
port 26 nsew default input
rlabel metal3 s 0 3680 480 3800 6 chanx_left_in[6]
port 27 nsew default input
rlabel metal3 s 0 4360 480 4480 6 chanx_left_in[7]
port 28 nsew default input
rlabel metal3 s 0 4904 480 5024 6 chanx_left_in[8]
port 29 nsew default input
rlabel metal3 s 0 5448 480 5568 6 chanx_left_in[9]
port 30 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_out[0]
port 31 nsew default tristate
rlabel metal3 s 0 17688 480 17808 6 chanx_left_out[10]
port 32 nsew default tristate
rlabel metal3 s 0 18368 480 18488 6 chanx_left_out[11]
port 33 nsew default tristate
rlabel metal3 s 0 18912 480 19032 6 chanx_left_out[12]
port 34 nsew default tristate
rlabel metal3 s 0 19456 480 19576 6 chanx_left_out[13]
port 35 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 chanx_left_out[14]
port 36 nsew default tristate
rlabel metal3 s 0 20680 480 20800 6 chanx_left_out[15]
port 37 nsew default tristate
rlabel metal3 s 0 21224 480 21344 6 chanx_left_out[16]
port 38 nsew default tristate
rlabel metal3 s 0 21768 480 21888 6 chanx_left_out[17]
port 39 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[18]
port 40 nsew default tristate
rlabel metal3 s 0 22992 480 23112 6 chanx_left_out[19]
port 41 nsew default tristate
rlabel metal3 s 0 12520 480 12640 6 chanx_left_out[1]
port 42 nsew default tristate
rlabel metal3 s 0 13064 480 13184 6 chanx_left_out[2]
port 43 nsew default tristate
rlabel metal3 s 0 13608 480 13728 6 chanx_left_out[3]
port 44 nsew default tristate
rlabel metal3 s 0 14288 480 14408 6 chanx_left_out[4]
port 45 nsew default tristate
rlabel metal3 s 0 14832 480 14952 6 chanx_left_out[5]
port 46 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 chanx_left_out[6]
port 47 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[7]
port 48 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 chanx_left_out[8]
port 49 nsew default tristate
rlabel metal3 s 0 17144 480 17264 6 chanx_left_out[9]
port 50 nsew default tristate
rlabel metal2 s 4802 0 4858 480 6 chany_bottom_in[0]
port 51 nsew default input
rlabel metal2 s 10506 0 10562 480 6 chany_bottom_in[10]
port 52 nsew default input
rlabel metal2 s 11058 0 11114 480 6 chany_bottom_in[11]
port 53 nsew default input
rlabel metal2 s 11702 0 11758 480 6 chany_bottom_in[12]
port 54 nsew default input
rlabel metal2 s 12254 0 12310 480 6 chany_bottom_in[13]
port 55 nsew default input
rlabel metal2 s 12806 0 12862 480 6 chany_bottom_in[14]
port 56 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[15]
port 57 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_in[16]
port 58 nsew default input
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_in[17]
port 59 nsew default input
rlabel metal2 s 15106 0 15162 480 6 chany_bottom_in[18]
port 60 nsew default input
rlabel metal2 s 15658 0 15714 480 6 chany_bottom_in[19]
port 61 nsew default input
rlabel metal2 s 5354 0 5410 480 6 chany_bottom_in[1]
port 62 nsew default input
rlabel metal2 s 5998 0 6054 480 6 chany_bottom_in[2]
port 63 nsew default input
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_in[3]
port 64 nsew default input
rlabel metal2 s 7102 0 7158 480 6 chany_bottom_in[4]
port 65 nsew default input
rlabel metal2 s 7654 0 7710 480 6 chany_bottom_in[5]
port 66 nsew default input
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[6]
port 67 nsew default input
rlabel metal2 s 8850 0 8906 480 6 chany_bottom_in[7]
port 68 nsew default input
rlabel metal2 s 9402 0 9458 480 6 chany_bottom_in[8]
port 69 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[9]
port 70 nsew default input
rlabel metal2 s 16210 0 16266 480 6 chany_bottom_out[0]
port 71 nsew default tristate
rlabel metal2 s 21914 0 21970 480 6 chany_bottom_out[10]
port 72 nsew default tristate
rlabel metal2 s 22466 0 22522 480 6 chany_bottom_out[11]
port 73 nsew default tristate
rlabel metal2 s 23110 0 23166 480 6 chany_bottom_out[12]
port 74 nsew default tristate
rlabel metal2 s 23662 0 23718 480 6 chany_bottom_out[13]
port 75 nsew default tristate
rlabel metal2 s 24214 0 24270 480 6 chany_bottom_out[14]
port 76 nsew default tristate
rlabel metal2 s 24766 0 24822 480 6 chany_bottom_out[15]
port 77 nsew default tristate
rlabel metal2 s 25318 0 25374 480 6 chany_bottom_out[16]
port 78 nsew default tristate
rlabel metal2 s 25962 0 26018 480 6 chany_bottom_out[17]
port 79 nsew default tristate
rlabel metal2 s 26514 0 26570 480 6 chany_bottom_out[18]
port 80 nsew default tristate
rlabel metal2 s 27066 0 27122 480 6 chany_bottom_out[19]
port 81 nsew default tristate
rlabel metal2 s 16762 0 16818 480 6 chany_bottom_out[1]
port 82 nsew default tristate
rlabel metal2 s 17406 0 17462 480 6 chany_bottom_out[2]
port 83 nsew default tristate
rlabel metal2 s 17958 0 18014 480 6 chany_bottom_out[3]
port 84 nsew default tristate
rlabel metal2 s 18510 0 18566 480 6 chany_bottom_out[4]
port 85 nsew default tristate
rlabel metal2 s 19062 0 19118 480 6 chany_bottom_out[5]
port 86 nsew default tristate
rlabel metal2 s 19614 0 19670 480 6 chany_bottom_out[6]
port 87 nsew default tristate
rlabel metal2 s 20258 0 20314 480 6 chany_bottom_out[7]
port 88 nsew default tristate
rlabel metal2 s 20810 0 20866 480 6 chany_bottom_out[8]
port 89 nsew default tristate
rlabel metal2 s 21362 0 21418 480 6 chany_bottom_out[9]
port 90 nsew default tristate
rlabel metal2 s 4802 27520 4858 28000 6 chany_top_in[0]
port 91 nsew default input
rlabel metal2 s 10506 27520 10562 28000 6 chany_top_in[10]
port 92 nsew default input
rlabel metal2 s 11058 27520 11114 28000 6 chany_top_in[11]
port 93 nsew default input
rlabel metal2 s 11702 27520 11758 28000 6 chany_top_in[12]
port 94 nsew default input
rlabel metal2 s 12254 27520 12310 28000 6 chany_top_in[13]
port 95 nsew default input
rlabel metal2 s 12806 27520 12862 28000 6 chany_top_in[14]
port 96 nsew default input
rlabel metal2 s 13358 27520 13414 28000 6 chany_top_in[15]
port 97 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_in[16]
port 98 nsew default input
rlabel metal2 s 14554 27520 14610 28000 6 chany_top_in[17]
port 99 nsew default input
rlabel metal2 s 15106 27520 15162 28000 6 chany_top_in[18]
port 100 nsew default input
rlabel metal2 s 15658 27520 15714 28000 6 chany_top_in[19]
port 101 nsew default input
rlabel metal2 s 5354 27520 5410 28000 6 chany_top_in[1]
port 102 nsew default input
rlabel metal2 s 5998 27520 6054 28000 6 chany_top_in[2]
port 103 nsew default input
rlabel metal2 s 6550 27520 6606 28000 6 chany_top_in[3]
port 104 nsew default input
rlabel metal2 s 7102 27520 7158 28000 6 chany_top_in[4]
port 105 nsew default input
rlabel metal2 s 7654 27520 7710 28000 6 chany_top_in[5]
port 106 nsew default input
rlabel metal2 s 8206 27520 8262 28000 6 chany_top_in[6]
port 107 nsew default input
rlabel metal2 s 8850 27520 8906 28000 6 chany_top_in[7]
port 108 nsew default input
rlabel metal2 s 9402 27520 9458 28000 6 chany_top_in[8]
port 109 nsew default input
rlabel metal2 s 9954 27520 10010 28000 6 chany_top_in[9]
port 110 nsew default input
rlabel metal2 s 16210 27520 16266 28000 6 chany_top_out[0]
port 111 nsew default tristate
rlabel metal2 s 21914 27520 21970 28000 6 chany_top_out[10]
port 112 nsew default tristate
rlabel metal2 s 22466 27520 22522 28000 6 chany_top_out[11]
port 113 nsew default tristate
rlabel metal2 s 23110 27520 23166 28000 6 chany_top_out[12]
port 114 nsew default tristate
rlabel metal2 s 23662 27520 23718 28000 6 chany_top_out[13]
port 115 nsew default tristate
rlabel metal2 s 24214 27520 24270 28000 6 chany_top_out[14]
port 116 nsew default tristate
rlabel metal2 s 24766 27520 24822 28000 6 chany_top_out[15]
port 117 nsew default tristate
rlabel metal2 s 25318 27520 25374 28000 6 chany_top_out[16]
port 118 nsew default tristate
rlabel metal2 s 25962 27520 26018 28000 6 chany_top_out[17]
port 119 nsew default tristate
rlabel metal2 s 26514 27520 26570 28000 6 chany_top_out[18]
port 120 nsew default tristate
rlabel metal2 s 27066 27520 27122 28000 6 chany_top_out[19]
port 121 nsew default tristate
rlabel metal2 s 16762 27520 16818 28000 6 chany_top_out[1]
port 122 nsew default tristate
rlabel metal2 s 17406 27520 17462 28000 6 chany_top_out[2]
port 123 nsew default tristate
rlabel metal2 s 17958 27520 18014 28000 6 chany_top_out[3]
port 124 nsew default tristate
rlabel metal2 s 18510 27520 18566 28000 6 chany_top_out[4]
port 125 nsew default tristate
rlabel metal2 s 19062 27520 19118 28000 6 chany_top_out[5]
port 126 nsew default tristate
rlabel metal2 s 19614 27520 19670 28000 6 chany_top_out[6]
port 127 nsew default tristate
rlabel metal2 s 20258 27520 20314 28000 6 chany_top_out[7]
port 128 nsew default tristate
rlabel metal2 s 20810 27520 20866 28000 6 chany_top_out[8]
port 129 nsew default tristate
rlabel metal2 s 21362 27520 21418 28000 6 chany_top_out[9]
port 130 nsew default tristate
rlabel metal3 s 0 23536 480 23656 6 left_top_grid_pin_42_
port 131 nsew default input
rlabel metal3 s 0 24080 480 24200 6 left_top_grid_pin_43_
port 132 nsew default input
rlabel metal3 s 0 24760 480 24880 6 left_top_grid_pin_44_
port 133 nsew default input
rlabel metal3 s 0 25304 480 25424 6 left_top_grid_pin_45_
port 134 nsew default input
rlabel metal3 s 0 25848 480 25968 6 left_top_grid_pin_46_
port 135 nsew default input
rlabel metal3 s 0 26528 480 26648 6 left_top_grid_pin_47_
port 136 nsew default input
rlabel metal3 s 0 27072 480 27192 6 left_top_grid_pin_48_
port 137 nsew default input
rlabel metal3 s 0 27616 480 27736 6 left_top_grid_pin_49_
port 138 nsew default input
rlabel metal3 s 27520 4632 28000 4752 6 prog_clk
port 139 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_34_
port 140 nsew default input
rlabel metal2 s 846 27520 902 28000 6 top_left_grid_pin_35_
port 141 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 top_left_grid_pin_36_
port 142 nsew default input
rlabel metal2 s 1950 27520 2006 28000 6 top_left_grid_pin_37_
port 143 nsew default input
rlabel metal2 s 2502 27520 2558 28000 6 top_left_grid_pin_38_
port 144 nsew default input
rlabel metal2 s 3146 27520 3202 28000 6 top_left_grid_pin_39_
port 145 nsew default input
rlabel metal2 s 3698 27520 3754 28000 6 top_left_grid_pin_40_
port 146 nsew default input
rlabel metal2 s 4250 27520 4306 28000 6 top_left_grid_pin_41_
port 147 nsew default input
rlabel metal2 s 27618 27520 27674 28000 6 top_right_grid_pin_1_
port 148 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 149 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 150 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
