VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cby_1__1_
  CLASS BLOCK ;
  FOREIGN cby_1__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 200.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 2.400 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 2.400 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 2.400 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 2.400 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 2.400 ;
    END
  END address[5]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.930 197.600 2.210 200.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.070 197.600 6.350 200.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.670 197.600 10.950 200.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.270 197.600 15.550 200.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.410 197.600 19.690 200.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 197.600 24.290 200.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 197.600 28.890 200.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.750 197.600 33.030 200.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.350 197.600 37.630 200.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.950 197.600 42.230 200.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 46.090 197.600 46.370 200.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 50.690 197.600 50.970 200.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 55.290 197.600 55.570 200.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.430 197.600 59.710 200.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.030 197.600 64.310 200.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.630 197.600 68.910 200.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.770 197.600 73.050 200.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.370 197.600 77.650 200.000 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 2.400 ;
    END
  END enable
  PIN left_grid_pin_1_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.400 33.960 ;
    END
  END left_grid_pin_1_
  PIN left_grid_pin_5_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END left_grid_pin_5_
  PIN left_grid_pin_9_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 2.400 167.240 ;
    END
  END left_grid_pin_9_
  PIN right_grid_pin_3_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 49.680 80.000 50.280 ;
    END
  END right_grid_pin_3_
  PIN right_grid_pin_7_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 149.640 80.000 150.240 ;
    END
  END right_grid_pin_7_
  PIN vpwr
    USE POWER ;
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 18.055 10.640 19.655 187.920 ;
    END
  END vpwr
  PIN vgnd
    USE GROUND ;
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 31.385 10.640 32.985 187.920 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 74.060 187.765 ;
      LAYER met1 ;
        RECT 0.070 0.040 79.050 198.520 ;
      LAYER met2 ;
        RECT 0.100 197.320 1.650 198.550 ;
        RECT 2.490 197.320 5.790 198.550 ;
        RECT 6.630 197.320 10.390 198.550 ;
        RECT 11.230 197.320 14.990 198.550 ;
        RECT 15.830 197.320 19.130 198.550 ;
        RECT 19.970 197.320 23.730 198.550 ;
        RECT 24.570 197.320 28.330 198.550 ;
        RECT 29.170 197.320 32.470 198.550 ;
        RECT 33.310 197.320 37.070 198.550 ;
        RECT 37.910 197.320 41.670 198.550 ;
        RECT 42.510 197.320 45.810 198.550 ;
        RECT 46.650 197.320 50.410 198.550 ;
        RECT 51.250 197.320 55.010 198.550 ;
        RECT 55.850 197.320 59.150 198.550 ;
        RECT 59.990 197.320 63.750 198.550 ;
        RECT 64.590 197.320 68.350 198.550 ;
        RECT 69.190 197.320 72.490 198.550 ;
        RECT 73.330 197.320 77.090 198.550 ;
        RECT 77.930 197.320 79.020 198.550 ;
        RECT 0.100 2.680 79.020 197.320 ;
        RECT 0.100 0.010 1.190 2.680 ;
        RECT 2.030 0.010 3.950 2.680 ;
        RECT 4.790 0.010 7.170 2.680 ;
        RECT 8.010 0.010 10.390 2.680 ;
        RECT 11.230 0.010 13.150 2.680 ;
        RECT 13.990 0.010 16.370 2.680 ;
        RECT 17.210 0.010 19.590 2.680 ;
        RECT 20.430 0.010 22.350 2.680 ;
        RECT 23.190 0.010 25.570 2.680 ;
        RECT 26.410 0.010 28.790 2.680 ;
        RECT 29.630 0.010 31.550 2.680 ;
        RECT 32.390 0.010 34.770 2.680 ;
        RECT 35.610 0.010 37.990 2.680 ;
        RECT 38.830 0.010 41.210 2.680 ;
        RECT 42.050 0.010 43.970 2.680 ;
        RECT 44.810 0.010 47.190 2.680 ;
        RECT 48.030 0.010 50.410 2.680 ;
        RECT 51.250 0.010 53.170 2.680 ;
        RECT 54.010 0.010 56.390 2.680 ;
        RECT 57.230 0.010 59.610 2.680 ;
        RECT 60.450 0.010 62.370 2.680 ;
        RECT 63.210 0.010 65.590 2.680 ;
        RECT 66.430 0.010 68.810 2.680 ;
        RECT 69.650 0.010 71.570 2.680 ;
        RECT 72.410 0.010 74.790 2.680 ;
        RECT 75.630 0.010 78.010 2.680 ;
        RECT 78.850 0.010 79.020 2.680 ;
      LAYER met3 ;
        RECT 0.270 167.640 77.890 187.845 ;
        RECT 2.800 166.240 77.890 167.640 ;
        RECT 0.270 150.640 77.890 166.240 ;
        RECT 0.270 149.240 77.200 150.640 ;
        RECT 0.270 101.000 77.890 149.240 ;
        RECT 2.800 99.600 77.890 101.000 ;
        RECT 0.270 50.680 77.890 99.600 ;
        RECT 0.270 49.280 77.200 50.680 ;
        RECT 0.270 34.360 77.890 49.280 ;
        RECT 2.800 32.960 77.890 34.360 ;
        RECT 0.270 6.295 77.890 32.960 ;
      LAYER met4 ;
        RECT 0.295 10.640 17.655 187.920 ;
        RECT 20.055 10.640 30.985 187.920 ;
        RECT 33.385 10.640 72.985 187.920 ;
  END
END cby_1__1_
END LIBRARY

