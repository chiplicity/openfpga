VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tie_array
  CLASS BLOCK ;
  FOREIGN tie_array ;
  ORIGIN 0.000 0.000 ;
  SIZE 52.300 BY 57.360 ;
  PIN x[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.020 0.000 0.300 4.000 ;
    END
  END x[0]
  PIN x[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.380 0.000 7.660 4.000 ;
    END
  END x[1]
  PIN x[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.740 0.000 15.020 4.000 ;
    END
  END x[2]
  PIN x[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.100 0.000 22.380 4.000 ;
    END
  END x[3]
  PIN x[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.920 0.000 30.200 4.000 ;
    END
  END x[4]
  PIN x[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.280 0.000 37.560 4.000 ;
    END
  END x[5]
  PIN x[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.640 0.000 44.920 4.000 ;
    END
  END x[6]
  PIN x[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.000 0.000 52.280 4.000 ;
    END
  END x[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 41.770 10.640 43.370 57.360 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 25.450 10.640 27.050 57.360 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.130 10.640 10.730 57.360 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 33.610 10.640 35.210 57.360 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 17.290 10.640 18.890 57.360 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.770 10.795 50.530 57.205 ;
      LAYER met1 ;
        RECT 0.000 10.640 52.300 57.360 ;
      LAYER met2 ;
        RECT 0.030 4.280 52.270 57.360 ;
        RECT 0.580 4.000 7.100 4.280 ;
        RECT 7.940 4.000 14.460 4.280 ;
        RECT 15.300 4.000 21.820 4.280 ;
        RECT 22.660 4.000 29.640 4.280 ;
        RECT 30.480 4.000 37.000 4.280 ;
        RECT 37.840 4.000 44.360 4.280 ;
        RECT 45.200 4.000 51.720 4.280 ;
      LAYER met3 ;
        RECT 9.130 10.715 43.370 57.285 ;
  END
END tie_array
END LIBRARY

