* NGSPICE file created from cbx_1__2_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 D Q CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VNB VPB VPWR
.ends

.subckt cbx_1__2_ SC_IN_BOT SC_IN_TOP SC_OUT_BOT SC_OUT_TOP bottom_grid_pin_0_ bottom_grid_pin_10_
+ bottom_grid_pin_11_ bottom_grid_pin_12_ bottom_grid_pin_13_ bottom_grid_pin_14_
+ bottom_grid_pin_15_ bottom_grid_pin_1_ bottom_grid_pin_2_ bottom_grid_pin_3_ bottom_grid_pin_4_
+ bottom_grid_pin_5_ bottom_grid_pin_6_ bottom_grid_pin_7_ bottom_grid_pin_8_ bottom_grid_pin_9_
+ bottom_width_0_height_0__pin_0_ bottom_width_0_height_0__pin_1_lower bottom_width_0_height_0__pin_1_upper
+ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11] chanx_left_in[12]
+ chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16] chanx_left_in[17]
+ chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3]
+ chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8]
+ chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11] chanx_left_out[12]
+ chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16] chanx_left_out[17]
+ chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3]
+ chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8]
+ chanx_left_out[9] chanx_right_in[0] chanx_right_in[10] chanx_right_in[11] chanx_right_in[12]
+ chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16] chanx_right_in[17]
+ chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11] chanx_right_out[12]
+ chanx_right_out[13] chanx_right_out[14] chanx_right_out[15] chanx_right_out[16]
+ chanx_right_out[17] chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chanx_right_out[9] gfpga_pad_EMBEDDED_IO_SOC_DIR gfpga_pad_EMBEDDED_IO_SOC_IN
+ gfpga_pad_EMBEDDED_IO_SOC_OUT prog_clk top_grid_pin_0_ VPWR VGND
XANTENNA_mux_top_ipin_7.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_7.mux_l4_in_0_/S mux_top_ipin_8.mux_l1_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_7_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_1__S mux_top_ipin_0.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_12.mux_l2_in_0__A1 mux_top_ipin_12.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_13.mux_l3_in_0_ mux_top_ipin_13.mux_l2_in_1_/X mux_top_ipin_13.mux_l2_in_0_/X
+ mux_top_ipin_13.mux_l3_in_1_/S mux_top_ipin_13.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_66_ chanx_left_in[12] chanx_right_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_2_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_10.mux_l2_in_2__A1 chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_6.mux_l2_in_0_ chanx_left_in[3] mux_top_ipin_6.mux_l1_in_0_/X mux_top_ipin_6.mux_l2_in_0_/S
+ mux_top_ipin_6.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_0.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_7.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_5.mux_l2_in_2__S mux_top_ipin_5.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l2_in_1__A1 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_1_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_49_ chanx_right_in[9] chanx_left_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xclkbuf_3_4_0_prog_clk clkbuf_2_2_0_prog_clk/X clkbuf_3_4_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_12.mux_l1_in_0__S mux_top_ipin_12.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_13.mux_l2_in_1_ chanx_left_in[10] chanx_right_in[2] mux_top_ipin_13.mux_l2_in_3_/S
+ mux_top_ipin_13.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_1_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_9.mux_l3_in_0__S mux_top_ipin_9.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_10.mux_l3_in_1__A1 mux_top_ipin_10.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_3.mux_l2_in_3__A1 chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_2.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l3_in_0__A1 mux_top_ipin_5.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D ccff_head VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_3_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_11.mux_l2_in_0__S mux_top_ipin_11.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_10.mux_l4_in_0__A1 mux_top_ipin_10.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_8.mux_l4_in_0__S mux_top_ipin_8.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_0.mux_l1_in_2__A0 chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_1.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_1.mux_l1_in_0_/S
+ mux_top_ipin_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_3.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_10.mux_l3_in_0__S mux_top_ipin_10.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_0.mux_l2_in_1__A0 chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_65_ chanx_left_in[13] chanx_right_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__D mux_bottom_ipin_0.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_48_ chanx_right_in[10] chanx_left_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_0.mux_l3_in_0__A0 mux_top_ipin_0.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_13.mux_l2_in_0_ chanx_left_in[2] mux_top_ipin_13.mux_l1_in_0_/X mux_top_ipin_13.mux_l2_in_3_/S
+ mux_top_ipin_13.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_11.mux_l2_in_3__S mux_top_ipin_11.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_15.mux_l3_in_1__S mux_top_ipin_15.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_6.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_6.mux_l1_in_0_/S
+ mux_top_ipin_6.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_2.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_6.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_14.mux_l2_in_1__A0 chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_9.mux_l2_in_0__A0 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ mux_bottom_ipin_0.mux_l3_in_1_/S mux_bottom_ipin_0.mux_l4_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_0.mux_l1_in_2__A1 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_12.mux_l2_in_3__A0 _26_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_14.mux_l3_in_0__A0 mux_top_ipin_14.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_7.mux_l2_in_2__A0 chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_0__S mux_top_ipin_7.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_14.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_1__A1 mux_top_ipin_0.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_64_ chanx_left_in[14] chanx_right_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_5_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_4.mux_l4_in_0_/X bottom_grid_pin_4_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_23_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_7.mux_l3_in_1__A0 mux_top_ipin_7.mux_l2_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_9.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0__S mux_top_ipin_6.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_47_ chanx_right_in[11] chanx_left_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_0.mux_l3_in_0__A1 mux_top_ipin_0.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0__S mux_bottom_ipin_0.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_7.mux_l4_in_0__A0 mux_top_ipin_7.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_1.mux_l2_in_2__S mux_top_ipin_1.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_7_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l2_in_1__A1 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_5.mux_l3_in_0__S mux_top_ipin_5.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_13.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_13.mux_l1_in_0_/S
+ mux_top_ipin_13.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_9.mux_l2_in_0__A1 mux_top_ipin_9.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ mux_bottom_ipin_0.mux_l2_in_3_/S mux_bottom_ipin_0.mux_l3_in_1_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_1_0_prog_clk clkbuf_0_prog_clk/X clkbuf_3_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_top_ipin_12.mux_l2_in_3__A1 chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_11.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_14.mux_l3_in_0__A1 mux_top_ipin_14.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_80_ bottom_width_0_height_0__pin_0_ gfpga_pad_EMBEDDED_IO_SOC_OUT VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__buf_2
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_7.mux_l2_in_2__A1 chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_6.mux_l2_in_3__S mux_top_ipin_6.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_4.mux_l4_in_0__S mux_top_ipin_4.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_63_ chanx_left_in[15] chanx_right_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_4.mux_l1_in_1__A0 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_7.mux_l3_in_1__A1 mux_top_ipin_7.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_1_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_46_ chanx_right_in[12] chanx_left_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_12.mux_l2_in_1__S mux_top_ipin_12.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29_ _29_/HI _29_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_ipin_7.mux_l4_in_0__A1 mux_top_ipin_7.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_4.mux_l2_in_0__A0 mux_top_ipin_4.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_6_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_11.mux_l4_in_0_/X bottom_grid_pin_11_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xclkbuf_3_3_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_3_3_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_10.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_bottom_ipin_0.mux_l4_in_0_/X top_grid_pin_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_2.mux_l2_in_2__A0 chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_11.mux_l3_in_1__S mux_top_ipin_11.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_11.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_ipin_0.mux_l1_in_1_/S mux_bottom_ipin_0.mux_l2_in_3_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_11.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_2.mux_l2_in_3_ _30_/HI chanx_right_in[15] mux_top_ipin_2.mux_l2_in_2_/S
+ mux_top_ipin_2.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_2.mux_l3_in_1__A0 mux_top_ipin_2.mux_l2_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_62_ chanx_left_in[16] chanx_right_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_3.mux_l1_in_0__S mux_top_ipin_3.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_5.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_4.mux_l1_in_1__A1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_2.mux_l4_in_0__A0 mux_top_ipin_2.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_13.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_45_ chanx_right_in[13] chanx_left_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_2.mux_l4_in_0_ mux_top_ipin_2.mux_l3_in_1_/X mux_top_ipin_2.mux_l3_in_0_/X
+ mux_top_ipin_2.mux_l4_in_0_/S mux_top_ipin_2.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28_ _28_/HI _28_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_ipin_4.mux_l2_in_0__A1 mux_top_ipin_4.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_7.mux_l2_in_3_ _18_/HI chanx_right_in[18] mux_top_ipin_7.mux_l2_in_2_/S
+ mux_top_ipin_7.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_2.mux_l2_in_0__S mux_top_ipin_2.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_2.mux_l3_in_1_ mux_top_ipin_2.mux_l2_in_3_/X mux_top_ipin_2.mux_l2_in_2_/X
+ mux_top_ipin_2.mux_l3_in_1_/S mux_top_ipin_2.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_9.mux_l2_in_3__A0 _20_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_8.mux_l1_in_1__S mux_top_ipin_8.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_2.mux_l2_in_2__A1 chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ ccff_head mux_bottom_ipin_0.mux_l1_in_1_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_1.mux_l3_in_0__S mux_top_ipin_1.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_6.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_2.mux_l2_in_2_ chanx_left_in[15] chanx_right_in[7] mux_top_ipin_2.mux_l2_in_2_/S
+ mux_top_ipin_2.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_7.mux_l4_in_0_ mux_top_ipin_7.mux_l3_in_1_/X mux_top_ipin_7.mux_l3_in_0_/X
+ mux_top_ipin_7.mux_l4_in_0_/S mux_top_ipin_7.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_7.mux_l2_in_1__S mux_top_ipin_7.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_2.mux_l3_in_1__A1 mux_top_ipin_2.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_5_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_61_ chanx_left_in[17] chanx_right_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_2.mux_l2_in_3__S mux_top_ipin_2.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_0.mux_l4_in_0__S mux_top_ipin_0.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_7.mux_l3_in_1_ mux_top_ipin_7.mux_l2_in_3_/X mux_top_ipin_7.mux_l2_in_2_/X
+ mux_top_ipin_7.mux_l3_in_1_/S mux_top_ipin_7.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_2.mux_l4_in_0__A1 mux_top_ipin_2.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_7_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_44_ chanx_right_in[14] chanx_left_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_6.mux_l3_in_1__S mux_top_ipin_6.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_3_0_prog_clk_A clkbuf_3_3_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_1__S mux_bottom_ipin_0.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_27_ _27_/HI _27_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_7.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[12] mux_top_ipin_7.mux_l2_in_2_/S
+ mux_top_ipin_7.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__34__A SC_IN_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_2.mux_l3_in_0_ mux_top_ipin_2.mux_l2_in_1_/X mux_top_ipin_2.mux_l2_in_0_/X
+ mux_top_ipin_2.mux_l3_in_1_/S mux_top_ipin_2.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_9.mux_l2_in_3__A1 chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_8.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_14.mux_l2_in_3_ _28_/HI chanx_right_in[19] mux_top_ipin_14.mux_l2_in_1_/S
+ mux_top_ipin_14.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_13.mux_l2_in_0__A0 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_2.mux_l2_in_1_ chanx_left_in[7] chanx_right_in[3] mux_top_ipin_2.mux_l2_in_2_/S
+ mux_top_ipin_2.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_13.mux_l2_in_2__S mux_top_ipin_13.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_11.mux_l2_in_2__A0 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__42__A chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
X_60_ chanx_left_in[18] chanx_right_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_14.mux_l4_in_0_ mux_top_ipin_14.mux_l3_in_1_/X mux_top_ipin_14.mux_l3_in_0_/X
+ mux_top_ipin_14.mux_l4_in_0_/S mux_top_ipin_14.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_6.mux_l2_in_1__A0 chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_2_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_7.mux_l3_in_0_ mux_top_ipin_7.mux_l2_in_1_/X mux_top_ipin_7.mux_l2_in_0_/X
+ mux_top_ipin_7.mux_l3_in_1_/S mux_top_ipin_7.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA__37__A gfpga_pad_EMBEDDED_IO_SOC_IN VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_11.mux_l3_in_1__A0 mux_top_ipin_11.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_43_ chanx_right_in[15] chanx_left_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_7.mux_l4_in_0_/X bottom_grid_pin_7_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_ipin_4.mux_l2_in_3__A0 _32_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_14.mux_l3_in_1_ mux_top_ipin_14.mux_l2_in_3_/X mux_top_ipin_14.mux_l2_in_2_/X
+ mux_top_ipin_14.mux_l3_in_1_/S mux_top_ipin_14.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_6.mux_l3_in_0__A0 mux_top_ipin_6.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_6_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26_ _26_/HI _26_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_top_ipin_7.mux_l2_in_1_ chanx_left_in[12] mux_top_ipin_7.mux_l1_in_2_/X mux_top_ipin_7.mux_l2_in_2_/S
+ mux_top_ipin_7.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_11.mux_l4_in_0__A0 mux_top_ipin_11.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__50__A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A0 mux_bottom_ipin_0.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_13.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_3.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_14.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[11] mux_top_ipin_14.mux_l2_in_1_/S
+ mux_top_ipin_14.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__45__A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_7.mux_l1_in_2_ chanx_right_in[8] chanx_left_in[8] mux_top_ipin_7.mux_l1_in_0_/S
+ mux_top_ipin_7.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_13.mux_l2_in_0__A1 mux_top_ipin_13.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_4.mux_l1_in_1__S mux_top_ipin_4.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_2_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_3_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_2.mux_l2_in_0_ chanx_left_in[3] mux_top_ipin_2.mux_l1_in_0_/X mux_top_ipin_2.mux_l2_in_2_/S
+ mux_top_ipin_2.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_11.mux_l2_in_2__A1 chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_6.mux_l2_in_1__A1 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_3.mux_l2_in_1__S mux_top_ipin_3.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_1.mux_l3_in_1_/S mux_top_ipin_1.mux_l4_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA__53__A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_11.mux_l3_in_1__A1 mux_top_ipin_11.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_42_ chanx_right_in[16] chanx_left_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_4.mux_l2_in_3__A1 chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_14.mux_l3_in_0_ mux_top_ipin_14.mux_l2_in_1_/X mux_top_ipin_14.mux_l2_in_0_/X
+ mux_top_ipin_14.mux_l3_in_1_/S mux_top_ipin_14.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA__48__A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l3_in_0__A1 mux_top_ipin_6.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_11.mux_l3_in_1_/S mux_top_ipin_11.mux_l4_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_25_ _25_/HI _25_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_top_ipin_7.mux_l2_in_0_ mux_top_ipin_7.mux_l1_in_1_/X mux_top_ipin_7.mux_l1_in_0_/X
+ mux_top_ipin_7.mux_l2_in_2_/S mux_top_ipin_7.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_2.mux_l3_in_1__S mux_top_ipin_2.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_11.mux_l4_in_0__A1 mux_top_ipin_11.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A1 mux_bottom_ipin_0.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_2_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l2_in_2__S mux_top_ipin_8.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_15.mux_l1_in_0__S mux_top_ipin_15.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_14.mux_l2_in_1_ chanx_left_in[11] chanx_right_in[3] mux_top_ipin_14.mux_l2_in_1_/S
+ mux_top_ipin_14.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_14.mux_l4_in_0_/X bottom_grid_pin_14_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__61__A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_7.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_7.mux_l1_in_0_/S
+ mux_top_ipin_7.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_1.mux_l2_in_1__A0 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__56__A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_5_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_4.mux_l3_in_0_/S mux_top_ipin_4.mux_l4_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_16_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_14.mux_l2_in_0__S mux_top_ipin_14.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_14.mux_l3_in_1_/S mux_top_ipin_14.mux_l4_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_4_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_2.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_2.mux_l1_in_0_/S
+ mux_top_ipin_2.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_1.mux_l3_in_0__A0 mux_top_ipin_1.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_7_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_15.mux_l1_in_2__A0 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_1.mux_l2_in_0_/S mux_top_ipin_1.mux_l3_in_1_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_41_ chanx_right_in[17] chanx_left_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_9_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_13.mux_l3_in_0__S mux_top_ipin_13.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__64__A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_11.mux_l2_in_3_/S mux_top_ipin_11.mux_l3_in_1_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_6_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_15.mux_l2_in_1__A0 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24_ _24_/HI _24_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__59__A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_7.mux_l3_in_1_/S mux_top_ipin_7.mux_l4_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_13.mux_l2_in_3__A0 _27_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_14.mux_l2_in_0_ chanx_left_in[3] mux_top_ipin_14.mux_l1_in_0_/X mux_top_ipin_14.mux_l2_in_1_/S
+ mux_top_ipin_14.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_14.mux_l2_in_3__S mux_top_ipin_14.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_0.mux_l4_in_0_/X bottom_grid_pin_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_ipin_12.mux_l4_in_0__S mux_top_ipin_12.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_15.mux_l3_in_0__A0 mux_top_ipin_15.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_7.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_7.mux_l1_in_0_/S
+ mux_top_ipin_7.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_8.mux_l2_in_2__A0 chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_2_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_14.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_4.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_1.mux_l2_in_1__A1 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_4.mux_l2_in_0_/S mux_top_ipin_4.mux_l3_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA__72__A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_0.mux_l1_in_1__S mux_top_ipin_0.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l3_in_1__A0 mux_top_ipin_8.mux_l2_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__67__A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_14.mux_l2_in_1_/S mux_top_ipin_14.mux_l3_in_1_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_1.mux_l3_in_0__A1 mux_top_ipin_1.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_15.mux_l1_in_2__A1 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_1.mux_l1_in_0_/S mux_top_ipin_1.mux_l2_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_40_ chanx_right_in[18] chanx_left_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_4_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l4_in_0__A0 mux_top_ipin_8.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__80__A bottom_width_0_height_0__pin_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A0 _21_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_11.mux_l1_in_2_/S mux_top_ipin_11.mux_l2_in_3_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_15.mux_l2_in_1__A1 mux_top_ipin_15.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23_ _23_/HI _23_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_15.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_5.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__75__A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_7.mux_l2_in_2_/S mux_top_ipin_7.mux_l3_in_1_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_9.mux_l2_in_0__S mux_top_ipin_9.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_13.mux_l2_in_3__A1 chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_12.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_15.mux_l3_in_0__A1 mux_top_ipin_15.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_8.mux_l2_in_2__A1 chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_4.mux_l2_in_2__S mux_top_ipin_4.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_11.mux_l1_in_0__S mux_top_ipin_11.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_4.mux_l1_in_2_/S mux_top_ipin_4.mux_l2_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_8_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_14.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_14.mux_l1_in_0_/S
+ mux_top_ipin_14.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_8.mux_l3_in_0__S mux_top_ipin_8.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_8.mux_l3_in_1__A1 mux_top_ipin_8.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_14.mux_l1_in_0_/S mux_top_ipin_14.mux_l2_in_1_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_1_0_prog_clk clkbuf_2_0_0_prog_clk/X clkbuf_3_1_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_10.mux_l2_in_1__A0 chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_0.mux_l4_in_0_/S mux_top_ipin_1.mux_l1_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_10.mux_l2_in_0__S mux_top_ipin_10.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__78__A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_9.mux_l2_in_3__S mux_top_ipin_9.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_7.mux_l4_in_0__S mux_top_ipin_7.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_5.mux_l2_in_0__A0 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l4_in_0__A1 mux_top_ipin_8.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1 chanx_right_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_10.mux_l4_in_0_/S mux_top_ipin_11.mux_l1_in_2_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_6_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22_ _22_/HI _22_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_ipin_10.mux_l3_in_0__A0 mux_top_ipin_10.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_3.mux_l2_in_2__A0 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_7.mux_l1_in_0_/S mux_top_ipin_7.mux_l2_in_2_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_15.mux_l2_in_1__S mux_top_ipin_15.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_12.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_0.mux_l4_in_0__S mux_bottom_ipin_0.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_6_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l3_in_1__A0 mux_top_ipin_3.mux_l2_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_10.mux_l2_in_3__S mux_top_ipin_10.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_3.mux_l4_in_0_/S mux_top_ipin_4.mux_l1_in_2_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_32_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_14.mux_l3_in_1__S mux_top_ipin_14.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_3.mux_l4_in_0__A0 mux_top_ipin_3.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_13.mux_l4_in_0_/S mux_top_ipin_14.mux_l1_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_4_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_10.mux_l2_in_1__A1 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_3.mux_l2_in_3_ _31_/HI chanx_right_in[14] mux_top_ipin_3.mux_l2_in_2_/S
+ mux_top_ipin_3.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_2_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_12.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_2.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0__A1 mux_top_ipin_5.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21_ _21_/HI _21_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_ipin_10.mux_l3_in_0__A1 mux_top_ipin_10.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_1_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0__S mux_top_ipin_6.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l2_in_2__A1 chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_6.mux_l4_in_0_/S mux_top_ipin_7.mux_l1_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_3.mux_l4_in_0_ mux_top_ipin_3.mux_l3_in_1_/X mux_top_ipin_3.mux_l3_in_0_/X
+ mux_top_ipin_3.mux_l4_in_0_/S mux_top_ipin_3.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_7.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_3_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1__A0 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_3.mux_l3_in_1__A1 mux_top_ipin_3.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0__S mux_top_ipin_5.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_8.mux_l2_in_3_ _19_/HI chanx_right_in[19] mux_top_ipin_8.mux_l2_in_1_/S
+ mux_top_ipin_8.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_3.mux_l3_in_1_ mux_top_ipin_3.mux_l2_in_3_/X mux_top_ipin_3.mux_l2_in_2_/X
+ mux_top_ipin_3.mux_l3_in_1_/S mux_top_ipin_3.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_4_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_0.mux_l2_in_2__S mux_top_ipin_0.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0__A0 mux_top_ipin_0.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l4_in_0__A1 mux_top_ipin_3.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_4.mux_l3_in_0__S mux_top_ipin_4.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_3.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[8] mux_top_ipin_3.mux_l2_in_2_/S
+ mux_top_ipin_3.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_8.mux_l4_in_0_ mux_top_ipin_8.mux_l3_in_1_/X mux_top_ipin_8.mux_l3_in_0_/X
+ mux_top_ipin_8.mux_l4_in_0_/S mux_top_ipin_8.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_10.mux_l2_in_3_ _24_/HI chanx_right_in[15] mux_top_ipin_10.mux_l2_in_3_/S
+ mux_top_ipin_10.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20_ _20_/HI _20_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_5.mux_l2_in_3__S mux_top_ipin_5.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_9.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l4_in_0__S mux_top_ipin_3.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_12.mux_l1_in_1__S mux_top_ipin_12.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_8.mux_l3_in_1_ mux_top_ipin_8.mux_l2_in_3_/X mux_top_ipin_8.mux_l2_in_2_/X
+ mux_top_ipin_8.mux_l3_in_0_/S mux_top_ipin_8.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_0_prog_clk prog_clk clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_10_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_9.mux_l3_in_1__S mux_top_ipin_9.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l2_in_0__A0 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_2.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_7.mux_l1_in_2__A0 chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_4_0_prog_clk_A clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_10.mux_l4_in_0_ mux_top_ipin_10.mux_l3_in_1_/X mux_top_ipin_10.mux_l3_in_0_/X
+ mux_top_ipin_10.mux_l4_in_0_/S mux_top_ipin_10.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_0.mux_l1_in_1__A1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__D mux_bottom_ipin_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_3.mux_l4_in_0_/X bottom_grid_pin_3_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_top_ipin_8.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[13] mux_top_ipin_8.mux_l2_in_1_/S
+ mux_top_ipin_8.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_12.mux_l2_in_2__A0 chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_11.mux_l2_in_1__S mux_top_ipin_11.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_3.mux_l3_in_0_ mux_top_ipin_3.mux_l2_in_1_/X mux_top_ipin_3.mux_l2_in_0_/X
+ mux_top_ipin_3.mux_l3_in_1_/S mux_top_ipin_3.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_7.mux_l2_in_1__A0 chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_15.mux_l2_in_3_ _29_/HI chanx_right_in[16] mux_top_ipin_15.mux_l2_in_3_/S
+ mux_top_ipin_15.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_0.mux_l2_in_0__A1 mux_top_ipin_0.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_10.mux_l3_in_1_ mux_top_ipin_10.mux_l2_in_3_/X mux_top_ipin_10.mux_l2_in_2_/X
+ mux_top_ipin_10.mux_l3_in_1_/S mux_top_ipin_10.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_12.mux_l3_in_1__A0 mux_top_ipin_12.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_5.mux_l2_in_3__A0 _33_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_3.mux_l2_in_1_ chanx_left_in[8] mux_top_ipin_3.mux_l1_in_2_/X mux_top_ipin_3.mux_l2_in_2_/S
+ mux_top_ipin_3.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_10.mux_l3_in_1__S mux_top_ipin_10.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_5_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_7.mux_l3_in_0__A0 mux_top_ipin_7.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_5.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_10.mux_l2_in_2_ chanx_left_in[15] chanx_right_in[7] mux_top_ipin_10.mux_l2_in_3_/S
+ mux_top_ipin_10.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_3_0_0_prog_clk clkbuf_2_0_0_prog_clk/X clkbuf_3_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_top_ipin_12.mux_l4_in_0__A0 mux_top_ipin_12.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_15.mux_l4_in_0_ mux_top_ipin_15.mux_l3_in_1_/X mux_top_ipin_15.mux_l3_in_0_/X
+ mux_top_ipin_15.mux_l4_in_0_/S mux_top_ipin_15.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_7_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_3.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_top_ipin_3.mux_l1_in_2_/S
+ mux_top_ipin_3.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_13.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_9.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_3.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_79_ ccff_tail gfpga_pad_EMBEDDED_IO_SOC_DIR VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_28_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_8.mux_l3_in_0_ mux_top_ipin_8.mux_l2_in_1_/X mux_top_ipin_8.mux_l2_in_0_/X
+ mux_top_ipin_8.mux_l3_in_0_/S mux_top_ipin_8.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_14.mux_l2_in_0__A1 mux_top_ipin_14.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_15.mux_l3_in_1_ mux_top_ipin_15.mux_l2_in_3_/X mux_top_ipin_15.mux_l2_in_2_/X
+ mux_top_ipin_15.mux_l3_in_1_/S mux_top_ipin_15.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_7.mux_l1_in_2__A1 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0__S mux_top_ipin_2.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_8.mux_l2_in_1_ chanx_left_in[13] mux_top_ipin_8.mux_l1_in_2_/X mux_top_ipin_8.mux_l2_in_1_/S
+ mux_top_ipin_8.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_12.mux_l2_in_2__A1 chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_7.mux_l2_in_1__A1 mux_top_ipin_7.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_15.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[10] mux_top_ipin_15.mux_l2_in_3_/S
+ mux_top_ipin_15.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_8.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0__S mux_top_ipin_1.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_10.mux_l3_in_0_ mux_top_ipin_10.mux_l2_in_1_/X mux_top_ipin_10.mux_l2_in_0_/X
+ mux_top_ipin_10.mux_l3_in_1_/S mux_top_ipin_10.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_12.mux_l3_in_1__A1 mux_top_ipin_12.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_8.mux_l1_in_2_ chanx_right_in[9] chanx_left_in[9] mux_top_ipin_8.mux_l1_in_0_/S
+ mux_top_ipin_8.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_7.mux_l1_in_1__S mux_top_ipin_7.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_14.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_4.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l2_in_3__A1 chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_10.mux_l4_in_0_/X bottom_grid_pin_10_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_top_ipin_3.mux_l2_in_0_ mux_top_ipin_3.mux_l1_in_1_/X mux_top_ipin_3.mux_l1_in_0_/X
+ mux_top_ipin_3.mux_l2_in_2_/S mux_top_ipin_3.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_7.mux_l3_in_0__A1 mux_top_ipin_7.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_4.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_10.mux_l2_in_1_ chanx_left_in[7] chanx_right_in[3] mux_top_ipin_10.mux_l2_in_3_/S
+ mux_top_ipin_10.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_1_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_12.mux_l4_in_0__A1 mux_top_ipin_12.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_0.mux_l3_in_0__S mux_top_ipin_0.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_3.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_3.mux_l1_in_2_/S
+ mux_top_ipin_3.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_6.mux_l2_in_1__S mux_top_ipin_6.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_78_ chanx_left_in[0] chanx_right_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1__S mux_bottom_ipin_0.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_6_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_9.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_15.mux_l3_in_0_ mux_top_ipin_15.mux_l2_in_1_/X mux_top_ipin_15.mux_l2_in_0_/X
+ mux_top_ipin_15.mux_l3_in_1_/S mux_top_ipin_15.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_2.mux_l2_in_1__A0 chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_1.mux_l2_in_3__S mux_top_ipin_1.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_8.mux_l2_in_0_ mux_top_ipin_8.mux_l1_in_1_/X mux_top_ipin_8.mux_l1_in_0_/X
+ mux_top_ipin_8.mux_l2_in_1_/S mux_top_ipin_8.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_5.mux_l3_in_1__S mux_top_ipin_5.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_2_3_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_0.mux_l2_in_3__A0 _22_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_15.mux_l2_in_1_ chanx_left_in[10] mux_top_ipin_15.mux_l1_in_2_/X mux_top_ipin_15.mux_l2_in_3_/S
+ mux_top_ipin_15.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_2.mux_l3_in_0__A0 mux_top_ipin_2.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_8.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_8.mux_l1_in_0_/S
+ mux_top_ipin_8.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_4.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_15.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_top_ipin_15.mux_l1_in_2_/S
+ mux_top_ipin_15.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_10.mux_l2_in_0_ chanx_left_in[3] mux_top_ipin_10.mux_l1_in_0_/X mux_top_ipin_10.mux_l2_in_3_/S
+ mux_top_ipin_10.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_3.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_3.mux_l1_in_2_/S
+ mux_top_ipin_3.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_14.mux_l2_in_3__A0 _28_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_77_ chanx_left_in[1] chanx_right_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_12.mux_l2_in_2__S mux_top_ipin_12.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_9.mux_l2_in_2__A0 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_2.mux_l2_in_1__A1 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_9.mux_l3_in_1__A0 mux_top_ipin_9.mux_l2_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_3__A1 chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_11.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_15.mux_l2_in_0_ mux_top_ipin_15.mux_l1_in_1_/X mux_top_ipin_15.mux_l1_in_0_/X
+ mux_top_ipin_15.mux_l2_in_3_/S mux_top_ipin_15.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_2.mux_l3_in_0__A1 mux_top_ipin_2.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_15.mux_l4_in_0__S mux_top_ipin_15.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_12.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_8.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_8.mux_l1_in_0_/S
+ mux_top_ipin_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_5_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_9.mux_l4_in_0__A0 mux_top_ipin_9.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_15.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_15.mux_l1_in_2_/S
+ mux_top_ipin_15.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_7_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_1__S mux_top_ipin_3.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_6.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_76_ chanx_left_in[2] chanx_right_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_14.mux_l2_in_3__A1 chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_13.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_10.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_10.mux_l1_in_0_/S
+ mux_top_ipin_10.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_9.mux_l2_in_2__A1 chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_59_ chanx_left_in[19] chanx_right_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_2.mux_l2_in_1__S mux_top_ipin_2.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_15.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_11.mux_l1_in_2__A0 chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l1_in_2__S mux_top_ipin_8.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_9.mux_l3_in_1__A1 mux_top_ipin_9.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_6.mux_l4_in_0_/X bottom_grid_pin_6_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_7_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_11.mux_l2_in_1__A0 chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_1.mux_l3_in_1__S mux_top_ipin_1.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_7.mux_l2_in_2__S mux_top_ipin_7.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0__A0 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_9.mux_l4_in_0__A1 mux_top_ipin_9.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ mux_top_ipin_15.mux_l4_in_0_/S ccff_tail clkbuf_3_7_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_22_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_14.mux_l1_in_0__S mux_top_ipin_14.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_15.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_15.mux_l1_in_2_/S
+ mux_top_ipin_15.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_11.mux_l3_in_0__A0 mux_top_ipin_11.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_4.mux_l2_in_2__A0 chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_75_ chanx_left_in[3] chanx_right_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_6_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_13.mux_l2_in_0__S mux_top_ipin_13.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_13.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__40__A chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_2__S mux_bottom_ipin_0.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_4.mux_l3_in_1__A0 mux_top_ipin_4.mux_l2_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_58_ chanx_right_in[0] chanx_left_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_21_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_11.mux_l1_in_2__A1 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_12.mux_l3_in_0__S mux_top_ipin_12.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_4.mux_l4_in_0__A0 mux_top_ipin_4.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_11.mux_l2_in_1__A1 mux_top_ipin_11.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_12.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_2.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0__A1 mux_top_ipin_6.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_13.mux_l2_in_3__S mux_top_ipin_13.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_11.mux_l4_in_0__S mux_top_ipin_11.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__43__A chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_13.mux_l4_in_0_/X bottom_grid_pin_13_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_ipin_11.mux_l3_in_0__A1 mux_top_ipin_11.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_4.mux_l2_in_2__A1 chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__38__A gfpga_pad_EMBEDDED_IO_SOC_IN VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_74_ chanx_left_in[4] chanx_right_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_4.mux_l2_in_3_ _32_/HI chanx_right_in[15] mux_top_ipin_4.mux_l2_in_0_/S
+ mux_top_ipin_4.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_4.mux_l3_in_1__A1 mux_top_ipin_4.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_ipin_0.mux_l2_in_3_ _21_/HI chanx_right_in[16] mux_bottom_ipin_0.mux_l2_in_3_/S
+ mux_bottom_ipin_0.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_57_ chanx_right_in[1] chanx_left_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_21_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__51__A chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_13.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_3.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_9.mux_l1_in_0__S mux_top_ipin_9.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_1.mux_l2_in_0__A0 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_4.mux_l4_in_0__A1 mux_top_ipin_4.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__46__A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_4.mux_l4_in_0_ mux_top_ipin_4.mux_l3_in_1_/X mux_top_ipin_4.mux_l3_in_0_/X
+ mux_top_ipin_4.mux_l4_in_0_/S mux_top_ipin_4.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_0.mux_l3_in_0_/S mux_top_ipin_0.mux_l4_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_19_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_5_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_4.mux_l1_in_2__S mux_top_ipin_4.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_0.mux_l4_in_0_ mux_bottom_ipin_0.mux_l3_in_1_/X mux_bottom_ipin_0.mux_l3_in_0_/X
+ mux_bottom_ipin_0.mux_l4_in_0_/S mux_bottom_ipin_0.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_9.mux_l2_in_3_ _20_/HI chanx_right_in[14] mux_top_ipin_9.mux_l2_in_0_/S
+ mux_top_ipin_9.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_8.mux_l2_in_0__S mux_top_ipin_8.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_10.mux_l3_in_1_/S mux_top_ipin_10.mux_l4_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_15.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_4.mux_l3_in_1_ mux_top_ipin_4.mux_l2_in_3_/X mux_top_ipin_4.mux_l2_in_2_/X
+ mux_top_ipin_4.mux_l3_in_0_/S mux_top_ipin_4.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_7_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_8.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_3.mux_l2_in_2__S mux_top_ipin_3.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_0.mux_l3_in_1_ mux_bottom_ipin_0.mux_l2_in_3_/X mux_bottom_ipin_0.mux_l2_in_2_/X
+ mux_bottom_ipin_0.mux_l3_in_1_/S mux_bottom_ipin_0.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_0_0_prog_clk_A clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_10.mux_l1_in_0__S mux_top_ipin_10.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__54__A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_15.mux_l2_in_0__A0 mux_top_ipin_15.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_73_ chanx_left_in[5] chanx_right_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_7.mux_l3_in_0__S mux_top_ipin_7.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_4.mux_l2_in_2_ chanx_left_in[15] chanx_right_in[9] mux_top_ipin_4.mux_l2_in_0_/S
+ mux_top_ipin_4.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_8.mux_l1_in_2__A0 chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_9.mux_l4_in_0_ mux_top_ipin_9.mux_l3_in_1_/X mux_top_ipin_9.mux_l3_in_0_/X
+ mux_top_ipin_9.mux_l4_in_0_/S mux_top_ipin_9.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__49__A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_3.mux_l3_in_1_/S mux_top_ipin_3.mux_l4_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_ipin_0.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[10] mux_bottom_ipin_0.mux_l2_in_3_/S
+ mux_bottom_ipin_0.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_56_ chanx_right_in[2] chanx_left_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_13.mux_l2_in_2__A0 chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_11.mux_l2_in_3_ _25_/HI chanx_right_in[16] mux_top_ipin_11.mux_l2_in_3_/S
+ mux_top_ipin_11.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_8.mux_l2_in_1__A0 chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l2_in_3__S mux_top_ipin_8.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l4_in_0__S mux_top_ipin_6.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_15.mux_l1_in_1__S mux_top_ipin_15.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_9.mux_l3_in_1_ mux_top_ipin_9.mux_l2_in_3_/X mux_top_ipin_9.mux_l2_in_2_/X
+ mux_top_ipin_9.mux_l3_in_1_/S mux_top_ipin_9.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_39_ chanx_right_in[19] chanx_left_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_13.mux_l3_in_1_/S mux_top_ipin_13.mux_l4_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_20_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_1.mux_l2_in_0__A1 mux_top_ipin_1.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_2_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l3_in_0__S mux_bottom_ipin_0.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_13.mux_l3_in_1__A0 mux_top_ipin_13.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_0.mux_l2_in_3_/S mux_top_ipin_0.mux_l3_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__62__A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_5_0_prog_clk_A clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_3__A0 _17_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_8.mux_l3_in_0__A0 mux_top_ipin_8.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__57__A chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_11.mux_l4_in_0_ mux_top_ipin_11.mux_l3_in_1_/X mux_top_ipin_11.mux_l3_in_0_/X
+ mux_top_ipin_11.mux_l4_in_0_/S mux_top_ipin_11.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_9.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[6] mux_top_ipin_9.mux_l2_in_0_/S
+ mux_top_ipin_9.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_10.mux_l2_in_3_/S mux_top_ipin_10.mux_l3_in_1_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_1_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_15.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l2_in_1__S mux_top_ipin_14.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_4.mux_l3_in_0_ mux_top_ipin_4.mux_l2_in_1_/X mux_top_ipin_4.mux_l2_in_0_/X
+ mux_top_ipin_4.mux_l3_in_0_/S mux_top_ipin_4.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_13.mux_l4_in_0__A0 mux_top_ipin_13.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_6.mux_l3_in_1_/S mux_top_ipin_6.mux_l4_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_ipin_0.mux_l3_in_0_ mux_bottom_ipin_0.mux_l2_in_1_/X mux_bottom_ipin_0.mux_l2_in_0_/X
+ mux_bottom_ipin_0.mux_l3_in_1_/S mux_bottom_ipin_0.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_11.mux_l3_in_1_ mux_top_ipin_11.mux_l2_in_3_/X mux_top_ipin_11.mux_l2_in_2_/X
+ mux_top_ipin_11.mux_l3_in_1_/S mux_top_ipin_11.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA__70__A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_15.mux_l2_in_0__A1 mux_top_ipin_15.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_72_ chanx_left_in[6] chanx_right_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_4.mux_l2_in_1_ chanx_left_in[9] mux_top_ipin_4.mux_l1_in_2_/X mux_top_ipin_4.mux_l2_in_0_/S
+ mux_top_ipin_4.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_13.mux_l3_in_1__S mux_top_ipin_13.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l1_in_2__A1 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_10.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__65__A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_3.mux_l2_in_2_/S mux_top_ipin_3.mux_l3_in_1_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_ipin_0.mux_l2_in_1_ chanx_left_in[10] mux_bottom_ipin_0.mux_l1_in_2_/X
+ mux_bottom_ipin_0.mux_l2_in_3_/S mux_bottom_ipin_0.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_13.mux_l2_in_2__A1 chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_55_ chanx_right_in[3] chanx_left_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_11.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[12] mux_top_ipin_11.mux_l2_in_3_/S
+ mux_top_ipin_11.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A0 mux_bottom_ipin_0.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_4.mux_l1_in_2_ chanx_right_in[5] chanx_left_in[5] mux_top_ipin_4.mux_l1_in_2_/S
+ mux_top_ipin_4.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_8.mux_l2_in_1__A1 mux_top_ipin_8.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_9.mux_l3_in_0_ mux_top_ipin_9.mux_l2_in_1_/X mux_top_ipin_9.mux_l2_in_0_/X
+ mux_top_ipin_9.mux_l3_in_1_/S mux_top_ipin_9.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_13.mux_l2_in_3_/S mux_top_ipin_13.mux_l3_in_1_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_38_ gfpga_pad_EMBEDDED_IO_SOC_IN bottom_width_0_height_0__pin_1_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_13.mux_l3_in_1__A1 mux_top_ipin_13.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_0.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_bottom_ipin_0.mux_l1_in_1_/S
+ mux_bottom_ipin_0.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_0.mux_l1_in_2_/S mux_top_ipin_0.mux_l2_in_3_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_34_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A0 mux_bottom_ipin_0.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_5.mux_l1_in_0__S mux_top_ipin_5.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_3__A1 chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_15.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_9.mux_l4_in_0_/X bottom_grid_pin_9_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_9.mux_l3_in_1_/S mux_top_ipin_9.mux_l4_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_5.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_8.mux_l3_in_0__A1 mux_top_ipin_8.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__73__A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_9.mux_l2_in_1_ chanx_left_in[6] chanx_right_in[2] mux_top_ipin_9.mux_l2_in_0_/S
+ mux_top_ipin_9.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_10.mux_l1_in_0_/S mux_top_ipin_10.mux_l2_in_3_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_22_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_10.mux_l2_in_0__A0 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_13.mux_l4_in_0__A1 mux_top_ipin_13.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_2__S mux_top_ipin_0.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__68__A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_2__A0 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_6.mux_l2_in_0_/S mux_top_ipin_6.mux_l3_in_1_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_4.mux_l2_in_0__S mux_top_ipin_4.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_11.mux_l3_in_0_ mux_top_ipin_11.mux_l2_in_1_/X mux_top_ipin_11.mux_l2_in_0_/X
+ mux_top_ipin_11.mux_l3_in_1_/S mux_top_ipin_11.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1 chanx_right_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_30_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_71_ chanx_left_in[7] chanx_right_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_4.mux_l2_in_0_ mux_top_ipin_4.mux_l1_in_1_/X mux_top_ipin_4.mux_l1_in_0_/X
+ mux_top_ipin_4.mux_l2_in_0_/S mux_top_ipin_4.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_3.mux_l2_in_1__A0 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_3.mux_l1_in_2_/S mux_top_ipin_3.mux_l2_in_2_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_ipin_0.mux_l2_in_0_ mux_bottom_ipin_0.mux_l1_in_1_/X mux_bottom_ipin_0.mux_l1_in_0_/X
+ mux_bottom_ipin_0.mux_l2_in_3_/S mux_bottom_ipin_0.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
X_54_ chanx_right_in[4] chanx_left_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_11.mux_l2_in_1_ chanx_left_in[12] mux_top_ipin_11.mux_l1_in_2_/X mux_top_ipin_11.mux_l2_in_3_/S
+ mux_top_ipin_11.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_6_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l3_in_0__S mux_top_ipin_3.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A1 mux_bottom_ipin_0.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_1.mux_l2_in_3__A0 _23_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_4.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_4.mux_l1_in_2_/S
+ mux_top_ipin_4.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__76__A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_9.mux_l2_in_1__S mux_top_ipin_9.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l3_in_0__A0 mux_top_ipin_3.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_13.mux_l1_in_0_/S mux_top_ipin_13.mux_l2_in_3_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_37_ gfpga_pad_EMBEDDED_IO_SOC_IN bottom_width_0_height_0__pin_1_lower VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_ipin_0.mux_l4_in_0_/S mux_top_ipin_0.mux_l1_in_2_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_ipin_0.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_bottom_ipin_0.mux_l1_in_1_/S
+ mux_bottom_ipin_0.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_11.mux_l1_in_2_ chanx_right_in[6] chanx_left_in[6] mux_top_ipin_11.mux_l1_in_2_/S
+ mux_top_ipin_11.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A1 mux_bottom_ipin_0.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_9.mux_l2_in_0_/S mux_top_ipin_9.mux_l3_in_1_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_4.mux_l2_in_3__S mux_top_ipin_4.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_2.mux_l4_in_0__S mux_top_ipin_2.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_11.mux_l1_in_1__S mux_top_ipin_11.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_9.mux_l2_in_0_ chanx_left_in[2] mux_top_ipin_9.mux_l1_in_0_/X mux_top_ipin_9.mux_l2_in_0_/S
+ mux_top_ipin_9.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_9.mux_l4_in_0_/S mux_top_ipin_10.mux_l1_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_8.mux_l3_in_1__S mux_top_ipin_8.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_10.mux_l2_in_0__A1 mux_top_ipin_10.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_3.mux_l1_in_2__A1 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_15.mux_l2_in_3__A0 _29_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_6.mux_l1_in_0_/S mux_top_ipin_6.mux_l2_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_10.mux_l2_in_1__S mux_top_ipin_10.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__79__A ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_70_ chanx_left_in[8] chanx_right_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_3.mux_l2_in_1__A1 mux_top_ipin_3.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_1_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_2.mux_l4_in_0_/S mux_top_ipin_3.mux_l1_in_2_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_53_ chanx_right_in[5] chanx_left_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_11.mux_l2_in_0_ mux_top_ipin_11.mux_l1_in_1_/X mux_top_ipin_11.mux_l1_in_0_/X
+ mux_top_ipin_11.mux_l2_in_3_/S mux_top_ipin_11.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_1.mux_l2_in_3__A1 chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_4.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_4.mux_l1_in_2_/S
+ mux_top_ipin_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_1.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_11.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_3_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l3_in_0__A1 mux_top_ipin_3.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_36_ _36_/A SC_OUT_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_15.mux_l2_in_2__S mux_top_ipin_15.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_12.mux_l4_in_0_/S mux_top_ipin_13.mux_l1_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_20_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_0.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_bottom_ipin_0.mux_l1_in_1_/S
+ mux_bottom_ipin_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_11.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_11.mux_l1_in_2_/S
+ mux_top_ipin_11.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_9.mux_l1_in_0_/S mux_top_ipin_9.mux_l2_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_19_ _19_/HI _19_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_4_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_1.mux_l1_in_0__S mux_top_ipin_1.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_15.mux_l2_in_3__A1 chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_5.mux_l4_in_0_/S mux_top_ipin_6.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_14.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_2.mux_l4_in_0_/X bottom_grid_pin_2_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_top_ipin_9.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_9.mux_l1_in_0_/S
+ mux_top_ipin_9.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_12.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_2.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_0.mux_l2_in_0__S mux_top_ipin_0.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_12.mux_l1_in_2__A0 chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_52_ chanx_right_in[6] chanx_left_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_7.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0__A mux_bottom_ipin_0.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35_ _35_/A SC_OUT_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_12.mux_l2_in_1__A0 chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_7.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_11.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_11.mux_l1_in_2_/S
+ mux_top_ipin_11.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_7.mux_l2_in_0__A0 mux_top_ipin_7.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18_ _18_/HI _18_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_ipin_5.mux_l2_in_1__S mux_top_ipin_5.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_8.mux_l4_in_0_/S mux_top_ipin_9.mux_l1_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_10.mux_l2_in_3__A0 _24_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_12.mux_l3_in_0__A0 mux_top_ipin_12.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_5.mux_l2_in_2__A0 chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_0.mux_l2_in_3__S mux_top_ipin_0.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_4_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_1.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_4.mux_l3_in_1__S mux_top_ipin_4.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_5.mux_l3_in_1__A0 mux_top_ipin_5.mux_l2_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_6_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_12.mux_l1_in_2__A1 chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_51_ chanx_right_in[7] chanx_left_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_12.mux_l1_in_2__S mux_top_ipin_12.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l4_in_0__A0 mux_top_ipin_5.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34_ SC_IN_BOT SC_IN_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_9_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_12.mux_l2_in_1__A1 mux_top_ipin_12.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0__A1 mux_top_ipin_7.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_2_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__D mux_bottom_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17_ _17_/HI _17_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_4.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_10.mux_l2_in_3__A1 chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_11.mux_l2_in_2__S mux_top_ipin_11.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_12.mux_l3_in_0__A1 mux_top_ipin_12.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_15.mux_l3_in_0__S mux_top_ipin_15.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l2_in_3_ _22_/HI chanx_right_in[17] mux_top_ipin_0.mux_l2_in_3_/S
+ mux_top_ipin_0.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_5.mux_l2_in_2__A1 chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_1_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_5.mux_l3_in_1__A1 mux_top_ipin_5.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l4_in_0__S mux_top_ipin_14.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_0.mux_l4_in_0_ mux_top_ipin_0.mux_l3_in_1_/X mux_top_ipin_0.mux_l3_in_0_/X
+ mux_top_ipin_0.mux_l4_in_0_/S mux_top_ipin_0.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_50_ chanx_right_in[8] chanx_left_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_3_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_2.mux_l2_in_0__A0 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l4_in_0__A1 mux_top_ipin_5.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_7.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_5.mux_l2_in_3_ _33_/HI chanx_right_in[18] mux_top_ipin_5.mux_l2_in_2_/S
+ mux_top_ipin_5.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_33_ _33_/HI _33_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_0.mux_l3_in_1_ mux_top_ipin_0.mux_l2_in_3_/X mux_top_ipin_0.mux_l2_in_2_/X
+ mux_top_ipin_0.mux_l3_in_0_/S mux_top_ipin_0.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_0.mux_l2_in_2__A0 chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_8.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[11] mux_top_ipin_0.mux_l2_in_3_/S
+ mux_top_ipin_0.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_0.mux_l3_in_1__A0 mux_top_ipin_0.mux_l2_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_5.mux_l4_in_0_ mux_top_ipin_5.mux_l3_in_1_/X mux_top_ipin_5.mux_l3_in_0_/X
+ mux_top_ipin_5.mux_l4_in_0_/S mux_top_ipin_5.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_1.mux_l2_in_1__S mux_top_ipin_1.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_7.mux_l1_in_2__S mux_top_ipin_7.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_7_0_prog_clk clkbuf_3_7_0_prog_clk/A clkbuf_3_7_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_29_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_0.mux_l4_in_0__A0 mux_top_ipin_0.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l2_in_2__A0 chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_5.mux_l3_in_1_ mux_top_ipin_5.mux_l2_in_3_/X mux_top_ipin_5.mux_l2_in_2_/X
+ mux_top_ipin_5.mux_l3_in_1_/S mux_top_ipin_5.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_0.mux_l3_in_1__S mux_top_ipin_0.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_9.mux_l2_in_1__A0 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_6.mux_l2_in_2__S mux_top_ipin_6.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_prog_clk_A clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_13.mux_l1_in_0__S mux_top_ipin_13.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0__A1 mux_top_ipin_2.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_14.mux_l3_in_1__A0 mux_top_ipin_14.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_2__S mux_bottom_ipin_0.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_5.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[10] mux_top_ipin_5.mux_l2_in_2_/S
+ mux_top_ipin_5.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32_ _32_/HI _32_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_9.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_7.mux_l2_in_3__A0 _18_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l3_in_0_ mux_top_ipin_0.mux_l2_in_1_/X mux_top_ipin_0.mux_l2_in_0_/X
+ mux_top_ipin_0.mux_l3_in_0_/S mux_top_ipin_0.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_9.mux_l3_in_0__A0 mux_top_ipin_9.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_2__A1 chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_12.mux_l2_in_3_ _26_/HI chanx_right_in[17] mux_top_ipin_12.mux_l2_in_2_/S
+ mux_top_ipin_12.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_12.mux_l2_in_0__S mux_top_ipin_12.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l4_in_0__A0 mux_top_ipin_14.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_9.mux_l4_in_0__S mux_top_ipin_9.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l2_in_1_ chanx_left_in[11] mux_top_ipin_0.mux_l1_in_2_/X mux_top_ipin_0.mux_l2_in_3_/S
+ mux_top_ipin_0.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_0.mux_l3_in_1__A1 mux_top_ipin_0.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_5_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_6_0_prog_clk_A clkbuf_3_7_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_11.mux_l3_in_0__S mux_top_ipin_11.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_12.mux_l4_in_0_ mux_top_ipin_12.mux_l3_in_1_/X mux_top_ipin_12.mux_l3_in_0_/X
+ mux_top_ipin_12.mux_l4_in_0_/S mux_top_ipin_12.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_10.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_7_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l1_in_2_ chanx_right_in[5] chanx_left_in[5] mux_top_ipin_0.mux_l1_in_2_/S
+ mux_top_ipin_0.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_0.mux_l4_in_0__A1 mux_top_ipin_0.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l2_in_2__A1 chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_5.mux_l3_in_0_ mux_top_ipin_5.mux_l2_in_1_/X mux_top_ipin_5.mux_l2_in_0_/X
+ mux_top_ipin_5.mux_l3_in_1_/S mux_top_ipin_5.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_5.mux_l4_in_0_/X bottom_grid_pin_5_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_6_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_9.mux_l2_in_1__A1 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_12.mux_l3_in_1_ mux_top_ipin_12.mux_l2_in_3_/X mux_top_ipin_12.mux_l2_in_2_/X
+ mux_top_ipin_12.mux_l3_in_1_/S mux_top_ipin_12.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_12.mux_l2_in_3__S mux_top_ipin_12.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_10.mux_l4_in_0__S mux_top_ipin_10.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_11.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_11.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l3_in_1__A1 mux_top_ipin_14.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_5.mux_l2_in_1_ chanx_left_in[10] chanx_right_in[2] mux_top_ipin_5.mux_l2_in_2_/S
+ mux_top_ipin_5.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_31_ _31_/HI _31_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_ipin_7.mux_l2_in_3__A1 chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_9.mux_l3_in_0__A1 mux_top_ipin_9.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_12.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[13] mux_top_ipin_12.mux_l2_in_2_/S
+ mux_top_ipin_12.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_11.mux_l2_in_0__A0 mux_top_ipin_11.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l4_in_0__A1 mux_top_ipin_14.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_1.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_11.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_4.mux_l1_in_2__A0 chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_0.mux_l2_in_0_ mux_top_ipin_0.mux_l1_in_1_/X mux_top_ipin_0.mux_l1_in_0_/X
+ mux_top_ipin_0.mux_l2_in_3_/S mux_top_ipin_0.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_8.mux_l1_in_0__S mux_top_ipin_8.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_3_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_4.mux_l2_in_1__A0 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_14.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_0.mux_l1_in_2_/S
+ mux_top_ipin_0.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_35_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_3.mux_l1_in_2__S mux_top_ipin_3.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_6.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_2.mux_l2_in_3__A0 _30_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_4.mux_l3_in_0__A0 mux_top_ipin_4.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0__S mux_top_ipin_7.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_12.mux_l3_in_0_ mux_top_ipin_12.mux_l2_in_1_/X mux_top_ipin_12.mux_l2_in_0_/X
+ mux_top_ipin_12.mux_l3_in_1_/S mux_top_ipin_12.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_11.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_5.mux_l2_in_0_ chanx_left_in[2] mux_top_ipin_5.mux_l1_in_0_/X mux_top_ipin_5.mux_l2_in_2_/S
+ mux_top_ipin_5.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_30_ _30_/HI _30_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_13_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_12.mux_l4_in_0_/X bottom_grid_pin_12_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_ipin_2.mux_l2_in_2__S mux_top_ipin_2.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_12.mux_l2_in_1_ chanx_left_in[13] mux_top_ipin_12.mux_l1_in_2_/X mux_top_ipin_12.mux_l2_in_2_/S
+ mux_top_ipin_12.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_6.mux_l3_in_0__S mux_top_ipin_6.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_11.mux_l2_in_0__A1 mux_top_ipin_11.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_4.mux_l1_in_2__A1 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0__S mux_bottom_ipin_0.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_12.mux_l1_in_2_ chanx_right_in[7] chanx_left_in[7] mux_top_ipin_12.mux_l1_in_2_/S
+ mux_top_ipin_12.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_7.mux_l2_in_3__S mux_top_ipin_7.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_5.mux_l4_in_0__S mux_top_ipin_5.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_4.mux_l2_in_1__A1 mux_top_ipin_4.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_0.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_0.mux_l1_in_2_/S
+ mux_top_ipin_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_35_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_2.mux_l2_in_3__A1 chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_4.mux_l3_in_0__A1 mux_top_ipin_4.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_6_0_prog_clk clkbuf_3_7_0_prog_clk/A clkbuf_3_6_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_23_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_13.mux_l2_in_1__S mux_top_ipin_13.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__41__A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_3__S mux_bottom_ipin_0.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_5_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_12.mux_l2_in_0_ mux_top_ipin_12.mux_l1_in_1_/X mux_top_ipin_12.mux_l1_in_0_/X
+ mux_top_ipin_12.mux_l2_in_2_/S mux_top_ipin_12.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_12.mux_l3_in_1__S mux_top_ipin_12.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_5.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_5.mux_l1_in_0_/S
+ mux_top_ipin_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_15.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_12.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_12.mux_l1_in_2_/S
+ mux_top_ipin_12.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_13.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_7_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__44__A chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_4.mux_l1_in_0__S mux_top_ipin_4.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l1_in_1__A0 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__39__A chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_13.mux_l2_in_1__A0 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_7.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_8.mux_l2_in_0__A0 mux_top_ipin_8.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_3.mux_l2_in_0__S mux_top_ipin_3.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_11.mux_l2_in_3__A0 _25_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__52__A chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_13.mux_l3_in_0__A0 mux_top_ipin_13.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_2_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_2__A0 chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__47__A chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_15.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_2.mux_l3_in_0__S mux_top_ipin_2.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_12.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_12.mux_l1_in_2_/S
+ mux_top_ipin_12.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_1_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_6.mux_l3_in_1__A0 mux_top_ipin_6.mux_l2_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_8.mux_l2_in_1__S mux_top_ipin_8.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_2.mux_l3_in_1_/S mux_top_ipin_2.mux_l4_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_14_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__60__A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_8.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_3.mux_l2_in_3__S mux_top_ipin_3.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l1_in_1__A1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_1.mux_l4_in_0__S mux_top_ipin_1.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_6.mux_l4_in_0__A0 mux_top_ipin_6.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_12.mux_l3_in_1_/S mux_top_ipin_12.mux_l4_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__55__A chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_8.mux_l4_in_0_/X bottom_grid_pin_8_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_15_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_7.mux_l3_in_1__S mux_top_ipin_7.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_13.mux_l2_in_1__A1 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A0 mux_bottom_ipin_0.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_8.mux_l2_in_0__A1 mux_top_ipin_8.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_11.mux_l2_in_3__A1 chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_10.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_13.mux_l3_in_0__A1 mux_top_ipin_13.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_6.mux_l2_in_2__A1 chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_15.mux_l1_in_2__S mux_top_ipin_15.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D mux_bottom_ipin_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_5.mux_l3_in_1_/S mux_top_ipin_5.mux_l4_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_9.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l3_in_1__S mux_bottom_ipin_0.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__63__A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_3_0_prog_clk clkbuf_0_prog_clk/X clkbuf_3_7_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_3.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__58__A chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_15.mux_l3_in_1_/S mux_top_ipin_15.mux_l4_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_6.mux_l3_in_1__A1 mux_top_ipin_6.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_2.mux_l2_in_2_/S mux_top_ipin_2.mux_l3_in_1_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_14.mux_l2_in_2__S mux_top_ipin_14.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A1 mux_bottom_ipin_0.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_1.mux_l2_in_3_ _23_/HI chanx_right_in[14] mux_top_ipin_1.mux_l2_in_0_/S
+ mux_top_ipin_1.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_3.mux_l2_in_0__A0 mux_top_ipin_3.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l4_in_0__A1 mux_top_ipin_6.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_12.mux_l2_in_2_/S mux_top_ipin_12.mux_l3_in_1_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__71__A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A1 mux_bottom_ipin_0.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_10.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_0.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0__S mux_top_ipin_0.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_7_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_1.mux_l2_in_2__A0 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_8.mux_l3_in_0_/S mux_top_ipin_8.mux_l4_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA__66__A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_1.mux_l4_in_0_ mux_top_ipin_1.mux_l3_in_1_/X mux_top_ipin_1.mux_l3_in_0_/X
+ mux_top_ipin_1.mux_l4_in_0_/S mux_top_ipin_1.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_10.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_5_0_prog_clk clkbuf_2_2_0_prog_clk/X clkbuf_3_5_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_33_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_15.mux_l4_in_0_/X bottom_grid_pin_15_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_18_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_7_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_1.mux_l3_in_1__A0 mux_top_ipin_1.mux_l2_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_69_ chanx_left_in[9] chanx_right_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_5.mux_l2_in_2_/S mux_top_ipin_5.mux_l3_in_1_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_15_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_6.mux_l2_in_3_ _17_/HI chanx_right_in[19] mux_top_ipin_6.mux_l2_in_0_/S
+ mux_top_ipin_6.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_1.mux_l3_in_1_ mux_top_ipin_1.mux_l2_in_3_/X mux_top_ipin_1.mux_l2_in_2_/X
+ mux_top_ipin_1.mux_l3_in_1_/S mux_top_ipin_1.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_15.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_5.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_15.mux_l2_in_3_/S mux_top_ipin_15.mux_l3_in_1_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA__74__A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_1.mux_l4_in_0__A0 mux_top_ipin_1.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_15.mux_l2_in_2__A0 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_2.mux_l1_in_0_/S mux_top_ipin_2.mux_l2_in_2_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_1_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__69__A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_1.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[6] mux_top_ipin_1.mux_l2_in_0_/S
+ mux_top_ipin_1.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_4.mux_l2_in_1__S mux_top_ipin_4.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_6.mux_l4_in_0_ mux_top_ipin_6.mux_l3_in_1_/X mux_top_ipin_6.mux_l3_in_0_/X
+ mux_top_ipin_6.mux_l4_in_0_/S mux_top_ipin_6.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_3.mux_l2_in_0__A1 mux_top_ipin_3.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_12.mux_l1_in_2_/S mux_top_ipin_12.mux_l2_in_2_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_15.mux_l3_in_1__A0 mux_top_ipin_15.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
+ mux_top_ipin_15.mux_l4_in_0_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l2_in_3__A0 _19_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_1.mux_l2_in_2__A1 chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_8.mux_l2_in_1_/S mux_top_ipin_8.mux_l3_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_6.mux_l3_in_1_ mux_top_ipin_6.mux_l2_in_3_/X mux_top_ipin_6.mux_l2_in_2_/X
+ mux_top_ipin_6.mux_l3_in_1_/S mux_top_ipin_6.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_15.mux_l4_in_0__A0 mux_top_ipin_15.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_2_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l3_in_1__S mux_top_ipin_3.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__77__A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_prog_clk_A clkbuf_3_3_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_1.mux_l4_in_0_/X bottom_grid_pin_1_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_ipin_9.mux_l2_in_2__S mux_top_ipin_9.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_68_ chanx_left_in[10] chanx_right_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_1.mux_l3_in_1__A1 mux_top_ipin_1.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_5.mux_l1_in_0_/S mux_top_ipin_5.mux_l2_in_2_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_3_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_6.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[11] mux_top_ipin_6.mux_l2_in_0_/S
+ mux_top_ipin_6.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_4_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_1.mux_l3_in_0_ mux_top_ipin_1.mux_l2_in_1_/X mux_top_ipin_1.mux_l2_in_0_/X
+ mux_top_ipin_1.mux_l3_in_1_/S mux_top_ipin_1.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_11.mux_l1_in_2__S mux_top_ipin_11.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_13.mux_l2_in_3_ _27_/HI chanx_right_in[18] mux_top_ipin_13.mux_l2_in_3_/S
+ mux_top_ipin_13.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_15.mux_l1_in_2_/S mux_top_ipin_15.mux_l2_in_3_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_1.mux_l4_in_0__A1 mux_top_ipin_1.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_15.mux_l2_in_2__A1 chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_15.mux_l2_in_0__S mux_top_ipin_15.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_1.mux_l4_in_0_/S mux_top_ipin_2.mux_l1_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_4_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_1.mux_l2_in_1_ chanx_left_in[6] chanx_right_in[2] mux_top_ipin_1.mux_l2_in_0_/S
+ mux_top_ipin_1.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_11.mux_l4_in_0_/S mux_top_ipin_12.mux_l1_in_2_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_10.mux_l2_in_2__S mux_top_ipin_10.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_12.mux_l1_in_1__A0 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_15.mux_l3_in_1__A1 mux_top_ipin_15.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_7_0_prog_clk_A clkbuf_3_7_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_8.mux_l2_in_3__A1 chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_13.mux_l4_in_0_ mux_top_ipin_13.mux_l3_in_1_/X mux_top_ipin_13.mux_l3_in_0_/X
+ mux_top_ipin_13.mux_l4_in_0_/S mux_top_ipin_13.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_14.mux_l3_in_0__S mux_top_ipin_14.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_8.mux_l1_in_0_/S mux_top_ipin_8.mux_l2_in_1_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_13_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_6.mux_l3_in_0_ mux_top_ipin_6.mux_l2_in_1_/X mux_top_ipin_6.mux_l2_in_0_/X
+ mux_top_ipin_6.mux_l3_in_1_/S mux_top_ipin_6.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_15.mux_l4_in_0__A1 mux_top_ipin_15.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_12.mux_l2_in_0__A0 mux_top_ipin_12.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_12.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_13.mux_l3_in_1_ mux_top_ipin_13.mux_l2_in_3_/X mux_top_ipin_13.mux_l2_in_2_/X
+ mux_top_ipin_13.mux_l3_in_1_/S mux_top_ipin_13.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_15.mux_l2_in_3__S mux_top_ipin_15.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_67_ chanx_left_in[11] chanx_right_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_13.mux_l4_in_0__S mux_top_ipin_13.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_4.mux_l4_in_0_/S mux_top_ipin_5.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_10.mux_l2_in_2__A0 chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_6.mux_l2_in_1_ chanx_left_in[11] chanx_right_in[3] mux_top_ipin_6.mux_l2_in_0_/S
+ mux_top_ipin_6.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_5.mux_l2_in_1__A0 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_13.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[10] mux_top_ipin_13.mux_l2_in_3_/S
+ mux_top_ipin_13.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_14.mux_l4_in_0_/S mux_top_ipin_15.mux_l1_in_2_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_10.mux_l3_in_1__A0 mux_top_ipin_10.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_4_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l2_in_3__A0 _31_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_6.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_2_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_1.mux_l2_in_0_ chanx_left_in[2] mux_top_ipin_1.mux_l1_in_0_/X mux_top_ipin_1.mux_l2_in_0_/S
+ mux_top_ipin_1.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_5.mux_l3_in_0__A0 mux_top_ipin_5.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_12.mux_l1_in_1__A1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_6_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_10.mux_l4_in_0__A0 mux_top_ipin_10.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

