magic
tech sky130A
magscale 1 2
timestamp 1605111277
<< locali >>
rect 7021 23103 7055 23273
rect 10241 13855 10275 14025
<< viali >>
rect 4261 25449 4295 25483
rect 1409 25313 1443 25347
rect 2513 25313 2547 25347
rect 4077 25313 4111 25347
rect 5181 25313 5215 25347
rect 6929 25313 6963 25347
rect 8033 25245 8067 25279
rect 9781 25245 9815 25279
rect 1593 25177 1627 25211
rect 5365 25177 5399 25211
rect 7113 25177 7147 25211
rect 2053 25109 2087 25143
rect 2421 25109 2455 25143
rect 2697 25109 2731 25143
rect 4721 25109 4755 25143
rect 10425 25109 10459 25143
rect 2697 24905 2731 24939
rect 4077 24905 4111 24939
rect 4629 24837 4663 24871
rect 10333 24837 10367 24871
rect 12449 24837 12483 24871
rect 1869 24769 1903 24803
rect 2329 24769 2363 24803
rect 5089 24769 5123 24803
rect 5181 24769 5215 24803
rect 5733 24769 5767 24803
rect 6561 24769 6595 24803
rect 7481 24769 7515 24803
rect 10793 24769 10827 24803
rect 10977 24769 11011 24803
rect 12265 24769 12299 24803
rect 12909 24769 12943 24803
rect 13093 24769 13127 24803
rect 1593 24701 1627 24735
rect 2881 24701 2915 24735
rect 3433 24701 3467 24735
rect 4537 24701 4571 24735
rect 4997 24701 5031 24735
rect 8309 24701 8343 24735
rect 11897 24701 11931 24735
rect 15209 24701 15243 24735
rect 7297 24633 7331 24667
rect 8493 24633 8527 24667
rect 10701 24633 10735 24667
rect 3065 24565 3099 24599
rect 6285 24565 6319 24599
rect 6929 24565 6963 24599
rect 7389 24565 7423 24599
rect 8033 24565 8067 24599
rect 10149 24565 10183 24599
rect 12817 24565 12851 24599
rect 15393 24565 15427 24599
rect 15761 24565 15795 24599
rect 4261 24361 4295 24395
rect 5549 24361 5583 24395
rect 6009 24361 6043 24395
rect 7021 24361 7055 24395
rect 8493 24361 8527 24395
rect 15485 24361 15519 24395
rect 16589 24361 16623 24395
rect 17693 24361 17727 24395
rect 19073 24361 19107 24395
rect 21097 24361 21131 24395
rect 1869 24293 1903 24327
rect 5089 24293 5123 24327
rect 10425 24293 10459 24327
rect 10876 24293 10910 24327
rect 1593 24225 1627 24259
rect 2881 24225 2915 24259
rect 4077 24225 4111 24259
rect 4721 24225 4755 24259
rect 5917 24225 5951 24259
rect 6653 24225 6687 24259
rect 7113 24225 7147 24259
rect 7380 24225 7414 24259
rect 10609 24225 10643 24259
rect 15301 24225 15335 24259
rect 16405 24225 16439 24259
rect 17509 24225 17543 24259
rect 18889 24225 18923 24259
rect 20913 24225 20947 24259
rect 6193 24157 6227 24191
rect 13277 24157 13311 24191
rect 2697 24021 2731 24055
rect 3065 24021 3099 24055
rect 3525 24021 3559 24055
rect 11989 24021 12023 24055
rect 12541 24021 12575 24055
rect 14933 24021 14967 24055
rect 2605 23817 2639 23851
rect 3617 23817 3651 23851
rect 6193 23817 6227 23851
rect 6561 23817 6595 23851
rect 9229 23817 9263 23851
rect 13829 23817 13863 23851
rect 18245 23817 18279 23851
rect 19349 23817 19383 23851
rect 20453 23817 20487 23851
rect 21557 23817 21591 23851
rect 22661 23817 22695 23851
rect 10701 23749 10735 23783
rect 3249 23681 3283 23715
rect 4169 23681 4203 23715
rect 7849 23681 7883 23715
rect 11253 23681 11287 23715
rect 11437 23681 11471 23715
rect 14933 23681 14967 23715
rect 1409 23613 1443 23647
rect 4261 23613 4295 23647
rect 4528 23613 4562 23647
rect 9965 23613 9999 23647
rect 12449 23613 12483 23647
rect 14749 23613 14783 23647
rect 18061 23613 18095 23647
rect 18613 23613 18647 23647
rect 19165 23613 19199 23647
rect 19717 23613 19751 23647
rect 20269 23613 20303 23647
rect 20821 23613 20855 23647
rect 21373 23613 21407 23647
rect 21925 23613 21959 23647
rect 22477 23613 22511 23647
rect 23029 23613 23063 23647
rect 2053 23545 2087 23579
rect 3065 23545 3099 23579
rect 7757 23545 7791 23579
rect 8094 23545 8128 23579
rect 11161 23545 11195 23579
rect 11897 23545 11931 23579
rect 12265 23545 12299 23579
rect 12716 23545 12750 23579
rect 15178 23545 15212 23579
rect 18981 23545 19015 23579
rect 1593 23477 1627 23511
rect 2513 23477 2547 23511
rect 2973 23477 3007 23511
rect 5641 23477 5675 23511
rect 6837 23477 6871 23511
rect 7389 23477 7423 23511
rect 10241 23477 10275 23511
rect 10793 23477 10827 23511
rect 14381 23477 14415 23511
rect 16313 23477 16347 23511
rect 16865 23477 16899 23511
rect 17509 23477 17543 23511
rect 21189 23477 21223 23511
rect 4261 23273 4295 23307
rect 5825 23273 5859 23307
rect 6469 23273 6503 23307
rect 7021 23273 7055 23307
rect 8493 23273 8527 23307
rect 9781 23273 9815 23307
rect 10701 23273 10735 23307
rect 13645 23273 13679 23307
rect 16773 23273 16807 23307
rect 19625 23273 19659 23307
rect 1869 23205 1903 23239
rect 4712 23205 4746 23239
rect 1593 23137 1627 23171
rect 2881 23137 2915 23171
rect 3893 23137 3927 23171
rect 4445 23137 4479 23171
rect 11060 23205 11094 23239
rect 15577 23205 15611 23239
rect 21189 23205 21223 23239
rect 7369 23137 7403 23171
rect 12817 23137 12851 23171
rect 15301 23137 15335 23171
rect 16589 23137 16623 23171
rect 17693 23137 17727 23171
rect 19441 23137 19475 23171
rect 20913 23137 20947 23171
rect 7021 23069 7055 23103
rect 7113 23069 7147 23103
rect 9505 23069 9539 23103
rect 10333 23069 10367 23103
rect 10793 23069 10827 23103
rect 13737 23069 13771 23103
rect 13829 23069 13863 23103
rect 2697 23001 2731 23035
rect 17877 23001 17911 23035
rect 3065 22933 3099 22967
rect 3525 22933 3559 22967
rect 6929 22933 6963 22967
rect 12173 22933 12207 22967
rect 13277 22933 13311 22967
rect 14289 22933 14323 22967
rect 14657 22933 14691 22967
rect 4997 22729 5031 22763
rect 5641 22729 5675 22763
rect 6285 22729 6319 22763
rect 6653 22729 6687 22763
rect 8401 22729 8435 22763
rect 11437 22729 11471 22763
rect 13277 22729 13311 22763
rect 13645 22729 13679 22763
rect 15485 22729 15519 22763
rect 10333 22661 10367 22695
rect 11713 22661 11747 22695
rect 1777 22593 1811 22627
rect 2881 22593 2915 22627
rect 7389 22593 7423 22627
rect 8309 22593 8343 22627
rect 8861 22593 8895 22627
rect 8953 22593 8987 22627
rect 9413 22593 9447 22627
rect 10793 22593 10827 22627
rect 10977 22593 11011 22627
rect 12725 22593 12759 22627
rect 1501 22525 1535 22559
rect 2973 22525 3007 22559
rect 3240 22525 3274 22559
rect 5457 22525 5491 22559
rect 7297 22525 7331 22559
rect 9873 22525 9907 22559
rect 12265 22525 12299 22559
rect 12541 22525 12575 22559
rect 14105 22525 14139 22559
rect 7205 22457 7239 22491
rect 14350 22457 14384 22491
rect 2421 22389 2455 22423
rect 4353 22389 4387 22423
rect 5273 22389 5307 22423
rect 6837 22389 6871 22423
rect 7941 22389 7975 22423
rect 8769 22389 8803 22423
rect 10149 22389 10183 22423
rect 10701 22389 10735 22423
rect 16037 22389 16071 22423
rect 16589 22389 16623 22423
rect 17693 22389 17727 22423
rect 19441 22389 19475 22423
rect 20913 22389 20947 22423
rect 2421 22185 2455 22219
rect 3801 22185 3835 22219
rect 8493 22185 8527 22219
rect 13369 22185 13403 22219
rect 13461 22185 13495 22219
rect 4721 22117 4755 22151
rect 11222 22117 11256 22151
rect 1409 22049 1443 22083
rect 2053 22049 2087 22083
rect 2513 22049 2547 22083
rect 5917 22049 5951 22083
rect 6929 22049 6963 22083
rect 7380 22049 7414 22083
rect 9689 22049 9723 22083
rect 13829 22049 13863 22083
rect 15301 22049 15335 22083
rect 15577 22049 15611 22083
rect 3157 21981 3191 22015
rect 4813 21981 4847 22015
rect 4997 21981 5031 22015
rect 6561 21981 6595 22015
rect 7113 21981 7147 22015
rect 9873 21981 9907 22015
rect 10977 21981 11011 22015
rect 13921 21981 13955 22015
rect 14105 21981 14139 22015
rect 1593 21913 1627 21947
rect 4353 21913 4387 21947
rect 6101 21913 6135 21947
rect 2697 21845 2731 21879
rect 3433 21845 3467 21879
rect 5365 21845 5399 21879
rect 5733 21845 5767 21879
rect 9045 21845 9079 21879
rect 9505 21845 9539 21879
rect 10609 21845 10643 21879
rect 12357 21845 12391 21879
rect 13001 21845 13035 21879
rect 14657 21845 14691 21879
rect 2329 21641 2363 21675
rect 2789 21641 2823 21675
rect 3893 21641 3927 21675
rect 5457 21641 5491 21675
rect 6101 21641 6135 21675
rect 7665 21641 7699 21675
rect 9965 21641 9999 21675
rect 11529 21641 11563 21675
rect 12081 21641 12115 21675
rect 13921 21641 13955 21675
rect 15945 21641 15979 21675
rect 4353 21573 4387 21607
rect 13001 21573 13035 21607
rect 3249 21505 3283 21539
rect 3341 21505 3375 21539
rect 4905 21505 4939 21539
rect 7573 21505 7607 21539
rect 8125 21505 8159 21539
rect 8309 21505 8343 21539
rect 9045 21505 9079 21539
rect 9505 21505 9539 21539
rect 10425 21505 10459 21539
rect 10977 21505 11011 21539
rect 11161 21505 11195 21539
rect 1501 21437 1535 21471
rect 4261 21437 4295 21471
rect 4813 21437 4847 21471
rect 6469 21437 6503 21471
rect 12265 21437 12299 21471
rect 13093 21437 13127 21471
rect 14565 21437 14599 21471
rect 1777 21369 1811 21403
rect 3157 21369 3191 21403
rect 13369 21369 13403 21403
rect 14810 21369 14844 21403
rect 2697 21301 2731 21335
rect 4721 21301 4755 21335
rect 5825 21301 5859 21335
rect 6285 21301 6319 21335
rect 7205 21301 7239 21335
rect 8033 21301 8067 21335
rect 8677 21301 8711 21335
rect 10517 21301 10551 21335
rect 10885 21301 10919 21335
rect 11989 21301 12023 21335
rect 14197 21301 14231 21335
rect 2513 21097 2547 21131
rect 3433 21097 3467 21131
rect 5457 21097 5491 21131
rect 6009 21097 6043 21131
rect 8493 21097 8527 21131
rect 13645 21097 13679 21131
rect 16313 21097 16347 21131
rect 1777 21029 1811 21063
rect 3801 21029 3835 21063
rect 4322 21029 4356 21063
rect 11222 21029 11256 21063
rect 1501 20961 1535 20995
rect 2789 20961 2823 20995
rect 4077 20961 4111 20995
rect 7021 20961 7055 20995
rect 7380 20961 7414 20995
rect 9689 20961 9723 20995
rect 10977 20961 11011 20995
rect 14013 20961 14047 20995
rect 15301 20961 15335 20995
rect 7113 20893 7147 20927
rect 9873 20893 9907 20927
rect 14105 20893 14139 20927
rect 14197 20893 14231 20927
rect 6377 20825 6411 20859
rect 6837 20825 6871 20859
rect 2973 20757 3007 20791
rect 9137 20757 9171 20791
rect 9505 20757 9539 20791
rect 10609 20757 10643 20791
rect 12357 20757 12391 20791
rect 13185 20757 13219 20791
rect 14749 20757 14783 20791
rect 15025 20757 15059 20791
rect 15761 20757 15795 20791
rect 2697 20553 2731 20587
rect 3801 20553 3835 20587
rect 4169 20553 4203 20587
rect 7205 20553 7239 20587
rect 9137 20553 9171 20587
rect 9781 20553 9815 20587
rect 11253 20553 11287 20587
rect 12265 20553 12299 20587
rect 13185 20553 13219 20587
rect 14289 20553 14323 20587
rect 16129 20553 16163 20587
rect 11621 20485 11655 20519
rect 1685 20417 1719 20451
rect 2605 20417 2639 20451
rect 3341 20417 3375 20451
rect 7757 20417 7791 20451
rect 10701 20417 10735 20451
rect 10885 20417 10919 20451
rect 13093 20417 13127 20451
rect 13645 20417 13679 20451
rect 13829 20417 13863 20451
rect 1409 20349 1443 20383
rect 4261 20349 4295 20383
rect 4517 20349 4551 20383
rect 12725 20349 12759 20383
rect 14749 20349 14783 20383
rect 2237 20281 2271 20315
rect 3065 20281 3099 20315
rect 6193 20281 6227 20315
rect 7665 20281 7699 20315
rect 8002 20281 8036 20315
rect 10149 20281 10183 20315
rect 10609 20281 10643 20315
rect 14657 20281 14691 20315
rect 15016 20281 15050 20315
rect 3157 20213 3191 20247
rect 5641 20213 5675 20247
rect 6653 20213 6687 20247
rect 10241 20213 10275 20247
rect 13553 20213 13587 20247
rect 3341 20009 3375 20043
rect 4077 20009 4111 20043
rect 7021 20009 7055 20043
rect 8493 20009 8527 20043
rect 9873 20009 9907 20043
rect 14013 20009 14047 20043
rect 16681 20009 16715 20043
rect 1777 19941 1811 19975
rect 9413 19941 9447 19975
rect 10333 19941 10367 19975
rect 10692 19941 10726 19975
rect 1501 19873 1535 19907
rect 2789 19873 2823 19907
rect 5356 19873 5390 19907
rect 7665 19873 7699 19907
rect 7941 19873 7975 19907
rect 8401 19873 8435 19907
rect 13277 19873 13311 19907
rect 14289 19873 14323 19907
rect 15557 19873 15591 19907
rect 5089 19805 5123 19839
rect 8677 19805 8711 19839
rect 10425 19805 10459 19839
rect 13369 19805 13403 19839
rect 13553 19805 13587 19839
rect 15301 19805 15335 19839
rect 2697 19737 2731 19771
rect 15117 19737 15151 19771
rect 2329 19669 2363 19703
rect 2973 19669 3007 19703
rect 3801 19669 3835 19703
rect 4813 19669 4847 19703
rect 6469 19669 6503 19703
rect 7757 19669 7791 19703
rect 8033 19669 8067 19703
rect 9045 19669 9079 19703
rect 11805 19669 11839 19703
rect 12541 19669 12575 19703
rect 12909 19669 12943 19703
rect 14657 19669 14691 19703
rect 7941 19465 7975 19499
rect 10977 19465 11011 19499
rect 12541 19465 12575 19499
rect 13553 19465 13587 19499
rect 15761 19465 15795 19499
rect 16313 19397 16347 19431
rect 4261 19329 4295 19363
rect 5549 19329 5583 19363
rect 6009 19329 6043 19363
rect 10517 19329 10551 19363
rect 13185 19329 13219 19363
rect 14381 19329 14415 19363
rect 2053 19261 2087 19295
rect 4629 19261 4663 19295
rect 4905 19261 4939 19295
rect 5457 19261 5491 19295
rect 8033 19261 8067 19295
rect 10333 19261 10367 19295
rect 11713 19261 11747 19295
rect 12173 19261 12207 19295
rect 12909 19261 12943 19295
rect 1961 19193 1995 19227
rect 2298 19193 2332 19227
rect 7481 19193 7515 19227
rect 8300 19193 8334 19227
rect 11437 19193 11471 19227
rect 14289 19193 14323 19227
rect 14648 19193 14682 19227
rect 3433 19125 3467 19159
rect 4721 19125 4755 19159
rect 4997 19125 5031 19159
rect 5365 19125 5399 19159
rect 6377 19125 6411 19159
rect 7021 19125 7055 19159
rect 9413 19125 9447 19159
rect 9965 19125 9999 19159
rect 11529 19125 11563 19159
rect 13001 19125 13035 19159
rect 1593 18921 1627 18955
rect 2053 18921 2087 18955
rect 4721 18921 4755 18955
rect 7757 18921 7791 18955
rect 8309 18921 8343 18955
rect 8953 18921 8987 18955
rect 11345 18921 11379 18955
rect 11437 18921 11471 18955
rect 12541 18921 12575 18955
rect 13001 18921 13035 18955
rect 13461 18921 13495 18955
rect 15577 18921 15611 18955
rect 8217 18853 8251 18887
rect 11897 18853 11931 18887
rect 2605 18785 2639 18819
rect 4077 18785 4111 18819
rect 5273 18785 5307 18819
rect 5540 18785 5574 18819
rect 7205 18785 7239 18819
rect 9965 18785 9999 18819
rect 11805 18785 11839 18819
rect 13369 18785 13403 18819
rect 2697 18717 2731 18751
rect 2881 18717 2915 18751
rect 8401 18717 8435 18751
rect 10149 18717 10183 18751
rect 11989 18717 12023 18751
rect 13553 18717 13587 18751
rect 3341 18649 3375 18683
rect 7849 18649 7883 18683
rect 14013 18649 14047 18683
rect 2237 18581 2271 18615
rect 3709 18581 3743 18615
rect 4261 18581 4295 18615
rect 4997 18581 5031 18615
rect 6653 18581 6687 18615
rect 9229 18581 9263 18615
rect 10701 18581 10735 18615
rect 12817 18581 12851 18615
rect 14381 18581 14415 18615
rect 14749 18581 14783 18615
rect 3617 18377 3651 18411
rect 4537 18377 4571 18411
rect 6561 18377 6595 18411
rect 7849 18377 7883 18411
rect 8217 18377 8251 18411
rect 9505 18377 9539 18411
rect 11437 18377 11471 18411
rect 12173 18377 12207 18411
rect 13093 18377 13127 18411
rect 14749 18377 14783 18411
rect 6837 18309 6871 18343
rect 11161 18309 11195 18343
rect 2237 18241 2271 18275
rect 4261 18241 4295 18275
rect 5181 18241 5215 18275
rect 5273 18241 5307 18275
rect 7389 18241 7423 18275
rect 8953 18241 8987 18275
rect 9873 18241 9907 18275
rect 10517 18241 10551 18275
rect 6193 18173 6227 18207
rect 8861 18173 8895 18207
rect 10333 18173 10367 18207
rect 11897 18173 11931 18207
rect 13369 18173 13403 18207
rect 13636 18173 13670 18207
rect 2145 18105 2179 18139
rect 2504 18105 2538 18139
rect 7205 18105 7239 18139
rect 1593 18037 1627 18071
rect 4721 18037 4755 18071
rect 5089 18037 5123 18071
rect 5825 18037 5859 18071
rect 7297 18037 7331 18071
rect 8401 18037 8435 18071
rect 8769 18037 8803 18071
rect 9965 18037 9999 18071
rect 10425 18037 10459 18071
rect 11713 18037 11747 18071
rect 12725 18037 12759 18071
rect 2329 17833 2363 17867
rect 2421 17833 2455 17867
rect 3433 17833 3467 17867
rect 4077 17833 4111 17867
rect 5181 17833 5215 17867
rect 7941 17833 7975 17867
rect 8493 17833 8527 17867
rect 13737 17833 13771 17867
rect 2789 17765 2823 17799
rect 6184 17765 6218 17799
rect 14197 17765 14231 17799
rect 14841 17765 14875 17799
rect 4445 17697 4479 17731
rect 5917 17697 5951 17731
rect 9137 17697 9171 17731
rect 10057 17697 10091 17731
rect 11253 17697 11287 17731
rect 11520 17697 11554 17731
rect 1409 17629 1443 17663
rect 1869 17629 1903 17663
rect 2881 17629 2915 17663
rect 3065 17629 3099 17663
rect 4537 17629 4571 17663
rect 4721 17629 4755 17663
rect 5549 17629 5583 17663
rect 8585 17629 8619 17663
rect 9505 17629 9539 17663
rect 10149 17629 10183 17663
rect 10241 17629 10275 17663
rect 12633 17561 12667 17595
rect 3801 17493 3835 17527
rect 7297 17493 7331 17527
rect 9689 17493 9723 17527
rect 10885 17493 10919 17527
rect 13369 17493 13403 17527
rect 1409 17289 1443 17323
rect 3341 17289 3375 17323
rect 6009 17289 6043 17323
rect 9781 17289 9815 17323
rect 11253 17289 11287 17323
rect 11805 17289 11839 17323
rect 12173 17289 12207 17323
rect 13277 17289 13311 17323
rect 14381 17289 14415 17323
rect 2421 17221 2455 17255
rect 3617 17221 3651 17255
rect 8769 17221 8803 17255
rect 2053 17153 2087 17187
rect 3801 17153 3835 17187
rect 7297 17153 7331 17187
rect 9873 17153 9907 17187
rect 13829 17153 13863 17187
rect 14657 17153 14691 17187
rect 1777 17085 1811 17119
rect 4068 17085 4102 17119
rect 7389 17085 7423 17119
rect 7656 17085 7690 17119
rect 13185 17085 13219 17119
rect 13737 17085 13771 17119
rect 14841 17085 14875 17119
rect 15097 17085 15131 17119
rect 9413 17017 9447 17051
rect 10140 17017 10174 17051
rect 1869 16949 1903 16983
rect 2789 16949 2823 16983
rect 5181 16949 5215 16983
rect 6285 16949 6319 16983
rect 12633 16949 12667 16983
rect 13645 16949 13679 16983
rect 16221 16949 16255 16983
rect 1685 16745 1719 16779
rect 2053 16745 2087 16779
rect 2145 16745 2179 16779
rect 3157 16745 3191 16779
rect 3893 16745 3927 16779
rect 4721 16745 4755 16779
rect 6745 16745 6779 16779
rect 7389 16745 7423 16779
rect 9965 16745 9999 16779
rect 10149 16745 10183 16779
rect 11253 16745 11287 16779
rect 11621 16745 11655 16779
rect 12449 16745 12483 16779
rect 2605 16677 2639 16711
rect 5825 16677 5859 16711
rect 8309 16677 8343 16711
rect 9137 16677 9171 16711
rect 10517 16677 10551 16711
rect 12541 16677 12575 16711
rect 13277 16677 13311 16711
rect 14197 16677 14231 16711
rect 2513 16609 2547 16643
rect 4353 16609 4387 16643
rect 5089 16609 5123 16643
rect 6653 16609 6687 16643
rect 7665 16609 7699 16643
rect 8217 16609 8251 16643
rect 9045 16609 9079 16643
rect 10609 16609 10643 16643
rect 13921 16609 13955 16643
rect 2697 16541 2731 16575
rect 5181 16541 5215 16575
rect 5273 16541 5307 16575
rect 6101 16541 6135 16575
rect 6837 16541 6871 16575
rect 8401 16541 8435 16575
rect 9229 16541 9263 16575
rect 10793 16541 10827 16575
rect 12725 16541 12759 16575
rect 6285 16473 6319 16507
rect 7849 16473 7883 16507
rect 8677 16473 8711 16507
rect 12081 16473 12115 16507
rect 11897 16405 11931 16439
rect 13737 16405 13771 16439
rect 14749 16405 14783 16439
rect 1593 16201 1627 16235
rect 5181 16201 5215 16235
rect 6377 16201 6411 16235
rect 7297 16201 7331 16235
rect 10793 16201 10827 16235
rect 12081 16201 12115 16235
rect 15209 16201 15243 16235
rect 5825 16065 5859 16099
rect 11253 16065 11287 16099
rect 11437 16065 11471 16099
rect 12633 16065 12667 16099
rect 13829 16065 13863 16099
rect 16589 16065 16623 16099
rect 1409 15997 1443 16031
rect 2697 15997 2731 16031
rect 4721 15997 4755 16031
rect 5641 15997 5675 16031
rect 10701 15997 10735 16031
rect 11161 15997 11195 16031
rect 12449 15997 12483 16031
rect 16313 15997 16347 16031
rect 17049 15997 17083 16031
rect 2942 15929 2976 15963
rect 5549 15929 5583 15963
rect 6837 15929 6871 15963
rect 8309 15929 8343 15963
rect 8401 15929 8435 15963
rect 14074 15929 14108 15963
rect 2053 15861 2087 15895
rect 2421 15861 2455 15895
rect 4077 15861 4111 15895
rect 7941 15861 7975 15895
rect 9689 15861 9723 15895
rect 13277 15861 13311 15895
rect 13645 15861 13679 15895
rect 3893 15657 3927 15691
rect 4261 15657 4295 15691
rect 5273 15657 5307 15691
rect 7389 15657 7423 15691
rect 10977 15657 11011 15691
rect 11437 15657 11471 15691
rect 14473 15657 14507 15691
rect 14841 15657 14875 15691
rect 15761 15657 15795 15691
rect 5632 15589 5666 15623
rect 7757 15589 7791 15623
rect 1501 15521 1535 15555
rect 1768 15521 1802 15555
rect 4077 15521 4111 15555
rect 5365 15521 5399 15555
rect 7849 15521 7883 15555
rect 8116 15521 8150 15555
rect 9689 15521 9723 15555
rect 11345 15521 11379 15555
rect 12541 15521 12575 15555
rect 12808 15521 12842 15555
rect 15669 15521 15703 15555
rect 9873 15453 9907 15487
rect 11621 15453 11655 15487
rect 15945 15453 15979 15487
rect 9229 15385 9263 15419
rect 10885 15385 10919 15419
rect 13921 15385 13955 15419
rect 2881 15317 2915 15351
rect 3433 15317 3467 15351
rect 4813 15317 4847 15351
rect 6745 15317 6779 15351
rect 10517 15317 10551 15351
rect 12173 15317 12207 15351
rect 15301 15317 15335 15351
rect 2237 15113 2271 15147
rect 3709 15113 3743 15147
rect 4077 15113 4111 15147
rect 6193 15113 6227 15147
rect 11897 15113 11931 15147
rect 12541 15113 12575 15147
rect 13645 15113 13679 15147
rect 15761 15113 15795 15147
rect 16681 15113 16715 15147
rect 7021 15045 7055 15079
rect 2881 14977 2915 15011
rect 8033 14977 8067 15011
rect 10333 14977 10367 15011
rect 11437 14977 11471 15011
rect 13001 14977 13035 15011
rect 13185 14977 13219 15011
rect 14381 14977 14415 15011
rect 4169 14909 4203 14943
rect 4425 14909 4459 14943
rect 6837 14909 6871 14943
rect 8289 14909 8323 14943
rect 11161 14909 11195 14943
rect 14648 14909 14682 14943
rect 2605 14841 2639 14875
rect 3341 14841 3375 14875
rect 7573 14841 7607 14875
rect 10609 14841 10643 14875
rect 11253 14841 11287 14875
rect 12909 14841 12943 14875
rect 14289 14841 14323 14875
rect 1593 14773 1627 14807
rect 2053 14773 2087 14807
rect 2697 14773 2731 14807
rect 5549 14773 5583 14807
rect 6653 14773 6687 14807
rect 7941 14773 7975 14807
rect 9413 14773 9447 14807
rect 10793 14773 10827 14807
rect 12265 14773 12299 14807
rect 16313 14773 16347 14807
rect 1409 14569 1443 14603
rect 2421 14569 2455 14603
rect 2881 14569 2915 14603
rect 7573 14569 7607 14603
rect 7941 14569 7975 14603
rect 9045 14569 9079 14603
rect 11805 14569 11839 14603
rect 12173 14569 12207 14603
rect 14105 14569 14139 14603
rect 14657 14569 14691 14603
rect 15025 14569 15059 14603
rect 15577 14569 15611 14603
rect 3801 14501 3835 14535
rect 4537 14501 4571 14535
rect 4905 14501 4939 14535
rect 5264 14501 5298 14535
rect 8033 14501 8067 14535
rect 11069 14501 11103 14535
rect 12970 14501 13004 14535
rect 16129 14501 16163 14535
rect 2789 14433 2823 14467
rect 4997 14433 5031 14467
rect 9321 14433 9355 14467
rect 12449 14433 12483 14467
rect 15853 14433 15887 14467
rect 2973 14365 3007 14399
rect 8125 14365 8159 14399
rect 8585 14365 8619 14399
rect 9689 14365 9723 14399
rect 11161 14365 11195 14399
rect 11345 14365 11379 14399
rect 12725 14365 12759 14399
rect 1869 14297 1903 14331
rect 2329 14297 2363 14331
rect 10517 14297 10551 14331
rect 12265 14297 12299 14331
rect 3433 14229 3467 14263
rect 6377 14229 6411 14263
rect 7021 14229 7055 14263
rect 7481 14229 7515 14263
rect 9137 14229 9171 14263
rect 10701 14229 10735 14263
rect 1501 14025 1535 14059
rect 3065 14025 3099 14059
rect 4169 14025 4203 14059
rect 4629 14025 4663 14059
rect 6285 14025 6319 14059
rect 9965 14025 9999 14059
rect 10241 14025 10275 14059
rect 11437 14025 11471 14059
rect 13829 14025 13863 14059
rect 14381 14025 14415 14059
rect 16313 14025 16347 14059
rect 2513 13957 2547 13991
rect 2973 13957 3007 13991
rect 4537 13957 4571 13991
rect 6837 13957 6871 13991
rect 7849 13957 7883 13991
rect 1961 13889 1995 13923
rect 2145 13889 2179 13923
rect 3709 13889 3743 13923
rect 5733 13889 5767 13923
rect 7435 13889 7469 13923
rect 8861 13889 8895 13923
rect 9045 13889 9079 13923
rect 9505 13889 9539 13923
rect 10425 13957 10459 13991
rect 10977 13889 11011 13923
rect 12173 13889 12207 13923
rect 12449 13889 12483 13923
rect 14841 13889 14875 13923
rect 1869 13821 1903 13855
rect 3525 13821 3559 13855
rect 4813 13821 4847 13855
rect 5641 13821 5675 13855
rect 7205 13821 7239 13855
rect 10149 13821 10183 13855
rect 10241 13821 10275 13855
rect 10793 13821 10827 13855
rect 12705 13821 12739 13855
rect 14933 13821 14967 13855
rect 15200 13821 15234 13855
rect 5549 13753 5583 13787
rect 8769 13753 8803 13787
rect 9873 13753 9907 13787
rect 10885 13753 10919 13787
rect 11805 13753 11839 13787
rect 3433 13685 3467 13719
rect 5181 13685 5215 13719
rect 6561 13685 6595 13719
rect 7297 13685 7331 13719
rect 8217 13685 8251 13719
rect 8401 13685 8435 13719
rect 1869 13481 1903 13515
rect 2421 13481 2455 13515
rect 3525 13481 3559 13515
rect 3801 13481 3835 13515
rect 4721 13481 4755 13515
rect 4813 13481 4847 13515
rect 5273 13481 5307 13515
rect 6837 13481 6871 13515
rect 7021 13481 7055 13515
rect 7481 13481 7515 13515
rect 8033 13481 8067 13515
rect 8493 13481 8527 13515
rect 9045 13481 9079 13515
rect 9413 13481 9447 13515
rect 10057 13481 10091 13515
rect 12817 13481 12851 13515
rect 13369 13481 13403 13515
rect 13921 13481 13955 13515
rect 15853 13481 15887 13515
rect 5181 13413 5215 13447
rect 7389 13413 7423 13447
rect 13829 13413 13863 13447
rect 14933 13413 14967 13447
rect 16957 13413 16991 13447
rect 1777 13345 1811 13379
rect 6285 13345 6319 13379
rect 6561 13345 6595 13379
rect 8585 13345 8619 13379
rect 11704 13345 11738 13379
rect 16681 13345 16715 13379
rect 2053 13277 2087 13311
rect 2973 13277 3007 13311
rect 5457 13277 5491 13311
rect 7573 13277 7607 13311
rect 10149 13277 10183 13311
rect 10241 13277 10275 13311
rect 11437 13277 11471 13311
rect 4353 13209 4387 13243
rect 9689 13209 9723 13243
rect 1409 13141 1443 13175
rect 2881 13141 2915 13175
rect 5917 13141 5951 13175
rect 6377 13141 6411 13175
rect 10793 13141 10827 13175
rect 11161 13141 11195 13175
rect 3433 12937 3467 12971
rect 4905 12937 4939 12971
rect 6285 12937 6319 12971
rect 9321 12937 9355 12971
rect 9689 12937 9723 12971
rect 10149 12937 10183 12971
rect 10701 12937 10735 12971
rect 12081 12937 12115 12971
rect 17049 12937 17083 12971
rect 6653 12869 6687 12903
rect 8677 12869 8711 12903
rect 10609 12869 10643 12903
rect 5825 12801 5859 12835
rect 11161 12801 11195 12835
rect 11345 12801 11379 12835
rect 12449 12801 12483 12835
rect 16221 12801 16255 12835
rect 18337 12801 18371 12835
rect 1409 12733 1443 12767
rect 1676 12733 1710 12767
rect 4537 12733 4571 12767
rect 5549 12733 5583 12767
rect 7297 12733 7331 12767
rect 15945 12733 15979 12767
rect 16681 12733 16715 12767
rect 18061 12733 18095 12767
rect 18797 12733 18831 12767
rect 3893 12665 3927 12699
rect 5641 12665 5675 12699
rect 7564 12665 7598 12699
rect 11069 12665 11103 12699
rect 2789 12597 2823 12631
rect 3985 12597 4019 12631
rect 5181 12597 5215 12631
rect 7113 12597 7147 12631
rect 11805 12597 11839 12631
rect 13001 12597 13035 12631
rect 1869 12393 1903 12427
rect 2421 12393 2455 12427
rect 2881 12393 2915 12427
rect 5641 12393 5675 12427
rect 8033 12393 8067 12427
rect 9229 12393 9263 12427
rect 11069 12393 11103 12427
rect 11621 12393 11655 12427
rect 3801 12325 3835 12359
rect 4537 12325 4571 12359
rect 6000 12325 6034 12359
rect 8217 12325 8251 12359
rect 10793 12325 10827 12359
rect 21189 12325 21223 12359
rect 1777 12257 1811 12291
rect 4445 12257 4479 12291
rect 5733 12257 5767 12291
rect 8677 12257 8711 12291
rect 10057 12257 10091 12291
rect 11437 12257 11471 12291
rect 11989 12257 12023 12291
rect 20913 12257 20947 12291
rect 2053 12189 2087 12223
rect 4629 12189 4663 12223
rect 10149 12189 10183 12223
rect 10241 12189 10275 12223
rect 12081 12189 12115 12223
rect 12265 12189 12299 12223
rect 12633 12189 12667 12223
rect 3249 12121 3283 12155
rect 4077 12121 4111 12155
rect 1409 12053 1443 12087
rect 5273 12053 5307 12087
rect 7113 12053 7147 12087
rect 7757 12053 7791 12087
rect 9689 12053 9723 12087
rect 11253 12053 11287 12087
rect 2053 11849 2087 11883
rect 4169 11849 4203 11883
rect 5181 11849 5215 11883
rect 6193 11849 6227 11883
rect 8217 11849 8251 11883
rect 8861 11849 8895 11883
rect 11345 11849 11379 11883
rect 12081 11849 12115 11883
rect 13829 11849 13863 11883
rect 4721 11781 4755 11815
rect 4905 11781 4939 11815
rect 9137 11781 9171 11815
rect 5825 11713 5859 11747
rect 6837 11713 6871 11747
rect 12449 11713 12483 11747
rect 2145 11645 2179 11679
rect 5089 11645 5123 11679
rect 5549 11645 5583 11679
rect 7104 11645 7138 11679
rect 9321 11645 9355 11679
rect 2412 11577 2446 11611
rect 6653 11577 6687 11611
rect 9588 11577 9622 11611
rect 12694 11577 12728 11611
rect 1593 11509 1627 11543
rect 3525 11509 3559 11543
rect 5641 11509 5675 11543
rect 10701 11509 10735 11543
rect 11713 11509 11747 11543
rect 20913 11509 20947 11543
rect 1409 11305 1443 11339
rect 1869 11305 1903 11339
rect 3433 11305 3467 11339
rect 3893 11305 3927 11339
rect 6101 11305 6135 11339
rect 6377 11305 6411 11339
rect 7297 11305 7331 11339
rect 8033 11305 8067 11339
rect 8493 11305 8527 11339
rect 10885 11305 10919 11339
rect 12449 11305 12483 11339
rect 13001 11305 13035 11339
rect 2881 11237 2915 11271
rect 4322 11237 4356 11271
rect 9965 11237 9999 11271
rect 18245 11237 18279 11271
rect 1777 11169 1811 11203
rect 2421 11169 2455 11203
rect 2973 11169 3007 11203
rect 4077 11169 4111 11203
rect 8401 11169 8435 11203
rect 9689 11169 9723 11203
rect 11069 11169 11103 11203
rect 11336 11169 11370 11203
rect 17969 11169 18003 11203
rect 1961 11101 1995 11135
rect 8677 11101 8711 11135
rect 7573 11033 7607 11067
rect 9413 11033 9447 11067
rect 10425 11033 10459 11067
rect 5457 10965 5491 10999
rect 6837 10965 6871 10999
rect 5641 10761 5675 10795
rect 8125 10761 8159 10795
rect 8953 10761 8987 10795
rect 9413 10761 9447 10795
rect 12265 10761 12299 10795
rect 18245 10761 18279 10795
rect 2145 10625 2179 10659
rect 2973 10625 3007 10659
rect 4261 10625 4295 10659
rect 7389 10625 7423 10659
rect 9781 10625 9815 10659
rect 12449 10625 12483 10659
rect 18705 10625 18739 10659
rect 19993 10625 20027 10659
rect 2697 10557 2731 10591
rect 4528 10557 4562 10591
rect 7205 10557 7239 10591
rect 9873 10557 9907 10591
rect 10140 10557 10174 10591
rect 18429 10557 18463 10591
rect 19165 10557 19199 10591
rect 19717 10557 19751 10591
rect 20453 10557 20487 10591
rect 1869 10489 1903 10523
rect 2789 10489 2823 10523
rect 3709 10489 3743 10523
rect 4169 10489 4203 10523
rect 6285 10489 6319 10523
rect 7297 10489 7331 10523
rect 2329 10421 2363 10455
rect 3341 10421 3375 10455
rect 6561 10421 6595 10455
rect 6837 10421 6871 10455
rect 8401 10421 8435 10455
rect 11253 10421 11287 10455
rect 11897 10421 11931 10455
rect 2789 10217 2823 10251
rect 3433 10217 3467 10251
rect 3801 10217 3835 10251
rect 4537 10217 4571 10251
rect 4905 10217 4939 10251
rect 7573 10217 7607 10251
rect 8217 10217 8251 10251
rect 10057 10217 10091 10251
rect 10793 10217 10827 10251
rect 11069 10217 11103 10251
rect 11253 10217 11287 10251
rect 1676 10149 1710 10183
rect 8769 10149 8803 10183
rect 19809 10149 19843 10183
rect 5273 10081 5307 10115
rect 5540 10081 5574 10115
rect 8125 10081 8159 10115
rect 11621 10081 11655 10115
rect 19533 10081 19567 10115
rect 1409 10013 1443 10047
rect 4077 10013 4111 10047
rect 8309 10013 8343 10047
rect 10149 10013 10183 10047
rect 10241 10013 10275 10047
rect 11713 10013 11747 10047
rect 11897 10013 11931 10047
rect 7757 9945 7791 9979
rect 9413 9945 9447 9979
rect 9689 9945 9723 9979
rect 6653 9877 6687 9911
rect 7297 9877 7331 9911
rect 3065 9673 3099 9707
rect 3985 9673 4019 9707
rect 6837 9673 6871 9707
rect 8217 9673 8251 9707
rect 10609 9673 10643 9707
rect 11713 9673 11747 9707
rect 11989 9673 12023 9707
rect 19533 9673 19567 9707
rect 1685 9537 1719 9571
rect 7389 9537 7423 9571
rect 3617 9469 3651 9503
rect 4169 9469 4203 9503
rect 4425 9469 4459 9503
rect 6561 9469 6595 9503
rect 7205 9469 7239 9503
rect 7849 9469 7883 9503
rect 8677 9469 8711 9503
rect 1952 9401 1986 9435
rect 6285 9401 6319 9435
rect 7297 9401 7331 9435
rect 8944 9401 8978 9435
rect 5549 9333 5583 9367
rect 10057 9333 10091 9367
rect 11253 9333 11287 9367
rect 1777 9129 1811 9163
rect 2053 9129 2087 9163
rect 3801 9129 3835 9163
rect 4537 9129 4571 9163
rect 5365 9129 5399 9163
rect 7757 9129 7791 9163
rect 8309 9129 8343 9163
rect 8769 9129 8803 9163
rect 9505 9129 9539 9163
rect 9689 9129 9723 9163
rect 2881 9061 2915 9095
rect 4445 9061 4479 9095
rect 5641 9061 5675 9095
rect 9045 9061 9079 9095
rect 2789 8993 2823 9027
rect 3525 8993 3559 9027
rect 6377 8993 6411 9027
rect 6633 8993 6667 9027
rect 10057 8993 10091 9027
rect 3065 8925 3099 8959
rect 4721 8925 4755 8959
rect 10149 8925 10183 8959
rect 10333 8925 10367 8959
rect 4077 8857 4111 8891
rect 2421 8789 2455 8823
rect 1593 8585 1627 8619
rect 1961 8585 1995 8619
rect 2513 8585 2547 8619
rect 2881 8585 2915 8619
rect 3985 8585 4019 8619
rect 5457 8585 5491 8619
rect 6469 8585 6503 8619
rect 7021 8585 7055 8619
rect 7573 8585 7607 8619
rect 9045 8585 9079 8619
rect 10609 8585 10643 8619
rect 3157 8517 3191 8551
rect 9689 8517 9723 8551
rect 3617 8449 3651 8483
rect 7665 8449 7699 8483
rect 10149 8449 10183 8483
rect 4077 8381 4111 8415
rect 4344 8381 4378 8415
rect 7932 8313 7966 8347
rect 3893 8041 3927 8075
rect 4537 8041 4571 8075
rect 5825 8041 5859 8075
rect 7665 8041 7699 8075
rect 9965 8041 9999 8075
rect 22477 8041 22511 8075
rect 3525 7973 3559 8007
rect 4445 7973 4479 8007
rect 22293 7905 22327 7939
rect 4721 7837 4755 7871
rect 4077 7769 4111 7803
rect 4169 7497 4203 7531
rect 4813 7497 4847 7531
rect 22293 7497 22327 7531
rect 23857 7497 23891 7531
rect 4537 7361 4571 7395
rect 23673 7293 23707 7327
rect 24225 7293 24259 7327
rect 23857 6409 23891 6443
rect 23673 6205 23707 6239
rect 24225 6205 24259 6239
rect 24225 5865 24259 5899
rect 24041 5729 24075 5763
rect 24041 5321 24075 5355
rect 24685 5321 24719 5355
rect 24501 5117 24535 5151
rect 25053 5117 25087 5151
rect 24777 4777 24811 4811
rect 24593 4641 24627 4675
rect 24685 4233 24719 4267
<< metal1 >>
rect 3878 26664 3884 26716
rect 3936 26704 3942 26716
rect 7098 26704 7104 26716
rect 3936 26676 7104 26704
rect 3936 26664 3942 26676
rect 7098 26664 7104 26676
rect 7156 26664 7162 26716
rect 4062 26392 4068 26444
rect 4120 26432 4126 26444
rect 5534 26432 5540 26444
rect 4120 26404 5540 26432
rect 4120 26392 4126 26404
rect 5534 26392 5540 26404
rect 5592 26392 5598 26444
rect 3510 26256 3516 26308
rect 3568 26296 3574 26308
rect 4890 26296 4896 26308
rect 3568 26268 4896 26296
rect 3568 26256 3574 26268
rect 4890 26256 4896 26268
rect 4948 26256 4954 26308
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 3326 25440 3332 25492
rect 3384 25480 3390 25492
rect 4249 25483 4307 25489
rect 4249 25480 4261 25483
rect 3384 25452 4261 25480
rect 3384 25440 3390 25452
rect 4249 25449 4261 25452
rect 4295 25449 4307 25483
rect 9950 25480 9956 25492
rect 4249 25443 4307 25449
rect 5276 25452 9956 25480
rect 2314 25412 2320 25424
rect 1412 25384 2320 25412
rect 1412 25353 1440 25384
rect 2314 25372 2320 25384
rect 2372 25412 2378 25424
rect 5276 25412 5304 25452
rect 9950 25440 9956 25452
rect 10008 25440 10014 25492
rect 2372 25384 5304 25412
rect 2372 25372 2378 25384
rect 5350 25372 5356 25424
rect 5408 25412 5414 25424
rect 6546 25412 6552 25424
rect 5408 25384 6552 25412
rect 5408 25372 5414 25384
rect 6546 25372 6552 25384
rect 6604 25412 6610 25424
rect 6604 25384 6960 25412
rect 6604 25372 6610 25384
rect 1397 25347 1455 25353
rect 1397 25313 1409 25347
rect 1443 25313 1455 25347
rect 2498 25344 2504 25356
rect 2459 25316 2504 25344
rect 1397 25307 1455 25313
rect 2498 25304 2504 25316
rect 2556 25304 2562 25356
rect 2590 25304 2596 25356
rect 2648 25344 2654 25356
rect 4065 25347 4123 25353
rect 4065 25344 4077 25347
rect 2648 25316 4077 25344
rect 2648 25304 2654 25316
rect 4065 25313 4077 25316
rect 4111 25344 4123 25347
rect 4154 25344 4160 25356
rect 4111 25316 4160 25344
rect 4111 25313 4123 25316
rect 4065 25307 4123 25313
rect 4154 25304 4160 25316
rect 4212 25304 4218 25356
rect 5169 25347 5227 25353
rect 5169 25313 5181 25347
rect 5215 25344 5227 25347
rect 5994 25344 6000 25356
rect 5215 25316 6000 25344
rect 5215 25313 5227 25316
rect 5169 25307 5227 25313
rect 5994 25304 6000 25316
rect 6052 25304 6058 25356
rect 6932 25353 6960 25384
rect 6917 25347 6975 25353
rect 6917 25313 6929 25347
rect 6963 25313 6975 25347
rect 6917 25307 6975 25313
rect 5258 25236 5264 25288
rect 5316 25276 5322 25288
rect 8021 25279 8079 25285
rect 8021 25276 8033 25279
rect 5316 25248 8033 25276
rect 5316 25236 5322 25248
rect 8021 25245 8033 25248
rect 8067 25245 8079 25279
rect 8021 25239 8079 25245
rect 9769 25279 9827 25285
rect 9769 25245 9781 25279
rect 9815 25245 9827 25279
rect 9769 25239 9827 25245
rect 1581 25211 1639 25217
rect 1581 25177 1593 25211
rect 1627 25208 1639 25211
rect 2866 25208 2872 25220
rect 1627 25180 2872 25208
rect 1627 25177 1639 25180
rect 1581 25171 1639 25177
rect 2866 25168 2872 25180
rect 2924 25168 2930 25220
rect 3786 25168 3792 25220
rect 3844 25208 3850 25220
rect 3844 25180 4844 25208
rect 3844 25168 3850 25180
rect 2038 25140 2044 25152
rect 1999 25112 2044 25140
rect 2038 25100 2044 25112
rect 2096 25100 2102 25152
rect 2406 25140 2412 25152
rect 2367 25112 2412 25140
rect 2406 25100 2412 25112
rect 2464 25100 2470 25152
rect 2685 25143 2743 25149
rect 2685 25109 2697 25143
rect 2731 25140 2743 25143
rect 2774 25140 2780 25152
rect 2731 25112 2780 25140
rect 2731 25109 2743 25112
rect 2685 25103 2743 25109
rect 2774 25100 2780 25112
rect 2832 25100 2838 25152
rect 4706 25140 4712 25152
rect 4667 25112 4712 25140
rect 4706 25100 4712 25112
rect 4764 25100 4770 25152
rect 4816 25140 4844 25180
rect 4890 25168 4896 25220
rect 4948 25208 4954 25220
rect 5353 25211 5411 25217
rect 5353 25208 5365 25211
rect 4948 25180 5365 25208
rect 4948 25168 4954 25180
rect 5353 25177 5365 25180
rect 5399 25177 5411 25211
rect 7098 25208 7104 25220
rect 7059 25180 7104 25208
rect 5353 25171 5411 25177
rect 7098 25168 7104 25180
rect 7156 25168 7162 25220
rect 9784 25140 9812 25239
rect 4816 25112 9812 25140
rect 10413 25143 10471 25149
rect 10413 25109 10425 25143
rect 10459 25140 10471 25143
rect 10778 25140 10784 25152
rect 10459 25112 10784 25140
rect 10459 25109 10471 25112
rect 10413 25103 10471 25109
rect 10778 25100 10784 25112
rect 10836 25100 10842 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 2498 24936 2504 24948
rect 1872 24908 2504 24936
rect 1872 24809 1900 24908
rect 2498 24896 2504 24908
rect 2556 24936 2562 24948
rect 2685 24939 2743 24945
rect 2685 24936 2697 24939
rect 2556 24908 2697 24936
rect 2556 24896 2562 24908
rect 2685 24905 2697 24908
rect 2731 24905 2743 24939
rect 2685 24899 2743 24905
rect 4065 24939 4123 24945
rect 4065 24905 4077 24939
rect 4111 24936 4123 24939
rect 4154 24936 4160 24948
rect 4111 24908 4160 24936
rect 4111 24905 4123 24908
rect 4065 24899 4123 24905
rect 4154 24896 4160 24908
rect 4212 24896 4218 24948
rect 2038 24828 2044 24880
rect 2096 24868 2102 24880
rect 4617 24871 4675 24877
rect 4617 24868 4629 24871
rect 2096 24840 4629 24868
rect 2096 24828 2102 24840
rect 4617 24837 4629 24840
rect 4663 24837 4675 24871
rect 10321 24871 10379 24877
rect 4617 24831 4675 24837
rect 6840 24840 8248 24868
rect 1857 24803 1915 24809
rect 1857 24769 1869 24803
rect 1903 24769 1915 24803
rect 1857 24763 1915 24769
rect 1581 24735 1639 24741
rect 1581 24701 1593 24735
rect 1627 24732 1639 24735
rect 2056 24732 2084 24828
rect 2314 24800 2320 24812
rect 2275 24772 2320 24800
rect 2314 24760 2320 24772
rect 2372 24760 2378 24812
rect 4706 24760 4712 24812
rect 4764 24800 4770 24812
rect 5077 24803 5135 24809
rect 5077 24800 5089 24803
rect 4764 24772 5089 24800
rect 4764 24760 4770 24772
rect 5077 24769 5089 24772
rect 5123 24769 5135 24803
rect 5077 24763 5135 24769
rect 5169 24803 5227 24809
rect 5169 24769 5181 24803
rect 5215 24800 5227 24803
rect 5350 24800 5356 24812
rect 5215 24772 5356 24800
rect 5215 24769 5227 24772
rect 5169 24763 5227 24769
rect 5350 24760 5356 24772
rect 5408 24760 5414 24812
rect 5721 24803 5779 24809
rect 5721 24769 5733 24803
rect 5767 24800 5779 24803
rect 5994 24800 6000 24812
rect 5767 24772 6000 24800
rect 5767 24769 5779 24772
rect 5721 24763 5779 24769
rect 5994 24760 6000 24772
rect 6052 24760 6058 24812
rect 6546 24800 6552 24812
rect 6507 24772 6552 24800
rect 6546 24760 6552 24772
rect 6604 24760 6610 24812
rect 1627 24704 2084 24732
rect 1627 24701 1639 24704
rect 1581 24695 1639 24701
rect 2682 24692 2688 24744
rect 2740 24732 2746 24744
rect 2869 24735 2927 24741
rect 2869 24732 2881 24735
rect 2740 24704 2881 24732
rect 2740 24692 2746 24704
rect 2869 24701 2881 24704
rect 2915 24732 2927 24735
rect 3421 24735 3479 24741
rect 3421 24732 3433 24735
rect 2915 24704 3433 24732
rect 2915 24701 2927 24704
rect 2869 24695 2927 24701
rect 3421 24701 3433 24704
rect 3467 24701 3479 24735
rect 3421 24695 3479 24701
rect 4525 24735 4583 24741
rect 4525 24701 4537 24735
rect 4571 24732 4583 24735
rect 4985 24735 5043 24741
rect 4985 24732 4997 24735
rect 4571 24704 4997 24732
rect 4571 24701 4583 24704
rect 4525 24695 4583 24701
rect 4985 24701 4997 24704
rect 5031 24732 5043 24735
rect 5258 24732 5264 24744
rect 5031 24704 5264 24732
rect 5031 24701 5043 24704
rect 4985 24695 5043 24701
rect 5258 24692 5264 24704
rect 5316 24692 5322 24744
rect 6840 24732 6868 24840
rect 7484 24809 7512 24840
rect 7469 24803 7527 24809
rect 7469 24769 7481 24803
rect 7515 24769 7527 24803
rect 8220 24800 8248 24840
rect 10321 24837 10333 24871
rect 10367 24837 10379 24871
rect 12437 24871 12495 24877
rect 12437 24868 12449 24871
rect 10321 24831 10379 24837
rect 10796 24840 12449 24868
rect 9214 24800 9220 24812
rect 8220 24772 9220 24800
rect 7469 24763 7527 24769
rect 9214 24760 9220 24772
rect 9272 24760 9278 24812
rect 9766 24760 9772 24812
rect 9824 24800 9830 24812
rect 10336 24800 10364 24831
rect 10796 24812 10824 24840
rect 12437 24837 12449 24840
rect 12483 24837 12495 24871
rect 12437 24831 12495 24837
rect 10778 24800 10784 24812
rect 9824 24772 10364 24800
rect 10739 24772 10784 24800
rect 9824 24760 9830 24772
rect 10778 24760 10784 24772
rect 10836 24760 10842 24812
rect 10962 24800 10968 24812
rect 10923 24772 10968 24800
rect 10962 24760 10968 24772
rect 11020 24760 11026 24812
rect 12253 24803 12311 24809
rect 12253 24769 12265 24803
rect 12299 24800 12311 24803
rect 12802 24800 12808 24812
rect 12299 24772 12808 24800
rect 12299 24769 12311 24772
rect 12253 24763 12311 24769
rect 12802 24760 12808 24772
rect 12860 24800 12866 24812
rect 12897 24803 12955 24809
rect 12897 24800 12909 24803
rect 12860 24772 12909 24800
rect 12860 24760 12866 24772
rect 12897 24769 12909 24772
rect 12943 24769 12955 24803
rect 13078 24800 13084 24812
rect 13039 24772 13084 24800
rect 12897 24763 12955 24769
rect 13078 24760 13084 24772
rect 13136 24760 13142 24812
rect 23842 24760 23848 24812
rect 23900 24800 23906 24812
rect 24762 24800 24768 24812
rect 23900 24772 24768 24800
rect 23900 24760 23906 24772
rect 24762 24760 24768 24772
rect 24820 24760 24826 24812
rect 6288 24704 6868 24732
rect 6288 24608 6316 24704
rect 7834 24692 7840 24744
rect 7892 24732 7898 24744
rect 8297 24735 8355 24741
rect 8297 24732 8309 24735
rect 7892 24704 8309 24732
rect 7892 24692 7898 24704
rect 8297 24701 8309 24704
rect 8343 24701 8355 24735
rect 8297 24695 8355 24701
rect 11885 24735 11943 24741
rect 11885 24701 11897 24735
rect 11931 24732 11943 24735
rect 13096 24732 13124 24760
rect 11931 24704 13124 24732
rect 15197 24735 15255 24741
rect 11931 24701 11943 24704
rect 11885 24695 11943 24701
rect 15197 24701 15209 24735
rect 15243 24732 15255 24735
rect 15562 24732 15568 24744
rect 15243 24704 15568 24732
rect 15243 24701 15255 24704
rect 15197 24695 15255 24701
rect 15562 24692 15568 24704
rect 15620 24692 15626 24744
rect 7006 24624 7012 24676
rect 7064 24664 7070 24676
rect 7285 24667 7343 24673
rect 7285 24664 7297 24667
rect 7064 24636 7297 24664
rect 7064 24624 7070 24636
rect 7285 24633 7297 24636
rect 7331 24664 7343 24667
rect 8481 24667 8539 24673
rect 8481 24664 8493 24667
rect 7331 24636 8493 24664
rect 7331 24633 7343 24636
rect 7285 24627 7343 24633
rect 8481 24633 8493 24636
rect 8527 24633 8539 24667
rect 10689 24667 10747 24673
rect 10689 24664 10701 24667
rect 8481 24627 8539 24633
rect 10152 24636 10701 24664
rect 10152 24608 10180 24636
rect 10689 24633 10701 24636
rect 10735 24633 10747 24667
rect 16482 24664 16488 24676
rect 10689 24627 10747 24633
rect 15396 24636 16488 24664
rect 3050 24596 3056 24608
rect 3011 24568 3056 24596
rect 3050 24556 3056 24568
rect 3108 24556 3114 24608
rect 6270 24596 6276 24608
rect 6231 24568 6276 24596
rect 6270 24556 6276 24568
rect 6328 24556 6334 24608
rect 6917 24599 6975 24605
rect 6917 24565 6929 24599
rect 6963 24596 6975 24599
rect 7098 24596 7104 24608
rect 6963 24568 7104 24596
rect 6963 24565 6975 24568
rect 6917 24559 6975 24565
rect 7098 24556 7104 24568
rect 7156 24556 7162 24608
rect 7377 24599 7435 24605
rect 7377 24565 7389 24599
rect 7423 24596 7435 24599
rect 8021 24599 8079 24605
rect 8021 24596 8033 24599
rect 7423 24568 8033 24596
rect 7423 24565 7435 24568
rect 7377 24559 7435 24565
rect 8021 24565 8033 24568
rect 8067 24596 8079 24599
rect 8202 24596 8208 24608
rect 8067 24568 8208 24596
rect 8067 24565 8079 24568
rect 8021 24559 8079 24565
rect 8202 24556 8208 24568
rect 8260 24556 8266 24608
rect 10134 24596 10140 24608
rect 10095 24568 10140 24596
rect 10134 24556 10140 24568
rect 10192 24556 10198 24608
rect 12526 24556 12532 24608
rect 12584 24596 12590 24608
rect 15396 24605 15424 24636
rect 16482 24624 16488 24636
rect 16540 24624 16546 24676
rect 12805 24599 12863 24605
rect 12805 24596 12817 24599
rect 12584 24568 12817 24596
rect 12584 24556 12590 24568
rect 12805 24565 12817 24568
rect 12851 24565 12863 24599
rect 12805 24559 12863 24565
rect 15381 24599 15439 24605
rect 15381 24565 15393 24599
rect 15427 24565 15439 24599
rect 15381 24559 15439 24565
rect 15562 24556 15568 24608
rect 15620 24596 15626 24608
rect 15749 24599 15807 24605
rect 15749 24596 15761 24599
rect 15620 24568 15761 24596
rect 15620 24556 15626 24568
rect 15749 24565 15761 24568
rect 15795 24565 15807 24599
rect 15749 24559 15807 24565
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 4154 24352 4160 24404
rect 4212 24392 4218 24404
rect 4249 24395 4307 24401
rect 4249 24392 4261 24395
rect 4212 24364 4261 24392
rect 4212 24352 4218 24364
rect 4249 24361 4261 24364
rect 4295 24361 4307 24395
rect 4249 24355 4307 24361
rect 4706 24352 4712 24404
rect 4764 24392 4770 24404
rect 5537 24395 5595 24401
rect 5537 24392 5549 24395
rect 4764 24364 5549 24392
rect 4764 24352 4770 24364
rect 5537 24361 5549 24364
rect 5583 24361 5595 24395
rect 5994 24392 6000 24404
rect 5955 24364 6000 24392
rect 5537 24355 5595 24361
rect 5994 24352 6000 24364
rect 6052 24352 6058 24404
rect 7006 24392 7012 24404
rect 6967 24364 7012 24392
rect 7006 24352 7012 24364
rect 7064 24352 7070 24404
rect 8478 24392 8484 24404
rect 8439 24364 8484 24392
rect 8478 24352 8484 24364
rect 8536 24352 8542 24404
rect 15473 24395 15531 24401
rect 15473 24361 15485 24395
rect 15519 24392 15531 24395
rect 16206 24392 16212 24404
rect 15519 24364 16212 24392
rect 15519 24361 15531 24364
rect 15473 24355 15531 24361
rect 16206 24352 16212 24364
rect 16264 24352 16270 24404
rect 16577 24395 16635 24401
rect 16577 24361 16589 24395
rect 16623 24392 16635 24395
rect 17402 24392 17408 24404
rect 16623 24364 17408 24392
rect 16623 24361 16635 24364
rect 16577 24355 16635 24361
rect 17402 24352 17408 24364
rect 17460 24352 17466 24404
rect 17681 24395 17739 24401
rect 17681 24361 17693 24395
rect 17727 24392 17739 24395
rect 18506 24392 18512 24404
rect 17727 24364 18512 24392
rect 17727 24361 17739 24364
rect 17681 24355 17739 24361
rect 18506 24352 18512 24364
rect 18564 24352 18570 24404
rect 19058 24392 19064 24404
rect 19019 24364 19064 24392
rect 19058 24352 19064 24364
rect 19116 24352 19122 24404
rect 21085 24395 21143 24401
rect 21085 24361 21097 24395
rect 21131 24392 21143 24395
rect 22462 24392 22468 24404
rect 21131 24364 22468 24392
rect 21131 24361 21143 24364
rect 21085 24355 21143 24361
rect 22462 24352 22468 24364
rect 22520 24352 22526 24404
rect 1857 24327 1915 24333
rect 1857 24293 1869 24327
rect 1903 24324 1915 24327
rect 1903 24296 4108 24324
rect 1903 24293 1915 24296
rect 1857 24287 1915 24293
rect 4080 24268 4108 24296
rect 4430 24284 4436 24336
rect 4488 24324 4494 24336
rect 5077 24327 5135 24333
rect 5077 24324 5089 24327
rect 4488 24296 5089 24324
rect 4488 24284 4494 24296
rect 5077 24293 5089 24296
rect 5123 24324 5135 24327
rect 7834 24324 7840 24336
rect 5123 24296 6684 24324
rect 5123 24293 5135 24296
rect 5077 24287 5135 24293
rect 1581 24259 1639 24265
rect 1581 24225 1593 24259
rect 1627 24256 1639 24259
rect 2406 24256 2412 24268
rect 1627 24228 2412 24256
rect 1627 24225 1639 24228
rect 1581 24219 1639 24225
rect 2406 24216 2412 24228
rect 2464 24216 2470 24268
rect 2498 24216 2504 24268
rect 2556 24256 2562 24268
rect 2866 24256 2872 24268
rect 2556 24228 2872 24256
rect 2556 24216 2562 24228
rect 2866 24216 2872 24228
rect 2924 24216 2930 24268
rect 4062 24256 4068 24268
rect 4023 24228 4068 24256
rect 4062 24216 4068 24228
rect 4120 24216 4126 24268
rect 4522 24216 4528 24268
rect 4580 24256 4586 24268
rect 4709 24259 4767 24265
rect 4709 24256 4721 24259
rect 4580 24228 4721 24256
rect 4580 24216 4586 24228
rect 4709 24225 4721 24228
rect 4755 24256 4767 24259
rect 5350 24256 5356 24268
rect 4755 24228 5356 24256
rect 4755 24225 4767 24228
rect 4709 24219 4767 24225
rect 5350 24216 5356 24228
rect 5408 24216 5414 24268
rect 5905 24259 5963 24265
rect 5905 24225 5917 24259
rect 5951 24256 5963 24259
rect 6546 24256 6552 24268
rect 5951 24228 6552 24256
rect 5951 24225 5963 24228
rect 5905 24219 5963 24225
rect 6546 24216 6552 24228
rect 6604 24216 6610 24268
rect 6656 24265 6684 24296
rect 7116 24296 7840 24324
rect 7116 24265 7144 24296
rect 7834 24284 7840 24296
rect 7892 24284 7898 24336
rect 10413 24327 10471 24333
rect 10413 24293 10425 24327
rect 10459 24324 10471 24327
rect 10864 24327 10922 24333
rect 10864 24324 10876 24327
rect 10459 24296 10876 24324
rect 10459 24293 10471 24296
rect 10413 24287 10471 24293
rect 10864 24293 10876 24296
rect 10910 24324 10922 24327
rect 10962 24324 10968 24336
rect 10910 24296 10968 24324
rect 10910 24293 10922 24296
rect 10864 24287 10922 24293
rect 10962 24284 10968 24296
rect 11020 24284 11026 24336
rect 7374 24265 7380 24268
rect 6641 24259 6699 24265
rect 6641 24225 6653 24259
rect 6687 24256 6699 24259
rect 7101 24259 7159 24265
rect 7101 24256 7113 24259
rect 6687 24228 7113 24256
rect 6687 24225 6699 24228
rect 6641 24219 6699 24225
rect 7101 24225 7113 24228
rect 7147 24225 7159 24259
rect 7368 24256 7380 24265
rect 7335 24228 7380 24256
rect 7101 24219 7159 24225
rect 7368 24219 7380 24228
rect 7374 24216 7380 24219
rect 7432 24216 7438 24268
rect 10597 24259 10655 24265
rect 10597 24225 10609 24259
rect 10643 24256 10655 24259
rect 10686 24256 10692 24268
rect 10643 24228 10692 24256
rect 10643 24225 10655 24228
rect 10597 24219 10655 24225
rect 10686 24216 10692 24228
rect 10744 24216 10750 24268
rect 14182 24216 14188 24268
rect 14240 24256 14246 24268
rect 15289 24259 15347 24265
rect 15289 24256 15301 24259
rect 14240 24228 15301 24256
rect 14240 24216 14246 24228
rect 15289 24225 15301 24228
rect 15335 24225 15347 24259
rect 16390 24256 16396 24268
rect 16351 24228 16396 24256
rect 15289 24219 15347 24225
rect 16390 24216 16396 24228
rect 16448 24216 16454 24268
rect 17494 24256 17500 24268
rect 17455 24228 17500 24256
rect 17494 24216 17500 24228
rect 17552 24216 17558 24268
rect 18874 24256 18880 24268
rect 18835 24228 18880 24256
rect 18874 24216 18880 24228
rect 18932 24216 18938 24268
rect 20901 24259 20959 24265
rect 20901 24225 20913 24259
rect 20947 24256 20959 24259
rect 21174 24256 21180 24268
rect 20947 24228 21180 24256
rect 20947 24225 20959 24228
rect 20901 24219 20959 24225
rect 21174 24216 21180 24228
rect 21232 24216 21238 24268
rect 6181 24191 6239 24197
rect 6181 24157 6193 24191
rect 6227 24188 6239 24191
rect 6454 24188 6460 24200
rect 6227 24160 6460 24188
rect 6227 24157 6239 24160
rect 6181 24151 6239 24157
rect 6454 24148 6460 24160
rect 6512 24148 6518 24200
rect 13262 24188 13268 24200
rect 13223 24160 13268 24188
rect 13262 24148 13268 24160
rect 13320 24148 13326 24200
rect 3326 24120 3332 24132
rect 2884 24092 3332 24120
rect 2685 24055 2743 24061
rect 2685 24021 2697 24055
rect 2731 24052 2743 24055
rect 2884 24052 2912 24092
rect 3326 24080 3332 24092
rect 3384 24080 3390 24132
rect 2731 24024 2912 24052
rect 2731 24021 2743 24024
rect 2685 24015 2743 24021
rect 2958 24012 2964 24064
rect 3016 24052 3022 24064
rect 3053 24055 3111 24061
rect 3053 24052 3065 24055
rect 3016 24024 3065 24052
rect 3016 24012 3022 24024
rect 3053 24021 3065 24024
rect 3099 24021 3111 24055
rect 3053 24015 3111 24021
rect 3513 24055 3571 24061
rect 3513 24021 3525 24055
rect 3559 24052 3571 24055
rect 4430 24052 4436 24064
rect 3559 24024 4436 24052
rect 3559 24021 3571 24024
rect 3513 24015 3571 24021
rect 4430 24012 4436 24024
rect 4488 24012 4494 24064
rect 11974 24052 11980 24064
rect 11935 24024 11980 24052
rect 11974 24012 11980 24024
rect 12032 24012 12038 24064
rect 12526 24052 12532 24064
rect 12487 24024 12532 24052
rect 12526 24012 12532 24024
rect 12584 24012 12590 24064
rect 14642 24012 14648 24064
rect 14700 24052 14706 24064
rect 14921 24055 14979 24061
rect 14921 24052 14933 24055
rect 14700 24024 14933 24052
rect 14700 24012 14706 24024
rect 14921 24021 14933 24024
rect 14967 24021 14979 24055
rect 14921 24015 14979 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 2406 23808 2412 23860
rect 2464 23848 2470 23860
rect 2593 23851 2651 23857
rect 2593 23848 2605 23851
rect 2464 23820 2605 23848
rect 2464 23808 2470 23820
rect 2593 23817 2605 23820
rect 2639 23817 2651 23851
rect 2593 23811 2651 23817
rect 2866 23808 2872 23860
rect 2924 23848 2930 23860
rect 3605 23851 3663 23857
rect 3605 23848 3617 23851
rect 2924 23820 3617 23848
rect 2924 23808 2930 23820
rect 3605 23817 3617 23820
rect 3651 23817 3663 23851
rect 3605 23811 3663 23817
rect 5994 23808 6000 23860
rect 6052 23848 6058 23860
rect 6181 23851 6239 23857
rect 6181 23848 6193 23851
rect 6052 23820 6193 23848
rect 6052 23808 6058 23820
rect 6181 23817 6193 23820
rect 6227 23817 6239 23851
rect 6546 23848 6552 23860
rect 6507 23820 6552 23848
rect 6181 23811 6239 23817
rect 6546 23808 6552 23820
rect 6604 23808 6610 23860
rect 9214 23848 9220 23860
rect 9175 23820 9220 23848
rect 9214 23808 9220 23820
rect 9272 23808 9278 23860
rect 10962 23808 10968 23860
rect 11020 23848 11026 23860
rect 13817 23851 13875 23857
rect 13817 23848 13829 23851
rect 11020 23820 13829 23848
rect 11020 23808 11026 23820
rect 13817 23817 13829 23820
rect 13863 23817 13875 23851
rect 13817 23811 13875 23817
rect 18233 23851 18291 23857
rect 18233 23817 18245 23851
rect 18279 23848 18291 23851
rect 19150 23848 19156 23860
rect 18279 23820 19156 23848
rect 18279 23817 18291 23820
rect 18233 23811 18291 23817
rect 19150 23808 19156 23820
rect 19208 23808 19214 23860
rect 19337 23851 19395 23857
rect 19337 23817 19349 23851
rect 19383 23848 19395 23851
rect 20254 23848 20260 23860
rect 19383 23820 20260 23848
rect 19383 23817 19395 23820
rect 19337 23811 19395 23817
rect 20254 23808 20260 23820
rect 20312 23808 20318 23860
rect 20438 23848 20444 23860
rect 20399 23820 20444 23848
rect 20438 23808 20444 23820
rect 20496 23808 20502 23860
rect 21542 23848 21548 23860
rect 21503 23820 21548 23848
rect 21542 23808 21548 23820
rect 21600 23808 21606 23860
rect 22649 23851 22707 23857
rect 22649 23817 22661 23851
rect 22695 23848 22707 23851
rect 23382 23848 23388 23860
rect 22695 23820 23388 23848
rect 22695 23817 22707 23820
rect 22649 23811 22707 23817
rect 23382 23808 23388 23820
rect 23440 23808 23446 23860
rect 10689 23783 10747 23789
rect 10689 23749 10701 23783
rect 10735 23780 10747 23783
rect 12250 23780 12256 23792
rect 10735 23752 12256 23780
rect 10735 23749 10747 23752
rect 10689 23743 10747 23749
rect 3234 23712 3240 23724
rect 3195 23684 3240 23712
rect 3234 23672 3240 23684
rect 3292 23672 3298 23724
rect 4157 23715 4215 23721
rect 4157 23681 4169 23715
rect 4203 23712 4215 23715
rect 7834 23712 7840 23724
rect 4203 23684 4384 23712
rect 7795 23684 7840 23712
rect 4203 23681 4215 23684
rect 4157 23675 4215 23681
rect 1397 23647 1455 23653
rect 1397 23613 1409 23647
rect 1443 23613 1455 23647
rect 1397 23607 1455 23613
rect 4249 23647 4307 23653
rect 4249 23613 4261 23647
rect 4295 23613 4307 23647
rect 4356 23644 4384 23684
rect 7834 23672 7840 23684
rect 7892 23672 7898 23724
rect 11256 23721 11284 23752
rect 12250 23740 12256 23752
rect 12308 23740 12314 23792
rect 11241 23715 11299 23721
rect 11241 23681 11253 23715
rect 11287 23681 11299 23715
rect 11422 23712 11428 23724
rect 11335 23684 11428 23712
rect 11241 23675 11299 23681
rect 11422 23672 11428 23684
rect 11480 23712 11486 23724
rect 11974 23712 11980 23724
rect 11480 23684 11980 23712
rect 11480 23672 11486 23684
rect 11974 23672 11980 23684
rect 12032 23672 12038 23724
rect 14642 23672 14648 23724
rect 14700 23712 14706 23724
rect 14921 23715 14979 23721
rect 14921 23712 14933 23715
rect 14700 23684 14933 23712
rect 14700 23672 14706 23684
rect 14921 23681 14933 23684
rect 14967 23681 14979 23715
rect 14921 23675 14979 23681
rect 18322 23672 18328 23724
rect 18380 23712 18386 23724
rect 18380 23684 19196 23712
rect 18380 23672 18386 23684
rect 4522 23653 4528 23656
rect 4516 23644 4528 23653
rect 4356 23616 4528 23644
rect 4249 23607 4307 23613
rect 4516 23607 4528 23616
rect 1412 23576 1440 23607
rect 2038 23576 2044 23588
rect 1412 23548 2044 23576
rect 2038 23536 2044 23548
rect 2096 23536 2102 23588
rect 3053 23579 3111 23585
rect 3053 23545 3065 23579
rect 3099 23576 3111 23579
rect 3326 23576 3332 23588
rect 3099 23548 3332 23576
rect 3099 23545 3111 23548
rect 3053 23539 3111 23545
rect 3326 23536 3332 23548
rect 3384 23576 3390 23588
rect 4062 23576 4068 23588
rect 3384 23548 4068 23576
rect 3384 23536 3390 23548
rect 4062 23536 4068 23548
rect 4120 23536 4126 23588
rect 4264 23576 4292 23607
rect 4522 23604 4528 23607
rect 4580 23604 4586 23656
rect 9953 23647 10011 23653
rect 9953 23613 9965 23647
rect 9999 23644 10011 23647
rect 11440 23644 11468 23672
rect 12434 23644 12440 23656
rect 9999 23616 11468 23644
rect 12395 23616 12440 23644
rect 9999 23613 10011 23616
rect 9953 23607 10011 23613
rect 12434 23604 12440 23616
rect 12492 23604 12498 23656
rect 13814 23604 13820 23656
rect 13872 23644 13878 23656
rect 14737 23647 14795 23653
rect 14737 23644 14749 23647
rect 13872 23616 14749 23644
rect 13872 23604 13878 23616
rect 14737 23613 14749 23616
rect 14783 23613 14795 23647
rect 14737 23607 14795 23613
rect 4430 23576 4436 23588
rect 4264 23548 4436 23576
rect 4430 23536 4436 23548
rect 4488 23536 4494 23588
rect 6454 23536 6460 23588
rect 6512 23576 6518 23588
rect 8110 23585 8116 23588
rect 7745 23579 7803 23585
rect 6512 23548 7420 23576
rect 6512 23536 6518 23548
rect 7392 23520 7420 23548
rect 7745 23545 7757 23579
rect 7791 23576 7803 23579
rect 8082 23579 8116 23585
rect 8082 23576 8094 23579
rect 7791 23548 8094 23576
rect 7791 23545 7803 23548
rect 7745 23539 7803 23545
rect 8082 23545 8094 23548
rect 8168 23576 8174 23588
rect 11149 23579 11207 23585
rect 11149 23576 11161 23579
rect 8168 23548 8230 23576
rect 10244 23548 11161 23576
rect 8082 23539 8116 23545
rect 8110 23536 8116 23539
rect 8168 23536 8174 23548
rect 1394 23468 1400 23520
rect 1452 23508 1458 23520
rect 1581 23511 1639 23517
rect 1581 23508 1593 23511
rect 1452 23480 1593 23508
rect 1452 23468 1458 23480
rect 1581 23477 1593 23480
rect 1627 23477 1639 23511
rect 1581 23471 1639 23477
rect 2501 23511 2559 23517
rect 2501 23477 2513 23511
rect 2547 23508 2559 23511
rect 2961 23511 3019 23517
rect 2961 23508 2973 23511
rect 2547 23480 2973 23508
rect 2547 23477 2559 23480
rect 2501 23471 2559 23477
rect 2961 23477 2973 23480
rect 3007 23508 3019 23511
rect 3418 23508 3424 23520
rect 3007 23480 3424 23508
rect 3007 23477 3019 23480
rect 2961 23471 3019 23477
rect 3418 23468 3424 23480
rect 3476 23468 3482 23520
rect 5534 23468 5540 23520
rect 5592 23508 5598 23520
rect 5629 23511 5687 23517
rect 5629 23508 5641 23511
rect 5592 23480 5641 23508
rect 5592 23468 5598 23480
rect 5629 23477 5641 23480
rect 5675 23477 5687 23511
rect 6822 23508 6828 23520
rect 6783 23480 6828 23508
rect 5629 23471 5687 23477
rect 6822 23468 6828 23480
rect 6880 23468 6886 23520
rect 7374 23508 7380 23520
rect 7287 23480 7380 23508
rect 7374 23468 7380 23480
rect 7432 23508 7438 23520
rect 8294 23508 8300 23520
rect 7432 23480 8300 23508
rect 7432 23468 7438 23480
rect 8294 23468 8300 23480
rect 8352 23468 8358 23520
rect 10042 23468 10048 23520
rect 10100 23508 10106 23520
rect 10244 23517 10272 23548
rect 11149 23545 11161 23548
rect 11195 23545 11207 23579
rect 11149 23539 11207 23545
rect 11885 23579 11943 23585
rect 11885 23545 11897 23579
rect 11931 23576 11943 23579
rect 12253 23579 12311 23585
rect 11931 23548 12112 23576
rect 11931 23545 11943 23548
rect 11885 23539 11943 23545
rect 10229 23511 10287 23517
rect 10229 23508 10241 23511
rect 10100 23480 10241 23508
rect 10100 23468 10106 23480
rect 10229 23477 10241 23480
rect 10275 23477 10287 23511
rect 10778 23508 10784 23520
rect 10739 23480 10784 23508
rect 10229 23471 10287 23477
rect 10778 23468 10784 23480
rect 10836 23468 10842 23520
rect 11164 23508 11192 23539
rect 11974 23508 11980 23520
rect 11164 23480 11980 23508
rect 11974 23468 11980 23480
rect 12032 23468 12038 23520
rect 12084 23508 12112 23548
rect 12253 23545 12265 23579
rect 12299 23576 12311 23579
rect 12704 23579 12762 23585
rect 12704 23576 12716 23579
rect 12299 23548 12716 23576
rect 12299 23545 12311 23548
rect 12253 23539 12311 23545
rect 12704 23545 12716 23548
rect 12750 23576 12762 23579
rect 13078 23576 13084 23588
rect 12750 23548 13084 23576
rect 12750 23545 12762 23548
rect 12704 23539 12762 23545
rect 13078 23536 13084 23548
rect 13136 23576 13142 23588
rect 14752 23576 14780 23607
rect 17954 23604 17960 23656
rect 18012 23644 18018 23656
rect 19168 23653 19196 23684
rect 18049 23647 18107 23653
rect 18049 23644 18061 23647
rect 18012 23616 18061 23644
rect 18012 23604 18018 23616
rect 18049 23613 18061 23616
rect 18095 23644 18107 23647
rect 18601 23647 18659 23653
rect 18601 23644 18613 23647
rect 18095 23616 18613 23644
rect 18095 23613 18107 23616
rect 18049 23607 18107 23613
rect 18601 23613 18613 23616
rect 18647 23613 18659 23647
rect 18601 23607 18659 23613
rect 19153 23647 19211 23653
rect 19153 23613 19165 23647
rect 19199 23644 19211 23647
rect 19705 23647 19763 23653
rect 19705 23644 19717 23647
rect 19199 23616 19717 23644
rect 19199 23613 19211 23616
rect 19153 23607 19211 23613
rect 19705 23613 19717 23616
rect 19751 23613 19763 23647
rect 19705 23607 19763 23613
rect 19978 23604 19984 23656
rect 20036 23644 20042 23656
rect 20257 23647 20315 23653
rect 20257 23644 20269 23647
rect 20036 23616 20269 23644
rect 20036 23604 20042 23616
rect 20257 23613 20269 23616
rect 20303 23644 20315 23647
rect 20809 23647 20867 23653
rect 20809 23644 20821 23647
rect 20303 23616 20821 23644
rect 20303 23613 20315 23616
rect 20257 23607 20315 23613
rect 20809 23613 20821 23616
rect 20855 23613 20867 23647
rect 20809 23607 20867 23613
rect 20990 23604 20996 23656
rect 21048 23644 21054 23656
rect 21361 23647 21419 23653
rect 21361 23644 21373 23647
rect 21048 23616 21373 23644
rect 21048 23604 21054 23616
rect 21361 23613 21373 23616
rect 21407 23644 21419 23647
rect 21913 23647 21971 23653
rect 21913 23644 21925 23647
rect 21407 23616 21925 23644
rect 21407 23613 21419 23616
rect 21361 23607 21419 23613
rect 21913 23613 21925 23616
rect 21959 23613 21971 23647
rect 21913 23607 21971 23613
rect 22094 23604 22100 23656
rect 22152 23644 22158 23656
rect 22465 23647 22523 23653
rect 22465 23644 22477 23647
rect 22152 23616 22477 23644
rect 22152 23604 22158 23616
rect 22465 23613 22477 23616
rect 22511 23644 22523 23647
rect 23017 23647 23075 23653
rect 23017 23644 23029 23647
rect 22511 23616 23029 23644
rect 22511 23613 22523 23616
rect 22465 23607 22523 23613
rect 23017 23613 23029 23616
rect 23063 23613 23075 23647
rect 23017 23607 23075 23613
rect 15166 23579 15224 23585
rect 15166 23576 15178 23579
rect 13136 23548 14596 23576
rect 14752 23548 15178 23576
rect 13136 23536 13142 23548
rect 12434 23508 12440 23520
rect 12084 23480 12440 23508
rect 12434 23468 12440 23480
rect 12492 23468 12498 23520
rect 14182 23468 14188 23520
rect 14240 23508 14246 23520
rect 14369 23511 14427 23517
rect 14369 23508 14381 23511
rect 14240 23480 14381 23508
rect 14240 23468 14246 23480
rect 14369 23477 14381 23480
rect 14415 23477 14427 23511
rect 14568 23508 14596 23548
rect 15166 23545 15178 23548
rect 15212 23576 15224 23579
rect 15470 23576 15476 23588
rect 15212 23548 15476 23576
rect 15212 23545 15224 23548
rect 15166 23539 15224 23545
rect 15470 23536 15476 23548
rect 15528 23536 15534 23588
rect 18138 23536 18144 23588
rect 18196 23576 18202 23588
rect 18874 23576 18880 23588
rect 18196 23548 18880 23576
rect 18196 23536 18202 23548
rect 18874 23536 18880 23548
rect 18932 23576 18938 23588
rect 18969 23579 19027 23585
rect 18969 23576 18981 23579
rect 18932 23548 18981 23576
rect 18932 23536 18938 23548
rect 18969 23545 18981 23548
rect 19015 23545 19027 23579
rect 18969 23539 19027 23545
rect 16301 23511 16359 23517
rect 16301 23508 16313 23511
rect 14568 23480 16313 23508
rect 14369 23471 14427 23477
rect 16301 23477 16313 23480
rect 16347 23477 16359 23511
rect 16301 23471 16359 23477
rect 16390 23468 16396 23520
rect 16448 23508 16454 23520
rect 16853 23511 16911 23517
rect 16853 23508 16865 23511
rect 16448 23480 16865 23508
rect 16448 23468 16454 23480
rect 16853 23477 16865 23480
rect 16899 23477 16911 23511
rect 17494 23508 17500 23520
rect 17455 23480 17500 23508
rect 16853 23471 16911 23477
rect 17494 23468 17500 23480
rect 17552 23468 17558 23520
rect 21174 23508 21180 23520
rect 21135 23480 21180 23508
rect 21174 23468 21180 23480
rect 21232 23468 21238 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 4154 23264 4160 23316
rect 4212 23304 4218 23316
rect 4249 23307 4307 23313
rect 4249 23304 4261 23307
rect 4212 23276 4261 23304
rect 4212 23264 4218 23276
rect 4249 23273 4261 23276
rect 4295 23273 4307 23307
rect 5810 23304 5816 23316
rect 5771 23276 5816 23304
rect 4249 23267 4307 23273
rect 5810 23264 5816 23276
rect 5868 23264 5874 23316
rect 6454 23304 6460 23316
rect 6415 23276 6460 23304
rect 6454 23264 6460 23276
rect 6512 23264 6518 23316
rect 7009 23307 7067 23313
rect 7009 23273 7021 23307
rect 7055 23304 7067 23307
rect 7834 23304 7840 23316
rect 7055 23276 7840 23304
rect 7055 23273 7067 23276
rect 7009 23267 7067 23273
rect 7834 23264 7840 23276
rect 7892 23264 7898 23316
rect 8294 23264 8300 23316
rect 8352 23304 8358 23316
rect 8481 23307 8539 23313
rect 8481 23304 8493 23307
rect 8352 23276 8493 23304
rect 8352 23264 8358 23276
rect 8481 23273 8493 23276
rect 8527 23273 8539 23307
rect 8481 23267 8539 23273
rect 9769 23307 9827 23313
rect 9769 23273 9781 23307
rect 9815 23304 9827 23307
rect 10134 23304 10140 23316
rect 9815 23276 10140 23304
rect 9815 23273 9827 23276
rect 9769 23267 9827 23273
rect 10134 23264 10140 23276
rect 10192 23264 10198 23316
rect 10689 23307 10747 23313
rect 10689 23273 10701 23307
rect 10735 23304 10747 23307
rect 10962 23304 10968 23316
rect 10735 23276 10968 23304
rect 10735 23273 10747 23276
rect 10689 23267 10747 23273
rect 10962 23264 10968 23276
rect 11020 23264 11026 23316
rect 13262 23264 13268 23316
rect 13320 23304 13326 23316
rect 13633 23307 13691 23313
rect 13633 23304 13645 23307
rect 13320 23276 13645 23304
rect 13320 23264 13326 23276
rect 13633 23273 13645 23276
rect 13679 23273 13691 23307
rect 13633 23267 13691 23273
rect 16761 23307 16819 23313
rect 16761 23273 16773 23307
rect 16807 23304 16819 23307
rect 17862 23304 17868 23316
rect 16807 23276 17868 23304
rect 16807 23273 16819 23276
rect 16761 23267 16819 23273
rect 17862 23264 17868 23276
rect 17920 23264 17926 23316
rect 19613 23307 19671 23313
rect 19613 23273 19625 23307
rect 19659 23304 19671 23307
rect 20070 23304 20076 23316
rect 19659 23276 20076 23304
rect 19659 23273 19671 23276
rect 19613 23267 19671 23273
rect 20070 23264 20076 23276
rect 20128 23264 20134 23316
rect 1857 23239 1915 23245
rect 1857 23205 1869 23239
rect 1903 23236 1915 23239
rect 2590 23236 2596 23248
rect 1903 23208 2596 23236
rect 1903 23205 1915 23208
rect 1857 23199 1915 23205
rect 2590 23196 2596 23208
rect 2648 23196 2654 23248
rect 4700 23239 4758 23245
rect 4700 23205 4712 23239
rect 4746 23236 4758 23239
rect 4982 23236 4988 23248
rect 4746 23208 4988 23236
rect 4746 23205 4758 23208
rect 4700 23199 4758 23205
rect 4982 23196 4988 23208
rect 5040 23236 5046 23248
rect 5442 23236 5448 23248
rect 5040 23208 5448 23236
rect 5040 23196 5046 23208
rect 5442 23196 5448 23208
rect 5500 23196 5506 23248
rect 11048 23239 11106 23245
rect 11048 23205 11060 23239
rect 11094 23236 11106 23239
rect 11422 23236 11428 23248
rect 11094 23208 11428 23236
rect 11094 23205 11106 23208
rect 11048 23199 11106 23205
rect 11422 23196 11428 23208
rect 11480 23196 11486 23248
rect 15565 23239 15623 23245
rect 15565 23205 15577 23239
rect 15611 23236 15623 23239
rect 16390 23236 16396 23248
rect 15611 23208 16396 23236
rect 15611 23205 15623 23208
rect 15565 23199 15623 23205
rect 16390 23196 16396 23208
rect 16448 23196 16454 23248
rect 21177 23239 21235 23245
rect 21177 23205 21189 23239
rect 21223 23236 21235 23239
rect 22002 23236 22008 23248
rect 21223 23208 22008 23236
rect 21223 23205 21235 23208
rect 21177 23199 21235 23205
rect 22002 23196 22008 23208
rect 22060 23196 22066 23248
rect 1581 23171 1639 23177
rect 1581 23137 1593 23171
rect 1627 23168 1639 23171
rect 1627 23140 2360 23168
rect 1627 23137 1639 23140
rect 1581 23131 1639 23137
rect 2332 23100 2360 23140
rect 2406 23128 2412 23180
rect 2464 23168 2470 23180
rect 2869 23171 2927 23177
rect 2869 23168 2881 23171
rect 2464 23140 2881 23168
rect 2464 23128 2470 23140
rect 2869 23137 2881 23140
rect 2915 23137 2927 23171
rect 3878 23168 3884 23180
rect 3791 23140 3884 23168
rect 2869 23131 2927 23137
rect 3878 23128 3884 23140
rect 3936 23168 3942 23180
rect 4430 23168 4436 23180
rect 3936 23140 4436 23168
rect 3936 23128 3942 23140
rect 4430 23128 4436 23140
rect 4488 23128 4494 23180
rect 6270 23128 6276 23180
rect 6328 23168 6334 23180
rect 7357 23171 7415 23177
rect 7357 23168 7369 23171
rect 6328 23140 7369 23168
rect 6328 23128 6334 23140
rect 7357 23137 7369 23140
rect 7403 23137 7415 23171
rect 7357 23131 7415 23137
rect 12434 23128 12440 23180
rect 12492 23168 12498 23180
rect 12805 23171 12863 23177
rect 12805 23168 12817 23171
rect 12492 23140 12817 23168
rect 12492 23128 12498 23140
rect 12805 23137 12817 23140
rect 12851 23168 12863 23171
rect 14550 23168 14556 23180
rect 12851 23140 14556 23168
rect 12851 23137 12863 23140
rect 12805 23131 12863 23137
rect 14550 23128 14556 23140
rect 14608 23128 14614 23180
rect 15289 23171 15347 23177
rect 15289 23137 15301 23171
rect 15335 23168 15347 23171
rect 16022 23168 16028 23180
rect 15335 23140 16028 23168
rect 15335 23137 15347 23140
rect 15289 23131 15347 23137
rect 16022 23128 16028 23140
rect 16080 23128 16086 23180
rect 16574 23128 16580 23180
rect 16632 23168 16638 23180
rect 17678 23168 17684 23180
rect 16632 23140 16677 23168
rect 17639 23140 17684 23168
rect 16632 23128 16638 23140
rect 17678 23128 17684 23140
rect 17736 23128 17742 23180
rect 19426 23168 19432 23180
rect 19387 23140 19432 23168
rect 19426 23128 19432 23140
rect 19484 23128 19490 23180
rect 20806 23128 20812 23180
rect 20864 23168 20870 23180
rect 20901 23171 20959 23177
rect 20901 23168 20913 23171
rect 20864 23140 20913 23168
rect 20864 23128 20870 23140
rect 20901 23137 20913 23140
rect 20947 23137 20959 23171
rect 20901 23131 20959 23137
rect 2774 23100 2780 23112
rect 2332 23072 2780 23100
rect 2774 23060 2780 23072
rect 2832 23060 2838 23112
rect 7006 23100 7012 23112
rect 6919 23072 7012 23100
rect 7006 23060 7012 23072
rect 7064 23100 7070 23112
rect 7101 23103 7159 23109
rect 7101 23100 7113 23103
rect 7064 23072 7113 23100
rect 7064 23060 7070 23072
rect 7101 23069 7113 23072
rect 7147 23069 7159 23103
rect 7101 23063 7159 23069
rect 9493 23103 9551 23109
rect 9493 23069 9505 23103
rect 9539 23100 9551 23103
rect 10321 23103 10379 23109
rect 10321 23100 10333 23103
rect 9539 23072 10333 23100
rect 9539 23069 9551 23072
rect 9493 23063 9551 23069
rect 10321 23069 10333 23072
rect 10367 23100 10379 23103
rect 10686 23100 10692 23112
rect 10367 23072 10692 23100
rect 10367 23069 10379 23072
rect 10321 23063 10379 23069
rect 10686 23060 10692 23072
rect 10744 23100 10750 23112
rect 10781 23103 10839 23109
rect 10781 23100 10793 23103
rect 10744 23072 10793 23100
rect 10744 23060 10750 23072
rect 10781 23069 10793 23072
rect 10827 23069 10839 23103
rect 13722 23100 13728 23112
rect 13683 23072 13728 23100
rect 10781 23063 10839 23069
rect 13722 23060 13728 23072
rect 13780 23060 13786 23112
rect 13817 23103 13875 23109
rect 13817 23069 13829 23103
rect 13863 23069 13875 23103
rect 13817 23063 13875 23069
rect 2685 23035 2743 23041
rect 2685 23001 2697 23035
rect 2731 23032 2743 23035
rect 3234 23032 3240 23044
rect 2731 23004 3240 23032
rect 2731 23001 2743 23004
rect 2685 22995 2743 23001
rect 3234 22992 3240 23004
rect 3292 22992 3298 23044
rect 13630 22992 13636 23044
rect 13688 23032 13694 23044
rect 13832 23032 13860 23063
rect 13688 23004 13860 23032
rect 13688 22992 13694 23004
rect 17770 22992 17776 23044
rect 17828 23032 17834 23044
rect 17865 23035 17923 23041
rect 17865 23032 17877 23035
rect 17828 23004 17877 23032
rect 17828 22992 17834 23004
rect 17865 23001 17877 23004
rect 17911 23001 17923 23035
rect 17865 22995 17923 23001
rect 3050 22964 3056 22976
rect 3011 22936 3056 22964
rect 3050 22924 3056 22936
rect 3108 22924 3114 22976
rect 3510 22964 3516 22976
rect 3471 22936 3516 22964
rect 3510 22924 3516 22936
rect 3568 22924 3574 22976
rect 6917 22967 6975 22973
rect 6917 22933 6929 22967
rect 6963 22964 6975 22967
rect 7282 22964 7288 22976
rect 6963 22936 7288 22964
rect 6963 22933 6975 22936
rect 6917 22927 6975 22933
rect 7282 22924 7288 22936
rect 7340 22924 7346 22976
rect 10962 22924 10968 22976
rect 11020 22964 11026 22976
rect 12161 22967 12219 22973
rect 12161 22964 12173 22967
rect 11020 22936 12173 22964
rect 11020 22924 11026 22936
rect 12161 22933 12173 22936
rect 12207 22933 12219 22967
rect 12161 22927 12219 22933
rect 12894 22924 12900 22976
rect 12952 22964 12958 22976
rect 13265 22967 13323 22973
rect 13265 22964 13277 22967
rect 12952 22936 13277 22964
rect 12952 22924 12958 22936
rect 13265 22933 13277 22936
rect 13311 22933 13323 22967
rect 13265 22927 13323 22933
rect 14090 22924 14096 22976
rect 14148 22964 14154 22976
rect 14277 22967 14335 22973
rect 14277 22964 14289 22967
rect 14148 22936 14289 22964
rect 14148 22924 14154 22936
rect 14277 22933 14289 22936
rect 14323 22933 14335 22967
rect 14277 22927 14335 22933
rect 14550 22924 14556 22976
rect 14608 22964 14614 22976
rect 14645 22967 14703 22973
rect 14645 22964 14657 22967
rect 14608 22936 14657 22964
rect 14608 22924 14614 22936
rect 14645 22933 14657 22936
rect 14691 22933 14703 22967
rect 14645 22927 14703 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 4982 22760 4988 22772
rect 4943 22732 4988 22760
rect 4982 22720 4988 22732
rect 5040 22720 5046 22772
rect 5534 22720 5540 22772
rect 5592 22760 5598 22772
rect 5629 22763 5687 22769
rect 5629 22760 5641 22763
rect 5592 22732 5641 22760
rect 5592 22720 5598 22732
rect 5629 22729 5641 22732
rect 5675 22729 5687 22763
rect 6270 22760 6276 22772
rect 6231 22732 6276 22760
rect 5629 22723 5687 22729
rect 6270 22720 6276 22732
rect 6328 22720 6334 22772
rect 6641 22763 6699 22769
rect 6641 22729 6653 22763
rect 6687 22760 6699 22763
rect 6822 22760 6828 22772
rect 6687 22732 6828 22760
rect 6687 22729 6699 22732
rect 6641 22723 6699 22729
rect 6822 22720 6828 22732
rect 6880 22720 6886 22772
rect 8202 22720 8208 22772
rect 8260 22760 8266 22772
rect 8389 22763 8447 22769
rect 8389 22760 8401 22763
rect 8260 22732 8401 22760
rect 8260 22720 8266 22732
rect 8389 22729 8401 22732
rect 8435 22729 8447 22763
rect 11422 22760 11428 22772
rect 11383 22732 11428 22760
rect 8389 22723 8447 22729
rect 11422 22720 11428 22732
rect 11480 22720 11486 22772
rect 13262 22760 13268 22772
rect 13223 22732 13268 22760
rect 13262 22720 13268 22732
rect 13320 22720 13326 22772
rect 13630 22760 13636 22772
rect 13591 22732 13636 22760
rect 13630 22720 13636 22732
rect 13688 22720 13694 22772
rect 15470 22760 15476 22772
rect 15431 22732 15476 22760
rect 15470 22720 15476 22732
rect 15528 22720 15534 22772
rect 9950 22652 9956 22704
rect 10008 22692 10014 22704
rect 10321 22695 10379 22701
rect 10321 22692 10333 22695
rect 10008 22664 10333 22692
rect 10008 22652 10014 22664
rect 10321 22661 10333 22664
rect 10367 22661 10379 22695
rect 11701 22695 11759 22701
rect 11701 22692 11713 22695
rect 10321 22655 10379 22661
rect 10796 22664 11713 22692
rect 10796 22636 10824 22664
rect 11701 22661 11713 22664
rect 11747 22661 11759 22695
rect 11701 22655 11759 22661
rect 1765 22627 1823 22633
rect 1765 22593 1777 22627
rect 1811 22624 1823 22627
rect 2682 22624 2688 22636
rect 1811 22596 2688 22624
rect 1811 22593 1823 22596
rect 1765 22587 1823 22593
rect 2682 22584 2688 22596
rect 2740 22584 2746 22636
rect 2869 22627 2927 22633
rect 2869 22593 2881 22627
rect 2915 22624 2927 22627
rect 7374 22624 7380 22636
rect 2915 22596 3096 22624
rect 7335 22596 7380 22624
rect 2915 22593 2927 22596
rect 2869 22587 2927 22593
rect 1489 22559 1547 22565
rect 1489 22525 1501 22559
rect 1535 22525 1547 22559
rect 1489 22519 1547 22525
rect 2961 22559 3019 22565
rect 2961 22525 2973 22559
rect 3007 22525 3019 22559
rect 3068 22556 3096 22596
rect 7374 22584 7380 22596
rect 7432 22584 7438 22636
rect 8297 22627 8355 22633
rect 8297 22593 8309 22627
rect 8343 22624 8355 22627
rect 8846 22624 8852 22636
rect 8343 22596 8852 22624
rect 8343 22593 8355 22596
rect 8297 22587 8355 22593
rect 8846 22584 8852 22596
rect 8904 22584 8910 22636
rect 8938 22584 8944 22636
rect 8996 22624 9002 22636
rect 9401 22627 9459 22633
rect 9401 22624 9413 22627
rect 8996 22596 9413 22624
rect 8996 22584 9002 22596
rect 9401 22593 9413 22596
rect 9447 22593 9459 22627
rect 10778 22624 10784 22636
rect 10739 22596 10784 22624
rect 9401 22587 9459 22593
rect 10778 22584 10784 22596
rect 10836 22584 10842 22636
rect 10962 22624 10968 22636
rect 10923 22596 10968 22624
rect 10962 22584 10968 22596
rect 11020 22584 11026 22636
rect 12710 22624 12716 22636
rect 12671 22596 12716 22624
rect 12710 22584 12716 22596
rect 12768 22584 12774 22636
rect 3234 22565 3240 22568
rect 3228 22556 3240 22565
rect 3068 22528 3240 22556
rect 2961 22519 3019 22525
rect 3228 22519 3240 22528
rect 1504 22488 1532 22519
rect 2682 22488 2688 22500
rect 1504 22460 2688 22488
rect 2682 22448 2688 22460
rect 2740 22448 2746 22500
rect 2976 22488 3004 22519
rect 3234 22516 3240 22519
rect 3292 22516 3298 22568
rect 5445 22559 5503 22565
rect 5445 22556 5457 22559
rect 5276 22528 5457 22556
rect 3878 22488 3884 22500
rect 2976 22460 3884 22488
rect 3878 22448 3884 22460
rect 3936 22448 3942 22500
rect 5276 22432 5304 22528
rect 5445 22525 5457 22528
rect 5491 22525 5503 22559
rect 5445 22519 5503 22525
rect 6822 22516 6828 22568
rect 6880 22516 6886 22568
rect 7282 22556 7288 22568
rect 7243 22528 7288 22556
rect 7282 22516 7288 22528
rect 7340 22516 7346 22568
rect 9861 22559 9919 22565
rect 9861 22525 9873 22559
rect 9907 22556 9919 22559
rect 10980 22556 11008 22584
rect 9907 22528 11008 22556
rect 12253 22559 12311 22565
rect 9907 22525 9919 22528
rect 9861 22519 9919 22525
rect 12253 22525 12265 22559
rect 12299 22556 12311 22559
rect 12529 22559 12587 22565
rect 12529 22556 12541 22559
rect 12299 22528 12541 22556
rect 12299 22525 12311 22528
rect 12253 22519 12311 22525
rect 12529 22525 12541 22528
rect 12575 22556 12587 22559
rect 12894 22556 12900 22568
rect 12575 22528 12900 22556
rect 12575 22525 12587 22528
rect 12529 22519 12587 22525
rect 12894 22516 12900 22528
rect 12952 22516 12958 22568
rect 14093 22559 14151 22565
rect 14093 22525 14105 22559
rect 14139 22556 14151 22559
rect 14139 22528 14596 22556
rect 14139 22525 14151 22528
rect 14093 22519 14151 22525
rect 6840 22488 6868 22516
rect 14568 22500 14596 22528
rect 7193 22491 7251 22497
rect 7193 22488 7205 22491
rect 6840 22460 7205 22488
rect 7193 22457 7205 22460
rect 7239 22457 7251 22491
rect 14338 22491 14396 22497
rect 14338 22488 14350 22491
rect 7193 22451 7251 22457
rect 14108 22460 14350 22488
rect 14108 22432 14136 22460
rect 14338 22457 14350 22460
rect 14384 22457 14396 22491
rect 14338 22451 14396 22457
rect 14550 22448 14556 22500
rect 14608 22448 14614 22500
rect 2406 22420 2412 22432
rect 2367 22392 2412 22420
rect 2406 22380 2412 22392
rect 2464 22380 2470 22432
rect 4246 22380 4252 22432
rect 4304 22420 4310 22432
rect 4341 22423 4399 22429
rect 4341 22420 4353 22423
rect 4304 22392 4353 22420
rect 4304 22380 4310 22392
rect 4341 22389 4353 22392
rect 4387 22389 4399 22423
rect 5258 22420 5264 22432
rect 5219 22392 5264 22420
rect 4341 22383 4399 22389
rect 5258 22380 5264 22392
rect 5316 22380 5322 22432
rect 6822 22420 6828 22432
rect 6783 22392 6828 22420
rect 6822 22380 6828 22392
rect 6880 22380 6886 22432
rect 7929 22423 7987 22429
rect 7929 22389 7941 22423
rect 7975 22420 7987 22423
rect 8754 22420 8760 22432
rect 7975 22392 8760 22420
rect 7975 22389 7987 22392
rect 7929 22383 7987 22389
rect 8754 22380 8760 22392
rect 8812 22380 8818 22432
rect 9674 22380 9680 22432
rect 9732 22420 9738 22432
rect 10137 22423 10195 22429
rect 10137 22420 10149 22423
rect 9732 22392 10149 22420
rect 9732 22380 9738 22392
rect 10137 22389 10149 22392
rect 10183 22420 10195 22423
rect 10689 22423 10747 22429
rect 10689 22420 10701 22423
rect 10183 22392 10701 22420
rect 10183 22389 10195 22392
rect 10137 22383 10195 22389
rect 10689 22389 10701 22392
rect 10735 22389 10747 22423
rect 10689 22383 10747 22389
rect 14090 22380 14096 22432
rect 14148 22380 14154 22432
rect 16022 22420 16028 22432
rect 15983 22392 16028 22420
rect 16022 22380 16028 22392
rect 16080 22380 16086 22432
rect 16574 22380 16580 22432
rect 16632 22420 16638 22432
rect 16632 22392 16677 22420
rect 16632 22380 16638 22392
rect 16850 22380 16856 22432
rect 16908 22420 16914 22432
rect 17678 22420 17684 22432
rect 16908 22392 17684 22420
rect 16908 22380 16914 22392
rect 17678 22380 17684 22392
rect 17736 22380 17742 22432
rect 19426 22420 19432 22432
rect 19387 22392 19432 22420
rect 19426 22380 19432 22392
rect 19484 22380 19490 22432
rect 20806 22380 20812 22432
rect 20864 22420 20870 22432
rect 20901 22423 20959 22429
rect 20901 22420 20913 22423
rect 20864 22392 20913 22420
rect 20864 22380 20870 22392
rect 20901 22389 20913 22392
rect 20947 22389 20959 22423
rect 20901 22383 20959 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 2409 22219 2467 22225
rect 2409 22185 2421 22219
rect 2455 22216 2467 22219
rect 2682 22216 2688 22228
rect 2455 22188 2688 22216
rect 2455 22185 2467 22188
rect 2409 22179 2467 22185
rect 2682 22176 2688 22188
rect 2740 22176 2746 22228
rect 3510 22176 3516 22228
rect 3568 22216 3574 22228
rect 3789 22219 3847 22225
rect 3789 22216 3801 22219
rect 3568 22188 3801 22216
rect 3568 22176 3574 22188
rect 3789 22185 3801 22188
rect 3835 22185 3847 22219
rect 3789 22179 3847 22185
rect 1397 22083 1455 22089
rect 1397 22049 1409 22083
rect 1443 22049 1455 22083
rect 2038 22080 2044 22092
rect 1999 22052 2044 22080
rect 1397 22043 1455 22049
rect 1412 22012 1440 22043
rect 2038 22040 2044 22052
rect 2096 22040 2102 22092
rect 2501 22083 2559 22089
rect 2501 22049 2513 22083
rect 2547 22080 2559 22083
rect 2682 22080 2688 22092
rect 2547 22052 2688 22080
rect 2547 22049 2559 22052
rect 2501 22043 2559 22049
rect 2682 22040 2688 22052
rect 2740 22040 2746 22092
rect 3804 22080 3832 22179
rect 8294 22176 8300 22228
rect 8352 22216 8358 22228
rect 8481 22219 8539 22225
rect 8481 22216 8493 22219
rect 8352 22188 8493 22216
rect 8352 22176 8358 22188
rect 8481 22185 8493 22188
rect 8527 22216 8539 22219
rect 8938 22216 8944 22228
rect 8527 22188 8944 22216
rect 8527 22185 8539 22188
rect 8481 22179 8539 22185
rect 8938 22176 8944 22188
rect 8996 22176 9002 22228
rect 13357 22219 13415 22225
rect 13357 22185 13369 22219
rect 13403 22216 13415 22219
rect 13449 22219 13507 22225
rect 13449 22216 13461 22219
rect 13403 22188 13461 22216
rect 13403 22185 13415 22188
rect 13357 22179 13415 22185
rect 13449 22185 13461 22188
rect 13495 22216 13507 22219
rect 13722 22216 13728 22228
rect 13495 22188 13728 22216
rect 13495 22185 13507 22188
rect 13449 22179 13507 22185
rect 13722 22176 13728 22188
rect 13780 22176 13786 22228
rect 4709 22151 4767 22157
rect 4709 22117 4721 22151
rect 4755 22148 4767 22151
rect 5442 22148 5448 22160
rect 4755 22120 5448 22148
rect 4755 22117 4767 22120
rect 4709 22111 4767 22117
rect 5442 22108 5448 22120
rect 5500 22108 5506 22160
rect 10962 22108 10968 22160
rect 11020 22148 11026 22160
rect 11210 22151 11268 22157
rect 11210 22148 11222 22151
rect 11020 22120 11222 22148
rect 11020 22108 11026 22120
rect 11210 22117 11222 22120
rect 11256 22148 11268 22151
rect 11514 22148 11520 22160
rect 11256 22120 11520 22148
rect 11256 22117 11268 22120
rect 11210 22111 11268 22117
rect 11514 22108 11520 22120
rect 11572 22108 11578 22160
rect 5258 22080 5264 22092
rect 3804 22052 5264 22080
rect 5258 22040 5264 22052
rect 5316 22040 5322 22092
rect 5905 22083 5963 22089
rect 5905 22049 5917 22083
rect 5951 22080 5963 22083
rect 5994 22080 6000 22092
rect 5951 22052 6000 22080
rect 5951 22049 5963 22052
rect 5905 22043 5963 22049
rect 5994 22040 6000 22052
rect 6052 22040 6058 22092
rect 7374 22089 7380 22092
rect 6917 22083 6975 22089
rect 6917 22049 6929 22083
rect 6963 22080 6975 22083
rect 7368 22080 7380 22089
rect 6963 22052 7380 22080
rect 6963 22049 6975 22052
rect 6917 22043 6975 22049
rect 7368 22043 7380 22052
rect 7374 22040 7380 22043
rect 7432 22040 7438 22092
rect 9677 22083 9735 22089
rect 9677 22049 9689 22083
rect 9723 22080 9735 22083
rect 9766 22080 9772 22092
rect 9723 22052 9772 22080
rect 9723 22049 9735 22052
rect 9677 22043 9735 22049
rect 9766 22040 9772 22052
rect 9824 22040 9830 22092
rect 10686 22040 10692 22092
rect 10744 22080 10750 22092
rect 12342 22080 12348 22092
rect 10744 22052 12348 22080
rect 10744 22040 10750 22052
rect 10980 22024 11008 22052
rect 12342 22040 12348 22052
rect 12400 22040 12406 22092
rect 13817 22083 13875 22089
rect 13817 22049 13829 22083
rect 13863 22080 13875 22083
rect 13998 22080 14004 22092
rect 13863 22052 14004 22080
rect 13863 22049 13875 22052
rect 13817 22043 13875 22049
rect 13998 22040 14004 22052
rect 14056 22040 14062 22092
rect 15289 22083 15347 22089
rect 15289 22049 15301 22083
rect 15335 22049 15347 22083
rect 15562 22080 15568 22092
rect 15523 22052 15568 22080
rect 15289 22043 15347 22049
rect 2314 22012 2320 22024
rect 1412 21984 2320 22012
rect 2314 21972 2320 21984
rect 2372 21972 2378 22024
rect 3145 22015 3203 22021
rect 3145 21981 3157 22015
rect 3191 22012 3203 22015
rect 3326 22012 3332 22024
rect 3191 21984 3332 22012
rect 3191 21981 3203 21984
rect 3145 21975 3203 21981
rect 3326 21972 3332 21984
rect 3384 21972 3390 22024
rect 4798 22012 4804 22024
rect 4759 21984 4804 22012
rect 4798 21972 4804 21984
rect 4856 21972 4862 22024
rect 4982 21972 4988 22024
rect 5040 22012 5046 22024
rect 5534 22012 5540 22024
rect 5040 21984 5540 22012
rect 5040 21972 5046 21984
rect 5534 21972 5540 21984
rect 5592 21972 5598 22024
rect 6549 22015 6607 22021
rect 6549 21981 6561 22015
rect 6595 22012 6607 22015
rect 7098 22012 7104 22024
rect 6595 21984 7104 22012
rect 6595 21981 6607 21984
rect 6549 21975 6607 21981
rect 7098 21972 7104 21984
rect 7156 21972 7162 22024
rect 9861 22015 9919 22021
rect 9861 21981 9873 22015
rect 9907 21981 9919 22015
rect 10962 22012 10968 22024
rect 10875 21984 10968 22012
rect 9861 21975 9919 21981
rect 1578 21944 1584 21956
rect 1539 21916 1584 21944
rect 1578 21904 1584 21916
rect 1636 21904 1642 21956
rect 4154 21904 4160 21956
rect 4212 21944 4218 21956
rect 4341 21947 4399 21953
rect 4341 21944 4353 21947
rect 4212 21916 4353 21944
rect 4212 21904 4218 21916
rect 4341 21913 4353 21916
rect 4387 21913 4399 21947
rect 6086 21944 6092 21956
rect 6047 21916 6092 21944
rect 4341 21907 4399 21913
rect 6086 21904 6092 21916
rect 6144 21904 6150 21956
rect 9674 21904 9680 21956
rect 9732 21944 9738 21956
rect 9876 21944 9904 21975
rect 10962 21972 10968 21984
rect 11020 21972 11026 22024
rect 13354 21972 13360 22024
rect 13412 22012 13418 22024
rect 13906 22012 13912 22024
rect 13412 21984 13912 22012
rect 13412 21972 13418 21984
rect 13906 21972 13912 21984
rect 13964 21972 13970 22024
rect 14090 22012 14096 22024
rect 14051 21984 14096 22012
rect 14090 21972 14096 21984
rect 14148 21972 14154 22024
rect 15304 22012 15332 22043
rect 15562 22040 15568 22052
rect 15620 22040 15626 22092
rect 15654 22012 15660 22024
rect 15304 21984 15660 22012
rect 15654 21972 15660 21984
rect 15712 21972 15718 22024
rect 9732 21916 9904 21944
rect 9732 21904 9738 21916
rect 2685 21879 2743 21885
rect 2685 21845 2697 21879
rect 2731 21876 2743 21879
rect 2866 21876 2872 21888
rect 2731 21848 2872 21876
rect 2731 21845 2743 21848
rect 2685 21839 2743 21845
rect 2866 21836 2872 21848
rect 2924 21836 2930 21888
rect 3142 21836 3148 21888
rect 3200 21876 3206 21888
rect 3421 21879 3479 21885
rect 3421 21876 3433 21879
rect 3200 21848 3433 21876
rect 3200 21836 3206 21848
rect 3421 21845 3433 21848
rect 3467 21845 3479 21879
rect 3421 21839 3479 21845
rect 5258 21836 5264 21888
rect 5316 21876 5322 21888
rect 5353 21879 5411 21885
rect 5353 21876 5365 21879
rect 5316 21848 5365 21876
rect 5316 21836 5322 21848
rect 5353 21845 5365 21848
rect 5399 21876 5411 21879
rect 5721 21879 5779 21885
rect 5721 21876 5733 21879
rect 5399 21848 5733 21876
rect 5399 21845 5411 21848
rect 5353 21839 5411 21845
rect 5721 21845 5733 21848
rect 5767 21845 5779 21879
rect 9030 21876 9036 21888
rect 8991 21848 9036 21876
rect 5721 21839 5779 21845
rect 9030 21836 9036 21848
rect 9088 21836 9094 21888
rect 9490 21876 9496 21888
rect 9451 21848 9496 21876
rect 9490 21836 9496 21848
rect 9548 21836 9554 21888
rect 10597 21879 10655 21885
rect 10597 21845 10609 21879
rect 10643 21876 10655 21879
rect 11146 21876 11152 21888
rect 10643 21848 11152 21876
rect 10643 21845 10655 21848
rect 10597 21839 10655 21845
rect 11146 21836 11152 21848
rect 11204 21876 11210 21888
rect 12345 21879 12403 21885
rect 12345 21876 12357 21879
rect 11204 21848 12357 21876
rect 11204 21836 11210 21848
rect 12345 21845 12357 21848
rect 12391 21845 12403 21879
rect 12345 21839 12403 21845
rect 12989 21879 13047 21885
rect 12989 21845 13001 21879
rect 13035 21876 13047 21879
rect 13078 21876 13084 21888
rect 13035 21848 13084 21876
rect 13035 21845 13047 21848
rect 12989 21839 13047 21845
rect 13078 21836 13084 21848
rect 13136 21836 13142 21888
rect 14645 21879 14703 21885
rect 14645 21845 14657 21879
rect 14691 21876 14703 21879
rect 14734 21876 14740 21888
rect 14691 21848 14740 21876
rect 14691 21845 14703 21848
rect 14645 21839 14703 21845
rect 14734 21836 14740 21848
rect 14792 21836 14798 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 2314 21672 2320 21684
rect 2275 21644 2320 21672
rect 2314 21632 2320 21644
rect 2372 21632 2378 21684
rect 2774 21632 2780 21684
rect 2832 21672 2838 21684
rect 3142 21672 3148 21684
rect 2832 21644 3148 21672
rect 2832 21632 2838 21644
rect 3142 21632 3148 21644
rect 3200 21632 3206 21684
rect 3881 21675 3939 21681
rect 3881 21641 3893 21675
rect 3927 21672 3939 21675
rect 4798 21672 4804 21684
rect 3927 21644 4804 21672
rect 3927 21641 3939 21644
rect 3881 21635 3939 21641
rect 4798 21632 4804 21644
rect 4856 21632 4862 21684
rect 5442 21672 5448 21684
rect 5403 21644 5448 21672
rect 5442 21632 5448 21644
rect 5500 21632 5506 21684
rect 5534 21632 5540 21684
rect 5592 21672 5598 21684
rect 6089 21675 6147 21681
rect 6089 21672 6101 21675
rect 5592 21644 6101 21672
rect 5592 21632 5598 21644
rect 6089 21641 6101 21644
rect 6135 21641 6147 21675
rect 6089 21635 6147 21641
rect 7282 21632 7288 21684
rect 7340 21672 7346 21684
rect 7653 21675 7711 21681
rect 7653 21672 7665 21675
rect 7340 21644 7665 21672
rect 7340 21632 7346 21644
rect 7653 21641 7665 21644
rect 7699 21641 7711 21675
rect 7653 21635 7711 21641
rect 9766 21632 9772 21684
rect 9824 21672 9830 21684
rect 9953 21675 10011 21681
rect 9953 21672 9965 21675
rect 9824 21644 9965 21672
rect 9824 21632 9830 21644
rect 9953 21641 9965 21644
rect 9999 21641 10011 21675
rect 11514 21672 11520 21684
rect 11475 21644 11520 21672
rect 9953 21635 10011 21641
rect 11514 21632 11520 21644
rect 11572 21632 11578 21684
rect 12069 21675 12127 21681
rect 12069 21641 12081 21675
rect 12115 21672 12127 21675
rect 12342 21672 12348 21684
rect 12115 21644 12348 21672
rect 12115 21641 12127 21644
rect 12069 21635 12127 21641
rect 12342 21632 12348 21644
rect 12400 21632 12406 21684
rect 13906 21672 13912 21684
rect 13867 21644 13912 21672
rect 13906 21632 13912 21644
rect 13964 21632 13970 21684
rect 14090 21632 14096 21684
rect 14148 21672 14154 21684
rect 15933 21675 15991 21681
rect 15933 21672 15945 21675
rect 14148 21644 15945 21672
rect 14148 21632 14154 21644
rect 15933 21641 15945 21644
rect 15979 21641 15991 21675
rect 15933 21635 15991 21641
rect 3418 21604 3424 21616
rect 3252 21576 3424 21604
rect 3252 21545 3280 21576
rect 3418 21564 3424 21576
rect 3476 21604 3482 21616
rect 4341 21607 4399 21613
rect 4341 21604 4353 21607
rect 3476 21576 4353 21604
rect 3476 21564 3482 21576
rect 4341 21573 4353 21576
rect 4387 21573 4399 21607
rect 4341 21567 4399 21573
rect 12989 21607 13047 21613
rect 12989 21573 13001 21607
rect 13035 21604 13047 21607
rect 14108 21604 14136 21632
rect 13035 21576 14136 21604
rect 13035 21573 13047 21576
rect 12989 21567 13047 21573
rect 3237 21539 3295 21545
rect 3237 21505 3249 21539
rect 3283 21505 3295 21539
rect 3237 21499 3295 21505
rect 3326 21496 3332 21548
rect 3384 21536 3390 21548
rect 4154 21536 4160 21548
rect 3384 21508 4160 21536
rect 3384 21496 3390 21508
rect 4154 21496 4160 21508
rect 4212 21496 4218 21548
rect 4890 21536 4896 21548
rect 4851 21508 4896 21536
rect 4890 21496 4896 21508
rect 4948 21496 4954 21548
rect 7561 21539 7619 21545
rect 7561 21505 7573 21539
rect 7607 21536 7619 21539
rect 8018 21536 8024 21548
rect 7607 21508 8024 21536
rect 7607 21505 7619 21508
rect 7561 21499 7619 21505
rect 8018 21496 8024 21508
rect 8076 21536 8082 21548
rect 8113 21539 8171 21545
rect 8113 21536 8125 21539
rect 8076 21508 8125 21536
rect 8076 21496 8082 21508
rect 8113 21505 8125 21508
rect 8159 21505 8171 21539
rect 8113 21499 8171 21505
rect 8297 21539 8355 21545
rect 8297 21505 8309 21539
rect 8343 21536 8355 21539
rect 9033 21539 9091 21545
rect 9033 21536 9045 21539
rect 8343 21508 9045 21536
rect 8343 21505 8355 21508
rect 8297 21499 8355 21505
rect 9033 21505 9045 21508
rect 9079 21536 9091 21539
rect 9122 21536 9128 21548
rect 9079 21508 9128 21536
rect 9079 21505 9091 21508
rect 9033 21499 9091 21505
rect 9122 21496 9128 21508
rect 9180 21496 9186 21548
rect 9493 21539 9551 21545
rect 9493 21505 9505 21539
rect 9539 21536 9551 21539
rect 9582 21536 9588 21548
rect 9539 21508 9588 21536
rect 9539 21505 9551 21508
rect 9493 21499 9551 21505
rect 9582 21496 9588 21508
rect 9640 21496 9646 21548
rect 10413 21539 10471 21545
rect 10413 21505 10425 21539
rect 10459 21536 10471 21539
rect 10870 21536 10876 21548
rect 10459 21508 10876 21536
rect 10459 21505 10471 21508
rect 10413 21499 10471 21505
rect 10870 21496 10876 21508
rect 10928 21536 10934 21548
rect 10965 21539 11023 21545
rect 10965 21536 10977 21539
rect 10928 21508 10977 21536
rect 10928 21496 10934 21508
rect 10965 21505 10977 21508
rect 11011 21505 11023 21539
rect 11146 21536 11152 21548
rect 11107 21508 11152 21536
rect 10965 21499 11023 21505
rect 11146 21496 11152 21508
rect 11204 21496 11210 21548
rect 1489 21471 1547 21477
rect 1489 21437 1501 21471
rect 1535 21468 1547 21471
rect 2038 21468 2044 21480
rect 1535 21440 2044 21468
rect 1535 21437 1547 21440
rect 1489 21431 1547 21437
rect 2038 21428 2044 21440
rect 2096 21428 2102 21480
rect 4249 21471 4307 21477
rect 4249 21437 4261 21471
rect 4295 21468 4307 21471
rect 4801 21471 4859 21477
rect 4801 21468 4813 21471
rect 4295 21440 4813 21468
rect 4295 21437 4307 21440
rect 4249 21431 4307 21437
rect 4801 21437 4813 21440
rect 4847 21468 4859 21471
rect 5074 21468 5080 21480
rect 4847 21440 5080 21468
rect 4847 21437 4859 21440
rect 4801 21431 4859 21437
rect 5074 21428 5080 21440
rect 5132 21428 5138 21480
rect 6454 21468 6460 21480
rect 6415 21440 6460 21468
rect 6454 21428 6460 21440
rect 6512 21428 6518 21480
rect 12253 21471 12311 21477
rect 12253 21468 12265 21471
rect 12176 21440 12265 21468
rect 1762 21400 1768 21412
rect 1723 21372 1768 21400
rect 1762 21360 1768 21372
rect 1820 21360 1826 21412
rect 3142 21400 3148 21412
rect 3103 21372 3148 21400
rect 3142 21360 3148 21372
rect 3200 21360 3206 21412
rect 7374 21360 7380 21412
rect 7432 21400 7438 21412
rect 7432 21372 8524 21400
rect 7432 21360 7438 21372
rect 2685 21335 2743 21341
rect 2685 21301 2697 21335
rect 2731 21332 2743 21335
rect 3160 21332 3188 21360
rect 8496 21344 8524 21372
rect 12176 21344 12204 21440
rect 12253 21437 12265 21440
rect 12299 21437 12311 21471
rect 13078 21468 13084 21480
rect 13039 21440 13084 21468
rect 12253 21431 12311 21437
rect 13078 21428 13084 21440
rect 13136 21428 13142 21480
rect 14550 21468 14556 21480
rect 14511 21440 14556 21468
rect 14550 21428 14556 21440
rect 14608 21428 14614 21480
rect 12802 21360 12808 21412
rect 12860 21400 12866 21412
rect 13357 21403 13415 21409
rect 13357 21400 13369 21403
rect 12860 21372 13369 21400
rect 12860 21360 12866 21372
rect 13357 21369 13369 21372
rect 13403 21369 13415 21403
rect 13357 21363 13415 21369
rect 14734 21360 14740 21412
rect 14792 21409 14798 21412
rect 14792 21403 14856 21409
rect 14792 21369 14810 21403
rect 14844 21369 14856 21403
rect 14792 21363 14856 21369
rect 14792 21360 14798 21363
rect 2731 21304 3188 21332
rect 4709 21335 4767 21341
rect 2731 21301 2743 21304
rect 2685 21295 2743 21301
rect 4709 21301 4721 21335
rect 4755 21332 4767 21335
rect 5810 21332 5816 21344
rect 4755 21304 5816 21332
rect 4755 21301 4767 21304
rect 4709 21295 4767 21301
rect 5810 21292 5816 21304
rect 5868 21292 5874 21344
rect 6273 21335 6331 21341
rect 6273 21301 6285 21335
rect 6319 21332 6331 21335
rect 7098 21332 7104 21344
rect 6319 21304 7104 21332
rect 6319 21301 6331 21304
rect 6273 21295 6331 21301
rect 7098 21292 7104 21304
rect 7156 21292 7162 21344
rect 7193 21335 7251 21341
rect 7193 21301 7205 21335
rect 7239 21332 7251 21335
rect 8018 21332 8024 21344
rect 7239 21304 8024 21332
rect 7239 21301 7251 21304
rect 7193 21295 7251 21301
rect 8018 21292 8024 21304
rect 8076 21292 8082 21344
rect 8478 21292 8484 21344
rect 8536 21332 8542 21344
rect 8665 21335 8723 21341
rect 8665 21332 8677 21335
rect 8536 21304 8677 21332
rect 8536 21292 8542 21304
rect 8665 21301 8677 21304
rect 8711 21301 8723 21335
rect 8665 21295 8723 21301
rect 10505 21335 10563 21341
rect 10505 21301 10517 21335
rect 10551 21332 10563 21335
rect 10686 21332 10692 21344
rect 10551 21304 10692 21332
rect 10551 21301 10563 21304
rect 10505 21295 10563 21301
rect 10686 21292 10692 21304
rect 10744 21292 10750 21344
rect 10870 21332 10876 21344
rect 10831 21304 10876 21332
rect 10870 21292 10876 21304
rect 10928 21292 10934 21344
rect 11977 21335 12035 21341
rect 11977 21301 11989 21335
rect 12023 21332 12035 21335
rect 12158 21332 12164 21344
rect 12023 21304 12164 21332
rect 12023 21301 12035 21304
rect 11977 21295 12035 21301
rect 12158 21292 12164 21304
rect 12216 21292 12222 21344
rect 13906 21292 13912 21344
rect 13964 21332 13970 21344
rect 14185 21335 14243 21341
rect 14185 21332 14197 21335
rect 13964 21304 14197 21332
rect 13964 21292 13970 21304
rect 14185 21301 14197 21304
rect 14231 21301 14243 21335
rect 14185 21295 14243 21301
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 2501 21131 2559 21137
rect 2501 21097 2513 21131
rect 2547 21128 2559 21131
rect 2682 21128 2688 21140
rect 2547 21100 2688 21128
rect 2547 21097 2559 21100
rect 2501 21091 2559 21097
rect 2682 21088 2688 21100
rect 2740 21088 2746 21140
rect 3418 21128 3424 21140
rect 3379 21100 3424 21128
rect 3418 21088 3424 21100
rect 3476 21088 3482 21140
rect 4154 21088 4160 21140
rect 4212 21128 4218 21140
rect 5445 21131 5503 21137
rect 5445 21128 5457 21131
rect 4212 21100 5457 21128
rect 4212 21088 4218 21100
rect 5445 21097 5457 21100
rect 5491 21097 5503 21131
rect 5994 21128 6000 21140
rect 5955 21100 6000 21128
rect 5445 21091 5503 21097
rect 5994 21088 6000 21100
rect 6052 21088 6058 21140
rect 8478 21128 8484 21140
rect 8439 21100 8484 21128
rect 8478 21088 8484 21100
rect 8536 21088 8542 21140
rect 13078 21088 13084 21140
rect 13136 21128 13142 21140
rect 13633 21131 13691 21137
rect 13633 21128 13645 21131
rect 13136 21100 13645 21128
rect 13136 21088 13142 21100
rect 13633 21097 13645 21100
rect 13679 21097 13691 21131
rect 16298 21128 16304 21140
rect 16259 21100 16304 21128
rect 13633 21091 13691 21097
rect 16298 21088 16304 21100
rect 16356 21088 16362 21140
rect 1765 21063 1823 21069
rect 1765 21029 1777 21063
rect 1811 21060 1823 21063
rect 2590 21060 2596 21072
rect 1811 21032 2596 21060
rect 1811 21029 1823 21032
rect 1765 21023 1823 21029
rect 2590 21020 2596 21032
rect 2648 21020 2654 21072
rect 3786 21060 3792 21072
rect 3699 21032 3792 21060
rect 3786 21020 3792 21032
rect 3844 21060 3850 21072
rect 4246 21060 4252 21072
rect 3844 21032 4252 21060
rect 3844 21020 3850 21032
rect 4246 21020 4252 21032
rect 4304 21069 4310 21072
rect 4304 21063 4368 21069
rect 4304 21029 4322 21063
rect 4356 21060 4368 21063
rect 4890 21060 4896 21072
rect 4356 21032 4896 21060
rect 4356 21029 4368 21032
rect 4304 21023 4368 21029
rect 4304 21020 4310 21023
rect 4890 21020 4896 21032
rect 4948 21020 4954 21072
rect 11146 21020 11152 21072
rect 11204 21069 11210 21072
rect 11204 21063 11268 21069
rect 11204 21029 11222 21063
rect 11256 21029 11268 21063
rect 11204 21023 11268 21029
rect 11204 21020 11210 21023
rect 1486 20992 1492 21004
rect 1447 20964 1492 20992
rect 1486 20952 1492 20964
rect 1544 20952 1550 21004
rect 2777 20995 2835 21001
rect 2777 20961 2789 20995
rect 2823 20961 2835 20995
rect 2777 20955 2835 20961
rect 2792 20924 2820 20955
rect 3878 20952 3884 21004
rect 3936 20992 3942 21004
rect 4065 20995 4123 21001
rect 4065 20992 4077 20995
rect 3936 20964 4077 20992
rect 3936 20952 3942 20964
rect 4065 20961 4077 20964
rect 4111 20961 4123 20995
rect 7006 20992 7012 21004
rect 6967 20964 7012 20992
rect 4065 20955 4123 20961
rect 7006 20952 7012 20964
rect 7064 20952 7070 21004
rect 7374 21001 7380 21004
rect 7368 20992 7380 21001
rect 7335 20964 7380 20992
rect 7368 20955 7380 20964
rect 7374 20952 7380 20955
rect 7432 20952 7438 21004
rect 9677 20995 9735 21001
rect 9677 20961 9689 20995
rect 9723 20992 9735 20995
rect 9950 20992 9956 21004
rect 9723 20964 9956 20992
rect 9723 20961 9735 20964
rect 9677 20955 9735 20961
rect 9950 20952 9956 20964
rect 10008 20952 10014 21004
rect 10962 20992 10968 21004
rect 10923 20964 10968 20992
rect 10962 20952 10968 20964
rect 11020 20952 11026 21004
rect 14001 20995 14059 21001
rect 14001 20961 14013 20995
rect 14047 20992 14059 20995
rect 14274 20992 14280 21004
rect 14047 20964 14280 20992
rect 14047 20961 14059 20964
rect 14001 20955 14059 20961
rect 14274 20952 14280 20964
rect 14332 20992 14338 21004
rect 15289 20995 15347 21001
rect 15289 20992 15301 20995
rect 14332 20964 15301 20992
rect 14332 20952 14338 20964
rect 15289 20961 15301 20964
rect 15335 20961 15347 20995
rect 15289 20955 15347 20961
rect 3326 20924 3332 20936
rect 2792 20896 3332 20924
rect 3326 20884 3332 20896
rect 3384 20924 3390 20936
rect 3970 20924 3976 20936
rect 3384 20896 3976 20924
rect 3384 20884 3390 20896
rect 3970 20884 3976 20896
rect 4028 20884 4034 20936
rect 7098 20924 7104 20936
rect 7011 20896 7104 20924
rect 7098 20884 7104 20896
rect 7156 20884 7162 20936
rect 9858 20924 9864 20936
rect 9819 20896 9864 20924
rect 9858 20884 9864 20896
rect 9916 20884 9922 20936
rect 13814 20884 13820 20936
rect 13872 20924 13878 20936
rect 14093 20927 14151 20933
rect 14093 20924 14105 20927
rect 13872 20896 14105 20924
rect 13872 20884 13878 20896
rect 14093 20893 14105 20896
rect 14139 20893 14151 20927
rect 14093 20887 14151 20893
rect 14185 20927 14243 20933
rect 14185 20893 14197 20927
rect 14231 20924 14243 20927
rect 14734 20924 14740 20936
rect 14231 20896 14740 20924
rect 14231 20893 14243 20896
rect 14185 20887 14243 20893
rect 14734 20884 14740 20896
rect 14792 20884 14798 20936
rect 5534 20816 5540 20868
rect 5592 20856 5598 20868
rect 6365 20859 6423 20865
rect 6365 20856 6377 20859
rect 5592 20828 6377 20856
rect 5592 20816 5598 20828
rect 6365 20825 6377 20828
rect 6411 20856 6423 20859
rect 6454 20856 6460 20868
rect 6411 20828 6460 20856
rect 6411 20825 6423 20828
rect 6365 20819 6423 20825
rect 6454 20816 6460 20828
rect 6512 20856 6518 20868
rect 6825 20859 6883 20865
rect 6825 20856 6837 20859
rect 6512 20828 6837 20856
rect 6512 20816 6518 20828
rect 6825 20825 6837 20828
rect 6871 20825 6883 20859
rect 6825 20819 6883 20825
rect 2958 20788 2964 20800
rect 2919 20760 2964 20788
rect 2958 20748 2964 20760
rect 3016 20748 3022 20800
rect 7116 20788 7144 20884
rect 7742 20788 7748 20800
rect 7116 20760 7748 20788
rect 7742 20748 7748 20760
rect 7800 20788 7806 20800
rect 9030 20788 9036 20800
rect 7800 20760 9036 20788
rect 7800 20748 7806 20760
rect 9030 20748 9036 20760
rect 9088 20788 9094 20800
rect 9125 20791 9183 20797
rect 9125 20788 9137 20791
rect 9088 20760 9137 20788
rect 9088 20748 9094 20760
rect 9125 20757 9137 20760
rect 9171 20788 9183 20791
rect 9493 20791 9551 20797
rect 9493 20788 9505 20791
rect 9171 20760 9505 20788
rect 9171 20757 9183 20760
rect 9125 20751 9183 20757
rect 9493 20757 9505 20760
rect 9539 20788 9551 20791
rect 9582 20788 9588 20800
rect 9539 20760 9588 20788
rect 9539 20757 9551 20760
rect 9493 20751 9551 20757
rect 9582 20748 9588 20760
rect 9640 20748 9646 20800
rect 10594 20788 10600 20800
rect 10555 20760 10600 20788
rect 10594 20748 10600 20760
rect 10652 20788 10658 20800
rect 10870 20788 10876 20800
rect 10652 20760 10876 20788
rect 10652 20748 10658 20760
rect 10870 20748 10876 20760
rect 10928 20748 10934 20800
rect 10962 20748 10968 20800
rect 11020 20788 11026 20800
rect 12345 20791 12403 20797
rect 12345 20788 12357 20791
rect 11020 20760 12357 20788
rect 11020 20748 11026 20760
rect 12345 20757 12357 20760
rect 12391 20757 12403 20791
rect 13170 20788 13176 20800
rect 13131 20760 13176 20788
rect 12345 20751 12403 20757
rect 13170 20748 13176 20760
rect 13228 20748 13234 20800
rect 14550 20748 14556 20800
rect 14608 20788 14614 20800
rect 14737 20791 14795 20797
rect 14737 20788 14749 20791
rect 14608 20760 14749 20788
rect 14608 20748 14614 20760
rect 14737 20757 14749 20760
rect 14783 20788 14795 20791
rect 14826 20788 14832 20800
rect 14783 20760 14832 20788
rect 14783 20757 14795 20760
rect 14737 20751 14795 20757
rect 14826 20748 14832 20760
rect 14884 20788 14890 20800
rect 15013 20791 15071 20797
rect 15013 20788 15025 20791
rect 14884 20760 15025 20788
rect 14884 20748 14890 20760
rect 15013 20757 15025 20760
rect 15059 20757 15071 20791
rect 15013 20751 15071 20757
rect 15654 20748 15660 20800
rect 15712 20788 15718 20800
rect 15749 20791 15807 20797
rect 15749 20788 15761 20791
rect 15712 20760 15761 20788
rect 15712 20748 15718 20760
rect 15749 20757 15761 20760
rect 15795 20757 15807 20791
rect 15749 20751 15807 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1486 20544 1492 20596
rect 1544 20584 1550 20596
rect 2038 20584 2044 20596
rect 1544 20556 2044 20584
rect 1544 20544 1550 20556
rect 2038 20544 2044 20556
rect 2096 20584 2102 20596
rect 2685 20587 2743 20593
rect 2685 20584 2697 20587
rect 2096 20556 2697 20584
rect 2096 20544 2102 20556
rect 2685 20553 2697 20556
rect 2731 20553 2743 20587
rect 3786 20584 3792 20596
rect 3747 20556 3792 20584
rect 2685 20547 2743 20553
rect 3786 20544 3792 20556
rect 3844 20544 3850 20596
rect 4154 20584 4160 20596
rect 4115 20556 4160 20584
rect 4154 20544 4160 20556
rect 4212 20544 4218 20596
rect 7193 20587 7251 20593
rect 7193 20553 7205 20587
rect 7239 20584 7251 20587
rect 7374 20584 7380 20596
rect 7239 20556 7380 20584
rect 7239 20553 7251 20556
rect 7193 20547 7251 20553
rect 7374 20544 7380 20556
rect 7432 20584 7438 20596
rect 9122 20584 9128 20596
rect 7432 20556 9128 20584
rect 7432 20544 7438 20556
rect 9122 20544 9128 20556
rect 9180 20544 9186 20596
rect 9769 20587 9827 20593
rect 9769 20553 9781 20587
rect 9815 20584 9827 20587
rect 9950 20584 9956 20596
rect 9815 20556 9956 20584
rect 9815 20553 9827 20556
rect 9769 20547 9827 20553
rect 9950 20544 9956 20556
rect 10008 20544 10014 20596
rect 11146 20544 11152 20596
rect 11204 20584 11210 20596
rect 11241 20587 11299 20593
rect 11241 20584 11253 20587
rect 11204 20556 11253 20584
rect 11204 20544 11210 20556
rect 11241 20553 11253 20556
rect 11287 20553 11299 20587
rect 11241 20547 11299 20553
rect 12253 20587 12311 20593
rect 12253 20553 12265 20587
rect 12299 20584 12311 20587
rect 13173 20587 13231 20593
rect 13173 20584 13185 20587
rect 12299 20556 13185 20584
rect 12299 20553 12311 20556
rect 12253 20547 12311 20553
rect 13173 20553 13185 20556
rect 13219 20584 13231 20587
rect 13722 20584 13728 20596
rect 13219 20556 13728 20584
rect 13219 20553 13231 20556
rect 13173 20547 13231 20553
rect 13722 20544 13728 20556
rect 13780 20544 13786 20596
rect 14274 20584 14280 20596
rect 14235 20556 14280 20584
rect 14274 20544 14280 20556
rect 14332 20544 14338 20596
rect 14734 20544 14740 20596
rect 14792 20584 14798 20596
rect 16117 20587 16175 20593
rect 16117 20584 16129 20587
rect 14792 20556 16129 20584
rect 14792 20544 14798 20556
rect 16117 20553 16129 20556
rect 16163 20553 16175 20587
rect 16117 20547 16175 20553
rect 1673 20451 1731 20457
rect 1673 20417 1685 20451
rect 1719 20448 1731 20451
rect 2498 20448 2504 20460
rect 1719 20420 2504 20448
rect 1719 20417 1731 20420
rect 1673 20411 1731 20417
rect 2498 20408 2504 20420
rect 2556 20408 2562 20460
rect 2593 20451 2651 20457
rect 2593 20417 2605 20451
rect 2639 20448 2651 20451
rect 3329 20451 3387 20457
rect 3329 20448 3341 20451
rect 2639 20420 3341 20448
rect 2639 20417 2651 20420
rect 2593 20411 2651 20417
rect 3329 20417 3341 20420
rect 3375 20448 3387 20451
rect 3418 20448 3424 20460
rect 3375 20420 3424 20448
rect 3375 20417 3387 20420
rect 3329 20411 3387 20417
rect 3418 20408 3424 20420
rect 3476 20408 3482 20460
rect 4172 20448 4200 20544
rect 11609 20519 11667 20525
rect 11609 20516 11621 20519
rect 10704 20488 11621 20516
rect 10704 20460 10732 20488
rect 11609 20485 11621 20488
rect 11655 20485 11667 20519
rect 11609 20479 11667 20485
rect 7742 20448 7748 20460
rect 4172 20420 4384 20448
rect 7703 20420 7748 20448
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20380 1455 20383
rect 2314 20380 2320 20392
rect 1443 20352 2320 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 2314 20340 2320 20352
rect 2372 20340 2378 20392
rect 4249 20383 4307 20389
rect 4249 20349 4261 20383
rect 4295 20349 4307 20383
rect 4356 20380 4384 20420
rect 7742 20408 7748 20420
rect 7800 20408 7806 20460
rect 10686 20448 10692 20460
rect 10647 20420 10692 20448
rect 10686 20408 10692 20420
rect 10744 20408 10750 20460
rect 10873 20451 10931 20457
rect 10873 20417 10885 20451
rect 10919 20448 10931 20451
rect 10962 20448 10968 20460
rect 10919 20420 10968 20448
rect 10919 20417 10931 20420
rect 10873 20411 10931 20417
rect 10962 20408 10968 20420
rect 11020 20408 11026 20460
rect 13081 20451 13139 20457
rect 13081 20417 13093 20451
rect 13127 20448 13139 20451
rect 13630 20448 13636 20460
rect 13127 20420 13636 20448
rect 13127 20417 13139 20420
rect 13081 20411 13139 20417
rect 13630 20408 13636 20420
rect 13688 20408 13694 20460
rect 13817 20451 13875 20457
rect 13817 20417 13829 20451
rect 13863 20448 13875 20451
rect 13863 20420 14688 20448
rect 13863 20417 13875 20420
rect 13817 20411 13875 20417
rect 4505 20383 4563 20389
rect 4505 20380 4517 20383
rect 4356 20352 4517 20380
rect 4249 20343 4307 20349
rect 4505 20349 4517 20352
rect 4551 20349 4563 20383
rect 4505 20343 4563 20349
rect 12713 20383 12771 20389
rect 12713 20349 12725 20383
rect 12759 20380 12771 20383
rect 13832 20380 13860 20411
rect 12759 20352 13860 20380
rect 12759 20349 12771 20352
rect 12713 20343 12771 20349
rect 2225 20315 2283 20321
rect 2225 20281 2237 20315
rect 2271 20312 2283 20315
rect 2682 20312 2688 20324
rect 2271 20284 2688 20312
rect 2271 20281 2283 20284
rect 2225 20275 2283 20281
rect 2682 20272 2688 20284
rect 2740 20272 2746 20324
rect 2774 20272 2780 20324
rect 2832 20312 2838 20324
rect 3053 20315 3111 20321
rect 3053 20312 3065 20315
rect 2832 20284 3065 20312
rect 2832 20272 2838 20284
rect 3053 20281 3065 20284
rect 3099 20312 3111 20315
rect 3694 20312 3700 20324
rect 3099 20284 3700 20312
rect 3099 20281 3111 20284
rect 3053 20275 3111 20281
rect 3694 20272 3700 20284
rect 3752 20272 3758 20324
rect 4264 20312 4292 20343
rect 4614 20312 4620 20324
rect 4264 20284 4620 20312
rect 4614 20272 4620 20284
rect 4672 20312 4678 20324
rect 5258 20312 5264 20324
rect 4672 20284 5264 20312
rect 4672 20272 4678 20284
rect 5258 20272 5264 20284
rect 5316 20312 5322 20324
rect 6178 20312 6184 20324
rect 5316 20284 6184 20312
rect 5316 20272 5322 20284
rect 6178 20272 6184 20284
rect 6236 20272 6242 20324
rect 7653 20315 7711 20321
rect 7653 20281 7665 20315
rect 7699 20312 7711 20315
rect 7990 20315 8048 20321
rect 7990 20312 8002 20315
rect 7699 20284 8002 20312
rect 7699 20281 7711 20284
rect 7653 20275 7711 20281
rect 7990 20281 8002 20284
rect 8036 20312 8048 20315
rect 8202 20312 8208 20324
rect 8036 20284 8208 20312
rect 8036 20281 8048 20284
rect 7990 20275 8048 20281
rect 8202 20272 8208 20284
rect 8260 20272 8266 20324
rect 10134 20312 10140 20324
rect 10047 20284 10140 20312
rect 10134 20272 10140 20284
rect 10192 20312 10198 20324
rect 14660 20321 14688 20420
rect 14737 20383 14795 20389
rect 14737 20349 14749 20383
rect 14783 20380 14795 20383
rect 14826 20380 14832 20392
rect 14783 20352 14832 20380
rect 14783 20349 14795 20352
rect 14737 20343 14795 20349
rect 14826 20340 14832 20352
rect 14884 20380 14890 20392
rect 15286 20380 15292 20392
rect 14884 20352 15292 20380
rect 14884 20340 14890 20352
rect 15286 20340 15292 20352
rect 15344 20340 15350 20392
rect 15010 20321 15016 20324
rect 10597 20315 10655 20321
rect 10597 20312 10609 20315
rect 10192 20284 10609 20312
rect 10192 20272 10198 20284
rect 10597 20281 10609 20284
rect 10643 20281 10655 20315
rect 10597 20275 10655 20281
rect 14645 20315 14703 20321
rect 14645 20281 14657 20315
rect 14691 20312 14703 20315
rect 15004 20312 15016 20321
rect 14691 20284 15016 20312
rect 14691 20281 14703 20284
rect 14645 20275 14703 20281
rect 15004 20275 15016 20284
rect 15010 20272 15016 20275
rect 15068 20272 15074 20324
rect 3142 20244 3148 20256
rect 3103 20216 3148 20244
rect 3142 20204 3148 20216
rect 3200 20204 3206 20256
rect 5350 20204 5356 20256
rect 5408 20244 5414 20256
rect 5629 20247 5687 20253
rect 5629 20244 5641 20247
rect 5408 20216 5641 20244
rect 5408 20204 5414 20216
rect 5629 20213 5641 20216
rect 5675 20213 5687 20247
rect 5629 20207 5687 20213
rect 6641 20247 6699 20253
rect 6641 20213 6653 20247
rect 6687 20244 6699 20247
rect 7006 20244 7012 20256
rect 6687 20216 7012 20244
rect 6687 20213 6699 20216
rect 6641 20207 6699 20213
rect 7006 20204 7012 20216
rect 7064 20244 7070 20256
rect 7742 20244 7748 20256
rect 7064 20216 7748 20244
rect 7064 20204 7070 20216
rect 7742 20204 7748 20216
rect 7800 20204 7806 20256
rect 9674 20204 9680 20256
rect 9732 20244 9738 20256
rect 10229 20247 10287 20253
rect 10229 20244 10241 20247
rect 9732 20216 10241 20244
rect 9732 20204 9738 20216
rect 10229 20213 10241 20216
rect 10275 20213 10287 20247
rect 10229 20207 10287 20213
rect 13170 20204 13176 20256
rect 13228 20244 13234 20256
rect 13541 20247 13599 20253
rect 13541 20244 13553 20247
rect 13228 20216 13553 20244
rect 13228 20204 13234 20216
rect 13541 20213 13553 20216
rect 13587 20213 13599 20247
rect 13541 20207 13599 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 3326 20040 3332 20052
rect 3287 20012 3332 20040
rect 3326 20000 3332 20012
rect 3384 20000 3390 20052
rect 3510 20000 3516 20052
rect 3568 20040 3574 20052
rect 4065 20043 4123 20049
rect 4065 20040 4077 20043
rect 3568 20012 4077 20040
rect 3568 20000 3574 20012
rect 4065 20009 4077 20012
rect 4111 20009 4123 20043
rect 4065 20003 4123 20009
rect 6178 20000 6184 20052
rect 6236 20040 6242 20052
rect 7009 20043 7067 20049
rect 7009 20040 7021 20043
rect 6236 20012 7021 20040
rect 6236 20000 6242 20012
rect 7009 20009 7021 20012
rect 7055 20009 7067 20043
rect 8478 20040 8484 20052
rect 8439 20012 8484 20040
rect 7009 20003 7067 20009
rect 1765 19975 1823 19981
rect 1765 19941 1777 19975
rect 1811 19972 1823 19975
rect 2406 19972 2412 19984
rect 1811 19944 2412 19972
rect 1811 19941 1823 19944
rect 1765 19935 1823 19941
rect 2406 19932 2412 19944
rect 2464 19932 2470 19984
rect 7024 19972 7052 20003
rect 8478 20000 8484 20012
rect 8536 20000 8542 20052
rect 9766 20000 9772 20052
rect 9824 20040 9830 20052
rect 9861 20043 9919 20049
rect 9861 20040 9873 20043
rect 9824 20012 9873 20040
rect 9824 20000 9830 20012
rect 9861 20009 9873 20012
rect 9907 20009 9919 20043
rect 9861 20003 9919 20009
rect 14001 20043 14059 20049
rect 14001 20009 14013 20043
rect 14047 20040 14059 20043
rect 14734 20040 14740 20052
rect 14047 20012 14740 20040
rect 14047 20009 14059 20012
rect 14001 20003 14059 20009
rect 14734 20000 14740 20012
rect 14792 20000 14798 20052
rect 16666 20040 16672 20052
rect 16627 20012 16672 20040
rect 16666 20000 16672 20012
rect 16724 20000 16730 20052
rect 9398 19972 9404 19984
rect 7024 19944 9404 19972
rect 9398 19932 9404 19944
rect 9456 19932 9462 19984
rect 10321 19975 10379 19981
rect 10321 19941 10333 19975
rect 10367 19972 10379 19975
rect 10680 19975 10738 19981
rect 10680 19972 10692 19975
rect 10367 19944 10692 19972
rect 10367 19941 10379 19944
rect 10321 19935 10379 19941
rect 10680 19941 10692 19944
rect 10726 19972 10738 19975
rect 10962 19972 10968 19984
rect 10726 19944 10968 19972
rect 10726 19941 10738 19944
rect 10680 19935 10738 19941
rect 10962 19932 10968 19944
rect 11020 19932 11026 19984
rect 1486 19904 1492 19916
rect 1447 19876 1492 19904
rect 1486 19864 1492 19876
rect 1544 19864 1550 19916
rect 2777 19907 2835 19913
rect 2777 19873 2789 19907
rect 2823 19904 2835 19907
rect 3326 19904 3332 19916
rect 2823 19876 3332 19904
rect 2823 19873 2835 19876
rect 2777 19867 2835 19873
rect 3326 19864 3332 19876
rect 3384 19864 3390 19916
rect 5350 19913 5356 19916
rect 5344 19904 5356 19913
rect 5311 19876 5356 19904
rect 5344 19867 5356 19876
rect 5350 19864 5356 19867
rect 5408 19864 5414 19916
rect 7653 19907 7711 19913
rect 7653 19873 7665 19907
rect 7699 19904 7711 19907
rect 7926 19904 7932 19916
rect 7699 19876 7932 19904
rect 7699 19873 7711 19876
rect 7653 19867 7711 19873
rect 7926 19864 7932 19876
rect 7984 19864 7990 19916
rect 8389 19907 8447 19913
rect 8389 19873 8401 19907
rect 8435 19904 8447 19907
rect 8570 19904 8576 19916
rect 8435 19876 8576 19904
rect 8435 19873 8447 19876
rect 8389 19867 8447 19873
rect 8570 19864 8576 19876
rect 8628 19864 8634 19916
rect 12434 19864 12440 19916
rect 12492 19904 12498 19916
rect 15562 19913 15568 19916
rect 13265 19907 13323 19913
rect 13265 19904 13277 19907
rect 12492 19876 13277 19904
rect 12492 19864 12498 19876
rect 13265 19873 13277 19876
rect 13311 19904 13323 19907
rect 14277 19907 14335 19913
rect 14277 19904 14289 19907
rect 13311 19876 14289 19904
rect 13311 19873 13323 19876
rect 13265 19867 13323 19873
rect 14277 19873 14289 19876
rect 14323 19873 14335 19907
rect 15545 19907 15568 19913
rect 15545 19904 15557 19907
rect 14277 19867 14335 19873
rect 15028 19876 15557 19904
rect 4614 19796 4620 19848
rect 4672 19836 4678 19848
rect 5077 19839 5135 19845
rect 5077 19836 5089 19839
rect 4672 19808 5089 19836
rect 4672 19796 4678 19808
rect 5077 19805 5089 19808
rect 5123 19805 5135 19839
rect 5077 19799 5135 19805
rect 8665 19839 8723 19845
rect 8665 19805 8677 19839
rect 8711 19805 8723 19839
rect 8665 19799 8723 19805
rect 2685 19771 2743 19777
rect 2685 19737 2697 19771
rect 2731 19768 2743 19771
rect 3142 19768 3148 19780
rect 2731 19740 3148 19768
rect 2731 19737 2743 19740
rect 2685 19731 2743 19737
rect 3142 19728 3148 19740
rect 3200 19728 3206 19780
rect 8680 19768 8708 19799
rect 9674 19796 9680 19848
rect 9732 19836 9738 19848
rect 10413 19839 10471 19845
rect 10413 19836 10425 19839
rect 9732 19808 10425 19836
rect 9732 19796 9738 19808
rect 10413 19805 10425 19808
rect 10459 19805 10471 19839
rect 10413 19799 10471 19805
rect 12526 19796 12532 19848
rect 12584 19836 12590 19848
rect 13357 19839 13415 19845
rect 13357 19836 13369 19839
rect 12584 19808 13369 19836
rect 12584 19796 12590 19808
rect 13357 19805 13369 19808
rect 13403 19805 13415 19839
rect 13538 19836 13544 19848
rect 13499 19808 13544 19836
rect 13357 19799 13415 19805
rect 13538 19796 13544 19808
rect 13596 19836 13602 19848
rect 15028 19836 15056 19876
rect 15545 19873 15557 19876
rect 15620 19904 15626 19916
rect 15620 19876 15693 19904
rect 15545 19867 15568 19873
rect 15562 19864 15568 19867
rect 15620 19864 15626 19876
rect 15286 19836 15292 19848
rect 13596 19808 15056 19836
rect 15247 19808 15292 19836
rect 13596 19796 13602 19808
rect 15286 19796 15292 19808
rect 15344 19796 15350 19848
rect 8938 19768 8944 19780
rect 8680 19740 8944 19768
rect 8938 19728 8944 19740
rect 8996 19768 9002 19780
rect 15105 19771 15163 19777
rect 8996 19740 9996 19768
rect 8996 19728 9002 19740
rect 2314 19700 2320 19712
rect 2275 19672 2320 19700
rect 2314 19660 2320 19672
rect 2372 19660 2378 19712
rect 2866 19660 2872 19712
rect 2924 19700 2930 19712
rect 2961 19703 3019 19709
rect 2961 19700 2973 19703
rect 2924 19672 2973 19700
rect 2924 19660 2930 19672
rect 2961 19669 2973 19672
rect 3007 19669 3019 19703
rect 2961 19663 3019 19669
rect 3789 19703 3847 19709
rect 3789 19669 3801 19703
rect 3835 19700 3847 19703
rect 4062 19700 4068 19712
rect 3835 19672 4068 19700
rect 3835 19669 3847 19672
rect 3789 19663 3847 19669
rect 4062 19660 4068 19672
rect 4120 19660 4126 19712
rect 4801 19703 4859 19709
rect 4801 19669 4813 19703
rect 4847 19700 4859 19703
rect 4890 19700 4896 19712
rect 4847 19672 4896 19700
rect 4847 19669 4859 19672
rect 4801 19663 4859 19669
rect 4890 19660 4896 19672
rect 4948 19700 4954 19712
rect 5442 19700 5448 19712
rect 4948 19672 5448 19700
rect 4948 19660 4954 19672
rect 5442 19660 5448 19672
rect 5500 19660 5506 19712
rect 6270 19660 6276 19712
rect 6328 19700 6334 19712
rect 6457 19703 6515 19709
rect 6457 19700 6469 19703
rect 6328 19672 6469 19700
rect 6328 19660 6334 19672
rect 6457 19669 6469 19672
rect 6503 19669 6515 19703
rect 7742 19700 7748 19712
rect 7703 19672 7748 19700
rect 6457 19663 6515 19669
rect 7742 19660 7748 19672
rect 7800 19660 7806 19712
rect 8018 19700 8024 19712
rect 7979 19672 8024 19700
rect 8018 19660 8024 19672
rect 8076 19660 8082 19712
rect 8754 19660 8760 19712
rect 8812 19700 8818 19712
rect 9033 19703 9091 19709
rect 9033 19700 9045 19703
rect 8812 19672 9045 19700
rect 8812 19660 8818 19672
rect 9033 19669 9045 19672
rect 9079 19669 9091 19703
rect 9968 19700 9996 19740
rect 15105 19737 15117 19771
rect 15151 19768 15163 19771
rect 15304 19768 15332 19796
rect 15151 19740 15332 19768
rect 15151 19737 15163 19740
rect 15105 19731 15163 19737
rect 11793 19703 11851 19709
rect 11793 19700 11805 19703
rect 9968 19672 11805 19700
rect 9033 19663 9091 19669
rect 11793 19669 11805 19672
rect 11839 19669 11851 19703
rect 11793 19663 11851 19669
rect 12434 19660 12440 19712
rect 12492 19700 12498 19712
rect 12529 19703 12587 19709
rect 12529 19700 12541 19703
rect 12492 19672 12541 19700
rect 12492 19660 12498 19672
rect 12529 19669 12541 19672
rect 12575 19669 12587 19703
rect 12894 19700 12900 19712
rect 12855 19672 12900 19700
rect 12529 19663 12587 19669
rect 12894 19660 12900 19672
rect 12952 19660 12958 19712
rect 14366 19660 14372 19712
rect 14424 19700 14430 19712
rect 14645 19703 14703 19709
rect 14645 19700 14657 19703
rect 14424 19672 14657 19700
rect 14424 19660 14430 19672
rect 14645 19669 14657 19672
rect 14691 19669 14703 19703
rect 14645 19663 14703 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 7929 19499 7987 19505
rect 7929 19465 7941 19499
rect 7975 19496 7987 19499
rect 8386 19496 8392 19508
rect 7975 19468 8392 19496
rect 7975 19465 7987 19468
rect 7929 19459 7987 19465
rect 8386 19456 8392 19468
rect 8444 19456 8450 19508
rect 10962 19496 10968 19508
rect 10923 19468 10968 19496
rect 10962 19456 10968 19468
rect 11020 19456 11026 19508
rect 12526 19496 12532 19508
rect 12487 19468 12532 19496
rect 12526 19456 12532 19468
rect 12584 19456 12590 19508
rect 13538 19496 13544 19508
rect 13499 19468 13544 19496
rect 13538 19456 13544 19468
rect 13596 19456 13602 19508
rect 15286 19456 15292 19508
rect 15344 19456 15350 19508
rect 15562 19456 15568 19508
rect 15620 19496 15626 19508
rect 15749 19499 15807 19505
rect 15749 19496 15761 19499
rect 15620 19468 15761 19496
rect 15620 19456 15626 19468
rect 15749 19465 15761 19468
rect 15795 19465 15807 19499
rect 15749 19459 15807 19465
rect 15304 19428 15332 19456
rect 16301 19431 16359 19437
rect 16301 19428 16313 19431
rect 15304 19400 16313 19428
rect 16301 19397 16313 19400
rect 16347 19397 16359 19431
rect 16301 19391 16359 19397
rect 3142 19320 3148 19372
rect 3200 19360 3206 19372
rect 4249 19363 4307 19369
rect 3200 19332 4108 19360
rect 3200 19320 3206 19332
rect 2041 19295 2099 19301
rect 2041 19261 2053 19295
rect 2087 19292 2099 19295
rect 2130 19292 2136 19304
rect 2087 19264 2136 19292
rect 2087 19261 2099 19264
rect 2041 19255 2099 19261
rect 2130 19252 2136 19264
rect 2188 19252 2194 19304
rect 4080 19292 4108 19332
rect 4249 19329 4261 19363
rect 4295 19360 4307 19363
rect 5350 19360 5356 19372
rect 4295 19332 5356 19360
rect 4295 19329 4307 19332
rect 4249 19323 4307 19329
rect 5350 19320 5356 19332
rect 5408 19360 5414 19372
rect 5537 19363 5595 19369
rect 5537 19360 5549 19363
rect 5408 19332 5549 19360
rect 5408 19320 5414 19332
rect 5537 19329 5549 19332
rect 5583 19360 5595 19363
rect 5997 19363 6055 19369
rect 5997 19360 6009 19363
rect 5583 19332 6009 19360
rect 5583 19329 5595 19332
rect 5537 19323 5595 19329
rect 5997 19329 6009 19332
rect 6043 19329 6055 19363
rect 5997 19323 6055 19329
rect 9398 19320 9404 19372
rect 9456 19360 9462 19372
rect 9456 19332 9628 19360
rect 9456 19320 9462 19332
rect 4617 19295 4675 19301
rect 4080 19264 4200 19292
rect 2314 19233 2320 19236
rect 1949 19227 2007 19233
rect 1949 19193 1961 19227
rect 1995 19224 2007 19227
rect 2286 19227 2320 19233
rect 2286 19224 2298 19227
rect 1995 19196 2298 19224
rect 1995 19193 2007 19196
rect 1949 19187 2007 19193
rect 2286 19193 2298 19196
rect 2372 19224 2378 19236
rect 2774 19224 2780 19236
rect 2372 19196 2780 19224
rect 2286 19187 2320 19193
rect 2314 19184 2320 19187
rect 2372 19184 2378 19196
rect 2774 19184 2780 19196
rect 2832 19184 2838 19236
rect 4172 19224 4200 19264
rect 4617 19261 4629 19295
rect 4663 19292 4675 19295
rect 4706 19292 4712 19304
rect 4663 19264 4712 19292
rect 4663 19261 4675 19264
rect 4617 19255 4675 19261
rect 4706 19252 4712 19264
rect 4764 19252 4770 19304
rect 4890 19292 4896 19304
rect 4851 19264 4896 19292
rect 4890 19252 4896 19264
rect 4948 19252 4954 19304
rect 4982 19252 4988 19304
rect 5040 19292 5046 19304
rect 5445 19295 5503 19301
rect 5445 19292 5457 19295
rect 5040 19264 5457 19292
rect 5040 19252 5046 19264
rect 5445 19261 5457 19264
rect 5491 19261 5503 19295
rect 5445 19255 5503 19261
rect 8021 19295 8079 19301
rect 8021 19261 8033 19295
rect 8067 19292 8079 19295
rect 8110 19292 8116 19304
rect 8067 19264 8116 19292
rect 8067 19261 8079 19264
rect 8021 19255 8079 19261
rect 8110 19252 8116 19264
rect 8168 19252 8174 19304
rect 9600 19292 9628 19332
rect 10134 19320 10140 19372
rect 10192 19360 10198 19372
rect 10505 19363 10563 19369
rect 10505 19360 10517 19363
rect 10192 19332 10517 19360
rect 10192 19320 10198 19332
rect 10505 19329 10517 19332
rect 10551 19329 10563 19363
rect 10505 19323 10563 19329
rect 12434 19320 12440 19372
rect 12492 19360 12498 19372
rect 13173 19363 13231 19369
rect 13173 19360 13185 19363
rect 12492 19332 13185 19360
rect 12492 19320 12498 19332
rect 13173 19329 13185 19332
rect 13219 19360 13231 19363
rect 14366 19360 14372 19372
rect 13219 19332 13768 19360
rect 14327 19332 14372 19360
rect 13219 19329 13231 19332
rect 13173 19323 13231 19329
rect 10321 19295 10379 19301
rect 10321 19292 10333 19295
rect 9600 19264 10333 19292
rect 10321 19261 10333 19264
rect 10367 19261 10379 19295
rect 10321 19255 10379 19261
rect 11330 19252 11336 19304
rect 11388 19292 11394 19304
rect 11701 19295 11759 19301
rect 11701 19292 11713 19295
rect 11388 19264 11713 19292
rect 11388 19252 11394 19264
rect 11701 19261 11713 19264
rect 11747 19261 11759 19295
rect 11701 19255 11759 19261
rect 11974 19252 11980 19304
rect 12032 19292 12038 19304
rect 12161 19295 12219 19301
rect 12161 19292 12173 19295
rect 12032 19264 12173 19292
rect 12032 19252 12038 19264
rect 12161 19261 12173 19264
rect 12207 19292 12219 19295
rect 12710 19292 12716 19304
rect 12207 19264 12716 19292
rect 12207 19261 12219 19264
rect 12161 19255 12219 19261
rect 12710 19252 12716 19264
rect 12768 19292 12774 19304
rect 12897 19295 12955 19301
rect 12897 19292 12909 19295
rect 12768 19264 12909 19292
rect 12768 19252 12774 19264
rect 12897 19261 12909 19264
rect 12943 19261 12955 19295
rect 13740 19292 13768 19332
rect 14366 19320 14372 19332
rect 14424 19320 14430 19372
rect 13740 19264 14320 19292
rect 12897 19255 12955 19261
rect 7466 19224 7472 19236
rect 4172 19196 5028 19224
rect 3421 19159 3479 19165
rect 3421 19125 3433 19159
rect 3467 19156 3479 19159
rect 4522 19156 4528 19168
rect 3467 19128 4528 19156
rect 3467 19125 3479 19128
rect 3421 19119 3479 19125
rect 4522 19116 4528 19128
rect 4580 19116 4586 19168
rect 4614 19116 4620 19168
rect 4672 19156 4678 19168
rect 5000 19165 5028 19196
rect 5368 19196 7472 19224
rect 4709 19159 4767 19165
rect 4709 19156 4721 19159
rect 4672 19128 4721 19156
rect 4672 19116 4678 19128
rect 4709 19125 4721 19128
rect 4755 19125 4767 19159
rect 4709 19119 4767 19125
rect 4985 19159 5043 19165
rect 4985 19125 4997 19159
rect 5031 19125 5043 19159
rect 4985 19119 5043 19125
rect 5258 19116 5264 19168
rect 5316 19156 5322 19168
rect 5368 19165 5396 19196
rect 7466 19184 7472 19196
rect 7524 19184 7530 19236
rect 7742 19184 7748 19236
rect 7800 19224 7806 19236
rect 8288 19227 8346 19233
rect 8288 19224 8300 19227
rect 7800 19196 8300 19224
rect 7800 19184 7806 19196
rect 8288 19193 8300 19196
rect 8334 19224 8346 19227
rect 8938 19224 8944 19236
rect 8334 19196 8944 19224
rect 8334 19193 8346 19196
rect 8288 19187 8346 19193
rect 8938 19184 8944 19196
rect 8996 19184 9002 19236
rect 11425 19227 11483 19233
rect 11425 19193 11437 19227
rect 11471 19224 11483 19227
rect 12526 19224 12532 19236
rect 11471 19196 12532 19224
rect 11471 19193 11483 19196
rect 11425 19187 11483 19193
rect 12526 19184 12532 19196
rect 12584 19184 12590 19236
rect 14292 19233 14320 19264
rect 14277 19227 14335 19233
rect 14277 19193 14289 19227
rect 14323 19224 14335 19227
rect 14636 19227 14694 19233
rect 14636 19224 14648 19227
rect 14323 19196 14648 19224
rect 14323 19193 14335 19196
rect 14277 19187 14335 19193
rect 14636 19193 14648 19196
rect 14682 19224 14694 19227
rect 14734 19224 14740 19236
rect 14682 19196 14740 19224
rect 14682 19193 14694 19196
rect 14636 19187 14694 19193
rect 14734 19184 14740 19196
rect 14792 19184 14798 19236
rect 5353 19159 5411 19165
rect 5353 19156 5365 19159
rect 5316 19128 5365 19156
rect 5316 19116 5322 19128
rect 5353 19125 5365 19128
rect 5399 19125 5411 19159
rect 6362 19156 6368 19168
rect 6323 19128 6368 19156
rect 5353 19119 5411 19125
rect 6362 19116 6368 19128
rect 6420 19116 6426 19168
rect 7006 19156 7012 19168
rect 6967 19128 7012 19156
rect 7006 19116 7012 19128
rect 7064 19116 7070 19168
rect 8386 19116 8392 19168
rect 8444 19156 8450 19168
rect 9401 19159 9459 19165
rect 9401 19156 9413 19159
rect 8444 19128 9413 19156
rect 8444 19116 8450 19128
rect 9401 19125 9413 19128
rect 9447 19125 9459 19159
rect 9401 19119 9459 19125
rect 9766 19116 9772 19168
rect 9824 19156 9830 19168
rect 9953 19159 10011 19165
rect 9953 19156 9965 19159
rect 9824 19128 9965 19156
rect 9824 19116 9830 19128
rect 9953 19125 9965 19128
rect 9999 19125 10011 19159
rect 9953 19119 10011 19125
rect 11517 19159 11575 19165
rect 11517 19125 11529 19159
rect 11563 19156 11575 19159
rect 12158 19156 12164 19168
rect 11563 19128 12164 19156
rect 11563 19125 11575 19128
rect 11517 19119 11575 19125
rect 12158 19116 12164 19128
rect 12216 19116 12222 19168
rect 12986 19116 12992 19168
rect 13044 19156 13050 19168
rect 13044 19128 13089 19156
rect 13044 19116 13050 19128
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1486 18912 1492 18964
rect 1544 18952 1550 18964
rect 1581 18955 1639 18961
rect 1581 18952 1593 18955
rect 1544 18924 1593 18952
rect 1544 18912 1550 18924
rect 1581 18921 1593 18924
rect 1627 18921 1639 18955
rect 2038 18952 2044 18964
rect 1999 18924 2044 18952
rect 1581 18915 1639 18921
rect 2038 18912 2044 18924
rect 2096 18912 2102 18964
rect 4062 18912 4068 18964
rect 4120 18952 4126 18964
rect 4709 18955 4767 18961
rect 4709 18952 4721 18955
rect 4120 18924 4721 18952
rect 4120 18912 4126 18924
rect 4709 18921 4721 18924
rect 4755 18952 4767 18955
rect 5350 18952 5356 18964
rect 4755 18924 5356 18952
rect 4755 18921 4767 18924
rect 4709 18915 4767 18921
rect 5350 18912 5356 18924
rect 5408 18952 5414 18964
rect 6362 18952 6368 18964
rect 5408 18924 6368 18952
rect 5408 18912 5414 18924
rect 6362 18912 6368 18924
rect 6420 18912 6426 18964
rect 7742 18952 7748 18964
rect 7703 18924 7748 18952
rect 7742 18912 7748 18924
rect 7800 18912 7806 18964
rect 8018 18912 8024 18964
rect 8076 18952 8082 18964
rect 8297 18955 8355 18961
rect 8297 18952 8309 18955
rect 8076 18924 8309 18952
rect 8076 18912 8082 18924
rect 8297 18921 8309 18924
rect 8343 18921 8355 18955
rect 8938 18952 8944 18964
rect 8899 18924 8944 18952
rect 8297 18915 8355 18921
rect 8938 18912 8944 18924
rect 8996 18912 9002 18964
rect 11330 18952 11336 18964
rect 11291 18924 11336 18952
rect 11330 18912 11336 18924
rect 11388 18912 11394 18964
rect 11425 18955 11483 18961
rect 11425 18921 11437 18955
rect 11471 18952 11483 18955
rect 12342 18952 12348 18964
rect 11471 18924 12348 18952
rect 11471 18921 11483 18924
rect 11425 18915 11483 18921
rect 12342 18912 12348 18924
rect 12400 18912 12406 18964
rect 12529 18955 12587 18961
rect 12529 18921 12541 18955
rect 12575 18952 12587 18955
rect 12986 18952 12992 18964
rect 12575 18924 12992 18952
rect 12575 18921 12587 18924
rect 12529 18915 12587 18921
rect 12986 18912 12992 18924
rect 13044 18912 13050 18964
rect 13446 18952 13452 18964
rect 13407 18924 13452 18952
rect 13446 18912 13452 18924
rect 13504 18912 13510 18964
rect 15562 18952 15568 18964
rect 15523 18924 15568 18952
rect 15562 18912 15568 18924
rect 15620 18912 15626 18964
rect 5442 18884 5448 18896
rect 5276 18856 5448 18884
rect 2038 18776 2044 18828
rect 2096 18816 2102 18828
rect 2222 18816 2228 18828
rect 2096 18788 2228 18816
rect 2096 18776 2102 18788
rect 2222 18776 2228 18788
rect 2280 18776 2286 18828
rect 2593 18819 2651 18825
rect 2593 18785 2605 18819
rect 2639 18816 2651 18819
rect 3694 18816 3700 18828
rect 2639 18788 3700 18816
rect 2639 18785 2651 18788
rect 2593 18779 2651 18785
rect 3694 18776 3700 18788
rect 3752 18776 3758 18828
rect 4065 18819 4123 18825
rect 4065 18785 4077 18819
rect 4111 18816 4123 18819
rect 4154 18816 4160 18828
rect 4111 18788 4160 18816
rect 4111 18785 4123 18788
rect 4065 18779 4123 18785
rect 4154 18776 4160 18788
rect 4212 18776 4218 18828
rect 4614 18776 4620 18828
rect 4672 18816 4678 18828
rect 5276 18825 5304 18856
rect 5442 18844 5448 18856
rect 5500 18844 5506 18896
rect 7006 18844 7012 18896
rect 7064 18884 7070 18896
rect 7834 18884 7840 18896
rect 7064 18856 7840 18884
rect 7064 18844 7070 18856
rect 7834 18844 7840 18856
rect 7892 18884 7898 18896
rect 8205 18887 8263 18893
rect 8205 18884 8217 18887
rect 7892 18856 8217 18884
rect 7892 18844 7898 18856
rect 8205 18853 8217 18856
rect 8251 18853 8263 18887
rect 11885 18887 11943 18893
rect 11885 18884 11897 18887
rect 8205 18847 8263 18853
rect 11440 18856 11897 18884
rect 11440 18828 11468 18856
rect 11885 18853 11897 18856
rect 11931 18853 11943 18887
rect 11885 18847 11943 18853
rect 5261 18819 5319 18825
rect 5261 18816 5273 18819
rect 4672 18788 5273 18816
rect 4672 18776 4678 18788
rect 5261 18785 5273 18788
rect 5307 18785 5319 18819
rect 5261 18779 5319 18785
rect 5528 18819 5586 18825
rect 5528 18785 5540 18819
rect 5574 18816 5586 18819
rect 6086 18816 6092 18828
rect 5574 18788 6092 18816
rect 5574 18785 5586 18788
rect 5528 18779 5586 18785
rect 6086 18776 6092 18788
rect 6144 18816 6150 18828
rect 7193 18819 7251 18825
rect 7193 18816 7205 18819
rect 6144 18788 7205 18816
rect 6144 18776 6150 18788
rect 7193 18785 7205 18788
rect 7239 18816 7251 18819
rect 7374 18816 7380 18828
rect 7239 18788 7380 18816
rect 7239 18785 7251 18788
rect 7193 18779 7251 18785
rect 7374 18776 7380 18788
rect 7432 18776 7438 18828
rect 9950 18816 9956 18828
rect 9911 18788 9956 18816
rect 9950 18776 9956 18788
rect 10008 18776 10014 18828
rect 11422 18776 11428 18828
rect 11480 18776 11486 18828
rect 11790 18816 11796 18828
rect 11751 18788 11796 18816
rect 11790 18776 11796 18788
rect 11848 18776 11854 18828
rect 13262 18776 13268 18828
rect 13320 18816 13326 18828
rect 13357 18819 13415 18825
rect 13357 18816 13369 18819
rect 13320 18788 13369 18816
rect 13320 18776 13326 18788
rect 13357 18785 13369 18788
rect 13403 18816 13415 18819
rect 13906 18816 13912 18828
rect 13403 18788 13912 18816
rect 13403 18785 13415 18788
rect 13357 18779 13415 18785
rect 13906 18776 13912 18788
rect 13964 18776 13970 18828
rect 2682 18748 2688 18760
rect 2643 18720 2688 18748
rect 2682 18708 2688 18720
rect 2740 18708 2746 18760
rect 2774 18708 2780 18760
rect 2832 18748 2838 18760
rect 2869 18751 2927 18757
rect 2869 18748 2881 18751
rect 2832 18720 2881 18748
rect 2832 18708 2838 18720
rect 2869 18717 2881 18720
rect 2915 18748 2927 18751
rect 3602 18748 3608 18760
rect 2915 18720 3608 18748
rect 2915 18717 2927 18720
rect 2869 18711 2927 18717
rect 3602 18708 3608 18720
rect 3660 18708 3666 18760
rect 8202 18708 8208 18760
rect 8260 18748 8266 18760
rect 8389 18751 8447 18757
rect 8389 18748 8401 18751
rect 8260 18720 8401 18748
rect 8260 18708 8266 18720
rect 8389 18717 8401 18720
rect 8435 18717 8447 18751
rect 10134 18748 10140 18760
rect 10095 18720 10140 18748
rect 8389 18711 8447 18717
rect 10134 18708 10140 18720
rect 10192 18708 10198 18760
rect 11974 18748 11980 18760
rect 11935 18720 11980 18748
rect 11974 18708 11980 18720
rect 12032 18748 12038 18760
rect 12434 18748 12440 18760
rect 12032 18720 12440 18748
rect 12032 18708 12038 18720
rect 12434 18708 12440 18720
rect 12492 18708 12498 18760
rect 13541 18751 13599 18757
rect 13541 18717 13553 18751
rect 13587 18717 13599 18751
rect 13541 18711 13599 18717
rect 3326 18680 3332 18692
rect 3287 18652 3332 18680
rect 3326 18640 3332 18652
rect 3384 18640 3390 18692
rect 6914 18640 6920 18692
rect 6972 18680 6978 18692
rect 7837 18683 7895 18689
rect 7837 18680 7849 18683
rect 6972 18652 7849 18680
rect 6972 18640 6978 18652
rect 7837 18649 7849 18652
rect 7883 18649 7895 18683
rect 13556 18680 13584 18711
rect 13630 18680 13636 18692
rect 7837 18643 7895 18649
rect 12820 18652 13636 18680
rect 2222 18612 2228 18624
rect 2183 18584 2228 18612
rect 2222 18572 2228 18584
rect 2280 18572 2286 18624
rect 3694 18612 3700 18624
rect 3655 18584 3700 18612
rect 3694 18572 3700 18584
rect 3752 18572 3758 18624
rect 4246 18612 4252 18624
rect 4207 18584 4252 18612
rect 4246 18572 4252 18584
rect 4304 18572 4310 18624
rect 4430 18572 4436 18624
rect 4488 18612 4494 18624
rect 4985 18615 5043 18621
rect 4985 18612 4997 18615
rect 4488 18584 4997 18612
rect 4488 18572 4494 18584
rect 4985 18581 4997 18584
rect 5031 18612 5043 18615
rect 5258 18612 5264 18624
rect 5031 18584 5264 18612
rect 5031 18581 5043 18584
rect 4985 18575 5043 18581
rect 5258 18572 5264 18584
rect 5316 18572 5322 18624
rect 6638 18612 6644 18624
rect 6599 18584 6644 18612
rect 6638 18572 6644 18584
rect 6696 18572 6702 18624
rect 9214 18612 9220 18624
rect 9175 18584 9220 18612
rect 9214 18572 9220 18584
rect 9272 18572 9278 18624
rect 10134 18572 10140 18624
rect 10192 18612 10198 18624
rect 10689 18615 10747 18621
rect 10689 18612 10701 18615
rect 10192 18584 10701 18612
rect 10192 18572 10198 18584
rect 10689 18581 10701 18584
rect 10735 18581 10747 18615
rect 10689 18575 10747 18581
rect 12618 18572 12624 18624
rect 12676 18612 12682 18624
rect 12820 18621 12848 18652
rect 13630 18640 13636 18652
rect 13688 18680 13694 18692
rect 14001 18683 14059 18689
rect 14001 18680 14013 18683
rect 13688 18652 14013 18680
rect 13688 18640 13694 18652
rect 14001 18649 14013 18652
rect 14047 18649 14059 18683
rect 14001 18643 14059 18649
rect 12805 18615 12863 18621
rect 12805 18612 12817 18615
rect 12676 18584 12817 18612
rect 12676 18572 12682 18584
rect 12805 18581 12817 18584
rect 12851 18581 12863 18615
rect 14366 18612 14372 18624
rect 14327 18584 14372 18612
rect 12805 18575 12863 18581
rect 14366 18572 14372 18584
rect 14424 18612 14430 18624
rect 14737 18615 14795 18621
rect 14737 18612 14749 18615
rect 14424 18584 14749 18612
rect 14424 18572 14430 18584
rect 14737 18581 14749 18584
rect 14783 18581 14795 18615
rect 14737 18575 14795 18581
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 3602 18408 3608 18420
rect 3563 18380 3608 18408
rect 3602 18368 3608 18380
rect 3660 18368 3666 18420
rect 4522 18408 4528 18420
rect 4483 18380 4528 18408
rect 4522 18368 4528 18380
rect 4580 18368 4586 18420
rect 6546 18408 6552 18420
rect 6507 18380 6552 18408
rect 6546 18368 6552 18380
rect 6604 18368 6610 18420
rect 7834 18408 7840 18420
rect 7795 18380 7840 18408
rect 7834 18368 7840 18380
rect 7892 18368 7898 18420
rect 8202 18408 8208 18420
rect 8163 18380 8208 18408
rect 8202 18368 8208 18380
rect 8260 18368 8266 18420
rect 9493 18411 9551 18417
rect 9493 18377 9505 18411
rect 9539 18408 9551 18411
rect 9950 18408 9956 18420
rect 9539 18380 9956 18408
rect 9539 18377 9551 18380
rect 9493 18371 9551 18377
rect 9950 18368 9956 18380
rect 10008 18368 10014 18420
rect 11422 18408 11428 18420
rect 11383 18380 11428 18408
rect 11422 18368 11428 18380
rect 11480 18368 11486 18420
rect 11790 18368 11796 18420
rect 11848 18408 11854 18420
rect 12161 18411 12219 18417
rect 12161 18408 12173 18411
rect 11848 18380 12173 18408
rect 11848 18368 11854 18380
rect 12161 18377 12173 18380
rect 12207 18408 12219 18411
rect 12342 18408 12348 18420
rect 12207 18380 12348 18408
rect 12207 18377 12219 18380
rect 12161 18371 12219 18377
rect 12342 18368 12348 18380
rect 12400 18368 12406 18420
rect 13081 18411 13139 18417
rect 13081 18377 13093 18411
rect 13127 18408 13139 18411
rect 13354 18408 13360 18420
rect 13127 18380 13360 18408
rect 13127 18377 13139 18380
rect 13081 18371 13139 18377
rect 13354 18368 13360 18380
rect 13412 18368 13418 18420
rect 14734 18408 14740 18420
rect 14695 18380 14740 18408
rect 14734 18368 14740 18380
rect 14792 18368 14798 18420
rect 4062 18300 4068 18352
rect 4120 18340 4126 18352
rect 4540 18340 4568 18368
rect 6825 18343 6883 18349
rect 4120 18312 5304 18340
rect 4120 18300 4126 18312
rect 2222 18272 2228 18284
rect 2183 18244 2228 18272
rect 2222 18232 2228 18244
rect 2280 18232 2286 18284
rect 4246 18272 4252 18284
rect 4207 18244 4252 18272
rect 4246 18232 4252 18244
rect 4304 18232 4310 18284
rect 5166 18272 5172 18284
rect 5127 18244 5172 18272
rect 5166 18232 5172 18244
rect 5224 18232 5230 18284
rect 5276 18281 5304 18312
rect 6825 18309 6837 18343
rect 6871 18309 6883 18343
rect 6825 18303 6883 18309
rect 11149 18343 11207 18349
rect 11149 18309 11161 18343
rect 11195 18340 11207 18343
rect 11974 18340 11980 18352
rect 11195 18312 11980 18340
rect 11195 18309 11207 18312
rect 11149 18303 11207 18309
rect 5261 18275 5319 18281
rect 5261 18241 5273 18275
rect 5307 18241 5319 18275
rect 5261 18235 5319 18241
rect 1578 18164 1584 18216
rect 1636 18204 1642 18216
rect 6181 18207 6239 18213
rect 6181 18204 6193 18207
rect 1636 18176 6193 18204
rect 1636 18164 1642 18176
rect 6181 18173 6193 18176
rect 6227 18173 6239 18207
rect 6840 18204 6868 18303
rect 11974 18300 11980 18312
rect 12032 18300 12038 18352
rect 7374 18272 7380 18284
rect 7335 18244 7380 18272
rect 7374 18232 7380 18244
rect 7432 18232 7438 18284
rect 8478 18232 8484 18284
rect 8536 18272 8542 18284
rect 8941 18275 8999 18281
rect 8941 18272 8953 18275
rect 8536 18244 8953 18272
rect 8536 18232 8542 18244
rect 8941 18241 8953 18244
rect 8987 18241 8999 18275
rect 8941 18235 8999 18241
rect 9674 18232 9680 18284
rect 9732 18272 9738 18284
rect 9861 18275 9919 18281
rect 9861 18272 9873 18275
rect 9732 18244 9873 18272
rect 9732 18232 9738 18244
rect 9861 18241 9873 18244
rect 9907 18272 9919 18275
rect 10505 18275 10563 18281
rect 10505 18272 10517 18275
rect 9907 18244 10517 18272
rect 9907 18241 9919 18244
rect 9861 18235 9919 18241
rect 10505 18241 10517 18244
rect 10551 18241 10563 18275
rect 10505 18235 10563 18241
rect 8849 18207 8907 18213
rect 8849 18204 8861 18207
rect 6840 18176 8861 18204
rect 6181 18167 6239 18173
rect 8849 18173 8861 18176
rect 8895 18204 8907 18207
rect 9214 18204 9220 18216
rect 8895 18176 9220 18204
rect 8895 18173 8907 18176
rect 8849 18167 8907 18173
rect 2133 18139 2191 18145
rect 2133 18105 2145 18139
rect 2179 18136 2191 18139
rect 2492 18139 2550 18145
rect 2492 18136 2504 18139
rect 2179 18108 2504 18136
rect 2179 18105 2191 18108
rect 2133 18099 2191 18105
rect 2492 18105 2504 18108
rect 2538 18136 2550 18139
rect 2590 18136 2596 18148
rect 2538 18108 2596 18136
rect 2538 18105 2550 18108
rect 2492 18099 2550 18105
rect 2590 18096 2596 18108
rect 2648 18096 2654 18148
rect 6196 18136 6224 18167
rect 9214 18164 9220 18176
rect 9272 18164 9278 18216
rect 9766 18164 9772 18216
rect 9824 18204 9830 18216
rect 10321 18207 10379 18213
rect 10321 18204 10333 18207
rect 9824 18176 10333 18204
rect 9824 18164 9830 18176
rect 10321 18173 10333 18176
rect 10367 18173 10379 18207
rect 10321 18167 10379 18173
rect 11885 18207 11943 18213
rect 11885 18173 11897 18207
rect 11931 18204 11943 18207
rect 12158 18204 12164 18216
rect 11931 18176 12164 18204
rect 11931 18173 11943 18176
rect 11885 18167 11943 18173
rect 12158 18164 12164 18176
rect 12216 18164 12222 18216
rect 13354 18204 13360 18216
rect 12360 18176 13360 18204
rect 7193 18139 7251 18145
rect 7193 18136 7205 18139
rect 6196 18108 7205 18136
rect 7193 18105 7205 18108
rect 7239 18136 7251 18139
rect 7742 18136 7748 18148
rect 7239 18108 7748 18136
rect 7239 18105 7251 18108
rect 7193 18099 7251 18105
rect 7742 18096 7748 18108
rect 7800 18096 7806 18148
rect 12360 18136 12388 18176
rect 13354 18164 13360 18176
rect 13412 18164 13418 18216
rect 13630 18213 13636 18216
rect 13624 18204 13636 18213
rect 13591 18176 13636 18204
rect 13624 18167 13636 18176
rect 13630 18164 13636 18167
rect 13688 18164 13694 18216
rect 11716 18108 12388 18136
rect 11716 18080 11744 18108
rect 1394 18028 1400 18080
rect 1452 18068 1458 18080
rect 1581 18071 1639 18077
rect 1581 18068 1593 18071
rect 1452 18040 1593 18068
rect 1452 18028 1458 18040
rect 1581 18037 1593 18040
rect 1627 18037 1639 18071
rect 1581 18031 1639 18037
rect 1946 18028 1952 18080
rect 2004 18068 2010 18080
rect 2774 18068 2780 18080
rect 2004 18040 2780 18068
rect 2004 18028 2010 18040
rect 2774 18028 2780 18040
rect 2832 18028 2838 18080
rect 4706 18068 4712 18080
rect 4667 18040 4712 18068
rect 4706 18028 4712 18040
rect 4764 18028 4770 18080
rect 5074 18068 5080 18080
rect 5035 18040 5080 18068
rect 5074 18028 5080 18040
rect 5132 18028 5138 18080
rect 5813 18071 5871 18077
rect 5813 18037 5825 18071
rect 5859 18068 5871 18071
rect 6086 18068 6092 18080
rect 5859 18040 6092 18068
rect 5859 18037 5871 18040
rect 5813 18031 5871 18037
rect 6086 18028 6092 18040
rect 6144 18028 6150 18080
rect 6546 18028 6552 18080
rect 6604 18068 6610 18080
rect 7098 18068 7104 18080
rect 6604 18040 7104 18068
rect 6604 18028 6610 18040
rect 7098 18028 7104 18040
rect 7156 18068 7162 18080
rect 7285 18071 7343 18077
rect 7285 18068 7297 18071
rect 7156 18040 7297 18068
rect 7156 18028 7162 18040
rect 7285 18037 7297 18040
rect 7331 18037 7343 18071
rect 8386 18068 8392 18080
rect 8347 18040 8392 18068
rect 7285 18031 7343 18037
rect 8386 18028 8392 18040
rect 8444 18028 8450 18080
rect 8754 18068 8760 18080
rect 8715 18040 8760 18068
rect 8754 18028 8760 18040
rect 8812 18028 8818 18080
rect 9950 18068 9956 18080
rect 9911 18040 9956 18068
rect 9950 18028 9956 18040
rect 10008 18028 10014 18080
rect 10134 18028 10140 18080
rect 10192 18068 10198 18080
rect 10413 18071 10471 18077
rect 10413 18068 10425 18071
rect 10192 18040 10425 18068
rect 10192 18028 10198 18040
rect 10413 18037 10425 18040
rect 10459 18037 10471 18071
rect 11698 18068 11704 18080
rect 11659 18040 11704 18068
rect 10413 18031 10471 18037
rect 11698 18028 11704 18040
rect 11756 18028 11762 18080
rect 12713 18071 12771 18077
rect 12713 18037 12725 18071
rect 12759 18068 12771 18071
rect 12802 18068 12808 18080
rect 12759 18040 12808 18068
rect 12759 18037 12771 18040
rect 12713 18031 12771 18037
rect 12802 18028 12808 18040
rect 12860 18028 12866 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 2314 17864 2320 17876
rect 2275 17836 2320 17864
rect 2314 17824 2320 17836
rect 2372 17824 2378 17876
rect 2409 17867 2467 17873
rect 2409 17833 2421 17867
rect 2455 17864 2467 17867
rect 2682 17864 2688 17876
rect 2455 17836 2688 17864
rect 2455 17833 2467 17836
rect 2409 17827 2467 17833
rect 2682 17824 2688 17836
rect 2740 17864 2746 17876
rect 3421 17867 3479 17873
rect 3421 17864 3433 17867
rect 2740 17836 3433 17864
rect 2740 17824 2746 17836
rect 3421 17833 3433 17836
rect 3467 17833 3479 17867
rect 3421 17827 3479 17833
rect 3694 17824 3700 17876
rect 3752 17864 3758 17876
rect 4065 17867 4123 17873
rect 4065 17864 4077 17867
rect 3752 17836 4077 17864
rect 3752 17824 3758 17836
rect 4065 17833 4077 17836
rect 4111 17833 4123 17867
rect 5166 17864 5172 17876
rect 5127 17836 5172 17864
rect 4065 17827 4123 17833
rect 5166 17824 5172 17836
rect 5224 17824 5230 17876
rect 7929 17867 7987 17873
rect 7929 17833 7941 17867
rect 7975 17864 7987 17867
rect 8018 17864 8024 17876
rect 7975 17836 8024 17864
rect 7975 17833 7987 17836
rect 7929 17827 7987 17833
rect 8018 17824 8024 17836
rect 8076 17824 8082 17876
rect 8478 17864 8484 17876
rect 8439 17836 8484 17864
rect 8478 17824 8484 17836
rect 8536 17824 8542 17876
rect 12434 17824 12440 17876
rect 12492 17864 12498 17876
rect 13725 17867 13783 17873
rect 13725 17864 13737 17867
rect 12492 17836 13737 17864
rect 12492 17824 12498 17836
rect 13725 17833 13737 17836
rect 13771 17833 13783 17867
rect 13725 17827 13783 17833
rect 2774 17756 2780 17808
rect 2832 17796 2838 17808
rect 2832 17768 2877 17796
rect 2832 17756 2838 17768
rect 5534 17756 5540 17808
rect 5592 17796 5598 17808
rect 5592 17768 5948 17796
rect 5592 17756 5598 17768
rect 4338 17688 4344 17740
rect 4396 17728 4402 17740
rect 5920 17737 5948 17768
rect 5994 17756 6000 17808
rect 6052 17796 6058 17808
rect 6172 17799 6230 17805
rect 6172 17796 6184 17799
rect 6052 17768 6184 17796
rect 6052 17756 6058 17768
rect 6172 17765 6184 17768
rect 6218 17796 6230 17799
rect 6638 17796 6644 17808
rect 6218 17768 6644 17796
rect 6218 17765 6230 17768
rect 6172 17759 6230 17765
rect 6638 17756 6644 17768
rect 6696 17756 6702 17808
rect 9858 17756 9864 17808
rect 9916 17796 9922 17808
rect 11698 17796 11704 17808
rect 9916 17768 11704 17796
rect 9916 17756 9922 17768
rect 4433 17731 4491 17737
rect 4433 17728 4445 17731
rect 4396 17700 4445 17728
rect 4396 17688 4402 17700
rect 4433 17697 4445 17700
rect 4479 17697 4491 17731
rect 4433 17691 4491 17697
rect 5905 17731 5963 17737
rect 5905 17697 5917 17731
rect 5951 17728 5963 17731
rect 7374 17728 7380 17740
rect 5951 17700 7380 17728
rect 5951 17697 5963 17700
rect 5905 17691 5963 17697
rect 7374 17688 7380 17700
rect 7432 17688 7438 17740
rect 9125 17731 9183 17737
rect 9125 17697 9137 17731
rect 9171 17728 9183 17731
rect 10042 17728 10048 17740
rect 9171 17700 10048 17728
rect 9171 17697 9183 17700
rect 9125 17691 9183 17697
rect 10042 17688 10048 17700
rect 10100 17688 10106 17740
rect 11256 17737 11284 17768
rect 11698 17756 11704 17768
rect 11756 17756 11762 17808
rect 13354 17756 13360 17808
rect 13412 17796 13418 17808
rect 14185 17799 14243 17805
rect 14185 17796 14197 17799
rect 13412 17768 14197 17796
rect 13412 17756 13418 17768
rect 14185 17765 14197 17768
rect 14231 17796 14243 17799
rect 14366 17796 14372 17808
rect 14231 17768 14372 17796
rect 14231 17765 14243 17768
rect 14185 17759 14243 17765
rect 14366 17756 14372 17768
rect 14424 17796 14430 17808
rect 14829 17799 14887 17805
rect 14829 17796 14841 17799
rect 14424 17768 14841 17796
rect 14424 17756 14430 17768
rect 14829 17765 14841 17768
rect 14875 17765 14887 17799
rect 14829 17759 14887 17765
rect 11514 17737 11520 17740
rect 11241 17731 11299 17737
rect 11241 17697 11253 17731
rect 11287 17697 11299 17731
rect 11508 17728 11520 17737
rect 11475 17700 11520 17728
rect 11241 17691 11299 17697
rect 11508 17691 11520 17700
rect 11514 17688 11520 17691
rect 11572 17688 11578 17740
rect 1397 17663 1455 17669
rect 1397 17629 1409 17663
rect 1443 17660 1455 17663
rect 1762 17660 1768 17672
rect 1443 17632 1768 17660
rect 1443 17629 1455 17632
rect 1397 17623 1455 17629
rect 1762 17620 1768 17632
rect 1820 17660 1826 17672
rect 1857 17663 1915 17669
rect 1857 17660 1869 17663
rect 1820 17632 1869 17660
rect 1820 17620 1826 17632
rect 1857 17629 1869 17632
rect 1903 17629 1915 17663
rect 1857 17623 1915 17629
rect 1946 17620 1952 17672
rect 2004 17660 2010 17672
rect 2869 17663 2927 17669
rect 2869 17660 2881 17663
rect 2004 17632 2881 17660
rect 2004 17620 2010 17632
rect 2869 17629 2881 17632
rect 2915 17629 2927 17663
rect 3050 17660 3056 17672
rect 3011 17632 3056 17660
rect 2869 17623 2927 17629
rect 3050 17620 3056 17632
rect 3108 17620 3114 17672
rect 3326 17620 3332 17672
rect 3384 17660 3390 17672
rect 4525 17663 4583 17669
rect 4525 17660 4537 17663
rect 3384 17632 4537 17660
rect 3384 17620 3390 17632
rect 4525 17629 4537 17632
rect 4571 17629 4583 17663
rect 4706 17660 4712 17672
rect 4667 17632 4712 17660
rect 4525 17623 4583 17629
rect 4706 17620 4712 17632
rect 4764 17620 4770 17672
rect 5534 17660 5540 17672
rect 5495 17632 5540 17660
rect 5534 17620 5540 17632
rect 5592 17620 5598 17672
rect 8570 17660 8576 17672
rect 8531 17632 8576 17660
rect 8570 17620 8576 17632
rect 8628 17620 8634 17672
rect 9493 17663 9551 17669
rect 9493 17629 9505 17663
rect 9539 17660 9551 17663
rect 10134 17660 10140 17672
rect 9539 17632 10140 17660
rect 9539 17629 9551 17632
rect 9493 17623 9551 17629
rect 10134 17620 10140 17632
rect 10192 17620 10198 17672
rect 10226 17620 10232 17672
rect 10284 17660 10290 17672
rect 10284 17632 10329 17660
rect 10284 17620 10290 17632
rect 2590 17552 2596 17604
rect 2648 17592 2654 17604
rect 3068 17592 3096 17620
rect 12618 17592 12624 17604
rect 2648 17564 3096 17592
rect 12579 17564 12624 17592
rect 2648 17552 2654 17564
rect 12618 17552 12624 17564
rect 12676 17552 12682 17604
rect 3786 17524 3792 17536
rect 3747 17496 3792 17524
rect 3786 17484 3792 17496
rect 3844 17484 3850 17536
rect 7282 17524 7288 17536
rect 7243 17496 7288 17524
rect 7282 17484 7288 17496
rect 7340 17484 7346 17536
rect 9674 17524 9680 17536
rect 9635 17496 9680 17524
rect 9674 17484 9680 17496
rect 9732 17484 9738 17536
rect 10870 17524 10876 17536
rect 10831 17496 10876 17524
rect 10870 17484 10876 17496
rect 10928 17484 10934 17536
rect 13357 17527 13415 17533
rect 13357 17493 13369 17527
rect 13403 17524 13415 17527
rect 13814 17524 13820 17536
rect 13403 17496 13820 17524
rect 13403 17493 13415 17496
rect 13357 17487 13415 17493
rect 13814 17484 13820 17496
rect 13872 17484 13878 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1397 17323 1455 17329
rect 1397 17289 1409 17323
rect 1443 17320 1455 17323
rect 2498 17320 2504 17332
rect 1443 17292 2504 17320
rect 1443 17289 1455 17292
rect 1397 17283 1455 17289
rect 2498 17280 2504 17292
rect 2556 17280 2562 17332
rect 3050 17280 3056 17332
rect 3108 17320 3114 17332
rect 3329 17323 3387 17329
rect 3329 17320 3341 17323
rect 3108 17292 3341 17320
rect 3108 17280 3114 17292
rect 3329 17289 3341 17292
rect 3375 17320 3387 17323
rect 4706 17320 4712 17332
rect 3375 17292 4712 17320
rect 3375 17289 3387 17292
rect 3329 17283 3387 17289
rect 4706 17280 4712 17292
rect 4764 17280 4770 17332
rect 5994 17320 6000 17332
rect 5955 17292 6000 17320
rect 5994 17280 6000 17292
rect 6052 17280 6058 17332
rect 9769 17323 9827 17329
rect 9769 17289 9781 17323
rect 9815 17320 9827 17323
rect 10226 17320 10232 17332
rect 9815 17292 10232 17320
rect 9815 17289 9827 17292
rect 9769 17283 9827 17289
rect 10226 17280 10232 17292
rect 10284 17320 10290 17332
rect 11241 17323 11299 17329
rect 11241 17320 11253 17323
rect 10284 17292 11253 17320
rect 10284 17280 10290 17292
rect 11241 17289 11253 17292
rect 11287 17320 11299 17323
rect 11514 17320 11520 17332
rect 11287 17292 11520 17320
rect 11287 17289 11299 17292
rect 11241 17283 11299 17289
rect 11514 17280 11520 17292
rect 11572 17320 11578 17332
rect 11793 17323 11851 17329
rect 11793 17320 11805 17323
rect 11572 17292 11805 17320
rect 11572 17280 11578 17292
rect 11793 17289 11805 17292
rect 11839 17289 11851 17323
rect 12158 17320 12164 17332
rect 12119 17292 12164 17320
rect 11793 17283 11851 17289
rect 12158 17280 12164 17292
rect 12216 17280 12222 17332
rect 13262 17320 13268 17332
rect 13223 17292 13268 17320
rect 13262 17280 13268 17292
rect 13320 17280 13326 17332
rect 14366 17320 14372 17332
rect 14327 17292 14372 17320
rect 14366 17280 14372 17292
rect 14424 17280 14430 17332
rect 1946 17212 1952 17264
rect 2004 17252 2010 17264
rect 2409 17255 2467 17261
rect 2409 17252 2421 17255
rect 2004 17224 2421 17252
rect 2004 17212 2010 17224
rect 2409 17221 2421 17224
rect 2455 17221 2467 17255
rect 2409 17215 2467 17221
rect 3234 17212 3240 17264
rect 3292 17252 3298 17264
rect 3605 17255 3663 17261
rect 3605 17252 3617 17255
rect 3292 17224 3617 17252
rect 3292 17212 3298 17224
rect 3605 17221 3617 17224
rect 3651 17221 3663 17255
rect 3605 17215 3663 17221
rect 8478 17212 8484 17264
rect 8536 17252 8542 17264
rect 8757 17255 8815 17261
rect 8757 17252 8769 17255
rect 8536 17224 8769 17252
rect 8536 17212 8542 17224
rect 8757 17221 8769 17224
rect 8803 17221 8815 17255
rect 8757 17215 8815 17221
rect 2038 17184 2044 17196
rect 1951 17156 2044 17184
rect 2038 17144 2044 17156
rect 2096 17184 2102 17196
rect 2314 17184 2320 17196
rect 2096 17156 2320 17184
rect 2096 17144 2102 17156
rect 2314 17144 2320 17156
rect 2372 17144 2378 17196
rect 3418 17144 3424 17196
rect 3476 17184 3482 17196
rect 3789 17187 3847 17193
rect 3789 17184 3801 17187
rect 3476 17156 3801 17184
rect 3476 17144 3482 17156
rect 3789 17153 3801 17156
rect 3835 17153 3847 17187
rect 3789 17147 3847 17153
rect 7285 17187 7343 17193
rect 7285 17153 7297 17187
rect 7331 17184 7343 17187
rect 9858 17184 9864 17196
rect 7331 17156 7512 17184
rect 9819 17156 9864 17184
rect 7331 17153 7343 17156
rect 7285 17147 7343 17153
rect 1762 17116 1768 17128
rect 1723 17088 1768 17116
rect 1762 17076 1768 17088
rect 1820 17076 1826 17128
rect 4062 17125 4068 17128
rect 4056 17116 4068 17125
rect 4023 17088 4068 17116
rect 4056 17079 4068 17088
rect 4062 17076 4068 17079
rect 4120 17076 4126 17128
rect 7374 17116 7380 17128
rect 7335 17088 7380 17116
rect 7374 17076 7380 17088
rect 7432 17076 7438 17128
rect 7484 17116 7512 17156
rect 9858 17144 9864 17156
rect 9916 17144 9922 17196
rect 13814 17184 13820 17196
rect 13775 17156 13820 17184
rect 13814 17144 13820 17156
rect 13872 17184 13878 17196
rect 14645 17187 14703 17193
rect 14645 17184 14657 17187
rect 13872 17156 14657 17184
rect 13872 17144 13878 17156
rect 14645 17153 14657 17156
rect 14691 17184 14703 17187
rect 14691 17156 14964 17184
rect 14691 17153 14703 17156
rect 14645 17147 14703 17153
rect 7650 17125 7656 17128
rect 7644 17116 7656 17125
rect 7484 17088 7656 17116
rect 7644 17079 7656 17088
rect 7650 17076 7656 17079
rect 7708 17076 7714 17128
rect 13173 17119 13231 17125
rect 13173 17085 13185 17119
rect 13219 17116 13231 17119
rect 13722 17116 13728 17128
rect 13219 17088 13728 17116
rect 13219 17085 13231 17088
rect 13173 17079 13231 17085
rect 13722 17076 13728 17088
rect 13780 17076 13786 17128
rect 14366 17076 14372 17128
rect 14424 17116 14430 17128
rect 14829 17119 14887 17125
rect 14829 17116 14841 17119
rect 14424 17088 14841 17116
rect 14424 17076 14430 17088
rect 14829 17085 14841 17088
rect 14875 17085 14887 17119
rect 14936 17116 14964 17156
rect 15085 17119 15143 17125
rect 15085 17116 15097 17119
rect 14936 17088 15097 17116
rect 14829 17079 14887 17085
rect 15085 17085 15097 17088
rect 15131 17116 15143 17119
rect 15131 17085 15148 17116
rect 15085 17079 15148 17085
rect 2130 17008 2136 17060
rect 2188 17048 2194 17060
rect 6730 17048 6736 17060
rect 2188 17020 6736 17048
rect 2188 17008 2194 17020
rect 6730 17008 6736 17020
rect 6788 17008 6794 17060
rect 9401 17051 9459 17057
rect 9401 17017 9413 17051
rect 9447 17048 9459 17051
rect 10128 17051 10186 17057
rect 10128 17048 10140 17051
rect 9447 17020 10140 17048
rect 9447 17017 9459 17020
rect 9401 17011 9459 17017
rect 10128 17017 10140 17020
rect 10174 17048 10186 17051
rect 10778 17048 10784 17060
rect 10174 17020 10784 17048
rect 10174 17017 10186 17020
rect 10128 17011 10186 17017
rect 10778 17008 10784 17020
rect 10836 17008 10842 17060
rect 15120 17048 15148 17079
rect 15286 17048 15292 17060
rect 15120 17020 15292 17048
rect 15286 17008 15292 17020
rect 15344 17008 15350 17060
rect 1854 16980 1860 16992
rect 1815 16952 1860 16980
rect 1854 16940 1860 16952
rect 1912 16940 1918 16992
rect 2774 16980 2780 16992
rect 2735 16952 2780 16980
rect 2774 16940 2780 16952
rect 2832 16940 2838 16992
rect 5169 16983 5227 16989
rect 5169 16949 5181 16983
rect 5215 16980 5227 16983
rect 5258 16980 5264 16992
rect 5215 16952 5264 16980
rect 5215 16949 5227 16952
rect 5169 16943 5227 16949
rect 5258 16940 5264 16952
rect 5316 16940 5322 16992
rect 6270 16980 6276 16992
rect 6231 16952 6276 16980
rect 6270 16940 6276 16952
rect 6328 16940 6334 16992
rect 12434 16940 12440 16992
rect 12492 16980 12498 16992
rect 12621 16983 12679 16989
rect 12621 16980 12633 16983
rect 12492 16952 12633 16980
rect 12492 16940 12498 16952
rect 12621 16949 12633 16952
rect 12667 16949 12679 16983
rect 12621 16943 12679 16949
rect 13170 16940 13176 16992
rect 13228 16980 13234 16992
rect 13633 16983 13691 16989
rect 13633 16980 13645 16983
rect 13228 16952 13645 16980
rect 13228 16940 13234 16952
rect 13633 16949 13645 16952
rect 13679 16949 13691 16983
rect 16206 16980 16212 16992
rect 16167 16952 16212 16980
rect 13633 16943 13691 16949
rect 16206 16940 16212 16952
rect 16264 16940 16270 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1486 16736 1492 16788
rect 1544 16776 1550 16788
rect 1673 16779 1731 16785
rect 1673 16776 1685 16779
rect 1544 16748 1685 16776
rect 1544 16736 1550 16748
rect 1673 16745 1685 16748
rect 1719 16776 1731 16779
rect 1854 16776 1860 16788
rect 1719 16748 1860 16776
rect 1719 16745 1731 16748
rect 1673 16739 1731 16745
rect 1854 16736 1860 16748
rect 1912 16736 1918 16788
rect 2038 16776 2044 16788
rect 1999 16748 2044 16776
rect 2038 16736 2044 16748
rect 2096 16736 2102 16788
rect 2133 16779 2191 16785
rect 2133 16745 2145 16779
rect 2179 16776 2191 16779
rect 2498 16776 2504 16788
rect 2179 16748 2504 16776
rect 2179 16745 2191 16748
rect 2133 16739 2191 16745
rect 2498 16736 2504 16748
rect 2556 16736 2562 16788
rect 3050 16736 3056 16788
rect 3108 16776 3114 16788
rect 3145 16779 3203 16785
rect 3145 16776 3157 16779
rect 3108 16748 3157 16776
rect 3108 16736 3114 16748
rect 3145 16745 3157 16748
rect 3191 16745 3203 16779
rect 3145 16739 3203 16745
rect 3881 16779 3939 16785
rect 3881 16745 3893 16779
rect 3927 16776 3939 16779
rect 4062 16776 4068 16788
rect 3927 16748 4068 16776
rect 3927 16745 3939 16748
rect 3881 16739 3939 16745
rect 4062 16736 4068 16748
rect 4120 16736 4126 16788
rect 4709 16779 4767 16785
rect 4709 16745 4721 16779
rect 4755 16776 4767 16779
rect 6270 16776 6276 16788
rect 4755 16748 6276 16776
rect 4755 16745 4767 16748
rect 4709 16739 4767 16745
rect 6270 16736 6276 16748
rect 6328 16736 6334 16788
rect 6730 16776 6736 16788
rect 6691 16748 6736 16776
rect 6730 16736 6736 16748
rect 6788 16736 6794 16788
rect 7377 16779 7435 16785
rect 7377 16745 7389 16779
rect 7423 16776 7435 16779
rect 8386 16776 8392 16788
rect 7423 16748 8392 16776
rect 7423 16745 7435 16748
rect 7377 16739 7435 16745
rect 8386 16736 8392 16748
rect 8444 16736 8450 16788
rect 8570 16736 8576 16788
rect 8628 16776 8634 16788
rect 9953 16779 10011 16785
rect 9953 16776 9965 16779
rect 8628 16748 9965 16776
rect 8628 16736 8634 16748
rect 9953 16745 9965 16748
rect 9999 16745 10011 16779
rect 9953 16739 10011 16745
rect 2222 16668 2228 16720
rect 2280 16708 2286 16720
rect 2593 16711 2651 16717
rect 2593 16708 2605 16711
rect 2280 16680 2605 16708
rect 2280 16668 2286 16680
rect 2593 16677 2605 16680
rect 2639 16677 2651 16711
rect 2593 16671 2651 16677
rect 5813 16711 5871 16717
rect 5813 16677 5825 16711
rect 5859 16708 5871 16711
rect 5994 16708 6000 16720
rect 5859 16680 6000 16708
rect 5859 16677 5871 16680
rect 5813 16671 5871 16677
rect 5994 16668 6000 16680
rect 6052 16668 6058 16720
rect 6086 16668 6092 16720
rect 6144 16708 6150 16720
rect 8297 16711 8355 16717
rect 8297 16708 8309 16711
rect 6144 16680 6776 16708
rect 6144 16668 6150 16680
rect 2406 16600 2412 16652
rect 2464 16640 2470 16652
rect 2501 16643 2559 16649
rect 2501 16640 2513 16643
rect 2464 16612 2513 16640
rect 2464 16600 2470 16612
rect 2501 16609 2513 16612
rect 2547 16640 2559 16643
rect 3786 16640 3792 16652
rect 2547 16612 3792 16640
rect 2547 16609 2559 16612
rect 2501 16603 2559 16609
rect 3786 16600 3792 16612
rect 3844 16600 3850 16652
rect 4338 16640 4344 16652
rect 4299 16612 4344 16640
rect 4338 16600 4344 16612
rect 4396 16600 4402 16652
rect 5074 16640 5080 16652
rect 5035 16612 5080 16640
rect 5074 16600 5080 16612
rect 5132 16600 5138 16652
rect 2590 16532 2596 16584
rect 2648 16572 2654 16584
rect 2685 16575 2743 16581
rect 2685 16572 2697 16575
rect 2648 16544 2697 16572
rect 2648 16532 2654 16544
rect 2685 16541 2697 16544
rect 2731 16541 2743 16575
rect 2685 16535 2743 16541
rect 4982 16532 4988 16584
rect 5040 16572 5046 16584
rect 5169 16575 5227 16581
rect 5169 16572 5181 16575
rect 5040 16544 5181 16572
rect 5040 16532 5046 16544
rect 5169 16541 5181 16544
rect 5215 16541 5227 16575
rect 5169 16535 5227 16541
rect 5258 16532 5264 16584
rect 5316 16572 5322 16584
rect 6104 16581 6132 16668
rect 6454 16640 6460 16652
rect 6288 16612 6460 16640
rect 6089 16575 6147 16581
rect 6089 16572 6101 16575
rect 5316 16544 6101 16572
rect 5316 16532 5322 16544
rect 6089 16541 6101 16544
rect 6135 16541 6147 16575
rect 6089 16535 6147 16541
rect 3878 16464 3884 16516
rect 3936 16504 3942 16516
rect 5276 16504 5304 16532
rect 6288 16513 6316 16612
rect 6454 16600 6460 16612
rect 6512 16600 6518 16652
rect 6641 16643 6699 16649
rect 6641 16609 6653 16643
rect 6687 16609 6699 16643
rect 6748 16640 6776 16680
rect 7668 16680 8309 16708
rect 7668 16652 7696 16680
rect 8297 16677 8309 16680
rect 8343 16677 8355 16711
rect 8404 16708 8432 16736
rect 9125 16711 9183 16717
rect 9125 16708 9137 16711
rect 8404 16680 9137 16708
rect 8297 16671 8355 16677
rect 9125 16677 9137 16680
rect 9171 16677 9183 16711
rect 9968 16708 9996 16739
rect 10042 16736 10048 16788
rect 10100 16776 10106 16788
rect 10137 16779 10195 16785
rect 10137 16776 10149 16779
rect 10100 16748 10149 16776
rect 10100 16736 10106 16748
rect 10137 16745 10149 16748
rect 10183 16745 10195 16779
rect 10137 16739 10195 16745
rect 11241 16779 11299 16785
rect 11241 16745 11253 16779
rect 11287 16776 11299 16779
rect 11606 16776 11612 16788
rect 11287 16748 11612 16776
rect 11287 16745 11299 16748
rect 11241 16739 11299 16745
rect 10505 16711 10563 16717
rect 10505 16708 10517 16711
rect 9968 16680 10517 16708
rect 9125 16671 9183 16677
rect 10505 16677 10517 16680
rect 10551 16677 10563 16711
rect 10505 16671 10563 16677
rect 7650 16640 7656 16652
rect 6748 16612 6868 16640
rect 7611 16612 7656 16640
rect 6641 16603 6699 16609
rect 3936 16476 5304 16504
rect 6273 16507 6331 16513
rect 3936 16464 3942 16476
rect 6273 16473 6285 16507
rect 6319 16473 6331 16507
rect 6273 16467 6331 16473
rect 3510 16396 3516 16448
rect 3568 16436 3574 16448
rect 6656 16436 6684 16603
rect 6840 16581 6868 16612
rect 7650 16600 7656 16612
rect 7708 16600 7714 16652
rect 7834 16600 7840 16652
rect 7892 16600 7898 16652
rect 8202 16640 8208 16652
rect 8163 16612 8208 16640
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 8754 16640 8760 16652
rect 8680 16612 8760 16640
rect 6825 16575 6883 16581
rect 6825 16541 6837 16575
rect 6871 16541 6883 16575
rect 6825 16535 6883 16541
rect 7852 16513 7880 16600
rect 8110 16532 8116 16584
rect 8168 16572 8174 16584
rect 8389 16575 8447 16581
rect 8389 16572 8401 16575
rect 8168 16544 8401 16572
rect 8168 16532 8174 16544
rect 8389 16541 8401 16544
rect 8435 16541 8447 16575
rect 8389 16535 8447 16541
rect 8680 16513 8708 16612
rect 8754 16600 8760 16612
rect 8812 16600 8818 16652
rect 9030 16640 9036 16652
rect 8991 16612 9036 16640
rect 9030 16600 9036 16612
rect 9088 16600 9094 16652
rect 10597 16643 10655 16649
rect 10597 16609 10609 16643
rect 10643 16640 10655 16643
rect 10686 16640 10692 16652
rect 10643 16612 10692 16640
rect 10643 16609 10655 16612
rect 10597 16603 10655 16609
rect 10686 16600 10692 16612
rect 10744 16600 10750 16652
rect 9214 16572 9220 16584
rect 9175 16544 9220 16572
rect 9214 16532 9220 16544
rect 9272 16532 9278 16584
rect 10778 16572 10784 16584
rect 10691 16544 10784 16572
rect 10778 16532 10784 16544
rect 10836 16572 10842 16584
rect 11256 16572 11284 16739
rect 11606 16736 11612 16748
rect 11664 16736 11670 16788
rect 12250 16736 12256 16788
rect 12308 16776 12314 16788
rect 12437 16779 12495 16785
rect 12437 16776 12449 16779
rect 12308 16748 12449 16776
rect 12308 16736 12314 16748
rect 12437 16745 12449 16748
rect 12483 16745 12495 16779
rect 12437 16739 12495 16745
rect 11422 16668 11428 16720
rect 11480 16708 11486 16720
rect 12529 16711 12587 16717
rect 12529 16708 12541 16711
rect 11480 16680 12541 16708
rect 11480 16668 11486 16680
rect 12529 16677 12541 16680
rect 12575 16677 12587 16711
rect 12529 16671 12587 16677
rect 13170 16668 13176 16720
rect 13228 16708 13234 16720
rect 13265 16711 13323 16717
rect 13265 16708 13277 16711
rect 13228 16680 13277 16708
rect 13228 16668 13234 16680
rect 13265 16677 13277 16680
rect 13311 16677 13323 16711
rect 14182 16708 14188 16720
rect 14143 16680 14188 16708
rect 13265 16671 13323 16677
rect 14182 16668 14188 16680
rect 14240 16668 14246 16720
rect 13906 16640 13912 16652
rect 13867 16612 13912 16640
rect 13906 16600 13912 16612
rect 13964 16600 13970 16652
rect 10836 16544 11284 16572
rect 12713 16575 12771 16581
rect 10836 16532 10842 16544
rect 12713 16541 12725 16575
rect 12759 16572 12771 16575
rect 13262 16572 13268 16584
rect 12759 16544 13268 16572
rect 12759 16541 12771 16544
rect 12713 16535 12771 16541
rect 13262 16532 13268 16544
rect 13320 16532 13326 16584
rect 7837 16507 7895 16513
rect 7837 16473 7849 16507
rect 7883 16473 7895 16507
rect 7837 16467 7895 16473
rect 8665 16507 8723 16513
rect 8665 16473 8677 16507
rect 8711 16473 8723 16507
rect 8665 16467 8723 16473
rect 11330 16464 11336 16516
rect 11388 16504 11394 16516
rect 12069 16507 12127 16513
rect 12069 16504 12081 16507
rect 11388 16476 12081 16504
rect 11388 16464 11394 16476
rect 12069 16473 12081 16476
rect 12115 16473 12127 16507
rect 12069 16467 12127 16473
rect 7190 16436 7196 16448
rect 3568 16408 7196 16436
rect 3568 16396 3574 16408
rect 7190 16396 7196 16408
rect 7248 16396 7254 16448
rect 11882 16436 11888 16448
rect 11843 16408 11888 16436
rect 11882 16396 11888 16408
rect 11940 16396 11946 16448
rect 13725 16439 13783 16445
rect 13725 16405 13737 16439
rect 13771 16436 13783 16439
rect 13814 16436 13820 16448
rect 13771 16408 13820 16436
rect 13771 16405 13783 16408
rect 13725 16399 13783 16405
rect 13814 16396 13820 16408
rect 13872 16436 13878 16448
rect 14734 16436 14740 16448
rect 13872 16408 14740 16436
rect 13872 16396 13878 16408
rect 14734 16396 14740 16408
rect 14792 16396 14798 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 1578 16232 1584 16244
rect 1539 16204 1584 16232
rect 1578 16192 1584 16204
rect 1636 16192 1642 16244
rect 5166 16232 5172 16244
rect 5127 16204 5172 16232
rect 5166 16192 5172 16204
rect 5224 16192 5230 16244
rect 6365 16235 6423 16241
rect 6365 16201 6377 16235
rect 6411 16232 6423 16235
rect 6730 16232 6736 16244
rect 6411 16204 6736 16232
rect 6411 16201 6423 16204
rect 6365 16195 6423 16201
rect 6730 16192 6736 16204
rect 6788 16192 6794 16244
rect 7190 16192 7196 16244
rect 7248 16232 7254 16244
rect 7285 16235 7343 16241
rect 7285 16232 7297 16235
rect 7248 16204 7297 16232
rect 7248 16192 7254 16204
rect 7285 16201 7297 16204
rect 7331 16201 7343 16235
rect 7285 16195 7343 16201
rect 10134 16192 10140 16244
rect 10192 16232 10198 16244
rect 10781 16235 10839 16241
rect 10781 16232 10793 16235
rect 10192 16204 10793 16232
rect 10192 16192 10198 16204
rect 10781 16201 10793 16204
rect 10827 16201 10839 16235
rect 10781 16195 10839 16201
rect 11422 16192 11428 16244
rect 11480 16232 11486 16244
rect 12069 16235 12127 16241
rect 12069 16232 12081 16235
rect 11480 16204 12081 16232
rect 11480 16192 11486 16204
rect 12069 16201 12081 16204
rect 12115 16201 12127 16235
rect 12069 16195 12127 16201
rect 15197 16235 15255 16241
rect 15197 16201 15209 16235
rect 15243 16232 15255 16235
rect 15286 16232 15292 16244
rect 15243 16204 15292 16232
rect 15243 16201 15255 16204
rect 15197 16195 15255 16201
rect 15286 16192 15292 16204
rect 15344 16192 15350 16244
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16096 5871 16099
rect 5994 16096 6000 16108
rect 5859 16068 6000 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 5994 16056 6000 16068
rect 6052 16056 6058 16108
rect 11238 16096 11244 16108
rect 11199 16068 11244 16096
rect 11238 16056 11244 16068
rect 11296 16056 11302 16108
rect 11425 16099 11483 16105
rect 11425 16065 11437 16099
rect 11471 16096 11483 16099
rect 11606 16096 11612 16108
rect 11471 16068 11612 16096
rect 11471 16065 11483 16068
rect 11425 16059 11483 16065
rect 11606 16056 11612 16068
rect 11664 16056 11670 16108
rect 12526 16056 12532 16108
rect 12584 16096 12590 16108
rect 12621 16099 12679 16105
rect 12621 16096 12633 16099
rect 12584 16068 12633 16096
rect 12584 16056 12590 16068
rect 12621 16065 12633 16068
rect 12667 16065 12679 16099
rect 13814 16096 13820 16108
rect 13775 16068 13820 16096
rect 12621 16059 12679 16065
rect 13814 16056 13820 16068
rect 13872 16056 13878 16108
rect 16574 16096 16580 16108
rect 16535 16068 16580 16096
rect 16574 16056 16580 16068
rect 16632 16056 16638 16108
rect 1394 16028 1400 16040
rect 1355 16000 1400 16028
rect 1394 15988 1400 16000
rect 1452 15988 1458 16040
rect 1578 15988 1584 16040
rect 1636 16028 1642 16040
rect 2685 16031 2743 16037
rect 2685 16028 2697 16031
rect 1636 16000 2697 16028
rect 1636 15988 1642 16000
rect 2685 15997 2697 16000
rect 2731 16028 2743 16031
rect 2731 16000 3096 16028
rect 2731 15997 2743 16000
rect 2685 15991 2743 15997
rect 2930 15963 2988 15969
rect 2930 15960 2942 15963
rect 2608 15932 2942 15960
rect 2608 15904 2636 15932
rect 2930 15929 2942 15932
rect 2976 15929 2988 15963
rect 3068 15960 3096 16000
rect 4154 15988 4160 16040
rect 4212 16028 4218 16040
rect 4709 16031 4767 16037
rect 4709 16028 4721 16031
rect 4212 16000 4721 16028
rect 4212 15988 4218 16000
rect 4709 15997 4721 16000
rect 4755 16028 4767 16031
rect 5074 16028 5080 16040
rect 4755 16000 5080 16028
rect 4755 15997 4767 16000
rect 4709 15991 4767 15997
rect 5074 15988 5080 16000
rect 5132 15988 5138 16040
rect 5629 16031 5687 16037
rect 5629 15997 5641 16031
rect 5675 16028 5687 16031
rect 6270 16028 6276 16040
rect 5675 16000 6276 16028
rect 5675 15997 5687 16000
rect 5629 15991 5687 15997
rect 6270 15988 6276 16000
rect 6328 15988 6334 16040
rect 7926 15988 7932 16040
rect 7984 16028 7990 16040
rect 10689 16031 10747 16037
rect 7984 16000 9352 16028
rect 7984 15988 7990 16000
rect 3068 15932 4200 15960
rect 2930 15923 2988 15929
rect 4172 15904 4200 15932
rect 5258 15920 5264 15972
rect 5316 15960 5322 15972
rect 5537 15963 5595 15969
rect 5537 15960 5549 15963
rect 5316 15932 5549 15960
rect 5316 15920 5322 15932
rect 5537 15929 5549 15932
rect 5583 15960 5595 15963
rect 6825 15963 6883 15969
rect 6825 15960 6837 15963
rect 5583 15932 6837 15960
rect 5583 15929 5595 15932
rect 5537 15923 5595 15929
rect 6825 15929 6837 15932
rect 6871 15929 6883 15963
rect 6825 15923 6883 15929
rect 8297 15963 8355 15969
rect 8297 15929 8309 15963
rect 8343 15960 8355 15963
rect 8389 15963 8447 15969
rect 8389 15960 8401 15963
rect 8343 15932 8401 15960
rect 8343 15929 8355 15932
rect 8297 15923 8355 15929
rect 8389 15929 8401 15932
rect 8435 15960 8447 15963
rect 8478 15960 8484 15972
rect 8435 15932 8484 15960
rect 8435 15929 8447 15932
rect 8389 15923 8447 15929
rect 8478 15920 8484 15932
rect 8536 15920 8542 15972
rect 9324 15904 9352 16000
rect 10689 15997 10701 16031
rect 10735 16028 10747 16031
rect 11149 16031 11207 16037
rect 11149 16028 11161 16031
rect 10735 16000 11161 16028
rect 10735 15997 10747 16000
rect 10689 15991 10747 15997
rect 11149 15997 11161 16000
rect 11195 16028 11207 16031
rect 11514 16028 11520 16040
rect 11195 16000 11520 16028
rect 11195 15997 11207 16000
rect 11149 15991 11207 15997
rect 11514 15988 11520 16000
rect 11572 15988 11578 16040
rect 12434 15988 12440 16040
rect 12492 16028 12498 16040
rect 16298 16028 16304 16040
rect 12492 16000 12537 16028
rect 16259 16000 16304 16028
rect 12492 15988 12498 16000
rect 16298 15988 16304 16000
rect 16356 16028 16362 16040
rect 17037 16031 17095 16037
rect 17037 16028 17049 16031
rect 16356 16000 17049 16028
rect 16356 15988 16362 16000
rect 17037 15997 17049 16000
rect 17083 15997 17095 16031
rect 17037 15991 17095 15997
rect 14062 15963 14120 15969
rect 14062 15960 14074 15963
rect 13648 15932 14074 15960
rect 13648 15904 13676 15932
rect 14062 15929 14074 15932
rect 14108 15929 14120 15963
rect 14062 15923 14120 15929
rect 2038 15892 2044 15904
rect 1999 15864 2044 15892
rect 2038 15852 2044 15864
rect 2096 15852 2102 15904
rect 2409 15895 2467 15901
rect 2409 15861 2421 15895
rect 2455 15892 2467 15895
rect 2590 15892 2596 15904
rect 2455 15864 2596 15892
rect 2455 15861 2467 15864
rect 2409 15855 2467 15861
rect 2590 15852 2596 15864
rect 2648 15852 2654 15904
rect 4062 15892 4068 15904
rect 4023 15864 4068 15892
rect 4062 15852 4068 15864
rect 4120 15852 4126 15904
rect 4154 15852 4160 15904
rect 4212 15852 4218 15904
rect 7929 15895 7987 15901
rect 7929 15861 7941 15895
rect 7975 15892 7987 15895
rect 8110 15892 8116 15904
rect 7975 15864 8116 15892
rect 7975 15861 7987 15864
rect 7929 15855 7987 15861
rect 8110 15852 8116 15864
rect 8168 15852 8174 15904
rect 9306 15852 9312 15904
rect 9364 15892 9370 15904
rect 9677 15895 9735 15901
rect 9677 15892 9689 15895
rect 9364 15864 9689 15892
rect 9364 15852 9370 15864
rect 9677 15861 9689 15864
rect 9723 15861 9735 15895
rect 13262 15892 13268 15904
rect 13223 15864 13268 15892
rect 9677 15855 9735 15861
rect 13262 15852 13268 15864
rect 13320 15852 13326 15904
rect 13630 15892 13636 15904
rect 13591 15864 13636 15892
rect 13630 15852 13636 15864
rect 13688 15852 13694 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 3878 15688 3884 15700
rect 3839 15660 3884 15688
rect 3878 15648 3884 15660
rect 3936 15648 3942 15700
rect 4246 15688 4252 15700
rect 4207 15660 4252 15688
rect 4246 15648 4252 15660
rect 4304 15648 4310 15700
rect 5258 15688 5264 15700
rect 5219 15660 5264 15688
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 7006 15648 7012 15700
rect 7064 15688 7070 15700
rect 7377 15691 7435 15697
rect 7377 15688 7389 15691
rect 7064 15660 7389 15688
rect 7064 15648 7070 15660
rect 7377 15657 7389 15660
rect 7423 15688 7435 15691
rect 8202 15688 8208 15700
rect 7423 15660 8208 15688
rect 7423 15657 7435 15660
rect 7377 15651 7435 15657
rect 8202 15648 8208 15660
rect 8260 15648 8266 15700
rect 10962 15688 10968 15700
rect 10923 15660 10968 15688
rect 10962 15648 10968 15660
rect 11020 15648 11026 15700
rect 11425 15691 11483 15697
rect 11425 15657 11437 15691
rect 11471 15688 11483 15691
rect 11882 15688 11888 15700
rect 11471 15660 11888 15688
rect 11471 15657 11483 15660
rect 11425 15651 11483 15657
rect 11882 15648 11888 15660
rect 11940 15688 11946 15700
rect 12342 15688 12348 15700
rect 11940 15660 12348 15688
rect 11940 15648 11946 15660
rect 12342 15648 12348 15660
rect 12400 15648 12406 15700
rect 13906 15648 13912 15700
rect 13964 15688 13970 15700
rect 14461 15691 14519 15697
rect 14461 15688 14473 15691
rect 13964 15660 14473 15688
rect 13964 15648 13970 15660
rect 14461 15657 14473 15660
rect 14507 15657 14519 15691
rect 14461 15651 14519 15657
rect 14734 15648 14740 15700
rect 14792 15688 14798 15700
rect 14829 15691 14887 15697
rect 14829 15688 14841 15691
rect 14792 15660 14841 15688
rect 14792 15648 14798 15660
rect 14829 15657 14841 15660
rect 14875 15657 14887 15691
rect 15746 15688 15752 15700
rect 15707 15660 15752 15688
rect 14829 15651 14887 15657
rect 15746 15648 15752 15660
rect 15804 15648 15810 15700
rect 5620 15623 5678 15629
rect 5620 15589 5632 15623
rect 5666 15620 5678 15623
rect 6178 15620 6184 15632
rect 5666 15592 6184 15620
rect 5666 15589 5678 15592
rect 5620 15583 5678 15589
rect 6178 15580 6184 15592
rect 6236 15620 6242 15632
rect 7282 15620 7288 15632
rect 6236 15592 7288 15620
rect 6236 15580 6242 15592
rect 7282 15580 7288 15592
rect 7340 15620 7346 15632
rect 7745 15623 7803 15629
rect 7745 15620 7757 15623
rect 7340 15592 7757 15620
rect 7340 15580 7346 15592
rect 7745 15589 7757 15592
rect 7791 15620 7803 15623
rect 9214 15620 9220 15632
rect 7791 15592 9220 15620
rect 7791 15589 7803 15592
rect 7745 15583 7803 15589
rect 9214 15580 9220 15592
rect 9272 15580 9278 15632
rect 13630 15620 13636 15632
rect 12452 15592 13636 15620
rect 1489 15555 1547 15561
rect 1489 15521 1501 15555
rect 1535 15552 1547 15555
rect 1578 15552 1584 15564
rect 1535 15524 1584 15552
rect 1535 15521 1547 15524
rect 1489 15515 1547 15521
rect 1578 15512 1584 15524
rect 1636 15512 1642 15564
rect 1756 15555 1814 15561
rect 1756 15521 1768 15555
rect 1802 15552 1814 15555
rect 2038 15552 2044 15564
rect 1802 15524 2044 15552
rect 1802 15521 1814 15524
rect 1756 15515 1814 15521
rect 2038 15512 2044 15524
rect 2096 15512 2102 15564
rect 3878 15512 3884 15564
rect 3936 15552 3942 15564
rect 4065 15555 4123 15561
rect 4065 15552 4077 15555
rect 3936 15524 4077 15552
rect 3936 15512 3942 15524
rect 4065 15521 4077 15524
rect 4111 15521 4123 15555
rect 4065 15515 4123 15521
rect 4154 15512 4160 15564
rect 4212 15552 4218 15564
rect 5350 15552 5356 15564
rect 4212 15524 5356 15552
rect 4212 15512 4218 15524
rect 5350 15512 5356 15524
rect 5408 15512 5414 15564
rect 7837 15555 7895 15561
rect 7837 15521 7849 15555
rect 7883 15552 7895 15555
rect 7926 15552 7932 15564
rect 7883 15524 7932 15552
rect 7883 15521 7895 15524
rect 7837 15515 7895 15521
rect 7926 15512 7932 15524
rect 7984 15512 7990 15564
rect 8110 15561 8116 15564
rect 8104 15552 8116 15561
rect 8071 15524 8116 15552
rect 8104 15515 8116 15524
rect 8110 15512 8116 15515
rect 8168 15512 8174 15564
rect 9674 15552 9680 15564
rect 9635 15524 9680 15552
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 11330 15552 11336 15564
rect 11291 15524 11336 15552
rect 11330 15512 11336 15524
rect 11388 15512 11394 15564
rect 9858 15484 9864 15496
rect 9819 15456 9864 15484
rect 9858 15444 9864 15456
rect 9916 15444 9922 15496
rect 11609 15487 11667 15493
rect 11609 15453 11621 15487
rect 11655 15484 11667 15487
rect 11882 15484 11888 15496
rect 11655 15456 11888 15484
rect 11655 15453 11667 15456
rect 11609 15447 11667 15453
rect 11882 15444 11888 15456
rect 11940 15484 11946 15496
rect 12452 15484 12480 15592
rect 13630 15580 13636 15592
rect 13688 15620 13694 15632
rect 13688 15592 13952 15620
rect 13688 15580 13694 15592
rect 12529 15555 12587 15561
rect 12529 15521 12541 15555
rect 12575 15552 12587 15555
rect 12618 15552 12624 15564
rect 12575 15524 12624 15552
rect 12575 15521 12587 15524
rect 12529 15515 12587 15521
rect 12618 15512 12624 15524
rect 12676 15512 12682 15564
rect 12796 15555 12854 15561
rect 12796 15521 12808 15555
rect 12842 15552 12854 15555
rect 13262 15552 13268 15564
rect 12842 15524 13268 15552
rect 12842 15521 12854 15524
rect 12796 15515 12854 15521
rect 13262 15512 13268 15524
rect 13320 15512 13326 15564
rect 11940 15456 12480 15484
rect 11940 15444 11946 15456
rect 9217 15419 9275 15425
rect 9217 15385 9229 15419
rect 9263 15416 9275 15419
rect 9490 15416 9496 15428
rect 9263 15388 9496 15416
rect 9263 15385 9275 15388
rect 9217 15379 9275 15385
rect 9490 15376 9496 15388
rect 9548 15376 9554 15428
rect 10870 15416 10876 15428
rect 10831 15388 10876 15416
rect 10870 15376 10876 15388
rect 10928 15376 10934 15428
rect 13924 15425 13952 15592
rect 14366 15580 14372 15632
rect 14424 15620 14430 15632
rect 14752 15620 14780 15648
rect 14424 15592 14780 15620
rect 14424 15580 14430 15592
rect 15654 15552 15660 15564
rect 15615 15524 15660 15552
rect 15654 15512 15660 15524
rect 15712 15512 15718 15564
rect 15378 15444 15384 15496
rect 15436 15484 15442 15496
rect 15933 15487 15991 15493
rect 15933 15484 15945 15487
rect 15436 15456 15945 15484
rect 15436 15444 15442 15456
rect 15933 15453 15945 15456
rect 15979 15484 15991 15487
rect 16482 15484 16488 15496
rect 15979 15456 16488 15484
rect 15979 15453 15991 15456
rect 15933 15447 15991 15453
rect 16482 15444 16488 15456
rect 16540 15444 16546 15496
rect 13909 15419 13967 15425
rect 13909 15385 13921 15419
rect 13955 15385 13967 15419
rect 13909 15379 13967 15385
rect 2590 15308 2596 15360
rect 2648 15348 2654 15360
rect 2869 15351 2927 15357
rect 2869 15348 2881 15351
rect 2648 15320 2881 15348
rect 2648 15308 2654 15320
rect 2869 15317 2881 15320
rect 2915 15348 2927 15351
rect 3421 15351 3479 15357
rect 3421 15348 3433 15351
rect 2915 15320 3433 15348
rect 2915 15317 2927 15320
rect 2869 15311 2927 15317
rect 3421 15317 3433 15320
rect 3467 15317 3479 15351
rect 3421 15311 3479 15317
rect 4801 15351 4859 15357
rect 4801 15317 4813 15351
rect 4847 15348 4859 15351
rect 4982 15348 4988 15360
rect 4847 15320 4988 15348
rect 4847 15317 4859 15320
rect 4801 15311 4859 15317
rect 4982 15308 4988 15320
rect 5040 15348 5046 15360
rect 5350 15348 5356 15360
rect 5040 15320 5356 15348
rect 5040 15308 5046 15320
rect 5350 15308 5356 15320
rect 5408 15308 5414 15360
rect 5534 15308 5540 15360
rect 5592 15348 5598 15360
rect 6733 15351 6791 15357
rect 6733 15348 6745 15351
rect 5592 15320 6745 15348
rect 5592 15308 5598 15320
rect 6733 15317 6745 15320
rect 6779 15317 6791 15351
rect 6733 15311 6791 15317
rect 10505 15351 10563 15357
rect 10505 15317 10517 15351
rect 10551 15348 10563 15351
rect 10686 15348 10692 15360
rect 10551 15320 10692 15348
rect 10551 15317 10563 15320
rect 10505 15311 10563 15317
rect 10686 15308 10692 15320
rect 10744 15308 10750 15360
rect 12161 15351 12219 15357
rect 12161 15317 12173 15351
rect 12207 15348 12219 15351
rect 12250 15348 12256 15360
rect 12207 15320 12256 15348
rect 12207 15317 12219 15320
rect 12161 15311 12219 15317
rect 12250 15308 12256 15320
rect 12308 15348 12314 15360
rect 13446 15348 13452 15360
rect 12308 15320 13452 15348
rect 12308 15308 12314 15320
rect 13446 15308 13452 15320
rect 13504 15308 13510 15360
rect 15286 15348 15292 15360
rect 15247 15320 15292 15348
rect 15286 15308 15292 15320
rect 15344 15308 15350 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 2222 15144 2228 15156
rect 2183 15116 2228 15144
rect 2222 15104 2228 15116
rect 2280 15104 2286 15156
rect 3697 15147 3755 15153
rect 3697 15113 3709 15147
rect 3743 15144 3755 15147
rect 3878 15144 3884 15156
rect 3743 15116 3884 15144
rect 3743 15113 3755 15116
rect 3697 15107 3755 15113
rect 3878 15104 3884 15116
rect 3936 15104 3942 15156
rect 4062 15144 4068 15156
rect 4023 15116 4068 15144
rect 4062 15104 4068 15116
rect 4120 15104 4126 15156
rect 6178 15144 6184 15156
rect 6139 15116 6184 15144
rect 6178 15104 6184 15116
rect 6236 15104 6242 15156
rect 11882 15144 11888 15156
rect 11843 15116 11888 15144
rect 11882 15104 11888 15116
rect 11940 15104 11946 15156
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 12529 15147 12587 15153
rect 12529 15144 12541 15147
rect 12492 15116 12541 15144
rect 12492 15104 12498 15116
rect 12529 15113 12541 15116
rect 12575 15113 12587 15147
rect 12529 15107 12587 15113
rect 13633 15147 13691 15153
rect 13633 15113 13645 15147
rect 13679 15144 13691 15147
rect 15749 15147 15807 15153
rect 15749 15144 15761 15147
rect 13679 15116 15761 15144
rect 13679 15113 13691 15116
rect 13633 15107 13691 15113
rect 15749 15113 15761 15116
rect 15795 15113 15807 15147
rect 15749 15107 15807 15113
rect 2038 14968 2044 15020
rect 2096 15008 2102 15020
rect 2869 15011 2927 15017
rect 2869 15008 2881 15011
rect 2096 14980 2881 15008
rect 2096 14968 2102 14980
rect 2869 14977 2881 14980
rect 2915 15008 2927 15011
rect 2958 15008 2964 15020
rect 2915 14980 2964 15008
rect 2915 14977 2927 14980
rect 2869 14971 2927 14977
rect 2958 14968 2964 14980
rect 3016 15008 3022 15020
rect 4080 15008 4108 15104
rect 6914 15036 6920 15088
rect 6972 15076 6978 15088
rect 7009 15079 7067 15085
rect 7009 15076 7021 15079
rect 6972 15048 7021 15076
rect 6972 15036 6978 15048
rect 7009 15045 7021 15048
rect 7055 15045 7067 15079
rect 7009 15039 7067 15045
rect 8018 15008 8024 15020
rect 3016 14980 3372 15008
rect 4080 14980 4292 15008
rect 7979 14980 8024 15008
rect 3016 14968 3022 14980
rect 2593 14875 2651 14881
rect 2593 14841 2605 14875
rect 2639 14872 2651 14875
rect 2774 14872 2780 14884
rect 2639 14844 2780 14872
rect 2639 14841 2651 14844
rect 2593 14835 2651 14841
rect 2774 14832 2780 14844
rect 2832 14872 2838 14884
rect 3050 14872 3056 14884
rect 2832 14844 3056 14872
rect 2832 14832 2838 14844
rect 3050 14832 3056 14844
rect 3108 14832 3114 14884
rect 3344 14881 3372 14980
rect 4154 14940 4160 14952
rect 4115 14912 4160 14940
rect 4154 14900 4160 14912
rect 4212 14900 4218 14952
rect 4264 14940 4292 14980
rect 8018 14968 8024 14980
rect 8076 14968 8082 15020
rect 10321 15011 10379 15017
rect 10321 14977 10333 15011
rect 10367 15008 10379 15011
rect 11425 15011 11483 15017
rect 11425 15008 11437 15011
rect 10367 14980 11437 15008
rect 10367 14977 10379 14980
rect 10321 14971 10379 14977
rect 11425 14977 11437 14980
rect 11471 15008 11483 15011
rect 11698 15008 11704 15020
rect 11471 14980 11704 15008
rect 11471 14977 11483 14980
rect 11425 14971 11483 14977
rect 11698 14968 11704 14980
rect 11756 14968 11762 15020
rect 11790 14968 11796 15020
rect 11848 15008 11854 15020
rect 12986 15008 12992 15020
rect 11848 14980 12992 15008
rect 11848 14968 11854 14980
rect 12986 14968 12992 14980
rect 13044 14968 13050 15020
rect 13173 15011 13231 15017
rect 13173 14977 13185 15011
rect 13219 15008 13231 15011
rect 13262 15008 13268 15020
rect 13219 14980 13268 15008
rect 13219 14977 13231 14980
rect 13173 14971 13231 14977
rect 13262 14968 13268 14980
rect 13320 15008 13326 15020
rect 13648 15008 13676 15107
rect 16482 15104 16488 15156
rect 16540 15144 16546 15156
rect 16669 15147 16727 15153
rect 16669 15144 16681 15147
rect 16540 15116 16681 15144
rect 16540 15104 16546 15116
rect 16669 15113 16681 15116
rect 16715 15113 16727 15147
rect 16669 15107 16727 15113
rect 14366 15008 14372 15020
rect 13320 14980 13676 15008
rect 14327 14980 14372 15008
rect 13320 14968 13326 14980
rect 14366 14968 14372 14980
rect 14424 14968 14430 15020
rect 4413 14943 4471 14949
rect 4413 14940 4425 14943
rect 4264 14912 4425 14940
rect 4413 14909 4425 14912
rect 4459 14909 4471 14943
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 4413 14903 4471 14909
rect 6748 14912 6837 14940
rect 3329 14875 3387 14881
rect 3329 14841 3341 14875
rect 3375 14872 3387 14875
rect 4246 14872 4252 14884
rect 3375 14844 4252 14872
rect 3375 14841 3387 14844
rect 3329 14835 3387 14841
rect 4246 14832 4252 14844
rect 4304 14872 4310 14884
rect 5442 14872 5448 14884
rect 4304 14844 5448 14872
rect 4304 14832 4310 14844
rect 5442 14832 5448 14844
rect 5500 14832 5506 14884
rect 6748 14816 6776 14912
rect 6825 14909 6837 14912
rect 6871 14909 6883 14943
rect 6825 14903 6883 14909
rect 7926 14900 7932 14952
rect 7984 14940 7990 14952
rect 8277 14943 8335 14949
rect 8277 14940 8289 14943
rect 7984 14912 8289 14940
rect 7984 14900 7990 14912
rect 8277 14909 8289 14912
rect 8323 14909 8335 14943
rect 11146 14940 11152 14952
rect 11107 14912 11152 14940
rect 8277 14903 8335 14909
rect 11146 14900 11152 14912
rect 11204 14940 11210 14952
rect 11514 14940 11520 14952
rect 11204 14912 11520 14940
rect 11204 14900 11210 14912
rect 11514 14900 11520 14912
rect 11572 14900 11578 14952
rect 14636 14943 14694 14949
rect 14636 14940 14648 14943
rect 14568 14912 14648 14940
rect 7561 14875 7619 14881
rect 7561 14841 7573 14875
rect 7607 14872 7619 14875
rect 8110 14872 8116 14884
rect 7607 14844 8116 14872
rect 7607 14841 7619 14844
rect 7561 14835 7619 14841
rect 8110 14832 8116 14844
rect 8168 14872 8174 14884
rect 8168 14844 8248 14872
rect 8168 14832 8174 14844
rect 1578 14804 1584 14816
rect 1539 14776 1584 14804
rect 1578 14764 1584 14776
rect 1636 14764 1642 14816
rect 2038 14804 2044 14816
rect 1999 14776 2044 14804
rect 2038 14764 2044 14776
rect 2096 14804 2102 14816
rect 2685 14807 2743 14813
rect 2685 14804 2697 14807
rect 2096 14776 2697 14804
rect 2096 14764 2102 14776
rect 2685 14773 2697 14776
rect 2731 14773 2743 14807
rect 5534 14804 5540 14816
rect 5495 14776 5540 14804
rect 2685 14767 2743 14773
rect 5534 14764 5540 14776
rect 5592 14764 5598 14816
rect 6641 14807 6699 14813
rect 6641 14773 6653 14807
rect 6687 14804 6699 14807
rect 6730 14804 6736 14816
rect 6687 14776 6736 14804
rect 6687 14773 6699 14776
rect 6641 14767 6699 14773
rect 6730 14764 6736 14776
rect 6788 14764 6794 14816
rect 7926 14804 7932 14816
rect 7887 14776 7932 14804
rect 7926 14764 7932 14776
rect 7984 14764 7990 14816
rect 8220 14804 8248 14844
rect 10042 14832 10048 14884
rect 10100 14872 10106 14884
rect 10597 14875 10655 14881
rect 10597 14872 10609 14875
rect 10100 14844 10609 14872
rect 10100 14832 10106 14844
rect 10597 14841 10609 14844
rect 10643 14872 10655 14875
rect 11241 14875 11299 14881
rect 11241 14872 11253 14875
rect 10643 14844 11253 14872
rect 10643 14841 10655 14844
rect 10597 14835 10655 14841
rect 11241 14841 11253 14844
rect 11287 14841 11299 14875
rect 11241 14835 11299 14841
rect 12710 14832 12716 14884
rect 12768 14872 12774 14884
rect 12897 14875 12955 14881
rect 12897 14872 12909 14875
rect 12768 14844 12909 14872
rect 12768 14832 12774 14844
rect 12897 14841 12909 14844
rect 12943 14841 12955 14875
rect 12897 14835 12955 14841
rect 14090 14832 14096 14884
rect 14148 14872 14154 14884
rect 14277 14875 14335 14881
rect 14277 14872 14289 14875
rect 14148 14844 14289 14872
rect 14148 14832 14154 14844
rect 14277 14841 14289 14844
rect 14323 14872 14335 14875
rect 14568 14872 14596 14912
rect 14636 14909 14648 14912
rect 14682 14940 14694 14943
rect 15378 14940 15384 14952
rect 14682 14912 15384 14940
rect 14682 14909 14694 14912
rect 14636 14903 14694 14909
rect 15378 14900 15384 14912
rect 15436 14900 15442 14952
rect 14323 14844 14596 14872
rect 14323 14841 14335 14844
rect 14277 14835 14335 14841
rect 9401 14807 9459 14813
rect 9401 14804 9413 14807
rect 8220 14776 9413 14804
rect 9401 14773 9413 14776
rect 9447 14804 9459 14807
rect 10134 14804 10140 14816
rect 9447 14776 10140 14804
rect 9447 14773 9459 14776
rect 9401 14767 9459 14773
rect 10134 14764 10140 14776
rect 10192 14764 10198 14816
rect 10781 14807 10839 14813
rect 10781 14773 10793 14807
rect 10827 14804 10839 14807
rect 11054 14804 11060 14816
rect 10827 14776 11060 14804
rect 10827 14773 10839 14776
rect 10781 14767 10839 14773
rect 11054 14764 11060 14776
rect 11112 14764 11118 14816
rect 12158 14764 12164 14816
rect 12216 14804 12222 14816
rect 12253 14807 12311 14813
rect 12253 14804 12265 14807
rect 12216 14776 12265 14804
rect 12216 14764 12222 14776
rect 12253 14773 12265 14776
rect 12299 14804 12311 14807
rect 12728 14804 12756 14832
rect 12299 14776 12756 14804
rect 12299 14773 12311 14776
rect 12253 14767 12311 14773
rect 15286 14764 15292 14816
rect 15344 14804 15350 14816
rect 15654 14804 15660 14816
rect 15344 14776 15660 14804
rect 15344 14764 15350 14776
rect 15654 14764 15660 14776
rect 15712 14804 15718 14816
rect 16301 14807 16359 14813
rect 16301 14804 16313 14807
rect 15712 14776 16313 14804
rect 15712 14764 15718 14776
rect 16301 14773 16313 14776
rect 16347 14773 16359 14807
rect 16301 14767 16359 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1397 14603 1455 14609
rect 1397 14569 1409 14603
rect 1443 14600 1455 14603
rect 1578 14600 1584 14612
rect 1443 14572 1584 14600
rect 1443 14569 1455 14572
rect 1397 14563 1455 14569
rect 1578 14560 1584 14572
rect 1636 14560 1642 14612
rect 2406 14600 2412 14612
rect 2367 14572 2412 14600
rect 2406 14560 2412 14572
rect 2464 14560 2470 14612
rect 2866 14600 2872 14612
rect 2779 14572 2872 14600
rect 2866 14560 2872 14572
rect 2924 14600 2930 14612
rect 3234 14600 3240 14612
rect 2924 14572 3240 14600
rect 2924 14560 2930 14572
rect 3234 14560 3240 14572
rect 3292 14560 3298 14612
rect 7561 14603 7619 14609
rect 7561 14569 7573 14603
rect 7607 14600 7619 14603
rect 7650 14600 7656 14612
rect 7607 14572 7656 14600
rect 7607 14569 7619 14572
rect 7561 14563 7619 14569
rect 7650 14560 7656 14572
rect 7708 14560 7714 14612
rect 7742 14560 7748 14612
rect 7800 14600 7806 14612
rect 7929 14603 7987 14609
rect 7929 14600 7941 14603
rect 7800 14572 7941 14600
rect 7800 14560 7806 14572
rect 7929 14569 7941 14572
rect 7975 14569 7987 14603
rect 9030 14600 9036 14612
rect 8991 14572 9036 14600
rect 7929 14563 7987 14569
rect 9030 14560 9036 14572
rect 9088 14560 9094 14612
rect 11790 14600 11796 14612
rect 11751 14572 11796 14600
rect 11790 14560 11796 14572
rect 11848 14560 11854 14612
rect 12161 14603 12219 14609
rect 12161 14569 12173 14603
rect 12207 14600 12219 14603
rect 13262 14600 13268 14612
rect 12207 14572 13268 14600
rect 12207 14569 12219 14572
rect 12161 14563 12219 14569
rect 13262 14560 13268 14572
rect 13320 14560 13326 14612
rect 14090 14600 14096 14612
rect 14051 14572 14096 14600
rect 14090 14560 14096 14572
rect 14148 14560 14154 14612
rect 14366 14560 14372 14612
rect 14424 14600 14430 14612
rect 14645 14603 14703 14609
rect 14645 14600 14657 14603
rect 14424 14572 14657 14600
rect 14424 14560 14430 14572
rect 14645 14569 14657 14572
rect 14691 14600 14703 14603
rect 15013 14603 15071 14609
rect 15013 14600 15025 14603
rect 14691 14572 15025 14600
rect 14691 14569 14703 14572
rect 14645 14563 14703 14569
rect 15013 14569 15025 14572
rect 15059 14569 15071 14603
rect 15013 14563 15071 14569
rect 15565 14603 15623 14609
rect 15565 14569 15577 14603
rect 15611 14600 15623 14603
rect 15746 14600 15752 14612
rect 15611 14572 15752 14600
rect 15611 14569 15623 14572
rect 15565 14563 15623 14569
rect 15746 14560 15752 14572
rect 15804 14560 15810 14612
rect 2222 14492 2228 14544
rect 2280 14532 2286 14544
rect 3789 14535 3847 14541
rect 3789 14532 3801 14535
rect 2280 14504 3801 14532
rect 2280 14492 2286 14504
rect 3789 14501 3801 14504
rect 3835 14501 3847 14535
rect 3789 14495 3847 14501
rect 4525 14535 4583 14541
rect 4525 14501 4537 14535
rect 4571 14532 4583 14535
rect 4706 14532 4712 14544
rect 4571 14504 4712 14532
rect 4571 14501 4583 14504
rect 4525 14495 4583 14501
rect 4706 14492 4712 14504
rect 4764 14532 4770 14544
rect 4893 14535 4951 14541
rect 4893 14532 4905 14535
rect 4764 14504 4905 14532
rect 4764 14492 4770 14504
rect 4893 14501 4905 14504
rect 4939 14532 4951 14535
rect 5252 14535 5310 14541
rect 5252 14532 5264 14535
rect 4939 14504 5264 14532
rect 4939 14501 4951 14504
rect 4893 14495 4951 14501
rect 5252 14501 5264 14504
rect 5298 14532 5310 14535
rect 5534 14532 5540 14544
rect 5298 14504 5540 14532
rect 5298 14501 5310 14504
rect 5252 14495 5310 14501
rect 5534 14492 5540 14504
rect 5592 14492 5598 14544
rect 7098 14492 7104 14544
rect 7156 14532 7162 14544
rect 8021 14535 8079 14541
rect 8021 14532 8033 14535
rect 7156 14504 8033 14532
rect 7156 14492 7162 14504
rect 8021 14501 8033 14504
rect 8067 14501 8079 14535
rect 8021 14495 8079 14501
rect 11057 14535 11115 14541
rect 11057 14501 11069 14535
rect 11103 14532 11115 14535
rect 11146 14532 11152 14544
rect 11103 14504 11152 14532
rect 11103 14501 11115 14504
rect 11057 14495 11115 14501
rect 11146 14492 11152 14504
rect 11204 14492 11210 14544
rect 12342 14492 12348 14544
rect 12400 14532 12406 14544
rect 12958 14535 13016 14541
rect 12958 14532 12970 14535
rect 12400 14504 12970 14532
rect 12400 14492 12406 14504
rect 12958 14501 12970 14504
rect 13004 14501 13016 14535
rect 16114 14532 16120 14544
rect 16075 14504 16120 14532
rect 12958 14495 13016 14501
rect 16114 14492 16120 14504
rect 16172 14492 16178 14544
rect 2777 14467 2835 14473
rect 2777 14433 2789 14467
rect 2823 14464 2835 14467
rect 3234 14464 3240 14476
rect 2823 14436 3240 14464
rect 2823 14433 2835 14436
rect 2777 14427 2835 14433
rect 3234 14424 3240 14436
rect 3292 14424 3298 14476
rect 4154 14424 4160 14476
rect 4212 14464 4218 14476
rect 4614 14464 4620 14476
rect 4212 14436 4620 14464
rect 4212 14424 4218 14436
rect 4614 14424 4620 14436
rect 4672 14464 4678 14476
rect 4985 14467 5043 14473
rect 4985 14464 4997 14467
rect 4672 14436 4997 14464
rect 4672 14424 4678 14436
rect 4985 14433 4997 14436
rect 5031 14433 5043 14467
rect 4985 14427 5043 14433
rect 9214 14424 9220 14476
rect 9272 14464 9278 14476
rect 9309 14467 9367 14473
rect 9309 14464 9321 14467
rect 9272 14436 9321 14464
rect 9272 14424 9278 14436
rect 9309 14433 9321 14436
rect 9355 14433 9367 14467
rect 9309 14427 9367 14433
rect 9950 14424 9956 14476
rect 10008 14464 10014 14476
rect 12437 14467 12495 14473
rect 12437 14464 12449 14467
rect 10008 14436 12449 14464
rect 10008 14424 10014 14436
rect 12437 14433 12449 14436
rect 12483 14464 12495 14467
rect 13354 14464 13360 14476
rect 12483 14436 13360 14464
rect 12483 14433 12495 14436
rect 12437 14427 12495 14433
rect 13354 14424 13360 14436
rect 13412 14424 13418 14476
rect 15838 14464 15844 14476
rect 15799 14436 15844 14464
rect 15838 14424 15844 14436
rect 15896 14424 15902 14476
rect 2406 14356 2412 14408
rect 2464 14396 2470 14408
rect 2866 14396 2872 14408
rect 2464 14368 2872 14396
rect 2464 14356 2470 14368
rect 2866 14356 2872 14368
rect 2924 14356 2930 14408
rect 2958 14356 2964 14408
rect 3016 14396 3022 14408
rect 7926 14396 7932 14408
rect 3016 14368 3061 14396
rect 7576 14368 7932 14396
rect 3016 14356 3022 14368
rect 1854 14328 1860 14340
rect 1815 14300 1860 14328
rect 1854 14288 1860 14300
rect 1912 14288 1918 14340
rect 2317 14331 2375 14337
rect 2317 14297 2329 14331
rect 2363 14328 2375 14331
rect 3050 14328 3056 14340
rect 2363 14300 3056 14328
rect 2363 14297 2375 14300
rect 2317 14291 2375 14297
rect 3050 14288 3056 14300
rect 3108 14288 3114 14340
rect 7374 14328 7380 14340
rect 6380 14300 7380 14328
rect 2590 14220 2596 14272
rect 2648 14260 2654 14272
rect 3421 14263 3479 14269
rect 3421 14260 3433 14263
rect 2648 14232 3433 14260
rect 2648 14220 2654 14232
rect 3421 14229 3433 14232
rect 3467 14229 3479 14263
rect 3421 14223 3479 14229
rect 6178 14220 6184 14272
rect 6236 14260 6242 14272
rect 6380 14269 6408 14300
rect 7374 14288 7380 14300
rect 7432 14288 7438 14340
rect 7576 14272 7604 14368
rect 7926 14356 7932 14368
rect 7984 14396 7990 14408
rect 8113 14399 8171 14405
rect 8113 14396 8125 14399
rect 7984 14368 8125 14396
rect 7984 14356 7990 14368
rect 8113 14365 8125 14368
rect 8159 14396 8171 14399
rect 8573 14399 8631 14405
rect 8573 14396 8585 14399
rect 8159 14368 8585 14396
rect 8159 14365 8171 14368
rect 8113 14359 8171 14365
rect 8573 14365 8585 14368
rect 8619 14396 8631 14399
rect 9030 14396 9036 14408
rect 8619 14368 9036 14396
rect 8619 14365 8631 14368
rect 8573 14359 8631 14365
rect 9030 14356 9036 14368
rect 9088 14356 9094 14408
rect 9674 14396 9680 14408
rect 9635 14368 9680 14396
rect 9674 14356 9680 14368
rect 9732 14356 9738 14408
rect 11149 14399 11207 14405
rect 11149 14365 11161 14399
rect 11195 14396 11207 14399
rect 11238 14396 11244 14408
rect 11195 14368 11244 14396
rect 11195 14365 11207 14368
rect 11149 14359 11207 14365
rect 11238 14356 11244 14368
rect 11296 14356 11302 14408
rect 11333 14399 11391 14405
rect 11333 14365 11345 14399
rect 11379 14365 11391 14399
rect 11333 14359 11391 14365
rect 12713 14399 12771 14405
rect 12713 14365 12725 14399
rect 12759 14365 12771 14399
rect 12713 14359 12771 14365
rect 10505 14331 10563 14337
rect 10505 14297 10517 14331
rect 10551 14328 10563 14331
rect 10962 14328 10968 14340
rect 10551 14300 10968 14328
rect 10551 14297 10563 14300
rect 10505 14291 10563 14297
rect 10962 14288 10968 14300
rect 11020 14288 11026 14340
rect 6365 14263 6423 14269
rect 6365 14260 6377 14263
rect 6236 14232 6377 14260
rect 6236 14220 6242 14232
rect 6365 14229 6377 14232
rect 6411 14229 6423 14263
rect 6365 14223 6423 14229
rect 7009 14263 7067 14269
rect 7009 14229 7021 14263
rect 7055 14260 7067 14263
rect 7190 14260 7196 14272
rect 7055 14232 7196 14260
rect 7055 14229 7067 14232
rect 7009 14223 7067 14229
rect 7190 14220 7196 14232
rect 7248 14220 7254 14272
rect 7469 14263 7527 14269
rect 7469 14229 7481 14263
rect 7515 14260 7527 14263
rect 7558 14260 7564 14272
rect 7515 14232 7564 14260
rect 7515 14229 7527 14232
rect 7469 14223 7527 14229
rect 7558 14220 7564 14232
rect 7616 14220 7622 14272
rect 9122 14260 9128 14272
rect 9035 14232 9128 14260
rect 9122 14220 9128 14232
rect 9180 14260 9186 14272
rect 10226 14260 10232 14272
rect 9180 14232 10232 14260
rect 9180 14220 9186 14232
rect 10226 14220 10232 14232
rect 10284 14220 10290 14272
rect 10686 14260 10692 14272
rect 10647 14232 10692 14260
rect 10686 14220 10692 14232
rect 10744 14220 10750 14272
rect 11238 14220 11244 14272
rect 11296 14260 11302 14272
rect 11348 14260 11376 14359
rect 12253 14331 12311 14337
rect 12253 14297 12265 14331
rect 12299 14328 12311 14331
rect 12434 14328 12440 14340
rect 12299 14300 12440 14328
rect 12299 14297 12311 14300
rect 12253 14291 12311 14297
rect 12434 14288 12440 14300
rect 12492 14328 12498 14340
rect 12728 14328 12756 14359
rect 12492 14300 12756 14328
rect 12492 14288 12498 14300
rect 11296 14232 11376 14260
rect 12728 14260 12756 14300
rect 14366 14260 14372 14272
rect 12728 14232 14372 14260
rect 11296 14220 11302 14232
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1489 14059 1547 14065
rect 1489 14025 1501 14059
rect 1535 14056 1547 14059
rect 3053 14059 3111 14065
rect 1535 14028 2728 14056
rect 1535 14025 1547 14028
rect 1489 14019 1547 14025
rect 1854 13948 1860 14000
rect 1912 13988 1918 14000
rect 1912 13960 1992 13988
rect 1912 13948 1918 13960
rect 1964 13929 1992 13960
rect 2406 13948 2412 14000
rect 2464 13988 2470 14000
rect 2501 13991 2559 13997
rect 2501 13988 2513 13991
rect 2464 13960 2513 13988
rect 2464 13948 2470 13960
rect 2501 13957 2513 13960
rect 2547 13957 2559 13991
rect 2501 13951 2559 13957
rect 1949 13923 2007 13929
rect 1949 13889 1961 13923
rect 1995 13889 2007 13923
rect 1949 13883 2007 13889
rect 2133 13923 2191 13929
rect 2133 13889 2145 13923
rect 2179 13920 2191 13923
rect 2590 13920 2596 13932
rect 2179 13892 2596 13920
rect 2179 13889 2191 13892
rect 2133 13883 2191 13889
rect 2590 13880 2596 13892
rect 2648 13880 2654 13932
rect 1578 13812 1584 13864
rect 1636 13852 1642 13864
rect 1857 13855 1915 13861
rect 1857 13852 1869 13855
rect 1636 13824 1869 13852
rect 1636 13812 1642 13824
rect 1857 13821 1869 13824
rect 1903 13821 1915 13855
rect 1857 13815 1915 13821
rect 2700 13784 2728 14028
rect 3053 14025 3065 14059
rect 3099 14056 3111 14059
rect 3142 14056 3148 14068
rect 3099 14028 3148 14056
rect 3099 14025 3111 14028
rect 3053 14019 3111 14025
rect 3142 14016 3148 14028
rect 3200 14016 3206 14068
rect 4157 14059 4215 14065
rect 4157 14025 4169 14059
rect 4203 14056 4215 14059
rect 4246 14056 4252 14068
rect 4203 14028 4252 14056
rect 4203 14025 4215 14028
rect 4157 14019 4215 14025
rect 4246 14016 4252 14028
rect 4304 14016 4310 14068
rect 4614 14056 4620 14068
rect 4575 14028 4620 14056
rect 4614 14016 4620 14028
rect 4672 14016 4678 14068
rect 6273 14059 6331 14065
rect 6273 14025 6285 14059
rect 6319 14056 6331 14059
rect 8846 14056 8852 14068
rect 6319 14028 8852 14056
rect 6319 14025 6331 14028
rect 6273 14019 6331 14025
rect 2958 13988 2964 14000
rect 2919 13960 2964 13988
rect 2958 13948 2964 13960
rect 3016 13948 3022 14000
rect 4522 13988 4528 14000
rect 4483 13960 4528 13988
rect 4522 13948 4528 13960
rect 4580 13948 4586 14000
rect 3602 13880 3608 13932
rect 3660 13920 3666 13932
rect 3697 13923 3755 13929
rect 3697 13920 3709 13923
rect 3660 13892 3709 13920
rect 3660 13880 3666 13892
rect 3697 13889 3709 13892
rect 3743 13920 3755 13923
rect 4062 13920 4068 13932
rect 3743 13892 4068 13920
rect 3743 13889 3755 13892
rect 3697 13883 3755 13889
rect 4062 13880 4068 13892
rect 4120 13880 4126 13932
rect 4540 13920 4568 13948
rect 4540 13892 5396 13920
rect 2774 13812 2780 13864
rect 2832 13852 2838 13864
rect 3513 13855 3571 13861
rect 3513 13852 3525 13855
rect 2832 13824 3525 13852
rect 2832 13812 2838 13824
rect 3513 13821 3525 13824
rect 3559 13852 3571 13855
rect 3786 13852 3792 13864
rect 3559 13824 3792 13852
rect 3559 13821 3571 13824
rect 3513 13815 3571 13821
rect 3786 13812 3792 13824
rect 3844 13812 3850 13864
rect 4801 13855 4859 13861
rect 4801 13821 4813 13855
rect 4847 13852 4859 13855
rect 4890 13852 4896 13864
rect 4847 13824 4896 13852
rect 4847 13821 4859 13824
rect 4801 13815 4859 13821
rect 4890 13812 4896 13824
rect 4948 13812 4954 13864
rect 5368 13852 5396 13892
rect 5534 13880 5540 13932
rect 5592 13920 5598 13932
rect 5721 13923 5779 13929
rect 5721 13920 5733 13923
rect 5592 13892 5733 13920
rect 5592 13880 5598 13892
rect 5721 13889 5733 13892
rect 5767 13889 5779 13923
rect 6288 13920 6316 14019
rect 8846 14016 8852 14028
rect 8904 14016 8910 14068
rect 9950 14056 9956 14068
rect 9911 14028 9956 14056
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 10226 14056 10232 14068
rect 10139 14028 10232 14056
rect 10226 14016 10232 14028
rect 10284 14056 10290 14068
rect 10870 14056 10876 14068
rect 10284 14028 10876 14056
rect 10284 14016 10290 14028
rect 10870 14016 10876 14028
rect 10928 14016 10934 14068
rect 11330 14016 11336 14068
rect 11388 14056 11394 14068
rect 11425 14059 11483 14065
rect 11425 14056 11437 14059
rect 11388 14028 11437 14056
rect 11388 14016 11394 14028
rect 11425 14025 11437 14028
rect 11471 14025 11483 14059
rect 12342 14056 12348 14068
rect 11425 14019 11483 14025
rect 12176 14028 12348 14056
rect 6825 13991 6883 13997
rect 6825 13957 6837 13991
rect 6871 13988 6883 13991
rect 6914 13988 6920 14000
rect 6871 13960 6920 13988
rect 6871 13957 6883 13960
rect 6825 13951 6883 13957
rect 6914 13948 6920 13960
rect 6972 13948 6978 14000
rect 7098 13948 7104 14000
rect 7156 13988 7162 14000
rect 7834 13988 7840 14000
rect 7156 13960 7840 13988
rect 7156 13948 7162 13960
rect 7834 13948 7840 13960
rect 7892 13948 7898 14000
rect 9858 13948 9864 14000
rect 9916 13988 9922 14000
rect 10413 13991 10471 13997
rect 10413 13988 10425 13991
rect 9916 13960 10425 13988
rect 9916 13948 9922 13960
rect 10413 13957 10425 13960
rect 10459 13957 10471 13991
rect 10413 13951 10471 13957
rect 5721 13883 5779 13889
rect 6104 13892 6316 13920
rect 5629 13855 5687 13861
rect 5629 13852 5641 13855
rect 5368 13824 5641 13852
rect 5629 13821 5641 13824
rect 5675 13821 5687 13855
rect 5629 13815 5687 13821
rect 2700 13756 3464 13784
rect 3436 13728 3464 13756
rect 5350 13744 5356 13796
rect 5408 13784 5414 13796
rect 5537 13787 5595 13793
rect 5537 13784 5549 13787
rect 5408 13756 5549 13784
rect 5408 13744 5414 13756
rect 5537 13753 5549 13756
rect 5583 13784 5595 13787
rect 6104 13784 6132 13892
rect 7374 13880 7380 13932
rect 7432 13929 7438 13932
rect 7432 13923 7481 13929
rect 7432 13889 7435 13923
rect 7469 13889 7481 13923
rect 8846 13920 8852 13932
rect 8807 13892 8852 13920
rect 7432 13883 7481 13889
rect 7432 13880 7438 13883
rect 8846 13880 8852 13892
rect 8904 13880 8910 13932
rect 9030 13920 9036 13932
rect 8991 13892 9036 13920
rect 9030 13880 9036 13892
rect 9088 13880 9094 13932
rect 9493 13923 9551 13929
rect 9493 13889 9505 13923
rect 9539 13920 9551 13923
rect 10962 13920 10968 13932
rect 9539 13892 10732 13920
rect 10923 13892 10968 13920
rect 9539 13889 9551 13892
rect 9493 13883 9551 13889
rect 10704 13864 10732 13892
rect 10962 13880 10968 13892
rect 11020 13920 11026 13932
rect 12176 13929 12204 14028
rect 12342 14016 12348 14028
rect 12400 14056 12406 14068
rect 13817 14059 13875 14065
rect 13817 14056 13829 14059
rect 12400 14028 13829 14056
rect 12400 14016 12406 14028
rect 13817 14025 13829 14028
rect 13863 14025 13875 14059
rect 14366 14056 14372 14068
rect 14327 14028 14372 14056
rect 13817 14019 13875 14025
rect 14366 14016 14372 14028
rect 14424 14016 14430 14068
rect 14458 14016 14464 14068
rect 14516 14056 14522 14068
rect 16301 14059 16359 14065
rect 16301 14056 16313 14059
rect 14516 14028 16313 14056
rect 14516 14016 14522 14028
rect 16301 14025 16313 14028
rect 16347 14025 16359 14059
rect 16301 14019 16359 14025
rect 12161 13923 12219 13929
rect 12161 13920 12173 13923
rect 11020 13892 12173 13920
rect 11020 13880 11026 13892
rect 12161 13889 12173 13892
rect 12207 13889 12219 13923
rect 12161 13883 12219 13889
rect 12434 13880 12440 13932
rect 12492 13920 12498 13932
rect 14829 13923 14887 13929
rect 12492 13892 12537 13920
rect 12492 13880 12498 13892
rect 14829 13889 14841 13923
rect 14875 13920 14887 13923
rect 14875 13892 15056 13920
rect 14875 13889 14887 13892
rect 14829 13883 14887 13889
rect 7190 13852 7196 13864
rect 7151 13824 7196 13852
rect 7190 13812 7196 13824
rect 7248 13812 7254 13864
rect 10137 13855 10195 13861
rect 10137 13821 10149 13855
rect 10183 13852 10195 13855
rect 10229 13855 10287 13861
rect 10229 13852 10241 13855
rect 10183 13824 10241 13852
rect 10183 13821 10195 13824
rect 10137 13815 10195 13821
rect 10229 13821 10241 13824
rect 10275 13821 10287 13855
rect 10229 13815 10287 13821
rect 10686 13812 10692 13864
rect 10744 13852 10750 13864
rect 12710 13861 12716 13864
rect 10781 13855 10839 13861
rect 10781 13852 10793 13855
rect 10744 13824 10793 13852
rect 10744 13812 10750 13824
rect 10781 13821 10793 13824
rect 10827 13821 10839 13855
rect 12693 13855 12716 13861
rect 12693 13852 12705 13855
rect 10781 13815 10839 13821
rect 11808 13824 12705 13852
rect 5583 13756 6132 13784
rect 5583 13753 5595 13756
rect 5537 13747 5595 13753
rect 6822 13744 6828 13796
rect 6880 13784 6886 13796
rect 8757 13787 8815 13793
rect 8757 13784 8769 13787
rect 6880 13756 7236 13784
rect 6880 13744 6886 13756
rect 3418 13716 3424 13728
rect 3379 13688 3424 13716
rect 3418 13676 3424 13688
rect 3476 13676 3482 13728
rect 5169 13719 5227 13725
rect 5169 13685 5181 13719
rect 5215 13716 5227 13719
rect 5994 13716 6000 13728
rect 5215 13688 6000 13716
rect 5215 13685 5227 13688
rect 5169 13679 5227 13685
rect 5994 13676 6000 13688
rect 6052 13676 6058 13728
rect 6178 13676 6184 13728
rect 6236 13716 6242 13728
rect 6549 13719 6607 13725
rect 6549 13716 6561 13719
rect 6236 13688 6561 13716
rect 6236 13676 6242 13688
rect 6549 13685 6561 13688
rect 6595 13685 6607 13719
rect 7208 13716 7236 13756
rect 8220 13756 8769 13784
rect 7285 13719 7343 13725
rect 7285 13716 7297 13719
rect 7208 13688 7297 13716
rect 6549 13679 6607 13685
rect 7285 13685 7297 13688
rect 7331 13685 7343 13719
rect 7285 13679 7343 13685
rect 7650 13676 7656 13728
rect 7708 13716 7714 13728
rect 8220 13725 8248 13756
rect 8757 13753 8769 13756
rect 8803 13753 8815 13787
rect 8757 13747 8815 13753
rect 9861 13787 9919 13793
rect 9861 13753 9873 13787
rect 9907 13784 9919 13787
rect 10873 13787 10931 13793
rect 10873 13784 10885 13787
rect 9907 13756 10885 13784
rect 9907 13753 9919 13756
rect 9861 13747 9919 13753
rect 10704 13728 10732 13756
rect 10873 13753 10885 13756
rect 10919 13753 10931 13787
rect 10873 13747 10931 13753
rect 11330 13744 11336 13796
rect 11388 13784 11394 13796
rect 11808 13793 11836 13824
rect 12693 13821 12705 13824
rect 12768 13852 12774 13864
rect 12768 13824 12841 13852
rect 12693 13815 12716 13821
rect 12710 13812 12716 13815
rect 12768 13812 12774 13824
rect 14366 13812 14372 13864
rect 14424 13852 14430 13864
rect 14921 13855 14979 13861
rect 14921 13852 14933 13855
rect 14424 13824 14933 13852
rect 14424 13812 14430 13824
rect 14921 13821 14933 13824
rect 14967 13821 14979 13855
rect 15028 13852 15056 13892
rect 15194 13861 15200 13864
rect 15188 13852 15200 13861
rect 15028 13824 15200 13852
rect 14921 13815 14979 13821
rect 15188 13815 15200 13824
rect 15194 13812 15200 13815
rect 15252 13812 15258 13864
rect 11793 13787 11851 13793
rect 11793 13784 11805 13787
rect 11388 13756 11805 13784
rect 11388 13744 11394 13756
rect 11793 13753 11805 13756
rect 11839 13753 11851 13787
rect 11793 13747 11851 13753
rect 8205 13719 8263 13725
rect 8205 13716 8217 13719
rect 7708 13688 8217 13716
rect 7708 13676 7714 13688
rect 8205 13685 8217 13688
rect 8251 13685 8263 13719
rect 8386 13716 8392 13728
rect 8347 13688 8392 13716
rect 8205 13679 8263 13685
rect 8386 13676 8392 13688
rect 8444 13676 8450 13728
rect 10686 13676 10692 13728
rect 10744 13676 10750 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1670 13472 1676 13524
rect 1728 13512 1734 13524
rect 1857 13515 1915 13521
rect 1857 13512 1869 13515
rect 1728 13484 1869 13512
rect 1728 13472 1734 13484
rect 1857 13481 1869 13484
rect 1903 13512 1915 13515
rect 2409 13515 2467 13521
rect 2409 13512 2421 13515
rect 1903 13484 2421 13512
rect 1903 13481 1915 13484
rect 1857 13475 1915 13481
rect 2409 13481 2421 13484
rect 2455 13481 2467 13515
rect 2409 13475 2467 13481
rect 3513 13515 3571 13521
rect 3513 13481 3525 13515
rect 3559 13512 3571 13515
rect 3602 13512 3608 13524
rect 3559 13484 3608 13512
rect 3559 13481 3571 13484
rect 3513 13475 3571 13481
rect 3602 13472 3608 13484
rect 3660 13472 3666 13524
rect 3786 13512 3792 13524
rect 3747 13484 3792 13512
rect 3786 13472 3792 13484
rect 3844 13472 3850 13524
rect 4706 13512 4712 13524
rect 4667 13484 4712 13512
rect 4706 13472 4712 13484
rect 4764 13472 4770 13524
rect 4801 13515 4859 13521
rect 4801 13481 4813 13515
rect 4847 13481 4859 13515
rect 5258 13512 5264 13524
rect 5219 13484 5264 13512
rect 4801 13475 4859 13481
rect 1762 13376 1768 13388
rect 1723 13348 1768 13376
rect 1762 13336 1768 13348
rect 1820 13336 1826 13388
rect 4816 13376 4844 13475
rect 5258 13472 5264 13484
rect 5316 13472 5322 13524
rect 5994 13472 6000 13524
rect 6052 13512 6058 13524
rect 6822 13512 6828 13524
rect 6052 13484 6828 13512
rect 6052 13472 6058 13484
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 7006 13472 7012 13524
rect 7064 13512 7070 13524
rect 7466 13512 7472 13524
rect 7064 13484 7109 13512
rect 7427 13484 7472 13512
rect 7064 13472 7070 13484
rect 7466 13472 7472 13484
rect 7524 13472 7530 13524
rect 7742 13472 7748 13524
rect 7800 13512 7806 13524
rect 8021 13515 8079 13521
rect 8021 13512 8033 13515
rect 7800 13484 8033 13512
rect 7800 13472 7806 13484
rect 8021 13481 8033 13484
rect 8067 13481 8079 13515
rect 8021 13475 8079 13481
rect 8481 13515 8539 13521
rect 8481 13481 8493 13515
rect 8527 13512 8539 13515
rect 8846 13512 8852 13524
rect 8527 13484 8852 13512
rect 8527 13481 8539 13484
rect 8481 13475 8539 13481
rect 8846 13472 8852 13484
rect 8904 13472 8910 13524
rect 8938 13472 8944 13524
rect 8996 13512 9002 13524
rect 9033 13515 9091 13521
rect 9033 13512 9045 13515
rect 8996 13484 9045 13512
rect 8996 13472 9002 13484
rect 9033 13481 9045 13484
rect 9079 13481 9091 13515
rect 9398 13512 9404 13524
rect 9359 13484 9404 13512
rect 9033 13475 9091 13481
rect 9398 13472 9404 13484
rect 9456 13472 9462 13524
rect 9674 13472 9680 13524
rect 9732 13512 9738 13524
rect 10045 13515 10103 13521
rect 10045 13512 10057 13515
rect 9732 13484 10057 13512
rect 9732 13472 9738 13484
rect 10045 13481 10057 13484
rect 10091 13481 10103 13515
rect 10045 13475 10103 13481
rect 12710 13472 12716 13524
rect 12768 13512 12774 13524
rect 12805 13515 12863 13521
rect 12805 13512 12817 13515
rect 12768 13484 12817 13512
rect 12768 13472 12774 13484
rect 12805 13481 12817 13484
rect 12851 13481 12863 13515
rect 13354 13512 13360 13524
rect 13315 13484 13360 13512
rect 12805 13475 12863 13481
rect 13354 13472 13360 13484
rect 13412 13472 13418 13524
rect 13446 13472 13452 13524
rect 13504 13512 13510 13524
rect 13909 13515 13967 13521
rect 13909 13512 13921 13515
rect 13504 13484 13921 13512
rect 13504 13472 13510 13484
rect 13909 13481 13921 13484
rect 13955 13481 13967 13515
rect 13909 13475 13967 13481
rect 15194 13472 15200 13524
rect 15252 13512 15258 13524
rect 15838 13512 15844 13524
rect 15252 13484 15844 13512
rect 15252 13472 15258 13484
rect 15838 13472 15844 13484
rect 15896 13472 15902 13524
rect 5169 13447 5227 13453
rect 5169 13413 5181 13447
rect 5215 13444 5227 13447
rect 5534 13444 5540 13456
rect 5215 13416 5540 13444
rect 5215 13413 5227 13416
rect 5169 13407 5227 13413
rect 5534 13404 5540 13416
rect 5592 13444 5598 13456
rect 5592 13416 6684 13444
rect 5592 13404 5598 13416
rect 6273 13379 6331 13385
rect 4816 13348 6224 13376
rect 2038 13308 2044 13320
rect 1951 13280 2044 13308
rect 2038 13268 2044 13280
rect 2096 13308 2102 13320
rect 2961 13311 3019 13317
rect 2096 13280 2912 13308
rect 2096 13268 2102 13280
rect 2884 13184 2912 13280
rect 2961 13277 2973 13311
rect 3007 13308 3019 13311
rect 4154 13308 4160 13320
rect 3007 13280 4160 13308
rect 3007 13277 3019 13280
rect 2961 13271 3019 13277
rect 4154 13268 4160 13280
rect 4212 13268 4218 13320
rect 5442 13308 5448 13320
rect 5403 13280 5448 13308
rect 5442 13268 5448 13280
rect 5500 13268 5506 13320
rect 6196 13308 6224 13348
rect 6273 13345 6285 13379
rect 6319 13376 6331 13379
rect 6546 13376 6552 13388
rect 6319 13348 6552 13376
rect 6319 13345 6331 13348
rect 6273 13339 6331 13345
rect 6546 13336 6552 13348
rect 6604 13336 6610 13388
rect 6656 13376 6684 13416
rect 7282 13404 7288 13456
rect 7340 13444 7346 13456
rect 7377 13447 7435 13453
rect 7377 13444 7389 13447
rect 7340 13416 7389 13444
rect 7340 13404 7346 13416
rect 7377 13413 7389 13416
rect 7423 13413 7435 13447
rect 7377 13407 7435 13413
rect 13817 13447 13875 13453
rect 13817 13413 13829 13447
rect 13863 13444 13875 13447
rect 14366 13444 14372 13456
rect 13863 13416 14372 13444
rect 13863 13413 13875 13416
rect 13817 13407 13875 13413
rect 14366 13404 14372 13416
rect 14424 13444 14430 13456
rect 14921 13447 14979 13453
rect 14921 13444 14933 13447
rect 14424 13416 14933 13444
rect 14424 13404 14430 13416
rect 14921 13413 14933 13416
rect 14967 13413 14979 13447
rect 14921 13407 14979 13413
rect 16850 13404 16856 13456
rect 16908 13444 16914 13456
rect 16945 13447 17003 13453
rect 16945 13444 16957 13447
rect 16908 13416 16957 13444
rect 16908 13404 16914 13416
rect 16945 13413 16957 13416
rect 16991 13413 17003 13447
rect 16945 13407 17003 13413
rect 11698 13385 11704 13388
rect 8573 13379 8631 13385
rect 8573 13376 8585 13379
rect 6656 13348 8585 13376
rect 8573 13345 8585 13348
rect 8619 13345 8631 13379
rect 11692 13376 11704 13385
rect 11659 13348 11704 13376
rect 8573 13339 8631 13345
rect 11692 13339 11704 13348
rect 11698 13336 11704 13339
rect 11756 13336 11762 13388
rect 16666 13376 16672 13388
rect 16627 13348 16672 13376
rect 16666 13336 16672 13348
rect 16724 13336 16730 13388
rect 7190 13308 7196 13320
rect 6196 13280 7196 13308
rect 7190 13268 7196 13280
rect 7248 13268 7254 13320
rect 7558 13308 7564 13320
rect 7519 13280 7564 13308
rect 7558 13268 7564 13280
rect 7616 13268 7622 13320
rect 9306 13268 9312 13320
rect 9364 13308 9370 13320
rect 10137 13311 10195 13317
rect 10137 13308 10149 13311
rect 9364 13280 10149 13308
rect 9364 13268 9370 13280
rect 10137 13277 10149 13280
rect 10183 13277 10195 13311
rect 10137 13271 10195 13277
rect 10226 13268 10232 13320
rect 10284 13308 10290 13320
rect 10284 13280 10329 13308
rect 10284 13268 10290 13280
rect 11238 13268 11244 13320
rect 11296 13308 11302 13320
rect 11425 13311 11483 13317
rect 11425 13308 11437 13311
rect 11296 13280 11437 13308
rect 11296 13268 11302 13280
rect 11425 13277 11437 13280
rect 11471 13277 11483 13311
rect 11425 13271 11483 13277
rect 4341 13243 4399 13249
rect 4341 13209 4353 13243
rect 4387 13240 4399 13243
rect 4890 13240 4896 13252
rect 4387 13212 4896 13240
rect 4387 13209 4399 13212
rect 4341 13203 4399 13209
rect 4890 13200 4896 13212
rect 4948 13240 4954 13252
rect 9677 13243 9735 13249
rect 4948 13212 6408 13240
rect 4948 13200 4954 13212
rect 6380 13184 6408 13212
rect 9677 13209 9689 13243
rect 9723 13240 9735 13243
rect 9766 13240 9772 13252
rect 9723 13212 9772 13240
rect 9723 13209 9735 13212
rect 9677 13203 9735 13209
rect 9766 13200 9772 13212
rect 9824 13200 9830 13252
rect 1397 13175 1455 13181
rect 1397 13141 1409 13175
rect 1443 13172 1455 13175
rect 2682 13172 2688 13184
rect 1443 13144 2688 13172
rect 1443 13141 1455 13144
rect 1397 13135 1455 13141
rect 2682 13132 2688 13144
rect 2740 13132 2746 13184
rect 2866 13172 2872 13184
rect 2827 13144 2872 13172
rect 2866 13132 2872 13144
rect 2924 13132 2930 13184
rect 5905 13175 5963 13181
rect 5905 13141 5917 13175
rect 5951 13172 5963 13175
rect 5994 13172 6000 13184
rect 5951 13144 6000 13172
rect 5951 13141 5963 13144
rect 5905 13135 5963 13141
rect 5994 13132 6000 13144
rect 6052 13132 6058 13184
rect 6362 13172 6368 13184
rect 6323 13144 6368 13172
rect 6362 13132 6368 13144
rect 6420 13132 6426 13184
rect 10778 13172 10784 13184
rect 10739 13144 10784 13172
rect 10778 13132 10784 13144
rect 10836 13132 10842 13184
rect 11149 13175 11207 13181
rect 11149 13141 11161 13175
rect 11195 13172 11207 13175
rect 11330 13172 11336 13184
rect 11195 13144 11336 13172
rect 11195 13141 11207 13144
rect 11149 13135 11207 13141
rect 11330 13132 11336 13144
rect 11388 13132 11394 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 3418 12968 3424 12980
rect 3379 12940 3424 12968
rect 3418 12928 3424 12940
rect 3476 12928 3482 12980
rect 4893 12971 4951 12977
rect 4893 12937 4905 12971
rect 4939 12968 4951 12971
rect 5258 12968 5264 12980
rect 4939 12940 5264 12968
rect 4939 12937 4951 12940
rect 4893 12931 4951 12937
rect 5258 12928 5264 12940
rect 5316 12928 5322 12980
rect 6273 12971 6331 12977
rect 6273 12937 6285 12971
rect 6319 12968 6331 12971
rect 7558 12968 7564 12980
rect 6319 12940 7564 12968
rect 6319 12937 6331 12940
rect 6273 12931 6331 12937
rect 7558 12928 7564 12940
rect 7616 12928 7622 12980
rect 8386 12928 8392 12980
rect 8444 12968 8450 12980
rect 9306 12968 9312 12980
rect 8444 12940 9312 12968
rect 8444 12928 8450 12940
rect 9306 12928 9312 12940
rect 9364 12928 9370 12980
rect 9674 12968 9680 12980
rect 9635 12940 9680 12968
rect 9674 12928 9680 12940
rect 9732 12928 9738 12980
rect 10137 12971 10195 12977
rect 10137 12937 10149 12971
rect 10183 12968 10195 12971
rect 10226 12968 10232 12980
rect 10183 12940 10232 12968
rect 10183 12937 10195 12940
rect 10137 12931 10195 12937
rect 10226 12928 10232 12940
rect 10284 12928 10290 12980
rect 10686 12968 10692 12980
rect 10647 12940 10692 12968
rect 10686 12928 10692 12940
rect 10744 12928 10750 12980
rect 10870 12928 10876 12980
rect 10928 12968 10934 12980
rect 12069 12971 12127 12977
rect 12069 12968 12081 12971
rect 10928 12940 12081 12968
rect 10928 12928 10934 12940
rect 12069 12937 12081 12940
rect 12115 12937 12127 12971
rect 12069 12931 12127 12937
rect 16666 12928 16672 12980
rect 16724 12968 16730 12980
rect 17034 12968 17040 12980
rect 16724 12940 17040 12968
rect 16724 12928 16730 12940
rect 17034 12928 17040 12940
rect 17092 12928 17098 12980
rect 6641 12903 6699 12909
rect 6641 12869 6653 12903
rect 6687 12900 6699 12903
rect 7006 12900 7012 12912
rect 6687 12872 7012 12900
rect 6687 12869 6699 12872
rect 6641 12863 6699 12869
rect 7006 12860 7012 12872
rect 7064 12900 7070 12912
rect 7282 12900 7288 12912
rect 7064 12872 7288 12900
rect 7064 12860 7070 12872
rect 7282 12860 7288 12872
rect 7340 12860 7346 12912
rect 8662 12900 8668 12912
rect 8623 12872 8668 12900
rect 8662 12860 8668 12872
rect 8720 12860 8726 12912
rect 10597 12903 10655 12909
rect 10597 12869 10609 12903
rect 10643 12900 10655 12903
rect 11422 12900 11428 12912
rect 10643 12872 11428 12900
rect 10643 12869 10655 12872
rect 10597 12863 10655 12869
rect 5813 12835 5871 12841
rect 5813 12801 5825 12835
rect 5859 12832 5871 12835
rect 5994 12832 6000 12844
rect 5859 12804 6000 12832
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 5994 12792 6000 12804
rect 6052 12832 6058 12844
rect 6052 12804 6960 12832
rect 6052 12792 6058 12804
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 1486 12764 1492 12776
rect 1443 12736 1492 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 1486 12724 1492 12736
rect 1544 12724 1550 12776
rect 1664 12767 1722 12773
rect 1664 12733 1676 12767
rect 1710 12764 1722 12767
rect 2038 12764 2044 12776
rect 1710 12736 2044 12764
rect 1710 12733 1722 12736
rect 1664 12727 1722 12733
rect 2038 12724 2044 12736
rect 2096 12724 2102 12776
rect 4525 12767 4583 12773
rect 4525 12733 4537 12767
rect 4571 12764 4583 12767
rect 5537 12767 5595 12773
rect 5537 12764 5549 12767
rect 4571 12736 5549 12764
rect 4571 12733 4583 12736
rect 4525 12727 4583 12733
rect 5537 12733 5549 12736
rect 5583 12764 5595 12767
rect 6822 12764 6828 12776
rect 5583 12736 6828 12764
rect 5583 12733 5595 12736
rect 5537 12727 5595 12733
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 3881 12699 3939 12705
rect 3881 12665 3893 12699
rect 3927 12696 3939 12699
rect 5074 12696 5080 12708
rect 3927 12668 5080 12696
rect 3927 12665 3939 12668
rect 3881 12659 3939 12665
rect 5074 12656 5080 12668
rect 5132 12696 5138 12708
rect 5629 12699 5687 12705
rect 5629 12696 5641 12699
rect 5132 12668 5641 12696
rect 5132 12656 5138 12668
rect 5629 12665 5641 12668
rect 5675 12665 5687 12699
rect 6932 12696 6960 12804
rect 7282 12764 7288 12776
rect 7243 12736 7288 12764
rect 7282 12724 7288 12736
rect 7340 12724 7346 12776
rect 7552 12699 7610 12705
rect 7552 12696 7564 12699
rect 6932 12668 7564 12696
rect 5629 12659 5687 12665
rect 7552 12665 7564 12668
rect 7598 12696 7610 12699
rect 7742 12696 7748 12708
rect 7598 12668 7748 12696
rect 7598 12665 7610 12668
rect 7552 12659 7610 12665
rect 7742 12656 7748 12668
rect 7800 12656 7806 12708
rect 10778 12656 10784 12708
rect 10836 12696 10842 12708
rect 10888 12696 10916 12872
rect 11422 12860 11428 12872
rect 11480 12860 11486 12912
rect 11054 12792 11060 12844
rect 11112 12832 11118 12844
rect 11149 12835 11207 12841
rect 11149 12832 11161 12835
rect 11112 12804 11161 12832
rect 11112 12792 11118 12804
rect 11149 12801 11161 12804
rect 11195 12801 11207 12835
rect 11330 12832 11336 12844
rect 11291 12804 11336 12832
rect 11149 12795 11207 12801
rect 11330 12792 11336 12804
rect 11388 12792 11394 12844
rect 12434 12792 12440 12844
rect 12492 12832 12498 12844
rect 16206 12832 16212 12844
rect 12492 12804 12537 12832
rect 16167 12804 16212 12832
rect 12492 12792 12498 12804
rect 16206 12792 16212 12804
rect 16264 12792 16270 12844
rect 18322 12832 18328 12844
rect 18283 12804 18328 12832
rect 18322 12792 18328 12804
rect 18380 12792 18386 12844
rect 15930 12764 15936 12776
rect 15891 12736 15936 12764
rect 15930 12724 15936 12736
rect 15988 12764 15994 12776
rect 16669 12767 16727 12773
rect 16669 12764 16681 12767
rect 15988 12736 16681 12764
rect 15988 12724 15994 12736
rect 16669 12733 16681 12736
rect 16715 12733 16727 12767
rect 18046 12764 18052 12776
rect 17959 12736 18052 12764
rect 16669 12727 16727 12733
rect 18046 12724 18052 12736
rect 18104 12764 18110 12776
rect 18785 12767 18843 12773
rect 18785 12764 18797 12767
rect 18104 12736 18797 12764
rect 18104 12724 18110 12736
rect 18785 12733 18797 12736
rect 18831 12733 18843 12767
rect 18785 12727 18843 12733
rect 11057 12699 11115 12705
rect 11057 12696 11069 12699
rect 10836 12668 11069 12696
rect 10836 12656 10842 12668
rect 11057 12665 11069 12668
rect 11103 12665 11115 12699
rect 11057 12659 11115 12665
rect 2777 12631 2835 12637
rect 2777 12597 2789 12631
rect 2823 12628 2835 12631
rect 2866 12628 2872 12640
rect 2823 12600 2872 12628
rect 2823 12597 2835 12600
rect 2777 12591 2835 12597
rect 2866 12588 2872 12600
rect 2924 12588 2930 12640
rect 3970 12628 3976 12640
rect 3931 12600 3976 12628
rect 3970 12588 3976 12600
rect 4028 12588 4034 12640
rect 5166 12628 5172 12640
rect 5127 12600 5172 12628
rect 5166 12588 5172 12600
rect 5224 12588 5230 12640
rect 7101 12631 7159 12637
rect 7101 12597 7113 12631
rect 7147 12628 7159 12631
rect 7466 12628 7472 12640
rect 7147 12600 7472 12628
rect 7147 12597 7159 12600
rect 7101 12591 7159 12597
rect 7466 12588 7472 12600
rect 7524 12588 7530 12640
rect 11790 12628 11796 12640
rect 11751 12600 11796 12628
rect 11790 12588 11796 12600
rect 11848 12588 11854 12640
rect 12986 12628 12992 12640
rect 12947 12600 12992 12628
rect 12986 12588 12992 12600
rect 13044 12588 13050 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1857 12427 1915 12433
rect 1857 12393 1869 12427
rect 1903 12424 1915 12427
rect 2130 12424 2136 12436
rect 1903 12396 2136 12424
rect 1903 12393 1915 12396
rect 1857 12387 1915 12393
rect 2130 12384 2136 12396
rect 2188 12384 2194 12436
rect 2406 12424 2412 12436
rect 2367 12396 2412 12424
rect 2406 12384 2412 12396
rect 2464 12384 2470 12436
rect 2869 12427 2927 12433
rect 2869 12393 2881 12427
rect 2915 12424 2927 12427
rect 2958 12424 2964 12436
rect 2915 12396 2964 12424
rect 2915 12393 2927 12396
rect 2869 12387 2927 12393
rect 2958 12384 2964 12396
rect 3016 12384 3022 12436
rect 3602 12384 3608 12436
rect 3660 12424 3666 12436
rect 4430 12424 4436 12436
rect 3660 12396 4436 12424
rect 3660 12384 3666 12396
rect 4430 12384 4436 12396
rect 4488 12384 4494 12436
rect 5626 12424 5632 12436
rect 5587 12396 5632 12424
rect 5626 12384 5632 12396
rect 5684 12384 5690 12436
rect 7282 12384 7288 12436
rect 7340 12424 7346 12436
rect 8021 12427 8079 12433
rect 8021 12424 8033 12427
rect 7340 12396 8033 12424
rect 7340 12384 7346 12396
rect 8021 12393 8033 12396
rect 8067 12393 8079 12427
rect 9214 12424 9220 12436
rect 9175 12396 9220 12424
rect 8021 12387 8079 12393
rect 9214 12384 9220 12396
rect 9272 12384 9278 12436
rect 11054 12424 11060 12436
rect 11015 12396 11060 12424
rect 11054 12384 11060 12396
rect 11112 12384 11118 12436
rect 11606 12424 11612 12436
rect 11567 12396 11612 12424
rect 11606 12384 11612 12396
rect 11664 12384 11670 12436
rect 2774 12316 2780 12368
rect 2832 12356 2838 12368
rect 3789 12359 3847 12365
rect 3789 12356 3801 12359
rect 2832 12328 3801 12356
rect 2832 12316 2838 12328
rect 3789 12325 3801 12328
rect 3835 12356 3847 12359
rect 4525 12359 4583 12365
rect 4525 12356 4537 12359
rect 3835 12328 4537 12356
rect 3835 12325 3847 12328
rect 3789 12319 3847 12325
rect 4525 12325 4537 12328
rect 4571 12325 4583 12359
rect 4525 12319 4583 12325
rect 5988 12359 6046 12365
rect 5988 12325 6000 12359
rect 6034 12356 6046 12359
rect 6178 12356 6184 12368
rect 6034 12328 6184 12356
rect 6034 12325 6046 12328
rect 5988 12319 6046 12325
rect 6178 12316 6184 12328
rect 6236 12316 6242 12368
rect 6914 12316 6920 12368
rect 6972 12356 6978 12368
rect 8205 12359 8263 12365
rect 8205 12356 8217 12359
rect 6972 12328 8217 12356
rect 6972 12316 6978 12328
rect 8205 12325 8217 12328
rect 8251 12325 8263 12359
rect 8205 12319 8263 12325
rect 9950 12316 9956 12368
rect 10008 12356 10014 12368
rect 10781 12359 10839 12365
rect 10008 12328 10732 12356
rect 10008 12316 10014 12328
rect 1578 12248 1584 12300
rect 1636 12288 1642 12300
rect 1765 12291 1823 12297
rect 1765 12288 1777 12291
rect 1636 12260 1777 12288
rect 1636 12248 1642 12260
rect 1765 12257 1777 12260
rect 1811 12257 1823 12291
rect 1765 12251 1823 12257
rect 4154 12248 4160 12300
rect 4212 12288 4218 12300
rect 4430 12288 4436 12300
rect 4212 12260 4436 12288
rect 4212 12248 4218 12260
rect 4430 12248 4436 12260
rect 4488 12248 4494 12300
rect 5718 12288 5724 12300
rect 5679 12260 5724 12288
rect 5718 12248 5724 12260
rect 5776 12288 5782 12300
rect 7558 12288 7564 12300
rect 5776 12260 7564 12288
rect 5776 12248 5782 12260
rect 7558 12248 7564 12260
rect 7616 12288 7622 12300
rect 8665 12291 8723 12297
rect 8665 12288 8677 12291
rect 7616 12260 8677 12288
rect 7616 12248 7622 12260
rect 8665 12257 8677 12260
rect 8711 12257 8723 12291
rect 8665 12251 8723 12257
rect 8846 12248 8852 12300
rect 8904 12288 8910 12300
rect 10045 12291 10103 12297
rect 10045 12288 10057 12291
rect 8904 12260 10057 12288
rect 8904 12248 8910 12260
rect 10045 12257 10057 12260
rect 10091 12257 10103 12291
rect 10704 12288 10732 12328
rect 10781 12325 10793 12359
rect 10827 12356 10839 12359
rect 11330 12356 11336 12368
rect 10827 12328 11336 12356
rect 10827 12325 10839 12328
rect 10781 12319 10839 12325
rect 11330 12316 11336 12328
rect 11388 12316 11394 12368
rect 20990 12316 20996 12368
rect 21048 12356 21054 12368
rect 21177 12359 21235 12365
rect 21177 12356 21189 12359
rect 21048 12328 21189 12356
rect 21048 12316 21054 12328
rect 21177 12325 21189 12328
rect 21223 12325 21235 12359
rect 21177 12319 21235 12325
rect 10870 12288 10876 12300
rect 10704 12260 10876 12288
rect 10045 12251 10103 12257
rect 10870 12248 10876 12260
rect 10928 12288 10934 12300
rect 11425 12291 11483 12297
rect 11425 12288 11437 12291
rect 10928 12260 11437 12288
rect 10928 12248 10934 12260
rect 11425 12257 11437 12260
rect 11471 12257 11483 12291
rect 11974 12288 11980 12300
rect 11935 12260 11980 12288
rect 11425 12251 11483 12257
rect 11974 12248 11980 12260
rect 12032 12248 12038 12300
rect 20898 12288 20904 12300
rect 20859 12260 20904 12288
rect 20898 12248 20904 12260
rect 20956 12248 20962 12300
rect 2041 12223 2099 12229
rect 2041 12189 2053 12223
rect 2087 12189 2099 12223
rect 4614 12220 4620 12232
rect 4575 12192 4620 12220
rect 2041 12183 2099 12189
rect 2056 12152 2084 12183
rect 4614 12180 4620 12192
rect 4672 12180 4678 12232
rect 9122 12180 9128 12232
rect 9180 12220 9186 12232
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 9180 12192 10149 12220
rect 9180 12180 9186 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 3237 12155 3295 12161
rect 3237 12152 3249 12155
rect 2056 12124 3249 12152
rect 3237 12121 3249 12124
rect 3283 12152 3295 12155
rect 3418 12152 3424 12164
rect 3283 12124 3424 12152
rect 3283 12121 3295 12124
rect 3237 12115 3295 12121
rect 3418 12112 3424 12124
rect 3476 12112 3482 12164
rect 4062 12152 4068 12164
rect 4023 12124 4068 12152
rect 4062 12112 4068 12124
rect 4120 12112 4126 12164
rect 9582 12112 9588 12164
rect 9640 12152 9646 12164
rect 10244 12152 10272 12183
rect 11330 12180 11336 12232
rect 11388 12220 11394 12232
rect 12069 12223 12127 12229
rect 12069 12220 12081 12223
rect 11388 12192 12081 12220
rect 11388 12180 11394 12192
rect 12069 12189 12081 12192
rect 12115 12189 12127 12223
rect 12250 12220 12256 12232
rect 12163 12192 12256 12220
rect 12069 12183 12127 12189
rect 12250 12180 12256 12192
rect 12308 12220 12314 12232
rect 12621 12223 12679 12229
rect 12621 12220 12633 12223
rect 12308 12192 12633 12220
rect 12308 12180 12314 12192
rect 12621 12189 12633 12192
rect 12667 12189 12679 12223
rect 12621 12183 12679 12189
rect 9640 12124 10272 12152
rect 9640 12112 9646 12124
rect 1397 12087 1455 12093
rect 1397 12053 1409 12087
rect 1443 12084 1455 12087
rect 1854 12084 1860 12096
rect 1443 12056 1860 12084
rect 1443 12053 1455 12056
rect 1397 12047 1455 12053
rect 1854 12044 1860 12056
rect 1912 12044 1918 12096
rect 5258 12084 5264 12096
rect 5219 12056 5264 12084
rect 5258 12044 5264 12056
rect 5316 12044 5322 12096
rect 7098 12084 7104 12096
rect 7059 12056 7104 12084
rect 7098 12044 7104 12056
rect 7156 12044 7162 12096
rect 7742 12084 7748 12096
rect 7703 12056 7748 12084
rect 7742 12044 7748 12056
rect 7800 12044 7806 12096
rect 9674 12084 9680 12096
rect 9635 12056 9680 12084
rect 9674 12044 9680 12056
rect 9732 12044 9738 12096
rect 11054 12044 11060 12096
rect 11112 12084 11118 12096
rect 11238 12084 11244 12096
rect 11112 12056 11244 12084
rect 11112 12044 11118 12056
rect 11238 12044 11244 12056
rect 11296 12084 11302 12096
rect 12986 12084 12992 12096
rect 11296 12056 12992 12084
rect 11296 12044 11302 12056
rect 12986 12044 12992 12056
rect 13044 12044 13050 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2041 11883 2099 11889
rect 2041 11849 2053 11883
rect 2087 11880 2099 11883
rect 2130 11880 2136 11892
rect 2087 11852 2136 11880
rect 2087 11849 2099 11852
rect 2041 11843 2099 11849
rect 2130 11840 2136 11852
rect 2188 11840 2194 11892
rect 4157 11883 4215 11889
rect 4157 11849 4169 11883
rect 4203 11880 4215 11883
rect 4430 11880 4436 11892
rect 4203 11852 4436 11880
rect 4203 11849 4215 11852
rect 4157 11843 4215 11849
rect 4430 11840 4436 11852
rect 4488 11840 4494 11892
rect 5074 11840 5080 11892
rect 5132 11880 5138 11892
rect 5169 11883 5227 11889
rect 5169 11880 5181 11883
rect 5132 11852 5181 11880
rect 5132 11840 5138 11852
rect 5169 11849 5181 11852
rect 5215 11849 5227 11883
rect 6178 11880 6184 11892
rect 6139 11852 6184 11880
rect 5169 11843 5227 11849
rect 6178 11840 6184 11852
rect 6236 11840 6242 11892
rect 7190 11880 7196 11892
rect 6840 11852 7196 11880
rect 3878 11772 3884 11824
rect 3936 11812 3942 11824
rect 4709 11815 4767 11821
rect 4709 11812 4721 11815
rect 3936 11784 4721 11812
rect 3936 11772 3942 11784
rect 4709 11781 4721 11784
rect 4755 11781 4767 11815
rect 4890 11812 4896 11824
rect 4803 11784 4896 11812
rect 4709 11775 4767 11781
rect 4724 11744 4752 11775
rect 4890 11772 4896 11784
rect 4948 11812 4954 11824
rect 6840 11812 6868 11852
rect 7190 11840 7196 11852
rect 7248 11840 7254 11892
rect 7742 11840 7748 11892
rect 7800 11880 7806 11892
rect 8205 11883 8263 11889
rect 8205 11880 8217 11883
rect 7800 11852 8217 11880
rect 7800 11840 7806 11852
rect 8205 11849 8217 11852
rect 8251 11849 8263 11883
rect 8846 11880 8852 11892
rect 8807 11852 8852 11880
rect 8205 11843 8263 11849
rect 8846 11840 8852 11852
rect 8904 11840 8910 11892
rect 11330 11880 11336 11892
rect 11291 11852 11336 11880
rect 11330 11840 11336 11852
rect 11388 11840 11394 11892
rect 12069 11883 12127 11889
rect 12069 11849 12081 11883
rect 12115 11880 12127 11883
rect 12250 11880 12256 11892
rect 12115 11852 12256 11880
rect 12115 11849 12127 11852
rect 12069 11843 12127 11849
rect 12250 11840 12256 11852
rect 12308 11840 12314 11892
rect 12802 11880 12808 11892
rect 12452 11852 12808 11880
rect 4948 11784 6868 11812
rect 4948 11772 4954 11784
rect 6840 11753 6868 11784
rect 7834 11772 7840 11824
rect 7892 11812 7898 11824
rect 9122 11812 9128 11824
rect 7892 11784 9128 11812
rect 7892 11772 7898 11784
rect 9122 11772 9128 11784
rect 9180 11772 9186 11824
rect 12452 11753 12480 11852
rect 12802 11840 12808 11852
rect 12860 11840 12866 11892
rect 13814 11880 13820 11892
rect 13775 11852 13820 11880
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 5813 11747 5871 11753
rect 4724 11716 5580 11744
rect 2133 11679 2191 11685
rect 2133 11645 2145 11679
rect 2179 11676 2191 11679
rect 4154 11676 4160 11688
rect 2179 11648 4160 11676
rect 2179 11645 2191 11648
rect 2133 11639 2191 11645
rect 4154 11636 4160 11648
rect 4212 11636 4218 11688
rect 5552 11685 5580 11716
rect 5813 11713 5825 11747
rect 5859 11744 5871 11747
rect 6825 11747 6883 11753
rect 5859 11716 6132 11744
rect 5859 11713 5871 11716
rect 5813 11707 5871 11713
rect 5077 11679 5135 11685
rect 5077 11645 5089 11679
rect 5123 11645 5135 11679
rect 5077 11639 5135 11645
rect 5537 11679 5595 11685
rect 5537 11645 5549 11679
rect 5583 11645 5595 11679
rect 5537 11639 5595 11645
rect 2400 11611 2458 11617
rect 2400 11577 2412 11611
rect 2446 11608 2458 11611
rect 2774 11608 2780 11620
rect 2446 11580 2780 11608
rect 2446 11577 2458 11580
rect 2400 11571 2458 11577
rect 2774 11568 2780 11580
rect 2832 11568 2838 11620
rect 5092 11608 5120 11639
rect 6104 11620 6132 11716
rect 6825 11713 6837 11747
rect 6871 11713 6883 11747
rect 6825 11707 6883 11713
rect 12437 11747 12495 11753
rect 12437 11713 12449 11747
rect 12483 11713 12495 11747
rect 12437 11707 12495 11713
rect 7098 11685 7104 11688
rect 7092 11676 7104 11685
rect 6932 11648 7104 11676
rect 5092 11580 5764 11608
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 3510 11540 3516 11552
rect 3471 11512 3516 11540
rect 3510 11500 3516 11512
rect 3568 11500 3574 11552
rect 5258 11500 5264 11552
rect 5316 11540 5322 11552
rect 5626 11540 5632 11552
rect 5316 11512 5632 11540
rect 5316 11500 5322 11512
rect 5626 11500 5632 11512
rect 5684 11500 5690 11552
rect 5736 11540 5764 11580
rect 6086 11568 6092 11620
rect 6144 11608 6150 11620
rect 6641 11611 6699 11617
rect 6641 11608 6653 11611
rect 6144 11580 6653 11608
rect 6144 11568 6150 11580
rect 6641 11577 6653 11580
rect 6687 11608 6699 11611
rect 6932 11608 6960 11648
rect 7092 11639 7104 11648
rect 7098 11636 7104 11639
rect 7156 11636 7162 11688
rect 9309 11679 9367 11685
rect 9309 11645 9321 11679
rect 9355 11676 9367 11679
rect 9398 11676 9404 11688
rect 9355 11648 9404 11676
rect 9355 11645 9367 11648
rect 9309 11639 9367 11645
rect 9398 11636 9404 11648
rect 9456 11636 9462 11688
rect 9582 11617 9588 11620
rect 9576 11608 9588 11617
rect 6687 11580 6960 11608
rect 9543 11580 9588 11608
rect 6687 11577 6699 11580
rect 6641 11571 6699 11577
rect 9576 11571 9588 11580
rect 9582 11568 9588 11571
rect 9640 11568 9646 11620
rect 12250 11568 12256 11620
rect 12308 11608 12314 11620
rect 12682 11611 12740 11617
rect 12682 11608 12694 11611
rect 12308 11580 12694 11608
rect 12308 11568 12314 11580
rect 12682 11577 12694 11580
rect 12728 11577 12740 11611
rect 12682 11571 12740 11577
rect 6362 11540 6368 11552
rect 5736 11512 6368 11540
rect 6362 11500 6368 11512
rect 6420 11500 6426 11552
rect 10686 11540 10692 11552
rect 10647 11512 10692 11540
rect 10686 11500 10692 11512
rect 10744 11500 10750 11552
rect 11701 11543 11759 11549
rect 11701 11509 11713 11543
rect 11747 11540 11759 11543
rect 11974 11540 11980 11552
rect 11747 11512 11980 11540
rect 11747 11509 11759 11512
rect 11701 11503 11759 11509
rect 11974 11500 11980 11512
rect 12032 11540 12038 11552
rect 12342 11540 12348 11552
rect 12032 11512 12348 11540
rect 12032 11500 12038 11512
rect 12342 11500 12348 11512
rect 12400 11500 12406 11552
rect 20898 11540 20904 11552
rect 20859 11512 20904 11540
rect 20898 11500 20904 11512
rect 20956 11500 20962 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1394 11336 1400 11348
rect 1355 11308 1400 11336
rect 1394 11296 1400 11308
rect 1452 11296 1458 11348
rect 1854 11336 1860 11348
rect 1815 11308 1860 11336
rect 1854 11296 1860 11308
rect 1912 11336 1918 11348
rect 3421 11339 3479 11345
rect 3421 11336 3433 11339
rect 1912 11308 3433 11336
rect 1912 11296 1918 11308
rect 3421 11305 3433 11308
rect 3467 11305 3479 11339
rect 3881 11339 3939 11345
rect 3881 11336 3893 11339
rect 3421 11299 3479 11305
rect 3620 11308 3893 11336
rect 2774 11228 2780 11280
rect 2832 11268 2838 11280
rect 2869 11271 2927 11277
rect 2869 11268 2881 11271
rect 2832 11240 2881 11268
rect 2832 11228 2838 11240
rect 2869 11237 2881 11240
rect 2915 11268 2927 11271
rect 3620 11268 3648 11308
rect 3881 11305 3893 11308
rect 3927 11336 3939 11339
rect 4614 11336 4620 11348
rect 3927 11308 4620 11336
rect 3927 11305 3939 11308
rect 3881 11299 3939 11305
rect 4614 11296 4620 11308
rect 4672 11296 4678 11348
rect 6086 11336 6092 11348
rect 6047 11308 6092 11336
rect 6086 11296 6092 11308
rect 6144 11296 6150 11348
rect 6362 11336 6368 11348
rect 6323 11308 6368 11336
rect 6362 11296 6368 11308
rect 6420 11296 6426 11348
rect 7282 11336 7288 11348
rect 7243 11308 7288 11336
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 8018 11336 8024 11348
rect 7979 11308 8024 11336
rect 8018 11296 8024 11308
rect 8076 11296 8082 11348
rect 8481 11339 8539 11345
rect 8481 11305 8493 11339
rect 8527 11336 8539 11339
rect 8938 11336 8944 11348
rect 8527 11308 8944 11336
rect 8527 11305 8539 11308
rect 8481 11299 8539 11305
rect 8938 11296 8944 11308
rect 8996 11336 9002 11348
rect 9674 11336 9680 11348
rect 8996 11308 9680 11336
rect 8996 11296 9002 11308
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 10870 11336 10876 11348
rect 10831 11308 10876 11336
rect 10870 11296 10876 11308
rect 10928 11296 10934 11348
rect 12250 11296 12256 11348
rect 12308 11336 12314 11348
rect 12437 11339 12495 11345
rect 12437 11336 12449 11339
rect 12308 11308 12449 11336
rect 12308 11296 12314 11308
rect 12437 11305 12449 11308
rect 12483 11305 12495 11339
rect 12986 11336 12992 11348
rect 12947 11308 12992 11336
rect 12437 11299 12495 11305
rect 12986 11296 12992 11308
rect 13044 11296 13050 11348
rect 4310 11271 4368 11277
rect 4310 11268 4322 11271
rect 2915 11240 3648 11268
rect 3712 11240 4322 11268
rect 2915 11237 2927 11240
rect 2869 11231 2927 11237
rect 1765 11203 1823 11209
rect 1765 11169 1777 11203
rect 1811 11200 1823 11203
rect 2409 11203 2467 11209
rect 2409 11200 2421 11203
rect 1811 11172 2421 11200
rect 1811 11169 1823 11172
rect 1765 11163 1823 11169
rect 2409 11169 2421 11172
rect 2455 11200 2467 11203
rect 2961 11203 3019 11209
rect 2961 11200 2973 11203
rect 2455 11172 2973 11200
rect 2455 11169 2467 11172
rect 2409 11163 2467 11169
rect 2961 11169 2973 11172
rect 3007 11169 3019 11203
rect 2961 11163 3019 11169
rect 3510 11160 3516 11212
rect 3568 11200 3574 11212
rect 3712 11200 3740 11240
rect 4310 11237 4322 11240
rect 4356 11237 4368 11271
rect 9950 11268 9956 11280
rect 9911 11240 9956 11268
rect 4310 11231 4368 11237
rect 9950 11228 9956 11240
rect 10008 11228 10014 11280
rect 18138 11228 18144 11280
rect 18196 11268 18202 11280
rect 18233 11271 18291 11277
rect 18233 11268 18245 11271
rect 18196 11240 18245 11268
rect 18196 11228 18202 11240
rect 18233 11237 18245 11240
rect 18279 11237 18291 11271
rect 18233 11231 18291 11237
rect 3568 11172 3740 11200
rect 4065 11203 4123 11209
rect 3568 11160 3574 11172
rect 4065 11169 4077 11203
rect 4111 11200 4123 11203
rect 4154 11200 4160 11212
rect 4111 11172 4160 11200
rect 4111 11169 4123 11172
rect 4065 11163 4123 11169
rect 4154 11160 4160 11172
rect 4212 11200 4218 11212
rect 4890 11200 4896 11212
rect 4212 11172 4896 11200
rect 4212 11160 4218 11172
rect 4890 11160 4896 11172
rect 4948 11160 4954 11212
rect 8389 11203 8447 11209
rect 8389 11169 8401 11203
rect 8435 11200 8447 11203
rect 8754 11200 8760 11212
rect 8435 11172 8760 11200
rect 8435 11169 8447 11172
rect 8389 11163 8447 11169
rect 8754 11160 8760 11172
rect 8812 11160 8818 11212
rect 9674 11200 9680 11212
rect 9587 11172 9680 11200
rect 9674 11160 9680 11172
rect 9732 11200 9738 11212
rect 9858 11200 9864 11212
rect 9732 11172 9864 11200
rect 9732 11160 9738 11172
rect 9858 11160 9864 11172
rect 9916 11160 9922 11212
rect 11054 11200 11060 11212
rect 11015 11172 11060 11200
rect 11054 11160 11060 11172
rect 11112 11160 11118 11212
rect 11330 11209 11336 11212
rect 11324 11200 11336 11209
rect 11291 11172 11336 11200
rect 11324 11163 11336 11172
rect 11330 11160 11336 11163
rect 11388 11160 11394 11212
rect 17954 11200 17960 11212
rect 17915 11172 17960 11200
rect 17954 11160 17960 11172
rect 18012 11160 18018 11212
rect 1949 11135 2007 11141
rect 1949 11101 1961 11135
rect 1995 11101 2007 11135
rect 1949 11095 2007 11101
rect 1964 11064 1992 11095
rect 8110 11092 8116 11144
rect 8168 11132 8174 11144
rect 8665 11135 8723 11141
rect 8665 11132 8677 11135
rect 8168 11104 8677 11132
rect 8168 11092 8174 11104
rect 8665 11101 8677 11104
rect 8711 11132 8723 11135
rect 9766 11132 9772 11144
rect 8711 11104 9772 11132
rect 8711 11101 8723 11104
rect 8665 11095 8723 11101
rect 9766 11092 9772 11104
rect 9824 11092 9830 11144
rect 7558 11064 7564 11076
rect 1964 11036 2728 11064
rect 7519 11036 7564 11064
rect 2700 10996 2728 11036
rect 7558 11024 7564 11036
rect 7616 11024 7622 11076
rect 9401 11067 9459 11073
rect 9401 11033 9413 11067
rect 9447 11064 9459 11067
rect 9582 11064 9588 11076
rect 9447 11036 9588 11064
rect 9447 11033 9459 11036
rect 9401 11027 9459 11033
rect 9582 11024 9588 11036
rect 9640 11064 9646 11076
rect 10134 11064 10140 11076
rect 9640 11036 10140 11064
rect 9640 11024 9646 11036
rect 10134 11024 10140 11036
rect 10192 11064 10198 11076
rect 10413 11067 10471 11073
rect 10413 11064 10425 11067
rect 10192 11036 10425 11064
rect 10192 11024 10198 11036
rect 10413 11033 10425 11036
rect 10459 11033 10471 11067
rect 10413 11027 10471 11033
rect 3326 10996 3332 11008
rect 2700 10968 3332 10996
rect 3326 10956 3332 10968
rect 3384 10956 3390 11008
rect 5442 10996 5448 11008
rect 5403 10968 5448 10996
rect 5442 10956 5448 10968
rect 5500 10956 5506 11008
rect 6454 10956 6460 11008
rect 6512 10996 6518 11008
rect 6825 10999 6883 11005
rect 6825 10996 6837 10999
rect 6512 10968 6837 10996
rect 6512 10956 6518 10968
rect 6825 10965 6837 10968
rect 6871 10965 6883 10999
rect 6825 10959 6883 10965
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 2038 10752 2044 10804
rect 2096 10792 2102 10804
rect 3418 10792 3424 10804
rect 2096 10764 3424 10792
rect 2096 10752 2102 10764
rect 3418 10752 3424 10764
rect 3476 10792 3482 10804
rect 5629 10795 5687 10801
rect 5629 10792 5641 10795
rect 3476 10764 5641 10792
rect 3476 10752 3482 10764
rect 5629 10761 5641 10764
rect 5675 10761 5687 10795
rect 8110 10792 8116 10804
rect 8071 10764 8116 10792
rect 5629 10755 5687 10761
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 8938 10792 8944 10804
rect 8899 10764 8944 10792
rect 8938 10752 8944 10764
rect 8996 10752 9002 10804
rect 9401 10795 9459 10801
rect 9401 10761 9413 10795
rect 9447 10792 9459 10795
rect 9582 10792 9588 10804
rect 9447 10764 9588 10792
rect 9447 10761 9459 10764
rect 9401 10755 9459 10761
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 12253 10795 12311 10801
rect 12253 10761 12265 10795
rect 12299 10792 12311 10795
rect 12986 10792 12992 10804
rect 12299 10764 12992 10792
rect 12299 10761 12311 10764
rect 12253 10755 12311 10761
rect 12986 10752 12992 10764
rect 13044 10752 13050 10804
rect 17954 10752 17960 10804
rect 18012 10792 18018 10804
rect 18233 10795 18291 10801
rect 18233 10792 18245 10795
rect 18012 10764 18245 10792
rect 18012 10752 18018 10764
rect 18233 10761 18245 10764
rect 18279 10761 18291 10795
rect 18233 10755 18291 10761
rect 2130 10656 2136 10668
rect 2091 10628 2136 10656
rect 2130 10616 2136 10628
rect 2188 10656 2194 10668
rect 2961 10659 3019 10665
rect 2188 10628 2728 10656
rect 2188 10616 2194 10628
rect 2700 10597 2728 10628
rect 2961 10625 2973 10659
rect 3007 10656 3019 10659
rect 3418 10656 3424 10668
rect 3007 10628 3424 10656
rect 3007 10625 3019 10628
rect 2961 10619 3019 10625
rect 3418 10616 3424 10628
rect 3476 10616 3482 10668
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4249 10659 4307 10665
rect 4249 10656 4261 10659
rect 4212 10628 4261 10656
rect 4212 10616 4218 10628
rect 4249 10625 4261 10628
rect 4295 10625 4307 10659
rect 4249 10619 4307 10625
rect 6454 10616 6460 10668
rect 6512 10656 6518 10668
rect 7377 10659 7435 10665
rect 7377 10656 7389 10659
rect 6512 10628 7389 10656
rect 6512 10616 6518 10628
rect 7377 10625 7389 10628
rect 7423 10625 7435 10659
rect 9766 10656 9772 10668
rect 9679 10628 9772 10656
rect 7377 10619 7435 10625
rect 9766 10616 9772 10628
rect 9824 10656 9830 10668
rect 9824 10628 9996 10656
rect 9824 10616 9830 10628
rect 2685 10591 2743 10597
rect 2685 10557 2697 10591
rect 2731 10557 2743 10591
rect 4516 10591 4574 10597
rect 4516 10588 4528 10591
rect 2685 10551 2743 10557
rect 4448 10560 4528 10588
rect 1857 10523 1915 10529
rect 1857 10489 1869 10523
rect 1903 10520 1915 10523
rect 2498 10520 2504 10532
rect 1903 10492 2504 10520
rect 1903 10489 1915 10492
rect 1857 10483 1915 10489
rect 2498 10480 2504 10492
rect 2556 10520 2562 10532
rect 2777 10523 2835 10529
rect 2777 10520 2789 10523
rect 2556 10492 2789 10520
rect 2556 10480 2562 10492
rect 2777 10489 2789 10492
rect 2823 10489 2835 10523
rect 2777 10483 2835 10489
rect 3142 10480 3148 10532
rect 3200 10520 3206 10532
rect 3510 10520 3516 10532
rect 3200 10492 3516 10520
rect 3200 10480 3206 10492
rect 3510 10480 3516 10492
rect 3568 10520 3574 10532
rect 3697 10523 3755 10529
rect 3697 10520 3709 10523
rect 3568 10492 3709 10520
rect 3568 10480 3574 10492
rect 3697 10489 3709 10492
rect 3743 10489 3755 10523
rect 3697 10483 3755 10489
rect 4157 10523 4215 10529
rect 4157 10489 4169 10523
rect 4203 10520 4215 10523
rect 4448 10520 4476 10560
rect 4516 10557 4528 10560
rect 4562 10588 4574 10591
rect 4798 10588 4804 10600
rect 4562 10560 4804 10588
rect 4562 10557 4574 10560
rect 4516 10551 4574 10557
rect 4798 10548 4804 10560
rect 4856 10588 4862 10600
rect 5442 10588 5448 10600
rect 4856 10560 5448 10588
rect 4856 10548 4862 10560
rect 5442 10548 5448 10560
rect 5500 10548 5506 10600
rect 6546 10548 6552 10600
rect 6604 10588 6610 10600
rect 7193 10591 7251 10597
rect 7193 10588 7205 10591
rect 6604 10560 7205 10588
rect 6604 10548 6610 10560
rect 7193 10557 7205 10560
rect 7239 10557 7251 10591
rect 7193 10551 7251 10557
rect 9674 10548 9680 10600
rect 9732 10588 9738 10600
rect 9861 10591 9919 10597
rect 9861 10588 9873 10591
rect 9732 10560 9873 10588
rect 9732 10548 9738 10560
rect 9861 10557 9873 10560
rect 9907 10557 9919 10591
rect 9968 10588 9996 10628
rect 12434 10616 12440 10668
rect 12492 10656 12498 10668
rect 18693 10659 18751 10665
rect 12492 10628 12537 10656
rect 12492 10616 12498 10628
rect 18693 10625 18705 10659
rect 18739 10656 18751 10659
rect 19426 10656 19432 10668
rect 18739 10628 19432 10656
rect 18739 10625 18751 10628
rect 18693 10619 18751 10625
rect 19426 10616 19432 10628
rect 19484 10616 19490 10668
rect 19978 10656 19984 10668
rect 19939 10628 19984 10656
rect 19978 10616 19984 10628
rect 20036 10616 20042 10668
rect 10128 10591 10186 10597
rect 10128 10588 10140 10591
rect 9968 10560 10140 10588
rect 9861 10551 9919 10557
rect 10128 10557 10140 10560
rect 10174 10588 10186 10591
rect 10686 10588 10692 10600
rect 10174 10560 10692 10588
rect 10174 10557 10186 10560
rect 10128 10551 10186 10557
rect 4203 10492 4476 10520
rect 6273 10523 6331 10529
rect 4203 10489 4215 10492
rect 4157 10483 4215 10489
rect 6273 10489 6285 10523
rect 6319 10520 6331 10523
rect 6730 10520 6736 10532
rect 6319 10492 6736 10520
rect 6319 10489 6331 10492
rect 6273 10483 6331 10489
rect 6730 10480 6736 10492
rect 6788 10520 6794 10532
rect 7285 10523 7343 10529
rect 7285 10520 7297 10523
rect 6788 10492 7297 10520
rect 6788 10480 6794 10492
rect 7285 10489 7297 10492
rect 7331 10489 7343 10523
rect 9876 10520 9904 10551
rect 10686 10548 10692 10560
rect 10744 10548 10750 10600
rect 18414 10588 18420 10600
rect 18375 10560 18420 10588
rect 18414 10548 18420 10560
rect 18472 10588 18478 10600
rect 19153 10591 19211 10597
rect 19153 10588 19165 10591
rect 18472 10560 19165 10588
rect 18472 10548 18478 10560
rect 19153 10557 19165 10560
rect 19199 10557 19211 10591
rect 19702 10588 19708 10600
rect 19663 10560 19708 10588
rect 19153 10551 19211 10557
rect 19702 10548 19708 10560
rect 19760 10588 19766 10600
rect 20441 10591 20499 10597
rect 20441 10588 20453 10591
rect 19760 10560 20453 10588
rect 19760 10548 19766 10560
rect 20441 10557 20453 10560
rect 20487 10557 20499 10591
rect 20441 10551 20499 10557
rect 11054 10520 11060 10532
rect 9876 10492 11060 10520
rect 7285 10483 7343 10489
rect 11054 10480 11060 10492
rect 11112 10480 11118 10532
rect 2317 10455 2375 10461
rect 2317 10421 2329 10455
rect 2363 10452 2375 10455
rect 2682 10452 2688 10464
rect 2363 10424 2688 10452
rect 2363 10421 2375 10424
rect 2317 10415 2375 10421
rect 2682 10412 2688 10424
rect 2740 10412 2746 10464
rect 3326 10452 3332 10464
rect 3287 10424 3332 10452
rect 3326 10412 3332 10424
rect 3384 10412 3390 10464
rect 6546 10452 6552 10464
rect 6507 10424 6552 10452
rect 6546 10412 6552 10424
rect 6604 10412 6610 10464
rect 6822 10452 6828 10464
rect 6783 10424 6828 10452
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 8386 10452 8392 10464
rect 8347 10424 8392 10452
rect 8386 10412 8392 10424
rect 8444 10412 8450 10464
rect 11241 10455 11299 10461
rect 11241 10421 11253 10455
rect 11287 10452 11299 10455
rect 11330 10452 11336 10464
rect 11287 10424 11336 10452
rect 11287 10421 11299 10424
rect 11241 10415 11299 10421
rect 11330 10412 11336 10424
rect 11388 10452 11394 10464
rect 11885 10455 11943 10461
rect 11885 10452 11897 10455
rect 11388 10424 11897 10452
rect 11388 10412 11394 10424
rect 11885 10421 11897 10424
rect 11931 10452 11943 10455
rect 11974 10452 11980 10464
rect 11931 10424 11980 10452
rect 11931 10421 11943 10424
rect 11885 10415 11943 10421
rect 11974 10412 11980 10424
rect 12032 10412 12038 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 2590 10208 2596 10260
rect 2648 10248 2654 10260
rect 2777 10251 2835 10257
rect 2777 10248 2789 10251
rect 2648 10220 2789 10248
rect 2648 10208 2654 10220
rect 2777 10217 2789 10220
rect 2823 10248 2835 10251
rect 3326 10248 3332 10260
rect 2823 10220 3332 10248
rect 2823 10217 2835 10220
rect 2777 10211 2835 10217
rect 3326 10208 3332 10220
rect 3384 10208 3390 10260
rect 3418 10208 3424 10260
rect 3476 10248 3482 10260
rect 3789 10251 3847 10257
rect 3476 10220 3521 10248
rect 3476 10208 3482 10220
rect 3789 10217 3801 10251
rect 3835 10248 3847 10251
rect 3878 10248 3884 10260
rect 3835 10220 3884 10248
rect 3835 10217 3847 10220
rect 3789 10211 3847 10217
rect 3878 10208 3884 10220
rect 3936 10248 3942 10260
rect 4154 10248 4160 10260
rect 3936 10220 4160 10248
rect 3936 10208 3942 10220
rect 4154 10208 4160 10220
rect 4212 10248 4218 10260
rect 4525 10251 4583 10257
rect 4525 10248 4537 10251
rect 4212 10220 4537 10248
rect 4212 10208 4218 10220
rect 4525 10217 4537 10220
rect 4571 10248 4583 10251
rect 4893 10251 4951 10257
rect 4893 10248 4905 10251
rect 4571 10220 4905 10248
rect 4571 10217 4583 10220
rect 4525 10211 4583 10217
rect 4893 10217 4905 10220
rect 4939 10217 4951 10251
rect 7558 10248 7564 10260
rect 7519 10220 7564 10248
rect 4893 10211 4951 10217
rect 1664 10183 1722 10189
rect 1664 10149 1676 10183
rect 1710 10180 1722 10183
rect 2038 10180 2044 10192
rect 1710 10152 2044 10180
rect 1710 10149 1722 10152
rect 1664 10143 1722 10149
rect 2038 10140 2044 10152
rect 2096 10140 2102 10192
rect 4908 10112 4936 10211
rect 7558 10208 7564 10220
rect 7616 10208 7622 10260
rect 8202 10248 8208 10260
rect 8163 10220 8208 10248
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 8386 10208 8392 10260
rect 8444 10248 8450 10260
rect 10042 10248 10048 10260
rect 8444 10220 10048 10248
rect 8444 10208 8450 10220
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 10781 10251 10839 10257
rect 10781 10217 10793 10251
rect 10827 10248 10839 10251
rect 11054 10248 11060 10260
rect 10827 10220 11060 10248
rect 10827 10217 10839 10220
rect 10781 10211 10839 10217
rect 11054 10208 11060 10220
rect 11112 10208 11118 10260
rect 11238 10248 11244 10260
rect 11199 10220 11244 10248
rect 11238 10208 11244 10220
rect 11296 10208 11302 10260
rect 8754 10180 8760 10192
rect 8715 10152 8760 10180
rect 8754 10140 8760 10152
rect 8812 10180 8818 10192
rect 9858 10180 9864 10192
rect 8812 10152 9864 10180
rect 8812 10140 8818 10152
rect 9858 10140 9864 10152
rect 9916 10140 9922 10192
rect 19797 10183 19855 10189
rect 19797 10149 19809 10183
rect 19843 10180 19855 10183
rect 21174 10180 21180 10192
rect 19843 10152 21180 10180
rect 19843 10149 19855 10152
rect 19797 10143 19855 10149
rect 21174 10140 21180 10152
rect 21232 10140 21238 10192
rect 5258 10112 5264 10124
rect 4908 10084 5264 10112
rect 5258 10072 5264 10084
rect 5316 10072 5322 10124
rect 5350 10072 5356 10124
rect 5408 10112 5414 10124
rect 5528 10115 5586 10121
rect 5528 10112 5540 10115
rect 5408 10084 5540 10112
rect 5408 10072 5414 10084
rect 5528 10081 5540 10084
rect 5574 10112 5586 10115
rect 7282 10112 7288 10124
rect 5574 10084 7288 10112
rect 5574 10081 5586 10084
rect 5528 10075 5586 10081
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 7834 10072 7840 10124
rect 7892 10112 7898 10124
rect 8113 10115 8171 10121
rect 8113 10112 8125 10115
rect 7892 10084 8125 10112
rect 7892 10072 7898 10084
rect 8113 10081 8125 10084
rect 8159 10081 8171 10115
rect 8113 10075 8171 10081
rect 11238 10072 11244 10124
rect 11296 10112 11302 10124
rect 11609 10115 11667 10121
rect 11609 10112 11621 10115
rect 11296 10084 11621 10112
rect 11296 10072 11302 10084
rect 11609 10081 11621 10084
rect 11655 10081 11667 10115
rect 19518 10112 19524 10124
rect 19479 10084 19524 10112
rect 11609 10075 11667 10081
rect 19518 10072 19524 10084
rect 19576 10072 19582 10124
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 4062 10044 4068 10056
rect 4023 10016 4068 10044
rect 4062 10004 4068 10016
rect 4120 10004 4126 10056
rect 8018 10004 8024 10056
rect 8076 10044 8082 10056
rect 8297 10047 8355 10053
rect 8297 10044 8309 10047
rect 8076 10016 8309 10044
rect 8076 10004 8082 10016
rect 8297 10013 8309 10016
rect 8343 10013 8355 10047
rect 10137 10047 10195 10053
rect 10137 10044 10149 10047
rect 8297 10007 8355 10013
rect 9416 10016 10149 10044
rect 7650 9976 7656 9988
rect 6380 9948 7656 9976
rect 3694 9868 3700 9920
rect 3752 9908 3758 9920
rect 6380 9908 6408 9948
rect 7650 9936 7656 9948
rect 7708 9936 7714 9988
rect 9416 9985 9444 10016
rect 10137 10013 10149 10016
rect 10183 10013 10195 10047
rect 10137 10007 10195 10013
rect 10229 10047 10287 10053
rect 10229 10013 10241 10047
rect 10275 10013 10287 10047
rect 11698 10044 11704 10056
rect 11659 10016 11704 10044
rect 10229 10007 10287 10013
rect 7745 9979 7803 9985
rect 7745 9945 7757 9979
rect 7791 9976 7803 9979
rect 9401 9979 9459 9985
rect 9401 9976 9413 9979
rect 7791 9948 9413 9976
rect 7791 9945 7803 9948
rect 7745 9939 7803 9945
rect 9401 9945 9413 9948
rect 9447 9945 9459 9979
rect 9674 9976 9680 9988
rect 9635 9948 9680 9976
rect 9401 9939 9459 9945
rect 9674 9936 9680 9948
rect 9732 9936 9738 9988
rect 9766 9936 9772 9988
rect 9824 9976 9830 9988
rect 10244 9976 10272 10007
rect 11698 10004 11704 10016
rect 11756 10004 11762 10056
rect 11885 10047 11943 10053
rect 11885 10013 11897 10047
rect 11931 10044 11943 10047
rect 11974 10044 11980 10056
rect 11931 10016 11980 10044
rect 11931 10013 11943 10016
rect 11885 10007 11943 10013
rect 11974 10004 11980 10016
rect 12032 10004 12038 10056
rect 9824 9948 10272 9976
rect 9824 9936 9830 9948
rect 3752 9880 6408 9908
rect 3752 9868 3758 9880
rect 6454 9868 6460 9920
rect 6512 9908 6518 9920
rect 6641 9911 6699 9917
rect 6641 9908 6653 9911
rect 6512 9880 6653 9908
rect 6512 9868 6518 9880
rect 6641 9877 6653 9880
rect 6687 9877 6699 9911
rect 7282 9908 7288 9920
rect 7243 9880 7288 9908
rect 6641 9871 6699 9877
rect 7282 9868 7288 9880
rect 7340 9868 7346 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 3053 9707 3111 9713
rect 3053 9673 3065 9707
rect 3099 9704 3111 9707
rect 3418 9704 3424 9716
rect 3099 9676 3424 9704
rect 3099 9673 3111 9676
rect 3053 9667 3111 9673
rect 3418 9664 3424 9676
rect 3476 9704 3482 9716
rect 3973 9707 4031 9713
rect 3973 9704 3985 9707
rect 3476 9676 3985 9704
rect 3476 9664 3482 9676
rect 3973 9673 3985 9676
rect 4019 9673 4031 9707
rect 3973 9667 4031 9673
rect 3326 9596 3332 9648
rect 3384 9636 3390 9648
rect 3694 9636 3700 9648
rect 3384 9608 3700 9636
rect 3384 9596 3390 9608
rect 3694 9596 3700 9608
rect 3752 9596 3758 9648
rect 1394 9528 1400 9580
rect 1452 9568 1458 9580
rect 1673 9571 1731 9577
rect 1673 9568 1685 9571
rect 1452 9540 1685 9568
rect 1452 9528 1458 9540
rect 1673 9537 1685 9540
rect 1719 9537 1731 9571
rect 3988 9568 4016 9667
rect 6730 9664 6736 9716
rect 6788 9704 6794 9716
rect 6825 9707 6883 9713
rect 6825 9704 6837 9707
rect 6788 9676 6837 9704
rect 6788 9664 6794 9676
rect 6825 9673 6837 9676
rect 6871 9673 6883 9707
rect 8202 9704 8208 9716
rect 8163 9676 8208 9704
rect 6825 9667 6883 9673
rect 8202 9664 8208 9676
rect 8260 9664 8266 9716
rect 10042 9664 10048 9716
rect 10100 9704 10106 9716
rect 10597 9707 10655 9713
rect 10597 9704 10609 9707
rect 10100 9676 10609 9704
rect 10100 9664 10106 9676
rect 10597 9673 10609 9676
rect 10643 9673 10655 9707
rect 11698 9704 11704 9716
rect 11659 9676 11704 9704
rect 10597 9667 10655 9673
rect 11698 9664 11704 9676
rect 11756 9664 11762 9716
rect 11974 9704 11980 9716
rect 11935 9676 11980 9704
rect 11974 9664 11980 9676
rect 12032 9664 12038 9716
rect 19518 9704 19524 9716
rect 19479 9676 19524 9704
rect 19518 9664 19524 9676
rect 19576 9664 19582 9716
rect 10686 9596 10692 9648
rect 10744 9636 10750 9648
rect 11514 9636 11520 9648
rect 10744 9608 11520 9636
rect 10744 9596 10750 9608
rect 11514 9596 11520 9608
rect 11572 9596 11578 9648
rect 12434 9596 12440 9648
rect 12492 9636 12498 9648
rect 15286 9636 15292 9648
rect 12492 9608 15292 9636
rect 12492 9596 12498 9608
rect 15286 9596 15292 9608
rect 15344 9596 15350 9648
rect 3988 9540 4292 9568
rect 1673 9531 1731 9537
rect 1688 9500 1716 9531
rect 3605 9503 3663 9509
rect 3605 9500 3617 9503
rect 1688 9472 3617 9500
rect 3605 9469 3617 9472
rect 3651 9500 3663 9503
rect 3878 9500 3884 9512
rect 3651 9472 3884 9500
rect 3651 9469 3663 9472
rect 3605 9463 3663 9469
rect 3878 9460 3884 9472
rect 3936 9500 3942 9512
rect 4157 9503 4215 9509
rect 4157 9500 4169 9503
rect 3936 9472 4169 9500
rect 3936 9460 3942 9472
rect 4157 9469 4169 9472
rect 4203 9469 4215 9503
rect 4264 9500 4292 9540
rect 7282 9528 7288 9580
rect 7340 9568 7346 9580
rect 7377 9571 7435 9577
rect 7377 9568 7389 9571
rect 7340 9540 7389 9568
rect 7340 9528 7346 9540
rect 7377 9537 7389 9540
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 4413 9503 4471 9509
rect 4413 9500 4425 9503
rect 4264 9472 4425 9500
rect 4157 9463 4215 9469
rect 4413 9469 4425 9472
rect 4459 9469 4471 9503
rect 6549 9503 6607 9509
rect 6549 9500 6561 9503
rect 4413 9463 4471 9469
rect 4632 9472 6561 9500
rect 1762 9392 1768 9444
rect 1820 9432 1826 9444
rect 1940 9435 1998 9441
rect 1940 9432 1952 9435
rect 1820 9404 1952 9432
rect 1820 9392 1826 9404
rect 1940 9401 1952 9404
rect 1986 9432 1998 9435
rect 2590 9432 2596 9444
rect 1986 9404 2596 9432
rect 1986 9401 1998 9404
rect 1940 9395 1998 9401
rect 2590 9392 2596 9404
rect 2648 9392 2654 9444
rect 2498 9324 2504 9376
rect 2556 9364 2562 9376
rect 4632 9364 4660 9472
rect 6549 9469 6561 9472
rect 6595 9500 6607 9503
rect 7193 9503 7251 9509
rect 7193 9500 7205 9503
rect 6595 9472 7205 9500
rect 6595 9469 6607 9472
rect 6549 9463 6607 9469
rect 7193 9469 7205 9472
rect 7239 9469 7251 9503
rect 7834 9500 7840 9512
rect 7795 9472 7840 9500
rect 7193 9463 7251 9469
rect 7834 9460 7840 9472
rect 7892 9460 7898 9512
rect 8662 9500 8668 9512
rect 8623 9472 8668 9500
rect 8662 9460 8668 9472
rect 8720 9500 8726 9512
rect 9490 9500 9496 9512
rect 8720 9472 9496 9500
rect 8720 9460 8726 9472
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 6273 9435 6331 9441
rect 6273 9401 6285 9435
rect 6319 9432 6331 9435
rect 7006 9432 7012 9444
rect 6319 9404 7012 9432
rect 6319 9401 6331 9404
rect 6273 9395 6331 9401
rect 7006 9392 7012 9404
rect 7064 9432 7070 9444
rect 8938 9441 8944 9444
rect 7285 9435 7343 9441
rect 7285 9432 7297 9435
rect 7064 9404 7297 9432
rect 7064 9392 7070 9404
rect 7285 9401 7297 9404
rect 7331 9401 7343 9435
rect 8932 9432 8944 9441
rect 8899 9404 8944 9432
rect 7285 9395 7343 9401
rect 8932 9395 8944 9404
rect 8938 9392 8944 9395
rect 8996 9392 9002 9444
rect 2556 9336 4660 9364
rect 2556 9324 2562 9336
rect 4706 9324 4712 9376
rect 4764 9364 4770 9376
rect 5537 9367 5595 9373
rect 5537 9364 5549 9367
rect 4764 9336 5549 9364
rect 4764 9324 4770 9336
rect 5537 9333 5549 9336
rect 5583 9333 5595 9367
rect 5537 9327 5595 9333
rect 10045 9367 10103 9373
rect 10045 9333 10057 9367
rect 10091 9364 10103 9367
rect 10134 9364 10140 9376
rect 10091 9336 10140 9364
rect 10091 9333 10103 9336
rect 10045 9327 10103 9333
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 11054 9324 11060 9376
rect 11112 9364 11118 9376
rect 11238 9364 11244 9376
rect 11112 9336 11244 9364
rect 11112 9324 11118 9336
rect 11238 9324 11244 9336
rect 11296 9324 11302 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1762 9160 1768 9172
rect 1723 9132 1768 9160
rect 1762 9120 1768 9132
rect 1820 9120 1826 9172
rect 2038 9160 2044 9172
rect 1999 9132 2044 9160
rect 2038 9120 2044 9132
rect 2096 9120 2102 9172
rect 2774 9120 2780 9172
rect 2832 9160 2838 9172
rect 3789 9163 3847 9169
rect 3789 9160 3801 9163
rect 2832 9132 3801 9160
rect 2832 9120 2838 9132
rect 3789 9129 3801 9132
rect 3835 9160 3847 9163
rect 4525 9163 4583 9169
rect 4525 9160 4537 9163
rect 3835 9132 4537 9160
rect 3835 9129 3847 9132
rect 3789 9123 3847 9129
rect 4525 9129 4537 9132
rect 4571 9129 4583 9163
rect 5350 9160 5356 9172
rect 5311 9132 5356 9160
rect 4525 9123 4583 9129
rect 5350 9120 5356 9132
rect 5408 9120 5414 9172
rect 7745 9163 7803 9169
rect 7745 9129 7757 9163
rect 7791 9160 7803 9163
rect 8018 9160 8024 9172
rect 7791 9132 8024 9160
rect 7791 9129 7803 9132
rect 7745 9123 7803 9129
rect 8018 9120 8024 9132
rect 8076 9160 8082 9172
rect 8297 9163 8355 9169
rect 8297 9160 8309 9163
rect 8076 9132 8309 9160
rect 8076 9120 8082 9132
rect 8297 9129 8309 9132
rect 8343 9129 8355 9163
rect 8297 9123 8355 9129
rect 8757 9163 8815 9169
rect 8757 9129 8769 9163
rect 8803 9160 8815 9163
rect 8938 9160 8944 9172
rect 8803 9132 8944 9160
rect 8803 9129 8815 9132
rect 8757 9123 8815 9129
rect 8938 9120 8944 9132
rect 8996 9160 9002 9172
rect 9493 9163 9551 9169
rect 9493 9160 9505 9163
rect 8996 9132 9505 9160
rect 8996 9120 9002 9132
rect 9493 9129 9505 9132
rect 9539 9160 9551 9163
rect 9582 9160 9588 9172
rect 9539 9132 9588 9160
rect 9539 9129 9551 9132
rect 9493 9123 9551 9129
rect 9582 9120 9588 9132
rect 9640 9120 9646 9172
rect 9677 9163 9735 9169
rect 9677 9129 9689 9163
rect 9723 9160 9735 9163
rect 9858 9160 9864 9172
rect 9723 9132 9864 9160
rect 9723 9129 9735 9132
rect 9677 9123 9735 9129
rect 9858 9120 9864 9132
rect 9916 9120 9922 9172
rect 2869 9095 2927 9101
rect 2869 9061 2881 9095
rect 2915 9092 2927 9095
rect 3050 9092 3056 9104
rect 2915 9064 3056 9092
rect 2915 9061 2927 9064
rect 2869 9055 2927 9061
rect 3050 9052 3056 9064
rect 3108 9052 3114 9104
rect 4062 9052 4068 9104
rect 4120 9092 4126 9104
rect 4433 9095 4491 9101
rect 4433 9092 4445 9095
rect 4120 9064 4445 9092
rect 4120 9052 4126 9064
rect 4433 9061 4445 9064
rect 4479 9061 4491 9095
rect 4433 9055 4491 9061
rect 5258 9052 5264 9104
rect 5316 9092 5322 9104
rect 5629 9095 5687 9101
rect 5629 9092 5641 9095
rect 5316 9064 5641 9092
rect 5316 9052 5322 9064
rect 5629 9061 5641 9064
rect 5675 9092 5687 9095
rect 7006 9092 7012 9104
rect 5675 9064 7012 9092
rect 5675 9061 5687 9064
rect 5629 9055 5687 9061
rect 2774 8984 2780 9036
rect 2832 9024 2838 9036
rect 3513 9027 3571 9033
rect 2832 8996 2877 9024
rect 2832 8984 2838 8996
rect 3513 8993 3525 9027
rect 3559 9024 3571 9027
rect 3786 9024 3792 9036
rect 3559 8996 3792 9024
rect 3559 8993 3571 8996
rect 3513 8987 3571 8993
rect 3786 8984 3792 8996
rect 3844 8984 3850 9036
rect 6380 9033 6408 9064
rect 7006 9052 7012 9064
rect 7064 9052 7070 9104
rect 8662 9052 8668 9104
rect 8720 9092 8726 9104
rect 9033 9095 9091 9101
rect 9033 9092 9045 9095
rect 8720 9064 9045 9092
rect 8720 9052 8726 9064
rect 9033 9061 9045 9064
rect 9079 9061 9091 9095
rect 9033 9055 9091 9061
rect 6365 9027 6423 9033
rect 6365 8993 6377 9027
rect 6411 8993 6423 9027
rect 6365 8987 6423 8993
rect 6454 8984 6460 9036
rect 6512 9024 6518 9036
rect 6621 9027 6679 9033
rect 6621 9024 6633 9027
rect 6512 8996 6633 9024
rect 6512 8984 6518 8996
rect 6621 8993 6633 8996
rect 6667 8993 6679 9027
rect 10042 9024 10048 9036
rect 10003 8996 10048 9024
rect 6621 8987 6679 8993
rect 10042 8984 10048 8996
rect 10100 8984 10106 9036
rect 3053 8959 3111 8965
rect 3053 8925 3065 8959
rect 3099 8956 3111 8959
rect 3142 8956 3148 8968
rect 3099 8928 3148 8956
rect 3099 8925 3111 8928
rect 3053 8919 3111 8925
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 4706 8956 4712 8968
rect 4667 8928 4712 8956
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 9674 8916 9680 8968
rect 9732 8956 9738 8968
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 9732 8928 10149 8956
rect 9732 8916 9738 8928
rect 10137 8925 10149 8928
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 10226 8916 10232 8968
rect 10284 8956 10290 8968
rect 10321 8959 10379 8965
rect 10321 8956 10333 8959
rect 10284 8928 10333 8956
rect 10284 8916 10290 8928
rect 10321 8925 10333 8928
rect 10367 8956 10379 8959
rect 10594 8956 10600 8968
rect 10367 8928 10600 8956
rect 10367 8925 10379 8928
rect 10321 8919 10379 8925
rect 10594 8916 10600 8928
rect 10652 8916 10658 8968
rect 3970 8848 3976 8900
rect 4028 8888 4034 8900
rect 4065 8891 4123 8897
rect 4065 8888 4077 8891
rect 4028 8860 4077 8888
rect 4028 8848 4034 8860
rect 4065 8857 4077 8860
rect 4111 8857 4123 8891
rect 4065 8851 4123 8857
rect 2406 8820 2412 8832
rect 2367 8792 2412 8820
rect 2406 8780 2412 8792
rect 2464 8780 2470 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1394 8576 1400 8628
rect 1452 8616 1458 8628
rect 1581 8619 1639 8625
rect 1581 8616 1593 8619
rect 1452 8588 1593 8616
rect 1452 8576 1458 8588
rect 1581 8585 1593 8588
rect 1627 8616 1639 8619
rect 1949 8619 2007 8625
rect 1949 8616 1961 8619
rect 1627 8588 1961 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 1949 8585 1961 8588
rect 1995 8585 2007 8619
rect 1949 8579 2007 8585
rect 2501 8619 2559 8625
rect 2501 8585 2513 8619
rect 2547 8616 2559 8619
rect 2774 8616 2780 8628
rect 2547 8588 2780 8616
rect 2547 8585 2559 8588
rect 2501 8579 2559 8585
rect 2774 8576 2780 8588
rect 2832 8576 2838 8628
rect 2869 8619 2927 8625
rect 2869 8585 2881 8619
rect 2915 8616 2927 8619
rect 3050 8616 3056 8628
rect 2915 8588 3056 8616
rect 2915 8585 2927 8588
rect 2869 8579 2927 8585
rect 3050 8576 3056 8588
rect 3108 8576 3114 8628
rect 3973 8619 4031 8625
rect 3973 8585 3985 8619
rect 4019 8616 4031 8619
rect 4062 8616 4068 8628
rect 4019 8588 4068 8616
rect 4019 8585 4031 8588
rect 3973 8579 4031 8585
rect 4062 8576 4068 8588
rect 4120 8576 4126 8628
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 5445 8619 5503 8625
rect 5445 8616 5457 8619
rect 5408 8588 5457 8616
rect 5408 8576 5414 8588
rect 5445 8585 5457 8588
rect 5491 8585 5503 8619
rect 6454 8616 6460 8628
rect 6415 8588 6460 8616
rect 5445 8579 5503 8585
rect 6454 8576 6460 8588
rect 6512 8576 6518 8628
rect 7006 8616 7012 8628
rect 6967 8588 7012 8616
rect 7006 8576 7012 8588
rect 7064 8576 7070 8628
rect 7561 8619 7619 8625
rect 7561 8585 7573 8619
rect 7607 8616 7619 8619
rect 8018 8616 8024 8628
rect 7607 8588 8024 8616
rect 7607 8585 7619 8588
rect 7561 8579 7619 8585
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 8938 8576 8944 8628
rect 8996 8616 9002 8628
rect 9033 8619 9091 8625
rect 9033 8616 9045 8619
rect 8996 8588 9045 8616
rect 8996 8576 9002 8588
rect 9033 8585 9045 8588
rect 9079 8585 9091 8619
rect 10594 8616 10600 8628
rect 10555 8588 10600 8616
rect 9033 8579 9091 8585
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 3142 8548 3148 8560
rect 3103 8520 3148 8548
rect 3142 8508 3148 8520
rect 3200 8508 3206 8560
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8480 3663 8483
rect 3878 8480 3884 8492
rect 3651 8452 3884 8480
rect 3651 8449 3663 8452
rect 3605 8443 3663 8449
rect 3878 8440 3884 8452
rect 3936 8480 3942 8492
rect 7024 8480 7052 8576
rect 9674 8548 9680 8560
rect 9635 8520 9680 8548
rect 9674 8508 9680 8520
rect 9732 8508 9738 8560
rect 7650 8480 7656 8492
rect 3936 8452 4200 8480
rect 7024 8452 7656 8480
rect 3936 8440 3942 8452
rect 3970 8372 3976 8424
rect 4028 8412 4034 8424
rect 4065 8415 4123 8421
rect 4065 8412 4077 8415
rect 4028 8384 4077 8412
rect 4028 8372 4034 8384
rect 4065 8381 4077 8384
rect 4111 8381 4123 8415
rect 4172 8412 4200 8452
rect 7650 8440 7656 8452
rect 7708 8440 7714 8492
rect 10042 8440 10048 8492
rect 10100 8480 10106 8492
rect 10137 8483 10195 8489
rect 10137 8480 10149 8483
rect 10100 8452 10149 8480
rect 10100 8440 10106 8452
rect 10137 8449 10149 8452
rect 10183 8449 10195 8483
rect 10137 8443 10195 8449
rect 4332 8415 4390 8421
rect 4332 8412 4344 8415
rect 4172 8384 4344 8412
rect 4065 8375 4123 8381
rect 4332 8381 4344 8384
rect 4378 8412 4390 8415
rect 4706 8412 4712 8424
rect 4378 8384 4712 8412
rect 4378 8381 4390 8384
rect 4332 8375 4390 8381
rect 4706 8372 4712 8384
rect 4764 8372 4770 8424
rect 7920 8347 7978 8353
rect 7920 8313 7932 8347
rect 7966 8344 7978 8347
rect 8018 8344 8024 8356
rect 7966 8316 8024 8344
rect 7966 8313 7978 8316
rect 7920 8307 7978 8313
rect 8018 8304 8024 8316
rect 8076 8304 8082 8356
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 3878 8072 3884 8084
rect 3839 8044 3884 8072
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 4522 8072 4528 8084
rect 4483 8044 4528 8072
rect 4522 8032 4528 8044
rect 4580 8032 4586 8084
rect 5813 8075 5871 8081
rect 5813 8041 5825 8075
rect 5859 8072 5871 8075
rect 6546 8072 6552 8084
rect 5859 8044 6552 8072
rect 5859 8041 5871 8044
rect 5813 8035 5871 8041
rect 6546 8032 6552 8044
rect 6604 8032 6610 8084
rect 7650 8072 7656 8084
rect 7611 8044 7656 8072
rect 7650 8032 7656 8044
rect 7708 8032 7714 8084
rect 9953 8075 10011 8081
rect 9953 8041 9965 8075
rect 9999 8072 10011 8075
rect 10042 8072 10048 8084
rect 9999 8044 10048 8072
rect 9999 8041 10011 8044
rect 9953 8035 10011 8041
rect 10042 8032 10048 8044
rect 10100 8032 10106 8084
rect 22465 8075 22523 8081
rect 22465 8041 22477 8075
rect 22511 8072 22523 8075
rect 23382 8072 23388 8084
rect 22511 8044 23388 8072
rect 22511 8041 22523 8044
rect 22465 8035 22523 8041
rect 23382 8032 23388 8044
rect 23440 8032 23446 8084
rect 3513 8007 3571 8013
rect 3513 7973 3525 8007
rect 3559 8004 3571 8007
rect 3970 8004 3976 8016
rect 3559 7976 3976 8004
rect 3559 7973 3571 7976
rect 3513 7967 3571 7973
rect 3970 7964 3976 7976
rect 4028 7964 4034 8016
rect 4154 7964 4160 8016
rect 4212 8004 4218 8016
rect 4433 8007 4491 8013
rect 4433 8004 4445 8007
rect 4212 7976 4445 8004
rect 4212 7964 4218 7976
rect 4433 7973 4445 7976
rect 4479 7973 4491 8007
rect 4433 7967 4491 7973
rect 22278 7936 22284 7948
rect 22239 7908 22284 7936
rect 22278 7896 22284 7908
rect 22336 7896 22342 7948
rect 4709 7871 4767 7877
rect 4709 7837 4721 7871
rect 4755 7868 4767 7871
rect 4798 7868 4804 7880
rect 4755 7840 4804 7868
rect 4755 7837 4767 7840
rect 4709 7831 4767 7837
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 4062 7800 4068 7812
rect 4023 7772 4068 7800
rect 4062 7760 4068 7772
rect 4120 7760 4126 7812
rect 566 7692 572 7744
rect 624 7732 630 7744
rect 4890 7732 4896 7744
rect 624 7704 4896 7732
rect 624 7692 630 7704
rect 4890 7692 4896 7704
rect 4948 7692 4954 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 4154 7528 4160 7540
rect 4115 7500 4160 7528
rect 4154 7488 4160 7500
rect 4212 7488 4218 7540
rect 4522 7488 4528 7540
rect 4580 7528 4586 7540
rect 4801 7531 4859 7537
rect 4801 7528 4813 7531
rect 4580 7500 4813 7528
rect 4580 7488 4586 7500
rect 4801 7497 4813 7500
rect 4847 7497 4859 7531
rect 22278 7528 22284 7540
rect 22239 7500 22284 7528
rect 4801 7491 4859 7497
rect 22278 7488 22284 7500
rect 22336 7488 22342 7540
rect 23842 7528 23848 7540
rect 23803 7500 23848 7528
rect 23842 7488 23848 7500
rect 23900 7488 23906 7540
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7392 4583 7395
rect 4798 7392 4804 7404
rect 4571 7364 4804 7392
rect 4571 7361 4583 7364
rect 4525 7355 4583 7361
rect 4798 7352 4804 7364
rect 4856 7352 4862 7404
rect 23658 7324 23664 7336
rect 23619 7296 23664 7324
rect 23658 7284 23664 7296
rect 23716 7324 23722 7336
rect 24213 7327 24271 7333
rect 24213 7324 24225 7327
rect 23716 7296 24225 7324
rect 23716 7284 23722 7296
rect 24213 7293 24225 7296
rect 24259 7293 24271 7327
rect 24213 7287 24271 7293
rect 566 7148 572 7200
rect 624 7188 630 7200
rect 3418 7188 3424 7200
rect 624 7160 3424 7188
rect 624 7148 630 7160
rect 3418 7148 3424 7160
rect 3476 7148 3482 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 23845 6443 23903 6449
rect 23845 6409 23857 6443
rect 23891 6440 23903 6443
rect 24762 6440 24768 6452
rect 23891 6412 24768 6440
rect 23891 6409 23903 6412
rect 23845 6403 23903 6409
rect 24762 6400 24768 6412
rect 24820 6400 24826 6452
rect 23658 6236 23664 6248
rect 23619 6208 23664 6236
rect 23658 6196 23664 6208
rect 23716 6236 23722 6248
rect 24213 6239 24271 6245
rect 24213 6236 24225 6239
rect 23716 6208 24225 6236
rect 23716 6196 23722 6208
rect 24213 6205 24225 6208
rect 24259 6205 24271 6239
rect 24213 6199 24271 6205
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 24213 5899 24271 5905
rect 24213 5865 24225 5899
rect 24259 5896 24271 5899
rect 24762 5896 24768 5908
rect 24259 5868 24768 5896
rect 24259 5865 24271 5868
rect 24213 5859 24271 5865
rect 24762 5856 24768 5868
rect 24820 5856 24826 5908
rect 24026 5760 24032 5772
rect 23987 5732 24032 5760
rect 24026 5720 24032 5732
rect 24084 5720 24090 5772
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 24026 5352 24032 5364
rect 23987 5324 24032 5352
rect 24026 5312 24032 5324
rect 24084 5312 24090 5364
rect 24670 5352 24676 5364
rect 24631 5324 24676 5352
rect 24670 5312 24676 5324
rect 24728 5312 24734 5364
rect 24486 5148 24492 5160
rect 24447 5120 24492 5148
rect 24486 5108 24492 5120
rect 24544 5148 24550 5160
rect 25041 5151 25099 5157
rect 25041 5148 25053 5151
rect 24544 5120 25053 5148
rect 24544 5108 24550 5120
rect 25041 5117 25053 5120
rect 25087 5117 25099 5151
rect 25041 5111 25099 5117
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 24762 4808 24768 4820
rect 24723 4780 24768 4808
rect 24762 4768 24768 4780
rect 24820 4768 24826 4820
rect 24578 4672 24584 4684
rect 24539 4644 24584 4672
rect 24578 4632 24584 4644
rect 24636 4632 24642 4684
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 24670 4264 24676 4276
rect 24631 4236 24676 4264
rect 24670 4224 24676 4236
rect 24728 4224 24734 4276
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 3884 26664 3936 26716
rect 7104 26664 7156 26716
rect 4068 26392 4120 26444
rect 5540 26392 5592 26444
rect 3516 26256 3568 26308
rect 4896 26256 4948 26308
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 3332 25440 3384 25492
rect 2320 25372 2372 25424
rect 9956 25440 10008 25492
rect 5356 25372 5408 25424
rect 6552 25372 6604 25424
rect 2504 25347 2556 25356
rect 2504 25313 2513 25347
rect 2513 25313 2547 25347
rect 2547 25313 2556 25347
rect 2504 25304 2556 25313
rect 2596 25304 2648 25356
rect 4160 25304 4212 25356
rect 6000 25304 6052 25356
rect 5264 25236 5316 25288
rect 2872 25168 2924 25220
rect 3792 25168 3844 25220
rect 2044 25143 2096 25152
rect 2044 25109 2053 25143
rect 2053 25109 2087 25143
rect 2087 25109 2096 25143
rect 2044 25100 2096 25109
rect 2412 25143 2464 25152
rect 2412 25109 2421 25143
rect 2421 25109 2455 25143
rect 2455 25109 2464 25143
rect 2412 25100 2464 25109
rect 2780 25100 2832 25152
rect 4712 25143 4764 25152
rect 4712 25109 4721 25143
rect 4721 25109 4755 25143
rect 4755 25109 4764 25143
rect 4712 25100 4764 25109
rect 4896 25168 4948 25220
rect 7104 25211 7156 25220
rect 7104 25177 7113 25211
rect 7113 25177 7147 25211
rect 7147 25177 7156 25211
rect 7104 25168 7156 25177
rect 10784 25100 10836 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 2504 24896 2556 24948
rect 4160 24896 4212 24948
rect 2044 24828 2096 24880
rect 2320 24803 2372 24812
rect 2320 24769 2329 24803
rect 2329 24769 2363 24803
rect 2363 24769 2372 24803
rect 2320 24760 2372 24769
rect 4712 24760 4764 24812
rect 5356 24760 5408 24812
rect 6000 24760 6052 24812
rect 6552 24803 6604 24812
rect 6552 24769 6561 24803
rect 6561 24769 6595 24803
rect 6595 24769 6604 24803
rect 6552 24760 6604 24769
rect 2688 24692 2740 24744
rect 5264 24692 5316 24744
rect 9220 24760 9272 24812
rect 9772 24760 9824 24812
rect 10784 24803 10836 24812
rect 10784 24769 10793 24803
rect 10793 24769 10827 24803
rect 10827 24769 10836 24803
rect 10784 24760 10836 24769
rect 10968 24803 11020 24812
rect 10968 24769 10977 24803
rect 10977 24769 11011 24803
rect 11011 24769 11020 24803
rect 10968 24760 11020 24769
rect 12808 24760 12860 24812
rect 13084 24803 13136 24812
rect 13084 24769 13093 24803
rect 13093 24769 13127 24803
rect 13127 24769 13136 24803
rect 13084 24760 13136 24769
rect 23848 24760 23900 24812
rect 24768 24760 24820 24812
rect 7840 24692 7892 24744
rect 15568 24692 15620 24744
rect 7012 24624 7064 24676
rect 3056 24599 3108 24608
rect 3056 24565 3065 24599
rect 3065 24565 3099 24599
rect 3099 24565 3108 24599
rect 3056 24556 3108 24565
rect 6276 24599 6328 24608
rect 6276 24565 6285 24599
rect 6285 24565 6319 24599
rect 6319 24565 6328 24599
rect 6276 24556 6328 24565
rect 7104 24556 7156 24608
rect 8208 24556 8260 24608
rect 10140 24599 10192 24608
rect 10140 24565 10149 24599
rect 10149 24565 10183 24599
rect 10183 24565 10192 24599
rect 10140 24556 10192 24565
rect 12532 24556 12584 24608
rect 16488 24624 16540 24676
rect 15568 24556 15620 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 4160 24352 4212 24404
rect 4712 24352 4764 24404
rect 6000 24395 6052 24404
rect 6000 24361 6009 24395
rect 6009 24361 6043 24395
rect 6043 24361 6052 24395
rect 6000 24352 6052 24361
rect 7012 24395 7064 24404
rect 7012 24361 7021 24395
rect 7021 24361 7055 24395
rect 7055 24361 7064 24395
rect 7012 24352 7064 24361
rect 8484 24395 8536 24404
rect 8484 24361 8493 24395
rect 8493 24361 8527 24395
rect 8527 24361 8536 24395
rect 8484 24352 8536 24361
rect 16212 24352 16264 24404
rect 17408 24352 17460 24404
rect 18512 24352 18564 24404
rect 19064 24395 19116 24404
rect 19064 24361 19073 24395
rect 19073 24361 19107 24395
rect 19107 24361 19116 24395
rect 19064 24352 19116 24361
rect 22468 24352 22520 24404
rect 4436 24284 4488 24336
rect 2412 24216 2464 24268
rect 2504 24216 2556 24268
rect 2872 24259 2924 24268
rect 2872 24225 2881 24259
rect 2881 24225 2915 24259
rect 2915 24225 2924 24259
rect 2872 24216 2924 24225
rect 4068 24259 4120 24268
rect 4068 24225 4077 24259
rect 4077 24225 4111 24259
rect 4111 24225 4120 24259
rect 4068 24216 4120 24225
rect 4528 24216 4580 24268
rect 5356 24216 5408 24268
rect 6552 24216 6604 24268
rect 7840 24284 7892 24336
rect 10968 24284 11020 24336
rect 7380 24259 7432 24268
rect 7380 24225 7414 24259
rect 7414 24225 7432 24259
rect 7380 24216 7432 24225
rect 10692 24216 10744 24268
rect 14188 24216 14240 24268
rect 16396 24259 16448 24268
rect 16396 24225 16405 24259
rect 16405 24225 16439 24259
rect 16439 24225 16448 24259
rect 16396 24216 16448 24225
rect 17500 24259 17552 24268
rect 17500 24225 17509 24259
rect 17509 24225 17543 24259
rect 17543 24225 17552 24259
rect 17500 24216 17552 24225
rect 18880 24259 18932 24268
rect 18880 24225 18889 24259
rect 18889 24225 18923 24259
rect 18923 24225 18932 24259
rect 18880 24216 18932 24225
rect 21180 24216 21232 24268
rect 6460 24148 6512 24200
rect 13268 24191 13320 24200
rect 13268 24157 13277 24191
rect 13277 24157 13311 24191
rect 13311 24157 13320 24191
rect 13268 24148 13320 24157
rect 3332 24080 3384 24132
rect 2964 24012 3016 24064
rect 4436 24012 4488 24064
rect 11980 24055 12032 24064
rect 11980 24021 11989 24055
rect 11989 24021 12023 24055
rect 12023 24021 12032 24055
rect 11980 24012 12032 24021
rect 12532 24055 12584 24064
rect 12532 24021 12541 24055
rect 12541 24021 12575 24055
rect 12575 24021 12584 24055
rect 12532 24012 12584 24021
rect 14648 24012 14700 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 2412 23808 2464 23860
rect 2872 23808 2924 23860
rect 6000 23808 6052 23860
rect 6552 23851 6604 23860
rect 6552 23817 6561 23851
rect 6561 23817 6595 23851
rect 6595 23817 6604 23851
rect 6552 23808 6604 23817
rect 9220 23851 9272 23860
rect 9220 23817 9229 23851
rect 9229 23817 9263 23851
rect 9263 23817 9272 23851
rect 9220 23808 9272 23817
rect 10968 23808 11020 23860
rect 19156 23808 19208 23860
rect 20260 23808 20312 23860
rect 20444 23851 20496 23860
rect 20444 23817 20453 23851
rect 20453 23817 20487 23851
rect 20487 23817 20496 23851
rect 20444 23808 20496 23817
rect 21548 23851 21600 23860
rect 21548 23817 21557 23851
rect 21557 23817 21591 23851
rect 21591 23817 21600 23851
rect 21548 23808 21600 23817
rect 23388 23808 23440 23860
rect 3240 23715 3292 23724
rect 3240 23681 3249 23715
rect 3249 23681 3283 23715
rect 3283 23681 3292 23715
rect 3240 23672 3292 23681
rect 7840 23715 7892 23724
rect 7840 23681 7849 23715
rect 7849 23681 7883 23715
rect 7883 23681 7892 23715
rect 7840 23672 7892 23681
rect 12256 23740 12308 23792
rect 11428 23715 11480 23724
rect 11428 23681 11437 23715
rect 11437 23681 11471 23715
rect 11471 23681 11480 23715
rect 11428 23672 11480 23681
rect 11980 23672 12032 23724
rect 14648 23672 14700 23724
rect 18328 23672 18380 23724
rect 4528 23647 4580 23656
rect 4528 23613 4562 23647
rect 4562 23613 4580 23647
rect 2044 23579 2096 23588
rect 2044 23545 2053 23579
rect 2053 23545 2087 23579
rect 2087 23545 2096 23579
rect 2044 23536 2096 23545
rect 3332 23536 3384 23588
rect 4068 23536 4120 23588
rect 4528 23604 4580 23613
rect 12440 23647 12492 23656
rect 12440 23613 12449 23647
rect 12449 23613 12483 23647
rect 12483 23613 12492 23647
rect 12440 23604 12492 23613
rect 13820 23604 13872 23656
rect 4436 23536 4488 23588
rect 6460 23536 6512 23588
rect 8116 23579 8168 23588
rect 8116 23545 8128 23579
rect 8128 23545 8168 23579
rect 8116 23536 8168 23545
rect 1400 23468 1452 23520
rect 3424 23468 3476 23520
rect 5540 23468 5592 23520
rect 6828 23511 6880 23520
rect 6828 23477 6837 23511
rect 6837 23477 6871 23511
rect 6871 23477 6880 23511
rect 6828 23468 6880 23477
rect 7380 23511 7432 23520
rect 7380 23477 7389 23511
rect 7389 23477 7423 23511
rect 7423 23477 7432 23511
rect 7380 23468 7432 23477
rect 8300 23468 8352 23520
rect 10048 23468 10100 23520
rect 10784 23511 10836 23520
rect 10784 23477 10793 23511
rect 10793 23477 10827 23511
rect 10827 23477 10836 23511
rect 10784 23468 10836 23477
rect 11980 23468 12032 23520
rect 13084 23536 13136 23588
rect 17960 23604 18012 23656
rect 19984 23604 20036 23656
rect 20996 23604 21048 23656
rect 22100 23604 22152 23656
rect 12440 23468 12492 23520
rect 14188 23468 14240 23520
rect 15476 23536 15528 23588
rect 18144 23536 18196 23588
rect 18880 23536 18932 23588
rect 16396 23468 16448 23520
rect 17500 23511 17552 23520
rect 17500 23477 17509 23511
rect 17509 23477 17543 23511
rect 17543 23477 17552 23511
rect 17500 23468 17552 23477
rect 21180 23511 21232 23520
rect 21180 23477 21189 23511
rect 21189 23477 21223 23511
rect 21223 23477 21232 23511
rect 21180 23468 21232 23477
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 4160 23264 4212 23316
rect 5816 23307 5868 23316
rect 5816 23273 5825 23307
rect 5825 23273 5859 23307
rect 5859 23273 5868 23307
rect 5816 23264 5868 23273
rect 6460 23307 6512 23316
rect 6460 23273 6469 23307
rect 6469 23273 6503 23307
rect 6503 23273 6512 23307
rect 6460 23264 6512 23273
rect 7840 23264 7892 23316
rect 8300 23264 8352 23316
rect 10140 23264 10192 23316
rect 10968 23264 11020 23316
rect 13268 23264 13320 23316
rect 17868 23264 17920 23316
rect 20076 23264 20128 23316
rect 2596 23196 2648 23248
rect 4988 23196 5040 23248
rect 5448 23196 5500 23248
rect 11428 23196 11480 23248
rect 16396 23196 16448 23248
rect 22008 23196 22060 23248
rect 2412 23128 2464 23180
rect 3884 23171 3936 23180
rect 3884 23137 3893 23171
rect 3893 23137 3927 23171
rect 3927 23137 3936 23171
rect 4436 23171 4488 23180
rect 3884 23128 3936 23137
rect 4436 23137 4445 23171
rect 4445 23137 4479 23171
rect 4479 23137 4488 23171
rect 4436 23128 4488 23137
rect 6276 23128 6328 23180
rect 12440 23128 12492 23180
rect 14556 23128 14608 23180
rect 16028 23128 16080 23180
rect 16580 23171 16632 23180
rect 16580 23137 16589 23171
rect 16589 23137 16623 23171
rect 16623 23137 16632 23171
rect 17684 23171 17736 23180
rect 16580 23128 16632 23137
rect 17684 23137 17693 23171
rect 17693 23137 17727 23171
rect 17727 23137 17736 23171
rect 17684 23128 17736 23137
rect 19432 23171 19484 23180
rect 19432 23137 19441 23171
rect 19441 23137 19475 23171
rect 19475 23137 19484 23171
rect 19432 23128 19484 23137
rect 20812 23128 20864 23180
rect 2780 23060 2832 23112
rect 7012 23103 7064 23112
rect 7012 23069 7021 23103
rect 7021 23069 7055 23103
rect 7055 23069 7064 23103
rect 7012 23060 7064 23069
rect 10692 23060 10744 23112
rect 13728 23103 13780 23112
rect 13728 23069 13737 23103
rect 13737 23069 13771 23103
rect 13771 23069 13780 23103
rect 13728 23060 13780 23069
rect 3240 22992 3292 23044
rect 13636 22992 13688 23044
rect 17776 22992 17828 23044
rect 3056 22967 3108 22976
rect 3056 22933 3065 22967
rect 3065 22933 3099 22967
rect 3099 22933 3108 22967
rect 3056 22924 3108 22933
rect 3516 22967 3568 22976
rect 3516 22933 3525 22967
rect 3525 22933 3559 22967
rect 3559 22933 3568 22967
rect 3516 22924 3568 22933
rect 7288 22924 7340 22976
rect 10968 22924 11020 22976
rect 12900 22924 12952 22976
rect 14096 22924 14148 22976
rect 14556 22924 14608 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 4988 22763 5040 22772
rect 4988 22729 4997 22763
rect 4997 22729 5031 22763
rect 5031 22729 5040 22763
rect 4988 22720 5040 22729
rect 5540 22720 5592 22772
rect 6276 22763 6328 22772
rect 6276 22729 6285 22763
rect 6285 22729 6319 22763
rect 6319 22729 6328 22763
rect 6276 22720 6328 22729
rect 6828 22720 6880 22772
rect 8208 22720 8260 22772
rect 11428 22763 11480 22772
rect 11428 22729 11437 22763
rect 11437 22729 11471 22763
rect 11471 22729 11480 22763
rect 11428 22720 11480 22729
rect 13268 22763 13320 22772
rect 13268 22729 13277 22763
rect 13277 22729 13311 22763
rect 13311 22729 13320 22763
rect 13268 22720 13320 22729
rect 13636 22763 13688 22772
rect 13636 22729 13645 22763
rect 13645 22729 13679 22763
rect 13679 22729 13688 22763
rect 13636 22720 13688 22729
rect 15476 22763 15528 22772
rect 15476 22729 15485 22763
rect 15485 22729 15519 22763
rect 15519 22729 15528 22763
rect 15476 22720 15528 22729
rect 9956 22652 10008 22704
rect 2688 22584 2740 22636
rect 7380 22627 7432 22636
rect 7380 22593 7389 22627
rect 7389 22593 7423 22627
rect 7423 22593 7432 22627
rect 7380 22584 7432 22593
rect 8852 22627 8904 22636
rect 8852 22593 8861 22627
rect 8861 22593 8895 22627
rect 8895 22593 8904 22627
rect 8852 22584 8904 22593
rect 8944 22627 8996 22636
rect 8944 22593 8953 22627
rect 8953 22593 8987 22627
rect 8987 22593 8996 22627
rect 8944 22584 8996 22593
rect 10784 22627 10836 22636
rect 10784 22593 10793 22627
rect 10793 22593 10827 22627
rect 10827 22593 10836 22627
rect 10784 22584 10836 22593
rect 10968 22627 11020 22636
rect 10968 22593 10977 22627
rect 10977 22593 11011 22627
rect 11011 22593 11020 22627
rect 10968 22584 11020 22593
rect 12716 22627 12768 22636
rect 12716 22593 12725 22627
rect 12725 22593 12759 22627
rect 12759 22593 12768 22627
rect 12716 22584 12768 22593
rect 3240 22559 3292 22568
rect 3240 22525 3274 22559
rect 3274 22525 3292 22559
rect 2688 22448 2740 22500
rect 3240 22516 3292 22525
rect 3884 22448 3936 22500
rect 6828 22516 6880 22568
rect 7288 22559 7340 22568
rect 7288 22525 7297 22559
rect 7297 22525 7331 22559
rect 7331 22525 7340 22559
rect 7288 22516 7340 22525
rect 12900 22516 12952 22568
rect 14556 22448 14608 22500
rect 2412 22423 2464 22432
rect 2412 22389 2421 22423
rect 2421 22389 2455 22423
rect 2455 22389 2464 22423
rect 2412 22380 2464 22389
rect 4252 22380 4304 22432
rect 5264 22423 5316 22432
rect 5264 22389 5273 22423
rect 5273 22389 5307 22423
rect 5307 22389 5316 22423
rect 5264 22380 5316 22389
rect 6828 22423 6880 22432
rect 6828 22389 6837 22423
rect 6837 22389 6871 22423
rect 6871 22389 6880 22423
rect 6828 22380 6880 22389
rect 8760 22423 8812 22432
rect 8760 22389 8769 22423
rect 8769 22389 8803 22423
rect 8803 22389 8812 22423
rect 8760 22380 8812 22389
rect 9680 22380 9732 22432
rect 14096 22380 14148 22432
rect 16028 22423 16080 22432
rect 16028 22389 16037 22423
rect 16037 22389 16071 22423
rect 16071 22389 16080 22423
rect 16028 22380 16080 22389
rect 16580 22423 16632 22432
rect 16580 22389 16589 22423
rect 16589 22389 16623 22423
rect 16623 22389 16632 22423
rect 16580 22380 16632 22389
rect 16856 22380 16908 22432
rect 17684 22423 17736 22432
rect 17684 22389 17693 22423
rect 17693 22389 17727 22423
rect 17727 22389 17736 22423
rect 17684 22380 17736 22389
rect 19432 22423 19484 22432
rect 19432 22389 19441 22423
rect 19441 22389 19475 22423
rect 19475 22389 19484 22423
rect 19432 22380 19484 22389
rect 20812 22380 20864 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 2688 22176 2740 22228
rect 3516 22176 3568 22228
rect 2044 22083 2096 22092
rect 2044 22049 2053 22083
rect 2053 22049 2087 22083
rect 2087 22049 2096 22083
rect 2044 22040 2096 22049
rect 2688 22040 2740 22092
rect 8300 22176 8352 22228
rect 8944 22176 8996 22228
rect 13728 22176 13780 22228
rect 5448 22108 5500 22160
rect 10968 22108 11020 22160
rect 11520 22108 11572 22160
rect 5264 22040 5316 22092
rect 6000 22040 6052 22092
rect 7380 22083 7432 22092
rect 7380 22049 7414 22083
rect 7414 22049 7432 22083
rect 7380 22040 7432 22049
rect 9772 22040 9824 22092
rect 10692 22040 10744 22092
rect 12348 22040 12400 22092
rect 14004 22040 14056 22092
rect 15568 22083 15620 22092
rect 2320 21972 2372 22024
rect 3332 21972 3384 22024
rect 4804 22015 4856 22024
rect 4804 21981 4813 22015
rect 4813 21981 4847 22015
rect 4847 21981 4856 22015
rect 4804 21972 4856 21981
rect 4988 22015 5040 22024
rect 4988 21981 4997 22015
rect 4997 21981 5031 22015
rect 5031 21981 5040 22015
rect 4988 21972 5040 21981
rect 5540 21972 5592 22024
rect 7104 22015 7156 22024
rect 7104 21981 7113 22015
rect 7113 21981 7147 22015
rect 7147 21981 7156 22015
rect 7104 21972 7156 21981
rect 10968 22015 11020 22024
rect 1584 21947 1636 21956
rect 1584 21913 1593 21947
rect 1593 21913 1627 21947
rect 1627 21913 1636 21947
rect 1584 21904 1636 21913
rect 4160 21904 4212 21956
rect 6092 21947 6144 21956
rect 6092 21913 6101 21947
rect 6101 21913 6135 21947
rect 6135 21913 6144 21947
rect 6092 21904 6144 21913
rect 9680 21904 9732 21956
rect 10968 21981 10977 22015
rect 10977 21981 11011 22015
rect 11011 21981 11020 22015
rect 10968 21972 11020 21981
rect 13360 21972 13412 22024
rect 13912 22015 13964 22024
rect 13912 21981 13921 22015
rect 13921 21981 13955 22015
rect 13955 21981 13964 22015
rect 13912 21972 13964 21981
rect 14096 22015 14148 22024
rect 14096 21981 14105 22015
rect 14105 21981 14139 22015
rect 14139 21981 14148 22015
rect 14096 21972 14148 21981
rect 15568 22049 15577 22083
rect 15577 22049 15611 22083
rect 15611 22049 15620 22083
rect 15568 22040 15620 22049
rect 15660 21972 15712 22024
rect 2872 21836 2924 21888
rect 3148 21836 3200 21888
rect 5264 21836 5316 21888
rect 9036 21879 9088 21888
rect 9036 21845 9045 21879
rect 9045 21845 9079 21879
rect 9079 21845 9088 21879
rect 9036 21836 9088 21845
rect 9496 21879 9548 21888
rect 9496 21845 9505 21879
rect 9505 21845 9539 21879
rect 9539 21845 9548 21879
rect 9496 21836 9548 21845
rect 11152 21836 11204 21888
rect 13084 21836 13136 21888
rect 14740 21836 14792 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 2320 21675 2372 21684
rect 2320 21641 2329 21675
rect 2329 21641 2363 21675
rect 2363 21641 2372 21675
rect 2320 21632 2372 21641
rect 2780 21675 2832 21684
rect 2780 21641 2789 21675
rect 2789 21641 2823 21675
rect 2823 21641 2832 21675
rect 2780 21632 2832 21641
rect 3148 21632 3200 21684
rect 4804 21632 4856 21684
rect 5448 21675 5500 21684
rect 5448 21641 5457 21675
rect 5457 21641 5491 21675
rect 5491 21641 5500 21675
rect 5448 21632 5500 21641
rect 5540 21632 5592 21684
rect 7288 21632 7340 21684
rect 9772 21632 9824 21684
rect 11520 21675 11572 21684
rect 11520 21641 11529 21675
rect 11529 21641 11563 21675
rect 11563 21641 11572 21675
rect 11520 21632 11572 21641
rect 12348 21632 12400 21684
rect 13912 21675 13964 21684
rect 13912 21641 13921 21675
rect 13921 21641 13955 21675
rect 13955 21641 13964 21675
rect 13912 21632 13964 21641
rect 14096 21632 14148 21684
rect 3424 21564 3476 21616
rect 3332 21539 3384 21548
rect 3332 21505 3341 21539
rect 3341 21505 3375 21539
rect 3375 21505 3384 21539
rect 3332 21496 3384 21505
rect 4160 21496 4212 21548
rect 4896 21539 4948 21548
rect 4896 21505 4905 21539
rect 4905 21505 4939 21539
rect 4939 21505 4948 21539
rect 4896 21496 4948 21505
rect 8024 21496 8076 21548
rect 9128 21496 9180 21548
rect 9588 21496 9640 21548
rect 10876 21496 10928 21548
rect 11152 21539 11204 21548
rect 11152 21505 11161 21539
rect 11161 21505 11195 21539
rect 11195 21505 11204 21539
rect 11152 21496 11204 21505
rect 2044 21428 2096 21480
rect 5080 21428 5132 21480
rect 6460 21471 6512 21480
rect 6460 21437 6469 21471
rect 6469 21437 6503 21471
rect 6503 21437 6512 21471
rect 6460 21428 6512 21437
rect 1768 21403 1820 21412
rect 1768 21369 1777 21403
rect 1777 21369 1811 21403
rect 1811 21369 1820 21403
rect 1768 21360 1820 21369
rect 3148 21403 3200 21412
rect 3148 21369 3157 21403
rect 3157 21369 3191 21403
rect 3191 21369 3200 21403
rect 3148 21360 3200 21369
rect 7380 21360 7432 21412
rect 13084 21471 13136 21480
rect 13084 21437 13093 21471
rect 13093 21437 13127 21471
rect 13127 21437 13136 21471
rect 13084 21428 13136 21437
rect 14556 21471 14608 21480
rect 14556 21437 14565 21471
rect 14565 21437 14599 21471
rect 14599 21437 14608 21471
rect 14556 21428 14608 21437
rect 12808 21360 12860 21412
rect 14740 21360 14792 21412
rect 5816 21335 5868 21344
rect 5816 21301 5825 21335
rect 5825 21301 5859 21335
rect 5859 21301 5868 21335
rect 5816 21292 5868 21301
rect 7104 21292 7156 21344
rect 8024 21335 8076 21344
rect 8024 21301 8033 21335
rect 8033 21301 8067 21335
rect 8067 21301 8076 21335
rect 8024 21292 8076 21301
rect 8484 21292 8536 21344
rect 10692 21292 10744 21344
rect 10876 21335 10928 21344
rect 10876 21301 10885 21335
rect 10885 21301 10919 21335
rect 10919 21301 10928 21335
rect 10876 21292 10928 21301
rect 12164 21292 12216 21344
rect 13912 21292 13964 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 2688 21088 2740 21140
rect 3424 21131 3476 21140
rect 3424 21097 3433 21131
rect 3433 21097 3467 21131
rect 3467 21097 3476 21131
rect 3424 21088 3476 21097
rect 4160 21088 4212 21140
rect 6000 21131 6052 21140
rect 6000 21097 6009 21131
rect 6009 21097 6043 21131
rect 6043 21097 6052 21131
rect 6000 21088 6052 21097
rect 8484 21131 8536 21140
rect 8484 21097 8493 21131
rect 8493 21097 8527 21131
rect 8527 21097 8536 21131
rect 8484 21088 8536 21097
rect 13084 21088 13136 21140
rect 16304 21131 16356 21140
rect 16304 21097 16313 21131
rect 16313 21097 16347 21131
rect 16347 21097 16356 21131
rect 16304 21088 16356 21097
rect 2596 21020 2648 21072
rect 3792 21063 3844 21072
rect 3792 21029 3801 21063
rect 3801 21029 3835 21063
rect 3835 21029 3844 21063
rect 3792 21020 3844 21029
rect 4252 21020 4304 21072
rect 4896 21020 4948 21072
rect 11152 21020 11204 21072
rect 1492 20995 1544 21004
rect 1492 20961 1501 20995
rect 1501 20961 1535 20995
rect 1535 20961 1544 20995
rect 1492 20952 1544 20961
rect 3884 20952 3936 21004
rect 7012 20995 7064 21004
rect 7012 20961 7021 20995
rect 7021 20961 7055 20995
rect 7055 20961 7064 20995
rect 7012 20952 7064 20961
rect 7380 20995 7432 21004
rect 7380 20961 7414 20995
rect 7414 20961 7432 20995
rect 7380 20952 7432 20961
rect 9956 20952 10008 21004
rect 10968 20995 11020 21004
rect 10968 20961 10977 20995
rect 10977 20961 11011 20995
rect 11011 20961 11020 20995
rect 10968 20952 11020 20961
rect 14280 20952 14332 21004
rect 3332 20884 3384 20936
rect 3976 20884 4028 20936
rect 7104 20927 7156 20936
rect 7104 20893 7113 20927
rect 7113 20893 7147 20927
rect 7147 20893 7156 20927
rect 7104 20884 7156 20893
rect 9864 20927 9916 20936
rect 9864 20893 9873 20927
rect 9873 20893 9907 20927
rect 9907 20893 9916 20927
rect 9864 20884 9916 20893
rect 13820 20884 13872 20936
rect 14740 20884 14792 20936
rect 5540 20816 5592 20868
rect 6460 20816 6512 20868
rect 2964 20791 3016 20800
rect 2964 20757 2973 20791
rect 2973 20757 3007 20791
rect 3007 20757 3016 20791
rect 2964 20748 3016 20757
rect 7748 20748 7800 20800
rect 9036 20748 9088 20800
rect 9588 20748 9640 20800
rect 10600 20791 10652 20800
rect 10600 20757 10609 20791
rect 10609 20757 10643 20791
rect 10643 20757 10652 20791
rect 10600 20748 10652 20757
rect 10876 20748 10928 20800
rect 10968 20748 11020 20800
rect 13176 20791 13228 20800
rect 13176 20757 13185 20791
rect 13185 20757 13219 20791
rect 13219 20757 13228 20791
rect 13176 20748 13228 20757
rect 14556 20748 14608 20800
rect 14832 20748 14884 20800
rect 15660 20748 15712 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1492 20544 1544 20596
rect 2044 20544 2096 20596
rect 3792 20587 3844 20596
rect 3792 20553 3801 20587
rect 3801 20553 3835 20587
rect 3835 20553 3844 20587
rect 3792 20544 3844 20553
rect 4160 20587 4212 20596
rect 4160 20553 4169 20587
rect 4169 20553 4203 20587
rect 4203 20553 4212 20587
rect 4160 20544 4212 20553
rect 7380 20544 7432 20596
rect 9128 20587 9180 20596
rect 9128 20553 9137 20587
rect 9137 20553 9171 20587
rect 9171 20553 9180 20587
rect 9128 20544 9180 20553
rect 9956 20544 10008 20596
rect 11152 20544 11204 20596
rect 13728 20544 13780 20596
rect 14280 20587 14332 20596
rect 14280 20553 14289 20587
rect 14289 20553 14323 20587
rect 14323 20553 14332 20587
rect 14280 20544 14332 20553
rect 14740 20544 14792 20596
rect 2504 20408 2556 20460
rect 3424 20408 3476 20460
rect 7748 20451 7800 20460
rect 2320 20340 2372 20392
rect 7748 20417 7757 20451
rect 7757 20417 7791 20451
rect 7791 20417 7800 20451
rect 7748 20408 7800 20417
rect 10692 20451 10744 20460
rect 10692 20417 10701 20451
rect 10701 20417 10735 20451
rect 10735 20417 10744 20451
rect 10692 20408 10744 20417
rect 10968 20408 11020 20460
rect 13636 20451 13688 20460
rect 13636 20417 13645 20451
rect 13645 20417 13679 20451
rect 13679 20417 13688 20451
rect 13636 20408 13688 20417
rect 2688 20272 2740 20324
rect 2780 20272 2832 20324
rect 3700 20272 3752 20324
rect 4620 20272 4672 20324
rect 5264 20272 5316 20324
rect 6184 20315 6236 20324
rect 6184 20281 6193 20315
rect 6193 20281 6227 20315
rect 6227 20281 6236 20315
rect 6184 20272 6236 20281
rect 8208 20272 8260 20324
rect 10140 20315 10192 20324
rect 10140 20281 10149 20315
rect 10149 20281 10183 20315
rect 10183 20281 10192 20315
rect 14832 20340 14884 20392
rect 15292 20340 15344 20392
rect 10140 20272 10192 20281
rect 15016 20315 15068 20324
rect 15016 20281 15050 20315
rect 15050 20281 15068 20315
rect 15016 20272 15068 20281
rect 3148 20247 3200 20256
rect 3148 20213 3157 20247
rect 3157 20213 3191 20247
rect 3191 20213 3200 20247
rect 3148 20204 3200 20213
rect 5356 20204 5408 20256
rect 7012 20204 7064 20256
rect 7748 20204 7800 20256
rect 9680 20204 9732 20256
rect 13176 20204 13228 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 3332 20043 3384 20052
rect 3332 20009 3341 20043
rect 3341 20009 3375 20043
rect 3375 20009 3384 20043
rect 3332 20000 3384 20009
rect 3516 20000 3568 20052
rect 6184 20000 6236 20052
rect 8484 20043 8536 20052
rect 2412 19932 2464 19984
rect 8484 20009 8493 20043
rect 8493 20009 8527 20043
rect 8527 20009 8536 20043
rect 8484 20000 8536 20009
rect 9772 20000 9824 20052
rect 14740 20000 14792 20052
rect 16672 20043 16724 20052
rect 16672 20009 16681 20043
rect 16681 20009 16715 20043
rect 16715 20009 16724 20043
rect 16672 20000 16724 20009
rect 9404 19975 9456 19984
rect 9404 19941 9413 19975
rect 9413 19941 9447 19975
rect 9447 19941 9456 19975
rect 9404 19932 9456 19941
rect 10968 19932 11020 19984
rect 1492 19907 1544 19916
rect 1492 19873 1501 19907
rect 1501 19873 1535 19907
rect 1535 19873 1544 19907
rect 1492 19864 1544 19873
rect 3332 19864 3384 19916
rect 5356 19907 5408 19916
rect 5356 19873 5390 19907
rect 5390 19873 5408 19907
rect 5356 19864 5408 19873
rect 7932 19907 7984 19916
rect 7932 19873 7941 19907
rect 7941 19873 7975 19907
rect 7975 19873 7984 19907
rect 7932 19864 7984 19873
rect 8576 19864 8628 19916
rect 12440 19864 12492 19916
rect 15568 19907 15620 19916
rect 4620 19796 4672 19848
rect 3148 19728 3200 19780
rect 9680 19796 9732 19848
rect 12532 19796 12584 19848
rect 13544 19839 13596 19848
rect 13544 19805 13553 19839
rect 13553 19805 13587 19839
rect 13587 19805 13596 19839
rect 15568 19873 15591 19907
rect 15591 19873 15620 19907
rect 15568 19864 15620 19873
rect 15292 19839 15344 19848
rect 13544 19796 13596 19805
rect 15292 19805 15301 19839
rect 15301 19805 15335 19839
rect 15335 19805 15344 19839
rect 15292 19796 15344 19805
rect 8944 19728 8996 19780
rect 2320 19703 2372 19712
rect 2320 19669 2329 19703
rect 2329 19669 2363 19703
rect 2363 19669 2372 19703
rect 2320 19660 2372 19669
rect 2872 19660 2924 19712
rect 4068 19660 4120 19712
rect 4896 19660 4948 19712
rect 5448 19660 5500 19712
rect 6276 19660 6328 19712
rect 7748 19703 7800 19712
rect 7748 19669 7757 19703
rect 7757 19669 7791 19703
rect 7791 19669 7800 19703
rect 7748 19660 7800 19669
rect 8024 19703 8076 19712
rect 8024 19669 8033 19703
rect 8033 19669 8067 19703
rect 8067 19669 8076 19703
rect 8024 19660 8076 19669
rect 8760 19660 8812 19712
rect 12440 19660 12492 19712
rect 12900 19703 12952 19712
rect 12900 19669 12909 19703
rect 12909 19669 12943 19703
rect 12943 19669 12952 19703
rect 12900 19660 12952 19669
rect 14372 19660 14424 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 8392 19456 8444 19508
rect 10968 19499 11020 19508
rect 10968 19465 10977 19499
rect 10977 19465 11011 19499
rect 11011 19465 11020 19499
rect 10968 19456 11020 19465
rect 12532 19499 12584 19508
rect 12532 19465 12541 19499
rect 12541 19465 12575 19499
rect 12575 19465 12584 19499
rect 12532 19456 12584 19465
rect 13544 19499 13596 19508
rect 13544 19465 13553 19499
rect 13553 19465 13587 19499
rect 13587 19465 13596 19499
rect 13544 19456 13596 19465
rect 15292 19456 15344 19508
rect 15568 19456 15620 19508
rect 3148 19320 3200 19372
rect 2136 19252 2188 19304
rect 5356 19320 5408 19372
rect 9404 19320 9456 19372
rect 2320 19227 2372 19236
rect 2320 19193 2332 19227
rect 2332 19193 2372 19227
rect 2320 19184 2372 19193
rect 2780 19184 2832 19236
rect 4712 19252 4764 19304
rect 4896 19295 4948 19304
rect 4896 19261 4905 19295
rect 4905 19261 4939 19295
rect 4939 19261 4948 19295
rect 4896 19252 4948 19261
rect 4988 19252 5040 19304
rect 8116 19252 8168 19304
rect 10140 19320 10192 19372
rect 12440 19320 12492 19372
rect 14372 19363 14424 19372
rect 11336 19252 11388 19304
rect 11980 19252 12032 19304
rect 12716 19252 12768 19304
rect 14372 19329 14381 19363
rect 14381 19329 14415 19363
rect 14415 19329 14424 19363
rect 14372 19320 14424 19329
rect 7472 19227 7524 19236
rect 4528 19116 4580 19168
rect 4620 19116 4672 19168
rect 5264 19116 5316 19168
rect 7472 19193 7481 19227
rect 7481 19193 7515 19227
rect 7515 19193 7524 19227
rect 7472 19184 7524 19193
rect 7748 19184 7800 19236
rect 8944 19184 8996 19236
rect 12532 19184 12584 19236
rect 14740 19184 14792 19236
rect 6368 19159 6420 19168
rect 6368 19125 6377 19159
rect 6377 19125 6411 19159
rect 6411 19125 6420 19159
rect 6368 19116 6420 19125
rect 7012 19159 7064 19168
rect 7012 19125 7021 19159
rect 7021 19125 7055 19159
rect 7055 19125 7064 19159
rect 7012 19116 7064 19125
rect 8392 19116 8444 19168
rect 9772 19116 9824 19168
rect 12164 19116 12216 19168
rect 12992 19159 13044 19168
rect 12992 19125 13001 19159
rect 13001 19125 13035 19159
rect 13035 19125 13044 19159
rect 12992 19116 13044 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1492 18912 1544 18964
rect 2044 18955 2096 18964
rect 2044 18921 2053 18955
rect 2053 18921 2087 18955
rect 2087 18921 2096 18955
rect 2044 18912 2096 18921
rect 4068 18912 4120 18964
rect 5356 18912 5408 18964
rect 6368 18912 6420 18964
rect 7748 18955 7800 18964
rect 7748 18921 7757 18955
rect 7757 18921 7791 18955
rect 7791 18921 7800 18955
rect 7748 18912 7800 18921
rect 8024 18912 8076 18964
rect 8944 18955 8996 18964
rect 8944 18921 8953 18955
rect 8953 18921 8987 18955
rect 8987 18921 8996 18955
rect 8944 18912 8996 18921
rect 11336 18955 11388 18964
rect 11336 18921 11345 18955
rect 11345 18921 11379 18955
rect 11379 18921 11388 18955
rect 11336 18912 11388 18921
rect 12348 18912 12400 18964
rect 12992 18955 13044 18964
rect 12992 18921 13001 18955
rect 13001 18921 13035 18955
rect 13035 18921 13044 18955
rect 12992 18912 13044 18921
rect 13452 18955 13504 18964
rect 13452 18921 13461 18955
rect 13461 18921 13495 18955
rect 13495 18921 13504 18955
rect 13452 18912 13504 18921
rect 15568 18955 15620 18964
rect 15568 18921 15577 18955
rect 15577 18921 15611 18955
rect 15611 18921 15620 18955
rect 15568 18912 15620 18921
rect 2044 18776 2096 18828
rect 2228 18776 2280 18828
rect 3700 18776 3752 18828
rect 4160 18776 4212 18828
rect 4620 18776 4672 18828
rect 5448 18844 5500 18896
rect 7012 18844 7064 18896
rect 7840 18844 7892 18896
rect 6092 18776 6144 18828
rect 7380 18776 7432 18828
rect 9956 18819 10008 18828
rect 9956 18785 9965 18819
rect 9965 18785 9999 18819
rect 9999 18785 10008 18819
rect 9956 18776 10008 18785
rect 11428 18776 11480 18828
rect 11796 18819 11848 18828
rect 11796 18785 11805 18819
rect 11805 18785 11839 18819
rect 11839 18785 11848 18819
rect 11796 18776 11848 18785
rect 13268 18776 13320 18828
rect 13912 18776 13964 18828
rect 2688 18751 2740 18760
rect 2688 18717 2697 18751
rect 2697 18717 2731 18751
rect 2731 18717 2740 18751
rect 2688 18708 2740 18717
rect 2780 18708 2832 18760
rect 3608 18708 3660 18760
rect 8208 18708 8260 18760
rect 10140 18751 10192 18760
rect 10140 18717 10149 18751
rect 10149 18717 10183 18751
rect 10183 18717 10192 18751
rect 10140 18708 10192 18717
rect 11980 18751 12032 18760
rect 11980 18717 11989 18751
rect 11989 18717 12023 18751
rect 12023 18717 12032 18751
rect 11980 18708 12032 18717
rect 12440 18708 12492 18760
rect 3332 18683 3384 18692
rect 3332 18649 3341 18683
rect 3341 18649 3375 18683
rect 3375 18649 3384 18683
rect 3332 18640 3384 18649
rect 6920 18640 6972 18692
rect 2228 18615 2280 18624
rect 2228 18581 2237 18615
rect 2237 18581 2271 18615
rect 2271 18581 2280 18615
rect 2228 18572 2280 18581
rect 3700 18615 3752 18624
rect 3700 18581 3709 18615
rect 3709 18581 3743 18615
rect 3743 18581 3752 18615
rect 3700 18572 3752 18581
rect 4252 18615 4304 18624
rect 4252 18581 4261 18615
rect 4261 18581 4295 18615
rect 4295 18581 4304 18615
rect 4252 18572 4304 18581
rect 4436 18572 4488 18624
rect 5264 18572 5316 18624
rect 6644 18615 6696 18624
rect 6644 18581 6653 18615
rect 6653 18581 6687 18615
rect 6687 18581 6696 18615
rect 6644 18572 6696 18581
rect 9220 18615 9272 18624
rect 9220 18581 9229 18615
rect 9229 18581 9263 18615
rect 9263 18581 9272 18615
rect 9220 18572 9272 18581
rect 10140 18572 10192 18624
rect 12624 18572 12676 18624
rect 13636 18640 13688 18692
rect 14372 18615 14424 18624
rect 14372 18581 14381 18615
rect 14381 18581 14415 18615
rect 14415 18581 14424 18615
rect 14372 18572 14424 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 3608 18411 3660 18420
rect 3608 18377 3617 18411
rect 3617 18377 3651 18411
rect 3651 18377 3660 18411
rect 3608 18368 3660 18377
rect 4528 18411 4580 18420
rect 4528 18377 4537 18411
rect 4537 18377 4571 18411
rect 4571 18377 4580 18411
rect 4528 18368 4580 18377
rect 6552 18411 6604 18420
rect 6552 18377 6561 18411
rect 6561 18377 6595 18411
rect 6595 18377 6604 18411
rect 6552 18368 6604 18377
rect 7840 18411 7892 18420
rect 7840 18377 7849 18411
rect 7849 18377 7883 18411
rect 7883 18377 7892 18411
rect 7840 18368 7892 18377
rect 8208 18411 8260 18420
rect 8208 18377 8217 18411
rect 8217 18377 8251 18411
rect 8251 18377 8260 18411
rect 8208 18368 8260 18377
rect 9956 18368 10008 18420
rect 11428 18411 11480 18420
rect 11428 18377 11437 18411
rect 11437 18377 11471 18411
rect 11471 18377 11480 18411
rect 11428 18368 11480 18377
rect 11796 18368 11848 18420
rect 12348 18368 12400 18420
rect 13360 18368 13412 18420
rect 14740 18411 14792 18420
rect 14740 18377 14749 18411
rect 14749 18377 14783 18411
rect 14783 18377 14792 18411
rect 14740 18368 14792 18377
rect 4068 18300 4120 18352
rect 2228 18275 2280 18284
rect 2228 18241 2237 18275
rect 2237 18241 2271 18275
rect 2271 18241 2280 18275
rect 2228 18232 2280 18241
rect 4252 18275 4304 18284
rect 4252 18241 4261 18275
rect 4261 18241 4295 18275
rect 4295 18241 4304 18275
rect 4252 18232 4304 18241
rect 5172 18275 5224 18284
rect 5172 18241 5181 18275
rect 5181 18241 5215 18275
rect 5215 18241 5224 18275
rect 5172 18232 5224 18241
rect 1584 18164 1636 18216
rect 11980 18300 12032 18352
rect 7380 18275 7432 18284
rect 7380 18241 7389 18275
rect 7389 18241 7423 18275
rect 7423 18241 7432 18275
rect 7380 18232 7432 18241
rect 8484 18232 8536 18284
rect 9680 18232 9732 18284
rect 2596 18096 2648 18148
rect 9220 18164 9272 18216
rect 9772 18164 9824 18216
rect 12164 18164 12216 18216
rect 13360 18207 13412 18216
rect 7748 18096 7800 18148
rect 13360 18173 13369 18207
rect 13369 18173 13403 18207
rect 13403 18173 13412 18207
rect 13360 18164 13412 18173
rect 13636 18207 13688 18216
rect 13636 18173 13670 18207
rect 13670 18173 13688 18207
rect 13636 18164 13688 18173
rect 1400 18028 1452 18080
rect 1952 18028 2004 18080
rect 2780 18028 2832 18080
rect 4712 18071 4764 18080
rect 4712 18037 4721 18071
rect 4721 18037 4755 18071
rect 4755 18037 4764 18071
rect 4712 18028 4764 18037
rect 5080 18071 5132 18080
rect 5080 18037 5089 18071
rect 5089 18037 5123 18071
rect 5123 18037 5132 18071
rect 5080 18028 5132 18037
rect 6092 18028 6144 18080
rect 6552 18028 6604 18080
rect 7104 18028 7156 18080
rect 8392 18071 8444 18080
rect 8392 18037 8401 18071
rect 8401 18037 8435 18071
rect 8435 18037 8444 18071
rect 8392 18028 8444 18037
rect 8760 18071 8812 18080
rect 8760 18037 8769 18071
rect 8769 18037 8803 18071
rect 8803 18037 8812 18071
rect 8760 18028 8812 18037
rect 9956 18071 10008 18080
rect 9956 18037 9965 18071
rect 9965 18037 9999 18071
rect 9999 18037 10008 18071
rect 9956 18028 10008 18037
rect 10140 18028 10192 18080
rect 11704 18071 11756 18080
rect 11704 18037 11713 18071
rect 11713 18037 11747 18071
rect 11747 18037 11756 18071
rect 11704 18028 11756 18037
rect 12808 18028 12860 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 2320 17867 2372 17876
rect 2320 17833 2329 17867
rect 2329 17833 2363 17867
rect 2363 17833 2372 17867
rect 2320 17824 2372 17833
rect 2688 17824 2740 17876
rect 3700 17824 3752 17876
rect 5172 17867 5224 17876
rect 5172 17833 5181 17867
rect 5181 17833 5215 17867
rect 5215 17833 5224 17867
rect 5172 17824 5224 17833
rect 8024 17824 8076 17876
rect 8484 17867 8536 17876
rect 8484 17833 8493 17867
rect 8493 17833 8527 17867
rect 8527 17833 8536 17867
rect 8484 17824 8536 17833
rect 12440 17824 12492 17876
rect 2780 17799 2832 17808
rect 2780 17765 2789 17799
rect 2789 17765 2823 17799
rect 2823 17765 2832 17799
rect 2780 17756 2832 17765
rect 5540 17756 5592 17808
rect 4344 17688 4396 17740
rect 6000 17756 6052 17808
rect 6644 17756 6696 17808
rect 9864 17756 9916 17808
rect 7380 17688 7432 17740
rect 10048 17731 10100 17740
rect 10048 17697 10057 17731
rect 10057 17697 10091 17731
rect 10091 17697 10100 17731
rect 10048 17688 10100 17697
rect 11704 17756 11756 17808
rect 13360 17756 13412 17808
rect 14372 17756 14424 17808
rect 11520 17731 11572 17740
rect 11520 17697 11554 17731
rect 11554 17697 11572 17731
rect 11520 17688 11572 17697
rect 1768 17620 1820 17672
rect 1952 17620 2004 17672
rect 3056 17663 3108 17672
rect 3056 17629 3065 17663
rect 3065 17629 3099 17663
rect 3099 17629 3108 17663
rect 3056 17620 3108 17629
rect 3332 17620 3384 17672
rect 4712 17663 4764 17672
rect 4712 17629 4721 17663
rect 4721 17629 4755 17663
rect 4755 17629 4764 17663
rect 4712 17620 4764 17629
rect 5540 17663 5592 17672
rect 5540 17629 5549 17663
rect 5549 17629 5583 17663
rect 5583 17629 5592 17663
rect 5540 17620 5592 17629
rect 8576 17663 8628 17672
rect 8576 17629 8585 17663
rect 8585 17629 8619 17663
rect 8619 17629 8628 17663
rect 8576 17620 8628 17629
rect 10140 17663 10192 17672
rect 10140 17629 10149 17663
rect 10149 17629 10183 17663
rect 10183 17629 10192 17663
rect 10140 17620 10192 17629
rect 10232 17663 10284 17672
rect 10232 17629 10241 17663
rect 10241 17629 10275 17663
rect 10275 17629 10284 17663
rect 10232 17620 10284 17629
rect 2596 17552 2648 17604
rect 12624 17595 12676 17604
rect 12624 17561 12633 17595
rect 12633 17561 12667 17595
rect 12667 17561 12676 17595
rect 12624 17552 12676 17561
rect 3792 17527 3844 17536
rect 3792 17493 3801 17527
rect 3801 17493 3835 17527
rect 3835 17493 3844 17527
rect 3792 17484 3844 17493
rect 7288 17527 7340 17536
rect 7288 17493 7297 17527
rect 7297 17493 7331 17527
rect 7331 17493 7340 17527
rect 7288 17484 7340 17493
rect 9680 17527 9732 17536
rect 9680 17493 9689 17527
rect 9689 17493 9723 17527
rect 9723 17493 9732 17527
rect 9680 17484 9732 17493
rect 10876 17527 10928 17536
rect 10876 17493 10885 17527
rect 10885 17493 10919 17527
rect 10919 17493 10928 17527
rect 10876 17484 10928 17493
rect 13820 17484 13872 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 2504 17280 2556 17332
rect 3056 17280 3108 17332
rect 4712 17280 4764 17332
rect 6000 17323 6052 17332
rect 6000 17289 6009 17323
rect 6009 17289 6043 17323
rect 6043 17289 6052 17323
rect 6000 17280 6052 17289
rect 10232 17280 10284 17332
rect 11520 17280 11572 17332
rect 12164 17323 12216 17332
rect 12164 17289 12173 17323
rect 12173 17289 12207 17323
rect 12207 17289 12216 17323
rect 12164 17280 12216 17289
rect 13268 17323 13320 17332
rect 13268 17289 13277 17323
rect 13277 17289 13311 17323
rect 13311 17289 13320 17323
rect 13268 17280 13320 17289
rect 14372 17323 14424 17332
rect 14372 17289 14381 17323
rect 14381 17289 14415 17323
rect 14415 17289 14424 17323
rect 14372 17280 14424 17289
rect 1952 17212 2004 17264
rect 3240 17212 3292 17264
rect 8484 17212 8536 17264
rect 2044 17187 2096 17196
rect 2044 17153 2053 17187
rect 2053 17153 2087 17187
rect 2087 17153 2096 17187
rect 2044 17144 2096 17153
rect 2320 17144 2372 17196
rect 3424 17144 3476 17196
rect 9864 17187 9916 17196
rect 1768 17119 1820 17128
rect 1768 17085 1777 17119
rect 1777 17085 1811 17119
rect 1811 17085 1820 17119
rect 1768 17076 1820 17085
rect 4068 17119 4120 17128
rect 4068 17085 4102 17119
rect 4102 17085 4120 17119
rect 4068 17076 4120 17085
rect 7380 17119 7432 17128
rect 7380 17085 7389 17119
rect 7389 17085 7423 17119
rect 7423 17085 7432 17119
rect 7380 17076 7432 17085
rect 9864 17153 9873 17187
rect 9873 17153 9907 17187
rect 9907 17153 9916 17187
rect 9864 17144 9916 17153
rect 13820 17187 13872 17196
rect 13820 17153 13829 17187
rect 13829 17153 13863 17187
rect 13863 17153 13872 17187
rect 13820 17144 13872 17153
rect 7656 17119 7708 17128
rect 7656 17085 7690 17119
rect 7690 17085 7708 17119
rect 7656 17076 7708 17085
rect 13728 17119 13780 17128
rect 13728 17085 13737 17119
rect 13737 17085 13771 17119
rect 13771 17085 13780 17119
rect 13728 17076 13780 17085
rect 14372 17076 14424 17128
rect 2136 17008 2188 17060
rect 6736 17008 6788 17060
rect 10784 17008 10836 17060
rect 15292 17008 15344 17060
rect 1860 16983 1912 16992
rect 1860 16949 1869 16983
rect 1869 16949 1903 16983
rect 1903 16949 1912 16983
rect 1860 16940 1912 16949
rect 2780 16983 2832 16992
rect 2780 16949 2789 16983
rect 2789 16949 2823 16983
rect 2823 16949 2832 16983
rect 2780 16940 2832 16949
rect 5264 16940 5316 16992
rect 6276 16983 6328 16992
rect 6276 16949 6285 16983
rect 6285 16949 6319 16983
rect 6319 16949 6328 16983
rect 6276 16940 6328 16949
rect 12440 16940 12492 16992
rect 13176 16940 13228 16992
rect 16212 16983 16264 16992
rect 16212 16949 16221 16983
rect 16221 16949 16255 16983
rect 16255 16949 16264 16983
rect 16212 16940 16264 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1492 16736 1544 16788
rect 1860 16736 1912 16788
rect 2044 16779 2096 16788
rect 2044 16745 2053 16779
rect 2053 16745 2087 16779
rect 2087 16745 2096 16779
rect 2044 16736 2096 16745
rect 2504 16736 2556 16788
rect 3056 16736 3108 16788
rect 4068 16736 4120 16788
rect 6276 16736 6328 16788
rect 6736 16779 6788 16788
rect 6736 16745 6745 16779
rect 6745 16745 6779 16779
rect 6779 16745 6788 16779
rect 6736 16736 6788 16745
rect 8392 16736 8444 16788
rect 8576 16736 8628 16788
rect 2228 16668 2280 16720
rect 6000 16668 6052 16720
rect 6092 16668 6144 16720
rect 2412 16600 2464 16652
rect 3792 16600 3844 16652
rect 4344 16643 4396 16652
rect 4344 16609 4353 16643
rect 4353 16609 4387 16643
rect 4387 16609 4396 16643
rect 4344 16600 4396 16609
rect 5080 16643 5132 16652
rect 5080 16609 5089 16643
rect 5089 16609 5123 16643
rect 5123 16609 5132 16643
rect 5080 16600 5132 16609
rect 2596 16532 2648 16584
rect 4988 16532 5040 16584
rect 5264 16575 5316 16584
rect 5264 16541 5273 16575
rect 5273 16541 5307 16575
rect 5307 16541 5316 16575
rect 5264 16532 5316 16541
rect 3884 16464 3936 16516
rect 6460 16600 6512 16652
rect 10048 16736 10100 16788
rect 11612 16779 11664 16788
rect 7656 16643 7708 16652
rect 3516 16396 3568 16448
rect 7656 16609 7665 16643
rect 7665 16609 7699 16643
rect 7699 16609 7708 16643
rect 7656 16600 7708 16609
rect 7840 16600 7892 16652
rect 8208 16643 8260 16652
rect 8208 16609 8217 16643
rect 8217 16609 8251 16643
rect 8251 16609 8260 16643
rect 8208 16600 8260 16609
rect 8116 16532 8168 16584
rect 8760 16600 8812 16652
rect 9036 16643 9088 16652
rect 9036 16609 9045 16643
rect 9045 16609 9079 16643
rect 9079 16609 9088 16643
rect 9036 16600 9088 16609
rect 10692 16600 10744 16652
rect 9220 16575 9272 16584
rect 9220 16541 9229 16575
rect 9229 16541 9263 16575
rect 9263 16541 9272 16575
rect 9220 16532 9272 16541
rect 10784 16575 10836 16584
rect 10784 16541 10793 16575
rect 10793 16541 10827 16575
rect 10827 16541 10836 16575
rect 11612 16745 11621 16779
rect 11621 16745 11655 16779
rect 11655 16745 11664 16779
rect 11612 16736 11664 16745
rect 12256 16736 12308 16788
rect 11428 16668 11480 16720
rect 13176 16668 13228 16720
rect 14188 16711 14240 16720
rect 14188 16677 14197 16711
rect 14197 16677 14231 16711
rect 14231 16677 14240 16711
rect 14188 16668 14240 16677
rect 13912 16643 13964 16652
rect 13912 16609 13921 16643
rect 13921 16609 13955 16643
rect 13955 16609 13964 16643
rect 13912 16600 13964 16609
rect 10784 16532 10836 16541
rect 13268 16532 13320 16584
rect 11336 16464 11388 16516
rect 7196 16396 7248 16448
rect 11888 16439 11940 16448
rect 11888 16405 11897 16439
rect 11897 16405 11931 16439
rect 11931 16405 11940 16439
rect 11888 16396 11940 16405
rect 13820 16396 13872 16448
rect 14740 16439 14792 16448
rect 14740 16405 14749 16439
rect 14749 16405 14783 16439
rect 14783 16405 14792 16439
rect 14740 16396 14792 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 5172 16235 5224 16244
rect 5172 16201 5181 16235
rect 5181 16201 5215 16235
rect 5215 16201 5224 16235
rect 5172 16192 5224 16201
rect 6736 16192 6788 16244
rect 7196 16192 7248 16244
rect 10140 16192 10192 16244
rect 11428 16192 11480 16244
rect 15292 16192 15344 16244
rect 6000 16056 6052 16108
rect 11244 16099 11296 16108
rect 11244 16065 11253 16099
rect 11253 16065 11287 16099
rect 11287 16065 11296 16099
rect 11244 16056 11296 16065
rect 11612 16056 11664 16108
rect 12532 16056 12584 16108
rect 13820 16099 13872 16108
rect 13820 16065 13829 16099
rect 13829 16065 13863 16099
rect 13863 16065 13872 16099
rect 13820 16056 13872 16065
rect 16580 16099 16632 16108
rect 16580 16065 16589 16099
rect 16589 16065 16623 16099
rect 16623 16065 16632 16099
rect 16580 16056 16632 16065
rect 1400 16031 1452 16040
rect 1400 15997 1409 16031
rect 1409 15997 1443 16031
rect 1443 15997 1452 16031
rect 1400 15988 1452 15997
rect 1584 15988 1636 16040
rect 4160 15988 4212 16040
rect 5080 15988 5132 16040
rect 6276 15988 6328 16040
rect 7932 15988 7984 16040
rect 5264 15920 5316 15972
rect 8484 15920 8536 15972
rect 11520 15988 11572 16040
rect 12440 16031 12492 16040
rect 12440 15997 12449 16031
rect 12449 15997 12483 16031
rect 12483 15997 12492 16031
rect 16304 16031 16356 16040
rect 12440 15988 12492 15997
rect 16304 15997 16313 16031
rect 16313 15997 16347 16031
rect 16347 15997 16356 16031
rect 16304 15988 16356 15997
rect 2044 15895 2096 15904
rect 2044 15861 2053 15895
rect 2053 15861 2087 15895
rect 2087 15861 2096 15895
rect 2044 15852 2096 15861
rect 2596 15852 2648 15904
rect 4068 15895 4120 15904
rect 4068 15861 4077 15895
rect 4077 15861 4111 15895
rect 4111 15861 4120 15895
rect 4068 15852 4120 15861
rect 4160 15852 4212 15904
rect 8116 15852 8168 15904
rect 9312 15852 9364 15904
rect 13268 15895 13320 15904
rect 13268 15861 13277 15895
rect 13277 15861 13311 15895
rect 13311 15861 13320 15895
rect 13268 15852 13320 15861
rect 13636 15895 13688 15904
rect 13636 15861 13645 15895
rect 13645 15861 13679 15895
rect 13679 15861 13688 15895
rect 13636 15852 13688 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 3884 15691 3936 15700
rect 3884 15657 3893 15691
rect 3893 15657 3927 15691
rect 3927 15657 3936 15691
rect 3884 15648 3936 15657
rect 4252 15691 4304 15700
rect 4252 15657 4261 15691
rect 4261 15657 4295 15691
rect 4295 15657 4304 15691
rect 4252 15648 4304 15657
rect 5264 15691 5316 15700
rect 5264 15657 5273 15691
rect 5273 15657 5307 15691
rect 5307 15657 5316 15691
rect 5264 15648 5316 15657
rect 7012 15648 7064 15700
rect 8208 15648 8260 15700
rect 10968 15691 11020 15700
rect 10968 15657 10977 15691
rect 10977 15657 11011 15691
rect 11011 15657 11020 15691
rect 10968 15648 11020 15657
rect 11888 15648 11940 15700
rect 12348 15648 12400 15700
rect 13912 15648 13964 15700
rect 14740 15648 14792 15700
rect 15752 15691 15804 15700
rect 15752 15657 15761 15691
rect 15761 15657 15795 15691
rect 15795 15657 15804 15691
rect 15752 15648 15804 15657
rect 6184 15580 6236 15632
rect 7288 15580 7340 15632
rect 9220 15580 9272 15632
rect 1584 15512 1636 15564
rect 2044 15512 2096 15564
rect 3884 15512 3936 15564
rect 4160 15512 4212 15564
rect 5356 15555 5408 15564
rect 5356 15521 5365 15555
rect 5365 15521 5399 15555
rect 5399 15521 5408 15555
rect 5356 15512 5408 15521
rect 7932 15512 7984 15564
rect 8116 15555 8168 15564
rect 8116 15521 8150 15555
rect 8150 15521 8168 15555
rect 8116 15512 8168 15521
rect 9680 15555 9732 15564
rect 9680 15521 9689 15555
rect 9689 15521 9723 15555
rect 9723 15521 9732 15555
rect 9680 15512 9732 15521
rect 11336 15555 11388 15564
rect 11336 15521 11345 15555
rect 11345 15521 11379 15555
rect 11379 15521 11388 15555
rect 11336 15512 11388 15521
rect 9864 15487 9916 15496
rect 9864 15453 9873 15487
rect 9873 15453 9907 15487
rect 9907 15453 9916 15487
rect 9864 15444 9916 15453
rect 11888 15444 11940 15496
rect 13636 15580 13688 15632
rect 12624 15512 12676 15564
rect 13268 15512 13320 15564
rect 9496 15376 9548 15428
rect 10876 15419 10928 15428
rect 10876 15385 10885 15419
rect 10885 15385 10919 15419
rect 10919 15385 10928 15419
rect 10876 15376 10928 15385
rect 14372 15580 14424 15632
rect 15660 15555 15712 15564
rect 15660 15521 15669 15555
rect 15669 15521 15703 15555
rect 15703 15521 15712 15555
rect 15660 15512 15712 15521
rect 15384 15444 15436 15496
rect 16488 15444 16540 15496
rect 2596 15308 2648 15360
rect 4988 15308 5040 15360
rect 5356 15308 5408 15360
rect 5540 15308 5592 15360
rect 10692 15308 10744 15360
rect 12256 15308 12308 15360
rect 13452 15308 13504 15360
rect 15292 15351 15344 15360
rect 15292 15317 15301 15351
rect 15301 15317 15335 15351
rect 15335 15317 15344 15351
rect 15292 15308 15344 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2228 15147 2280 15156
rect 2228 15113 2237 15147
rect 2237 15113 2271 15147
rect 2271 15113 2280 15147
rect 2228 15104 2280 15113
rect 3884 15104 3936 15156
rect 4068 15147 4120 15156
rect 4068 15113 4077 15147
rect 4077 15113 4111 15147
rect 4111 15113 4120 15147
rect 4068 15104 4120 15113
rect 6184 15147 6236 15156
rect 6184 15113 6193 15147
rect 6193 15113 6227 15147
rect 6227 15113 6236 15147
rect 6184 15104 6236 15113
rect 11888 15147 11940 15156
rect 11888 15113 11897 15147
rect 11897 15113 11931 15147
rect 11931 15113 11940 15147
rect 11888 15104 11940 15113
rect 12440 15104 12492 15156
rect 2044 14968 2096 15020
rect 2964 14968 3016 15020
rect 6920 15036 6972 15088
rect 8024 15011 8076 15020
rect 2780 14832 2832 14884
rect 3056 14832 3108 14884
rect 4160 14943 4212 14952
rect 4160 14909 4169 14943
rect 4169 14909 4203 14943
rect 4203 14909 4212 14943
rect 4160 14900 4212 14909
rect 8024 14977 8033 15011
rect 8033 14977 8067 15011
rect 8067 14977 8076 15011
rect 8024 14968 8076 14977
rect 11704 14968 11756 15020
rect 11796 14968 11848 15020
rect 12992 15011 13044 15020
rect 12992 14977 13001 15011
rect 13001 14977 13035 15011
rect 13035 14977 13044 15011
rect 12992 14968 13044 14977
rect 13268 14968 13320 15020
rect 16488 15104 16540 15156
rect 14372 15011 14424 15020
rect 14372 14977 14381 15011
rect 14381 14977 14415 15011
rect 14415 14977 14424 15011
rect 14372 14968 14424 14977
rect 4252 14832 4304 14884
rect 5448 14832 5500 14884
rect 7932 14900 7984 14952
rect 11152 14943 11204 14952
rect 11152 14909 11161 14943
rect 11161 14909 11195 14943
rect 11195 14909 11204 14943
rect 11152 14900 11204 14909
rect 11520 14900 11572 14952
rect 8116 14832 8168 14884
rect 1584 14807 1636 14816
rect 1584 14773 1593 14807
rect 1593 14773 1627 14807
rect 1627 14773 1636 14807
rect 1584 14764 1636 14773
rect 2044 14807 2096 14816
rect 2044 14773 2053 14807
rect 2053 14773 2087 14807
rect 2087 14773 2096 14807
rect 2044 14764 2096 14773
rect 5540 14807 5592 14816
rect 5540 14773 5549 14807
rect 5549 14773 5583 14807
rect 5583 14773 5592 14807
rect 5540 14764 5592 14773
rect 6736 14764 6788 14816
rect 7932 14807 7984 14816
rect 7932 14773 7941 14807
rect 7941 14773 7975 14807
rect 7975 14773 7984 14807
rect 7932 14764 7984 14773
rect 10048 14832 10100 14884
rect 12716 14832 12768 14884
rect 14096 14832 14148 14884
rect 15384 14900 15436 14952
rect 10140 14764 10192 14816
rect 11060 14764 11112 14816
rect 12164 14764 12216 14816
rect 15292 14764 15344 14816
rect 15660 14764 15712 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1584 14560 1636 14612
rect 2412 14603 2464 14612
rect 2412 14569 2421 14603
rect 2421 14569 2455 14603
rect 2455 14569 2464 14603
rect 2412 14560 2464 14569
rect 2872 14603 2924 14612
rect 2872 14569 2881 14603
rect 2881 14569 2915 14603
rect 2915 14569 2924 14603
rect 2872 14560 2924 14569
rect 3240 14560 3292 14612
rect 7656 14560 7708 14612
rect 7748 14560 7800 14612
rect 9036 14603 9088 14612
rect 9036 14569 9045 14603
rect 9045 14569 9079 14603
rect 9079 14569 9088 14603
rect 9036 14560 9088 14569
rect 11796 14603 11848 14612
rect 11796 14569 11805 14603
rect 11805 14569 11839 14603
rect 11839 14569 11848 14603
rect 11796 14560 11848 14569
rect 13268 14560 13320 14612
rect 14096 14603 14148 14612
rect 14096 14569 14105 14603
rect 14105 14569 14139 14603
rect 14139 14569 14148 14603
rect 14096 14560 14148 14569
rect 14372 14560 14424 14612
rect 15752 14560 15804 14612
rect 2228 14492 2280 14544
rect 4712 14492 4764 14544
rect 5540 14492 5592 14544
rect 7104 14492 7156 14544
rect 11152 14492 11204 14544
rect 12348 14492 12400 14544
rect 16120 14535 16172 14544
rect 16120 14501 16129 14535
rect 16129 14501 16163 14535
rect 16163 14501 16172 14535
rect 16120 14492 16172 14501
rect 3240 14424 3292 14476
rect 4160 14424 4212 14476
rect 4620 14424 4672 14476
rect 9220 14424 9272 14476
rect 9956 14424 10008 14476
rect 13360 14424 13412 14476
rect 15844 14467 15896 14476
rect 15844 14433 15853 14467
rect 15853 14433 15887 14467
rect 15887 14433 15896 14467
rect 15844 14424 15896 14433
rect 2412 14356 2464 14408
rect 2872 14356 2924 14408
rect 2964 14399 3016 14408
rect 2964 14365 2973 14399
rect 2973 14365 3007 14399
rect 3007 14365 3016 14399
rect 2964 14356 3016 14365
rect 1860 14331 1912 14340
rect 1860 14297 1869 14331
rect 1869 14297 1903 14331
rect 1903 14297 1912 14331
rect 1860 14288 1912 14297
rect 3056 14288 3108 14340
rect 2596 14220 2648 14272
rect 6184 14220 6236 14272
rect 7380 14288 7432 14340
rect 7932 14356 7984 14408
rect 9036 14356 9088 14408
rect 9680 14399 9732 14408
rect 9680 14365 9689 14399
rect 9689 14365 9723 14399
rect 9723 14365 9732 14399
rect 9680 14356 9732 14365
rect 11244 14356 11296 14408
rect 10968 14288 11020 14340
rect 7196 14220 7248 14272
rect 7564 14220 7616 14272
rect 9128 14263 9180 14272
rect 9128 14229 9137 14263
rect 9137 14229 9171 14263
rect 9171 14229 9180 14263
rect 9128 14220 9180 14229
rect 10232 14220 10284 14272
rect 10692 14263 10744 14272
rect 10692 14229 10701 14263
rect 10701 14229 10735 14263
rect 10735 14229 10744 14263
rect 10692 14220 10744 14229
rect 11244 14220 11296 14272
rect 12440 14288 12492 14340
rect 14372 14220 14424 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1860 13948 1912 14000
rect 2412 13948 2464 14000
rect 2596 13880 2648 13932
rect 1584 13812 1636 13864
rect 3148 14016 3200 14068
rect 4252 14016 4304 14068
rect 4620 14059 4672 14068
rect 4620 14025 4629 14059
rect 4629 14025 4663 14059
rect 4663 14025 4672 14059
rect 4620 14016 4672 14025
rect 2964 13991 3016 14000
rect 2964 13957 2973 13991
rect 2973 13957 3007 13991
rect 3007 13957 3016 13991
rect 2964 13948 3016 13957
rect 4528 13991 4580 14000
rect 4528 13957 4537 13991
rect 4537 13957 4571 13991
rect 4571 13957 4580 13991
rect 4528 13948 4580 13957
rect 3608 13880 3660 13932
rect 4068 13880 4120 13932
rect 2780 13812 2832 13864
rect 3792 13812 3844 13864
rect 4896 13812 4948 13864
rect 5540 13880 5592 13932
rect 8852 14016 8904 14068
rect 9956 14059 10008 14068
rect 9956 14025 9965 14059
rect 9965 14025 9999 14059
rect 9999 14025 10008 14059
rect 9956 14016 10008 14025
rect 10232 14059 10284 14068
rect 10232 14025 10241 14059
rect 10241 14025 10275 14059
rect 10275 14025 10284 14059
rect 10232 14016 10284 14025
rect 10876 14016 10928 14068
rect 11336 14016 11388 14068
rect 6920 13948 6972 14000
rect 7104 13948 7156 14000
rect 7840 13991 7892 14000
rect 7840 13957 7849 13991
rect 7849 13957 7883 13991
rect 7883 13957 7892 13991
rect 7840 13948 7892 13957
rect 9864 13948 9916 14000
rect 5356 13744 5408 13796
rect 7380 13880 7432 13932
rect 8852 13923 8904 13932
rect 8852 13889 8861 13923
rect 8861 13889 8895 13923
rect 8895 13889 8904 13923
rect 8852 13880 8904 13889
rect 9036 13923 9088 13932
rect 9036 13889 9045 13923
rect 9045 13889 9079 13923
rect 9079 13889 9088 13923
rect 9036 13880 9088 13889
rect 10968 13923 11020 13932
rect 10968 13889 10977 13923
rect 10977 13889 11011 13923
rect 11011 13889 11020 13923
rect 12348 14016 12400 14068
rect 14372 14059 14424 14068
rect 14372 14025 14381 14059
rect 14381 14025 14415 14059
rect 14415 14025 14424 14059
rect 14372 14016 14424 14025
rect 14464 14016 14516 14068
rect 10968 13880 11020 13889
rect 12440 13923 12492 13932
rect 12440 13889 12449 13923
rect 12449 13889 12483 13923
rect 12483 13889 12492 13923
rect 12440 13880 12492 13889
rect 7196 13855 7248 13864
rect 7196 13821 7205 13855
rect 7205 13821 7239 13855
rect 7239 13821 7248 13855
rect 7196 13812 7248 13821
rect 10692 13812 10744 13864
rect 12716 13855 12768 13864
rect 6828 13744 6880 13796
rect 3424 13719 3476 13728
rect 3424 13685 3433 13719
rect 3433 13685 3467 13719
rect 3467 13685 3476 13719
rect 3424 13676 3476 13685
rect 6000 13676 6052 13728
rect 6184 13676 6236 13728
rect 7656 13676 7708 13728
rect 11336 13744 11388 13796
rect 12716 13821 12739 13855
rect 12739 13821 12768 13855
rect 12716 13812 12768 13821
rect 14372 13812 14424 13864
rect 15200 13855 15252 13864
rect 15200 13821 15234 13855
rect 15234 13821 15252 13855
rect 15200 13812 15252 13821
rect 8392 13719 8444 13728
rect 8392 13685 8401 13719
rect 8401 13685 8435 13719
rect 8435 13685 8444 13719
rect 8392 13676 8444 13685
rect 10692 13676 10744 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1676 13472 1728 13524
rect 3608 13472 3660 13524
rect 3792 13515 3844 13524
rect 3792 13481 3801 13515
rect 3801 13481 3835 13515
rect 3835 13481 3844 13515
rect 3792 13472 3844 13481
rect 4712 13515 4764 13524
rect 4712 13481 4721 13515
rect 4721 13481 4755 13515
rect 4755 13481 4764 13515
rect 4712 13472 4764 13481
rect 5264 13515 5316 13524
rect 1768 13379 1820 13388
rect 1768 13345 1777 13379
rect 1777 13345 1811 13379
rect 1811 13345 1820 13379
rect 1768 13336 1820 13345
rect 5264 13481 5273 13515
rect 5273 13481 5307 13515
rect 5307 13481 5316 13515
rect 5264 13472 5316 13481
rect 6000 13472 6052 13524
rect 6828 13515 6880 13524
rect 6828 13481 6837 13515
rect 6837 13481 6871 13515
rect 6871 13481 6880 13515
rect 6828 13472 6880 13481
rect 7012 13515 7064 13524
rect 7012 13481 7021 13515
rect 7021 13481 7055 13515
rect 7055 13481 7064 13515
rect 7472 13515 7524 13524
rect 7012 13472 7064 13481
rect 7472 13481 7481 13515
rect 7481 13481 7515 13515
rect 7515 13481 7524 13515
rect 7472 13472 7524 13481
rect 7748 13472 7800 13524
rect 8852 13472 8904 13524
rect 8944 13472 8996 13524
rect 9404 13515 9456 13524
rect 9404 13481 9413 13515
rect 9413 13481 9447 13515
rect 9447 13481 9456 13515
rect 9404 13472 9456 13481
rect 9680 13472 9732 13524
rect 12716 13472 12768 13524
rect 13360 13515 13412 13524
rect 13360 13481 13369 13515
rect 13369 13481 13403 13515
rect 13403 13481 13412 13515
rect 13360 13472 13412 13481
rect 13452 13472 13504 13524
rect 15200 13472 15252 13524
rect 15844 13515 15896 13524
rect 15844 13481 15853 13515
rect 15853 13481 15887 13515
rect 15887 13481 15896 13515
rect 15844 13472 15896 13481
rect 5540 13404 5592 13456
rect 2044 13311 2096 13320
rect 2044 13277 2053 13311
rect 2053 13277 2087 13311
rect 2087 13277 2096 13311
rect 2044 13268 2096 13277
rect 4160 13268 4212 13320
rect 5448 13311 5500 13320
rect 5448 13277 5457 13311
rect 5457 13277 5491 13311
rect 5491 13277 5500 13311
rect 5448 13268 5500 13277
rect 6552 13379 6604 13388
rect 6552 13345 6561 13379
rect 6561 13345 6595 13379
rect 6595 13345 6604 13379
rect 6552 13336 6604 13345
rect 7288 13404 7340 13456
rect 14372 13404 14424 13456
rect 16856 13404 16908 13456
rect 11704 13379 11756 13388
rect 11704 13345 11738 13379
rect 11738 13345 11756 13379
rect 11704 13336 11756 13345
rect 16672 13379 16724 13388
rect 16672 13345 16681 13379
rect 16681 13345 16715 13379
rect 16715 13345 16724 13379
rect 16672 13336 16724 13345
rect 7196 13268 7248 13320
rect 7564 13311 7616 13320
rect 7564 13277 7573 13311
rect 7573 13277 7607 13311
rect 7607 13277 7616 13311
rect 7564 13268 7616 13277
rect 9312 13268 9364 13320
rect 10232 13311 10284 13320
rect 10232 13277 10241 13311
rect 10241 13277 10275 13311
rect 10275 13277 10284 13311
rect 10232 13268 10284 13277
rect 11244 13268 11296 13320
rect 4896 13200 4948 13252
rect 9772 13200 9824 13252
rect 2688 13132 2740 13184
rect 2872 13175 2924 13184
rect 2872 13141 2881 13175
rect 2881 13141 2915 13175
rect 2915 13141 2924 13175
rect 2872 13132 2924 13141
rect 6000 13132 6052 13184
rect 6368 13175 6420 13184
rect 6368 13141 6377 13175
rect 6377 13141 6411 13175
rect 6411 13141 6420 13175
rect 6368 13132 6420 13141
rect 10784 13175 10836 13184
rect 10784 13141 10793 13175
rect 10793 13141 10827 13175
rect 10827 13141 10836 13175
rect 10784 13132 10836 13141
rect 11336 13132 11388 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 3424 12971 3476 12980
rect 3424 12937 3433 12971
rect 3433 12937 3467 12971
rect 3467 12937 3476 12971
rect 3424 12928 3476 12937
rect 5264 12928 5316 12980
rect 7564 12928 7616 12980
rect 8392 12928 8444 12980
rect 9312 12971 9364 12980
rect 9312 12937 9321 12971
rect 9321 12937 9355 12971
rect 9355 12937 9364 12971
rect 9312 12928 9364 12937
rect 9680 12971 9732 12980
rect 9680 12937 9689 12971
rect 9689 12937 9723 12971
rect 9723 12937 9732 12971
rect 9680 12928 9732 12937
rect 10232 12928 10284 12980
rect 10692 12971 10744 12980
rect 10692 12937 10701 12971
rect 10701 12937 10735 12971
rect 10735 12937 10744 12971
rect 10692 12928 10744 12937
rect 10876 12928 10928 12980
rect 16672 12928 16724 12980
rect 17040 12971 17092 12980
rect 17040 12937 17049 12971
rect 17049 12937 17083 12971
rect 17083 12937 17092 12971
rect 17040 12928 17092 12937
rect 7012 12860 7064 12912
rect 7288 12860 7340 12912
rect 8668 12903 8720 12912
rect 8668 12869 8677 12903
rect 8677 12869 8711 12903
rect 8711 12869 8720 12903
rect 8668 12860 8720 12869
rect 6000 12792 6052 12844
rect 1492 12724 1544 12776
rect 2044 12724 2096 12776
rect 6828 12724 6880 12776
rect 5080 12656 5132 12708
rect 7288 12767 7340 12776
rect 7288 12733 7297 12767
rect 7297 12733 7331 12767
rect 7331 12733 7340 12767
rect 7288 12724 7340 12733
rect 7748 12656 7800 12708
rect 10784 12656 10836 12708
rect 11428 12860 11480 12912
rect 11060 12792 11112 12844
rect 11336 12835 11388 12844
rect 11336 12801 11345 12835
rect 11345 12801 11379 12835
rect 11379 12801 11388 12835
rect 11336 12792 11388 12801
rect 12440 12835 12492 12844
rect 12440 12801 12449 12835
rect 12449 12801 12483 12835
rect 12483 12801 12492 12835
rect 16212 12835 16264 12844
rect 12440 12792 12492 12801
rect 16212 12801 16221 12835
rect 16221 12801 16255 12835
rect 16255 12801 16264 12835
rect 16212 12792 16264 12801
rect 18328 12835 18380 12844
rect 18328 12801 18337 12835
rect 18337 12801 18371 12835
rect 18371 12801 18380 12835
rect 18328 12792 18380 12801
rect 15936 12767 15988 12776
rect 15936 12733 15945 12767
rect 15945 12733 15979 12767
rect 15979 12733 15988 12767
rect 15936 12724 15988 12733
rect 18052 12767 18104 12776
rect 18052 12733 18061 12767
rect 18061 12733 18095 12767
rect 18095 12733 18104 12767
rect 18052 12724 18104 12733
rect 2872 12588 2924 12640
rect 3976 12631 4028 12640
rect 3976 12597 3985 12631
rect 3985 12597 4019 12631
rect 4019 12597 4028 12631
rect 3976 12588 4028 12597
rect 5172 12631 5224 12640
rect 5172 12597 5181 12631
rect 5181 12597 5215 12631
rect 5215 12597 5224 12631
rect 5172 12588 5224 12597
rect 7472 12588 7524 12640
rect 11796 12631 11848 12640
rect 11796 12597 11805 12631
rect 11805 12597 11839 12631
rect 11839 12597 11848 12631
rect 11796 12588 11848 12597
rect 12992 12631 13044 12640
rect 12992 12597 13001 12631
rect 13001 12597 13035 12631
rect 13035 12597 13044 12631
rect 12992 12588 13044 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 2136 12384 2188 12436
rect 2412 12427 2464 12436
rect 2412 12393 2421 12427
rect 2421 12393 2455 12427
rect 2455 12393 2464 12427
rect 2412 12384 2464 12393
rect 2964 12384 3016 12436
rect 3608 12384 3660 12436
rect 4436 12384 4488 12436
rect 5632 12427 5684 12436
rect 5632 12393 5641 12427
rect 5641 12393 5675 12427
rect 5675 12393 5684 12427
rect 5632 12384 5684 12393
rect 7288 12384 7340 12436
rect 9220 12427 9272 12436
rect 9220 12393 9229 12427
rect 9229 12393 9263 12427
rect 9263 12393 9272 12427
rect 9220 12384 9272 12393
rect 11060 12427 11112 12436
rect 11060 12393 11069 12427
rect 11069 12393 11103 12427
rect 11103 12393 11112 12427
rect 11060 12384 11112 12393
rect 11612 12427 11664 12436
rect 11612 12393 11621 12427
rect 11621 12393 11655 12427
rect 11655 12393 11664 12427
rect 11612 12384 11664 12393
rect 2780 12316 2832 12368
rect 6184 12316 6236 12368
rect 6920 12316 6972 12368
rect 9956 12316 10008 12368
rect 1584 12248 1636 12300
rect 4160 12248 4212 12300
rect 4436 12291 4488 12300
rect 4436 12257 4445 12291
rect 4445 12257 4479 12291
rect 4479 12257 4488 12291
rect 4436 12248 4488 12257
rect 5724 12291 5776 12300
rect 5724 12257 5733 12291
rect 5733 12257 5767 12291
rect 5767 12257 5776 12291
rect 5724 12248 5776 12257
rect 7564 12248 7616 12300
rect 8852 12248 8904 12300
rect 11336 12316 11388 12368
rect 20996 12316 21048 12368
rect 10876 12248 10928 12300
rect 11980 12291 12032 12300
rect 11980 12257 11989 12291
rect 11989 12257 12023 12291
rect 12023 12257 12032 12291
rect 11980 12248 12032 12257
rect 20904 12291 20956 12300
rect 20904 12257 20913 12291
rect 20913 12257 20947 12291
rect 20947 12257 20956 12291
rect 20904 12248 20956 12257
rect 4620 12223 4672 12232
rect 4620 12189 4629 12223
rect 4629 12189 4663 12223
rect 4663 12189 4672 12223
rect 4620 12180 4672 12189
rect 9128 12180 9180 12232
rect 3424 12112 3476 12164
rect 4068 12155 4120 12164
rect 4068 12121 4077 12155
rect 4077 12121 4111 12155
rect 4111 12121 4120 12155
rect 4068 12112 4120 12121
rect 9588 12112 9640 12164
rect 11336 12180 11388 12232
rect 12256 12223 12308 12232
rect 12256 12189 12265 12223
rect 12265 12189 12299 12223
rect 12299 12189 12308 12223
rect 12256 12180 12308 12189
rect 1860 12044 1912 12096
rect 5264 12087 5316 12096
rect 5264 12053 5273 12087
rect 5273 12053 5307 12087
rect 5307 12053 5316 12087
rect 5264 12044 5316 12053
rect 7104 12087 7156 12096
rect 7104 12053 7113 12087
rect 7113 12053 7147 12087
rect 7147 12053 7156 12087
rect 7104 12044 7156 12053
rect 7748 12087 7800 12096
rect 7748 12053 7757 12087
rect 7757 12053 7791 12087
rect 7791 12053 7800 12087
rect 7748 12044 7800 12053
rect 9680 12087 9732 12096
rect 9680 12053 9689 12087
rect 9689 12053 9723 12087
rect 9723 12053 9732 12087
rect 9680 12044 9732 12053
rect 11060 12044 11112 12096
rect 11244 12087 11296 12096
rect 11244 12053 11253 12087
rect 11253 12053 11287 12087
rect 11287 12053 11296 12087
rect 11244 12044 11296 12053
rect 12992 12044 13044 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2136 11840 2188 11892
rect 4436 11840 4488 11892
rect 5080 11840 5132 11892
rect 6184 11883 6236 11892
rect 6184 11849 6193 11883
rect 6193 11849 6227 11883
rect 6227 11849 6236 11883
rect 6184 11840 6236 11849
rect 3884 11772 3936 11824
rect 4896 11815 4948 11824
rect 4896 11781 4905 11815
rect 4905 11781 4939 11815
rect 4939 11781 4948 11815
rect 7196 11840 7248 11892
rect 7748 11840 7800 11892
rect 8852 11883 8904 11892
rect 8852 11849 8861 11883
rect 8861 11849 8895 11883
rect 8895 11849 8904 11883
rect 8852 11840 8904 11849
rect 11336 11883 11388 11892
rect 11336 11849 11345 11883
rect 11345 11849 11379 11883
rect 11379 11849 11388 11883
rect 11336 11840 11388 11849
rect 12256 11840 12308 11892
rect 4896 11772 4948 11781
rect 7840 11772 7892 11824
rect 9128 11815 9180 11824
rect 9128 11781 9137 11815
rect 9137 11781 9171 11815
rect 9171 11781 9180 11815
rect 9128 11772 9180 11781
rect 12808 11840 12860 11892
rect 13820 11883 13872 11892
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 4160 11636 4212 11688
rect 2780 11568 2832 11620
rect 7104 11679 7156 11688
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 3516 11543 3568 11552
rect 3516 11509 3525 11543
rect 3525 11509 3559 11543
rect 3559 11509 3568 11543
rect 3516 11500 3568 11509
rect 5264 11500 5316 11552
rect 5632 11543 5684 11552
rect 5632 11509 5641 11543
rect 5641 11509 5675 11543
rect 5675 11509 5684 11543
rect 5632 11500 5684 11509
rect 6092 11568 6144 11620
rect 7104 11645 7138 11679
rect 7138 11645 7156 11679
rect 7104 11636 7156 11645
rect 9404 11636 9456 11688
rect 9588 11611 9640 11620
rect 9588 11577 9622 11611
rect 9622 11577 9640 11611
rect 9588 11568 9640 11577
rect 12256 11568 12308 11620
rect 6368 11500 6420 11552
rect 10692 11543 10744 11552
rect 10692 11509 10701 11543
rect 10701 11509 10735 11543
rect 10735 11509 10744 11543
rect 10692 11500 10744 11509
rect 11980 11500 12032 11552
rect 12348 11500 12400 11552
rect 20904 11543 20956 11552
rect 20904 11509 20913 11543
rect 20913 11509 20947 11543
rect 20947 11509 20956 11543
rect 20904 11500 20956 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1400 11339 1452 11348
rect 1400 11305 1409 11339
rect 1409 11305 1443 11339
rect 1443 11305 1452 11339
rect 1400 11296 1452 11305
rect 1860 11339 1912 11348
rect 1860 11305 1869 11339
rect 1869 11305 1903 11339
rect 1903 11305 1912 11339
rect 1860 11296 1912 11305
rect 2780 11228 2832 11280
rect 4620 11296 4672 11348
rect 6092 11339 6144 11348
rect 6092 11305 6101 11339
rect 6101 11305 6135 11339
rect 6135 11305 6144 11339
rect 6092 11296 6144 11305
rect 6368 11339 6420 11348
rect 6368 11305 6377 11339
rect 6377 11305 6411 11339
rect 6411 11305 6420 11339
rect 6368 11296 6420 11305
rect 7288 11339 7340 11348
rect 7288 11305 7297 11339
rect 7297 11305 7331 11339
rect 7331 11305 7340 11339
rect 7288 11296 7340 11305
rect 8024 11339 8076 11348
rect 8024 11305 8033 11339
rect 8033 11305 8067 11339
rect 8067 11305 8076 11339
rect 8024 11296 8076 11305
rect 8944 11296 8996 11348
rect 9680 11296 9732 11348
rect 10876 11339 10928 11348
rect 10876 11305 10885 11339
rect 10885 11305 10919 11339
rect 10919 11305 10928 11339
rect 10876 11296 10928 11305
rect 12256 11296 12308 11348
rect 12992 11339 13044 11348
rect 12992 11305 13001 11339
rect 13001 11305 13035 11339
rect 13035 11305 13044 11339
rect 12992 11296 13044 11305
rect 3516 11160 3568 11212
rect 9956 11271 10008 11280
rect 9956 11237 9965 11271
rect 9965 11237 9999 11271
rect 9999 11237 10008 11271
rect 9956 11228 10008 11237
rect 18144 11228 18196 11280
rect 4160 11160 4212 11212
rect 4896 11160 4948 11212
rect 8760 11160 8812 11212
rect 9680 11203 9732 11212
rect 9680 11169 9689 11203
rect 9689 11169 9723 11203
rect 9723 11169 9732 11203
rect 9680 11160 9732 11169
rect 9864 11160 9916 11212
rect 11060 11203 11112 11212
rect 11060 11169 11069 11203
rect 11069 11169 11103 11203
rect 11103 11169 11112 11203
rect 11060 11160 11112 11169
rect 11336 11203 11388 11212
rect 11336 11169 11370 11203
rect 11370 11169 11388 11203
rect 11336 11160 11388 11169
rect 17960 11203 18012 11212
rect 17960 11169 17969 11203
rect 17969 11169 18003 11203
rect 18003 11169 18012 11203
rect 17960 11160 18012 11169
rect 8116 11092 8168 11144
rect 9772 11092 9824 11144
rect 7564 11067 7616 11076
rect 7564 11033 7573 11067
rect 7573 11033 7607 11067
rect 7607 11033 7616 11067
rect 7564 11024 7616 11033
rect 9588 11024 9640 11076
rect 10140 11024 10192 11076
rect 3332 10956 3384 11008
rect 5448 10999 5500 11008
rect 5448 10965 5457 10999
rect 5457 10965 5491 10999
rect 5491 10965 5500 10999
rect 5448 10956 5500 10965
rect 6460 10956 6512 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 2044 10752 2096 10804
rect 3424 10752 3476 10804
rect 8116 10795 8168 10804
rect 8116 10761 8125 10795
rect 8125 10761 8159 10795
rect 8159 10761 8168 10795
rect 8116 10752 8168 10761
rect 8944 10795 8996 10804
rect 8944 10761 8953 10795
rect 8953 10761 8987 10795
rect 8987 10761 8996 10795
rect 8944 10752 8996 10761
rect 9588 10752 9640 10804
rect 12992 10752 13044 10804
rect 17960 10752 18012 10804
rect 2136 10659 2188 10668
rect 2136 10625 2145 10659
rect 2145 10625 2179 10659
rect 2179 10625 2188 10659
rect 2136 10616 2188 10625
rect 3424 10616 3476 10668
rect 4160 10616 4212 10668
rect 6460 10616 6512 10668
rect 9772 10659 9824 10668
rect 9772 10625 9781 10659
rect 9781 10625 9815 10659
rect 9815 10625 9824 10659
rect 9772 10616 9824 10625
rect 2504 10480 2556 10532
rect 3148 10480 3200 10532
rect 3516 10480 3568 10532
rect 4804 10548 4856 10600
rect 5448 10548 5500 10600
rect 6552 10548 6604 10600
rect 9680 10548 9732 10600
rect 12440 10659 12492 10668
rect 12440 10625 12449 10659
rect 12449 10625 12483 10659
rect 12483 10625 12492 10659
rect 12440 10616 12492 10625
rect 19432 10616 19484 10668
rect 19984 10659 20036 10668
rect 19984 10625 19993 10659
rect 19993 10625 20027 10659
rect 20027 10625 20036 10659
rect 19984 10616 20036 10625
rect 6736 10480 6788 10532
rect 10692 10548 10744 10600
rect 18420 10591 18472 10600
rect 18420 10557 18429 10591
rect 18429 10557 18463 10591
rect 18463 10557 18472 10591
rect 18420 10548 18472 10557
rect 19708 10591 19760 10600
rect 19708 10557 19717 10591
rect 19717 10557 19751 10591
rect 19751 10557 19760 10591
rect 19708 10548 19760 10557
rect 11060 10480 11112 10532
rect 2688 10412 2740 10464
rect 3332 10455 3384 10464
rect 3332 10421 3341 10455
rect 3341 10421 3375 10455
rect 3375 10421 3384 10455
rect 3332 10412 3384 10421
rect 6552 10455 6604 10464
rect 6552 10421 6561 10455
rect 6561 10421 6595 10455
rect 6595 10421 6604 10455
rect 6552 10412 6604 10421
rect 6828 10455 6880 10464
rect 6828 10421 6837 10455
rect 6837 10421 6871 10455
rect 6871 10421 6880 10455
rect 6828 10412 6880 10421
rect 8392 10455 8444 10464
rect 8392 10421 8401 10455
rect 8401 10421 8435 10455
rect 8435 10421 8444 10455
rect 8392 10412 8444 10421
rect 11336 10412 11388 10464
rect 11980 10412 12032 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2596 10208 2648 10260
rect 3332 10208 3384 10260
rect 3424 10251 3476 10260
rect 3424 10217 3433 10251
rect 3433 10217 3467 10251
rect 3467 10217 3476 10251
rect 3424 10208 3476 10217
rect 3884 10208 3936 10260
rect 4160 10208 4212 10260
rect 7564 10251 7616 10260
rect 2044 10140 2096 10192
rect 7564 10217 7573 10251
rect 7573 10217 7607 10251
rect 7607 10217 7616 10251
rect 7564 10208 7616 10217
rect 8208 10251 8260 10260
rect 8208 10217 8217 10251
rect 8217 10217 8251 10251
rect 8251 10217 8260 10251
rect 8208 10208 8260 10217
rect 8392 10208 8444 10260
rect 10048 10251 10100 10260
rect 10048 10217 10057 10251
rect 10057 10217 10091 10251
rect 10091 10217 10100 10251
rect 10048 10208 10100 10217
rect 11060 10251 11112 10260
rect 11060 10217 11069 10251
rect 11069 10217 11103 10251
rect 11103 10217 11112 10251
rect 11060 10208 11112 10217
rect 11244 10251 11296 10260
rect 11244 10217 11253 10251
rect 11253 10217 11287 10251
rect 11287 10217 11296 10251
rect 11244 10208 11296 10217
rect 8760 10183 8812 10192
rect 8760 10149 8769 10183
rect 8769 10149 8803 10183
rect 8803 10149 8812 10183
rect 8760 10140 8812 10149
rect 9864 10140 9916 10192
rect 21180 10140 21232 10192
rect 5264 10115 5316 10124
rect 5264 10081 5273 10115
rect 5273 10081 5307 10115
rect 5307 10081 5316 10115
rect 5264 10072 5316 10081
rect 5356 10072 5408 10124
rect 7288 10072 7340 10124
rect 7840 10072 7892 10124
rect 11244 10072 11296 10124
rect 19524 10115 19576 10124
rect 19524 10081 19533 10115
rect 19533 10081 19567 10115
rect 19567 10081 19576 10115
rect 19524 10072 19576 10081
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 4068 10047 4120 10056
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 8024 10004 8076 10056
rect 3700 9868 3752 9920
rect 7656 9936 7708 9988
rect 11704 10047 11756 10056
rect 9680 9979 9732 9988
rect 9680 9945 9689 9979
rect 9689 9945 9723 9979
rect 9723 9945 9732 9979
rect 9680 9936 9732 9945
rect 9772 9936 9824 9988
rect 11704 10013 11713 10047
rect 11713 10013 11747 10047
rect 11747 10013 11756 10047
rect 11704 10004 11756 10013
rect 11980 10004 12032 10056
rect 6460 9868 6512 9920
rect 7288 9911 7340 9920
rect 7288 9877 7297 9911
rect 7297 9877 7331 9911
rect 7331 9877 7340 9911
rect 7288 9868 7340 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 3424 9664 3476 9716
rect 3332 9596 3384 9648
rect 3700 9596 3752 9648
rect 1400 9528 1452 9580
rect 6736 9664 6788 9716
rect 8208 9707 8260 9716
rect 8208 9673 8217 9707
rect 8217 9673 8251 9707
rect 8251 9673 8260 9707
rect 8208 9664 8260 9673
rect 10048 9664 10100 9716
rect 11704 9707 11756 9716
rect 11704 9673 11713 9707
rect 11713 9673 11747 9707
rect 11747 9673 11756 9707
rect 11704 9664 11756 9673
rect 11980 9707 12032 9716
rect 11980 9673 11989 9707
rect 11989 9673 12023 9707
rect 12023 9673 12032 9707
rect 11980 9664 12032 9673
rect 19524 9707 19576 9716
rect 19524 9673 19533 9707
rect 19533 9673 19567 9707
rect 19567 9673 19576 9707
rect 19524 9664 19576 9673
rect 10692 9596 10744 9648
rect 11520 9596 11572 9648
rect 12440 9596 12492 9648
rect 15292 9596 15344 9648
rect 3884 9460 3936 9512
rect 7288 9528 7340 9580
rect 1768 9392 1820 9444
rect 2596 9392 2648 9444
rect 2504 9324 2556 9376
rect 7840 9503 7892 9512
rect 7840 9469 7849 9503
rect 7849 9469 7883 9503
rect 7883 9469 7892 9503
rect 7840 9460 7892 9469
rect 8668 9503 8720 9512
rect 8668 9469 8677 9503
rect 8677 9469 8711 9503
rect 8711 9469 8720 9503
rect 8668 9460 8720 9469
rect 9496 9460 9548 9512
rect 7012 9392 7064 9444
rect 8944 9435 8996 9444
rect 8944 9401 8978 9435
rect 8978 9401 8996 9435
rect 8944 9392 8996 9401
rect 4712 9324 4764 9376
rect 10140 9324 10192 9376
rect 11060 9324 11112 9376
rect 11244 9367 11296 9376
rect 11244 9333 11253 9367
rect 11253 9333 11287 9367
rect 11287 9333 11296 9367
rect 11244 9324 11296 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1768 9163 1820 9172
rect 1768 9129 1777 9163
rect 1777 9129 1811 9163
rect 1811 9129 1820 9163
rect 1768 9120 1820 9129
rect 2044 9163 2096 9172
rect 2044 9129 2053 9163
rect 2053 9129 2087 9163
rect 2087 9129 2096 9163
rect 2044 9120 2096 9129
rect 2780 9120 2832 9172
rect 5356 9163 5408 9172
rect 5356 9129 5365 9163
rect 5365 9129 5399 9163
rect 5399 9129 5408 9163
rect 5356 9120 5408 9129
rect 8024 9120 8076 9172
rect 8944 9120 8996 9172
rect 9588 9120 9640 9172
rect 9864 9120 9916 9172
rect 3056 9052 3108 9104
rect 4068 9052 4120 9104
rect 5264 9052 5316 9104
rect 2780 9027 2832 9036
rect 2780 8993 2789 9027
rect 2789 8993 2823 9027
rect 2823 8993 2832 9027
rect 2780 8984 2832 8993
rect 3792 8984 3844 9036
rect 7012 9052 7064 9104
rect 8668 9052 8720 9104
rect 6460 8984 6512 9036
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 3148 8916 3200 8968
rect 4712 8959 4764 8968
rect 4712 8925 4721 8959
rect 4721 8925 4755 8959
rect 4755 8925 4764 8959
rect 4712 8916 4764 8925
rect 9680 8916 9732 8968
rect 10232 8916 10284 8968
rect 10600 8916 10652 8968
rect 3976 8848 4028 8900
rect 2412 8823 2464 8832
rect 2412 8789 2421 8823
rect 2421 8789 2455 8823
rect 2455 8789 2464 8823
rect 2412 8780 2464 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 1400 8576 1452 8628
rect 2780 8576 2832 8628
rect 3056 8576 3108 8628
rect 4068 8576 4120 8628
rect 5356 8576 5408 8628
rect 6460 8619 6512 8628
rect 6460 8585 6469 8619
rect 6469 8585 6503 8619
rect 6503 8585 6512 8619
rect 6460 8576 6512 8585
rect 7012 8619 7064 8628
rect 7012 8585 7021 8619
rect 7021 8585 7055 8619
rect 7055 8585 7064 8619
rect 7012 8576 7064 8585
rect 8024 8576 8076 8628
rect 8944 8576 8996 8628
rect 10600 8619 10652 8628
rect 10600 8585 10609 8619
rect 10609 8585 10643 8619
rect 10643 8585 10652 8619
rect 10600 8576 10652 8585
rect 3148 8551 3200 8560
rect 3148 8517 3157 8551
rect 3157 8517 3191 8551
rect 3191 8517 3200 8551
rect 3148 8508 3200 8517
rect 3884 8440 3936 8492
rect 9680 8551 9732 8560
rect 9680 8517 9689 8551
rect 9689 8517 9723 8551
rect 9723 8517 9732 8551
rect 9680 8508 9732 8517
rect 7656 8483 7708 8492
rect 3976 8372 4028 8424
rect 7656 8449 7665 8483
rect 7665 8449 7699 8483
rect 7699 8449 7708 8483
rect 7656 8440 7708 8449
rect 10048 8440 10100 8492
rect 4712 8372 4764 8424
rect 8024 8304 8076 8356
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 3884 8075 3936 8084
rect 3884 8041 3893 8075
rect 3893 8041 3927 8075
rect 3927 8041 3936 8075
rect 3884 8032 3936 8041
rect 4528 8075 4580 8084
rect 4528 8041 4537 8075
rect 4537 8041 4571 8075
rect 4571 8041 4580 8075
rect 4528 8032 4580 8041
rect 6552 8032 6604 8084
rect 7656 8075 7708 8084
rect 7656 8041 7665 8075
rect 7665 8041 7699 8075
rect 7699 8041 7708 8075
rect 7656 8032 7708 8041
rect 10048 8032 10100 8084
rect 23388 8032 23440 8084
rect 3976 7964 4028 8016
rect 4160 7964 4212 8016
rect 22284 7939 22336 7948
rect 22284 7905 22293 7939
rect 22293 7905 22327 7939
rect 22327 7905 22336 7939
rect 22284 7896 22336 7905
rect 4804 7828 4856 7880
rect 4068 7803 4120 7812
rect 4068 7769 4077 7803
rect 4077 7769 4111 7803
rect 4111 7769 4120 7803
rect 4068 7760 4120 7769
rect 572 7692 624 7744
rect 4896 7692 4948 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 4160 7531 4212 7540
rect 4160 7497 4169 7531
rect 4169 7497 4203 7531
rect 4203 7497 4212 7531
rect 4160 7488 4212 7497
rect 4528 7488 4580 7540
rect 22284 7531 22336 7540
rect 22284 7497 22293 7531
rect 22293 7497 22327 7531
rect 22327 7497 22336 7531
rect 22284 7488 22336 7497
rect 23848 7531 23900 7540
rect 23848 7497 23857 7531
rect 23857 7497 23891 7531
rect 23891 7497 23900 7531
rect 23848 7488 23900 7497
rect 4804 7352 4856 7404
rect 23664 7327 23716 7336
rect 23664 7293 23673 7327
rect 23673 7293 23707 7327
rect 23707 7293 23716 7327
rect 23664 7284 23716 7293
rect 572 7148 624 7200
rect 3424 7148 3476 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 24768 6400 24820 6452
rect 23664 6239 23716 6248
rect 23664 6205 23673 6239
rect 23673 6205 23707 6239
rect 23707 6205 23716 6239
rect 23664 6196 23716 6205
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 24768 5856 24820 5908
rect 24032 5763 24084 5772
rect 24032 5729 24041 5763
rect 24041 5729 24075 5763
rect 24075 5729 24084 5763
rect 24032 5720 24084 5729
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 24032 5355 24084 5364
rect 24032 5321 24041 5355
rect 24041 5321 24075 5355
rect 24075 5321 24084 5355
rect 24032 5312 24084 5321
rect 24676 5355 24728 5364
rect 24676 5321 24685 5355
rect 24685 5321 24719 5355
rect 24719 5321 24728 5355
rect 24676 5312 24728 5321
rect 24492 5151 24544 5160
rect 24492 5117 24501 5151
rect 24501 5117 24535 5151
rect 24535 5117 24544 5151
rect 24492 5108 24544 5117
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 24768 4811 24820 4820
rect 24768 4777 24777 4811
rect 24777 4777 24811 4811
rect 24811 4777 24820 4811
rect 24768 4768 24820 4777
rect 24584 4675 24636 4684
rect 24584 4641 24593 4675
rect 24593 4641 24627 4675
rect 24627 4641 24636 4675
rect 24584 4632 24636 4641
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 24676 4267 24728 4276
rect 24676 4233 24685 4267
rect 24685 4233 24719 4267
rect 24719 4233 24728 4267
rect 24676 4224 24728 4233
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
<< metal2 >>
rect 294 27520 350 28000
rect 846 27520 902 28000
rect 1398 27520 1454 28000
rect 1950 27520 2006 28000
rect 2502 27520 2558 28000
rect 3146 27520 3202 28000
rect 3698 27520 3754 28000
rect 3882 27704 3938 27713
rect 3882 27639 3938 27648
rect 308 18873 336 27520
rect 294 18864 350 18873
rect 294 18799 350 18808
rect 860 17649 888 27520
rect 1412 23610 1440 27520
rect 1412 23582 1532 23610
rect 1400 23520 1452 23526
rect 1400 23462 1452 23468
rect 1412 20369 1440 23462
rect 1504 21162 1532 23582
rect 1582 22264 1638 22273
rect 1582 22199 1638 22208
rect 1596 21962 1624 22199
rect 1584 21956 1636 21962
rect 1584 21898 1636 21904
rect 1768 21412 1820 21418
rect 1768 21354 1820 21360
rect 1780 21185 1808 21354
rect 1766 21176 1822 21185
rect 1504 21134 1624 21162
rect 1492 21004 1544 21010
rect 1492 20946 1544 20952
rect 1504 20602 1532 20946
rect 1492 20596 1544 20602
rect 1492 20538 1544 20544
rect 1398 20360 1454 20369
rect 1398 20295 1454 20304
rect 1490 19952 1546 19961
rect 1490 19887 1492 19896
rect 1544 19887 1546 19896
rect 1492 19858 1544 19864
rect 1504 18970 1532 19858
rect 1492 18964 1544 18970
rect 1492 18906 1544 18912
rect 1596 18222 1624 21134
rect 1766 21111 1822 21120
rect 1584 18216 1636 18222
rect 1636 18176 1716 18204
rect 1584 18158 1636 18164
rect 1400 18080 1452 18086
rect 1400 18022 1452 18028
rect 846 17640 902 17649
rect 846 17575 902 17584
rect 1412 16046 1440 18022
rect 1492 16788 1544 16794
rect 1492 16730 1544 16736
rect 1400 16040 1452 16046
rect 1398 16008 1400 16017
rect 1452 16008 1454 16017
rect 1398 15943 1454 15952
rect 1504 15473 1532 16730
rect 1582 16688 1638 16697
rect 1582 16623 1638 16632
rect 1596 16250 1624 16623
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1584 16040 1636 16046
rect 1584 15982 1636 15988
rect 1596 15570 1624 15982
rect 1584 15564 1636 15570
rect 1584 15506 1636 15512
rect 1490 15464 1546 15473
rect 1490 15399 1546 15408
rect 1596 14906 1624 15506
rect 1504 14878 1624 14906
rect 1504 12782 1532 14878
rect 1584 14816 1636 14822
rect 1584 14758 1636 14764
rect 1596 14618 1624 14758
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 1596 13870 1624 14554
rect 1584 13864 1636 13870
rect 1584 13806 1636 13812
rect 1688 13530 1716 18176
rect 1964 18086 1992 27520
rect 2516 26874 2544 27520
rect 2332 26846 2544 26874
rect 2332 25514 2360 26846
rect 2240 25486 2360 25514
rect 2044 25152 2096 25158
rect 2044 25094 2096 25100
rect 2056 24886 2084 25094
rect 2044 24880 2096 24886
rect 2044 24822 2096 24828
rect 2042 23624 2098 23633
rect 2042 23559 2044 23568
rect 2096 23559 2098 23568
rect 2044 23530 2096 23536
rect 2042 22264 2098 22273
rect 2042 22199 2098 22208
rect 2056 22098 2084 22199
rect 2044 22092 2096 22098
rect 2044 22034 2096 22040
rect 2056 21486 2084 22034
rect 2044 21480 2096 21486
rect 2044 21422 2096 21428
rect 2044 20596 2096 20602
rect 2044 20538 2096 20544
rect 2056 18970 2084 20538
rect 2136 19304 2188 19310
rect 2136 19246 2188 19252
rect 2044 18964 2096 18970
rect 2044 18906 2096 18912
rect 2044 18828 2096 18834
rect 2044 18770 2096 18776
rect 2056 18170 2084 18770
rect 2148 18306 2176 19246
rect 2240 18834 2268 25486
rect 2320 25424 2372 25430
rect 2320 25366 2372 25372
rect 2332 24818 2360 25366
rect 2504 25356 2556 25362
rect 2504 25298 2556 25304
rect 2596 25356 2648 25362
rect 2596 25298 2648 25304
rect 2412 25152 2464 25158
rect 2412 25094 2464 25100
rect 2320 24812 2372 24818
rect 2320 24754 2372 24760
rect 2424 24274 2452 25094
rect 2516 24954 2544 25298
rect 2504 24948 2556 24954
rect 2504 24890 2556 24896
rect 2412 24268 2464 24274
rect 2412 24210 2464 24216
rect 2504 24268 2556 24274
rect 2504 24210 2556 24216
rect 2424 23866 2452 24210
rect 2412 23860 2464 23866
rect 2412 23802 2464 23808
rect 2412 23180 2464 23186
rect 2412 23122 2464 23128
rect 2318 22944 2374 22953
rect 2318 22879 2374 22888
rect 2332 22030 2360 22879
rect 2424 22438 2452 23122
rect 2412 22432 2464 22438
rect 2412 22374 2464 22380
rect 2320 22024 2372 22030
rect 2320 21966 2372 21972
rect 2332 21690 2360 21966
rect 2320 21684 2372 21690
rect 2320 21626 2372 21632
rect 2320 20392 2372 20398
rect 2320 20334 2372 20340
rect 2332 19718 2360 20334
rect 2424 19990 2452 22374
rect 2516 20466 2544 24210
rect 2608 23254 2636 25298
rect 2872 25220 2924 25226
rect 2872 25162 2924 25168
rect 2780 25152 2832 25158
rect 2780 25094 2832 25100
rect 2688 24744 2740 24750
rect 2792 24721 2820 25094
rect 2688 24686 2740 24692
rect 2778 24712 2834 24721
rect 2596 23248 2648 23254
rect 2596 23190 2648 23196
rect 2700 22642 2728 24686
rect 2778 24647 2834 24656
rect 2884 24426 2912 25162
rect 3056 24608 3108 24614
rect 3056 24550 3108 24556
rect 2792 24398 2912 24426
rect 2792 23202 2820 24398
rect 2872 24268 2924 24274
rect 2872 24210 2924 24216
rect 2884 23866 2912 24210
rect 2964 24064 3016 24070
rect 3068 24041 3096 24550
rect 2964 24006 3016 24012
rect 3054 24032 3110 24041
rect 2872 23860 2924 23866
rect 2872 23802 2924 23808
rect 2792 23174 2912 23202
rect 2780 23112 2832 23118
rect 2780 23054 2832 23060
rect 2688 22636 2740 22642
rect 2688 22578 2740 22584
rect 2686 22536 2742 22545
rect 2686 22471 2688 22480
rect 2740 22471 2742 22480
rect 2688 22442 2740 22448
rect 2594 22400 2650 22409
rect 2594 22335 2650 22344
rect 2608 21078 2636 22335
rect 2700 22234 2728 22442
rect 2688 22228 2740 22234
rect 2688 22170 2740 22176
rect 2688 22092 2740 22098
rect 2688 22034 2740 22040
rect 2700 21321 2728 22034
rect 2792 21690 2820 23054
rect 2884 22817 2912 23174
rect 2870 22808 2926 22817
rect 2870 22743 2926 22752
rect 2872 21888 2924 21894
rect 2872 21830 2924 21836
rect 2780 21684 2832 21690
rect 2780 21626 2832 21632
rect 2686 21312 2742 21321
rect 2686 21247 2742 21256
rect 2700 21146 2728 21247
rect 2688 21140 2740 21146
rect 2688 21082 2740 21088
rect 2596 21072 2648 21078
rect 2596 21014 2648 21020
rect 2504 20460 2556 20466
rect 2504 20402 2556 20408
rect 2688 20324 2740 20330
rect 2780 20324 2832 20330
rect 2740 20284 2780 20312
rect 2688 20266 2740 20272
rect 2780 20266 2832 20272
rect 2412 19984 2464 19990
rect 2412 19926 2464 19932
rect 2884 19825 2912 21830
rect 2976 21593 3004 24006
rect 3054 23967 3110 23976
rect 3056 22976 3108 22982
rect 3056 22918 3108 22924
rect 2962 21584 3018 21593
rect 2962 21519 3018 21528
rect 3068 21049 3096 22918
rect 3160 22420 3188 27520
rect 3514 27160 3570 27169
rect 3514 27095 3570 27104
rect 3528 26314 3556 27095
rect 3516 26308 3568 26314
rect 3516 26250 3568 26256
rect 3330 25936 3386 25945
rect 3330 25871 3386 25880
rect 3344 25498 3372 25871
rect 3332 25492 3384 25498
rect 3332 25434 3384 25440
rect 3712 24834 3740 27520
rect 3896 26722 3924 27639
rect 4250 27520 4306 28000
rect 4802 27520 4858 28000
rect 5354 27520 5410 28000
rect 5998 27520 6054 28000
rect 6550 27520 6606 28000
rect 7102 27520 7158 28000
rect 7654 27520 7710 28000
rect 8206 27520 8262 28000
rect 8850 27520 8906 28000
rect 9402 27520 9458 28000
rect 9954 27520 10010 28000
rect 10506 27520 10562 28000
rect 11058 27520 11114 28000
rect 11702 27520 11758 28000
rect 12254 27520 12310 28000
rect 12806 27520 12862 28000
rect 13358 27520 13414 28000
rect 13910 27520 13966 28000
rect 14554 27520 14610 28000
rect 15106 27520 15162 28000
rect 15658 27520 15714 28000
rect 16210 27520 16266 28000
rect 16762 27520 16818 28000
rect 17406 27520 17462 28000
rect 17958 27520 18014 28000
rect 18510 27520 18566 28000
rect 19062 27520 19118 28000
rect 19614 27520 19670 28000
rect 20258 27520 20314 28000
rect 20810 27520 20866 28000
rect 21362 27520 21418 28000
rect 21914 27520 21970 28000
rect 22466 27520 22522 28000
rect 23110 27520 23166 28000
rect 23662 27520 23718 28000
rect 24214 27520 24270 28000
rect 24766 27520 24822 28000
rect 25318 27520 25374 28000
rect 25962 27520 26018 28000
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 3884 26716 3936 26722
rect 3884 26658 3936 26664
rect 4066 26480 4122 26489
rect 4066 26415 4068 26424
rect 4120 26415 4122 26424
rect 4068 26386 4120 26392
rect 4160 25356 4212 25362
rect 4160 25298 4212 25304
rect 4066 25256 4122 25265
rect 3792 25220 3844 25226
rect 4066 25191 4122 25200
rect 3792 25162 3844 25168
rect 3620 24806 3740 24834
rect 3332 24132 3384 24138
rect 3332 24074 3384 24080
rect 3240 23724 3292 23730
rect 3240 23666 3292 23672
rect 3252 23361 3280 23666
rect 3344 23594 3372 24074
rect 3332 23588 3384 23594
rect 3332 23530 3384 23536
rect 3424 23520 3476 23526
rect 3424 23462 3476 23468
rect 3238 23352 3294 23361
rect 3238 23287 3294 23296
rect 3252 23050 3280 23287
rect 3240 23044 3292 23050
rect 3240 22986 3292 22992
rect 3252 22574 3280 22986
rect 3240 22568 3292 22574
rect 3240 22510 3292 22516
rect 3160 22392 3280 22420
rect 3148 21888 3200 21894
rect 3148 21830 3200 21836
rect 3160 21690 3188 21830
rect 3148 21684 3200 21690
rect 3148 21626 3200 21632
rect 3146 21584 3202 21593
rect 3146 21519 3202 21528
rect 3160 21418 3188 21519
rect 3148 21412 3200 21418
rect 3148 21354 3200 21360
rect 3054 21040 3110 21049
rect 3054 20975 3110 20984
rect 2964 20800 3016 20806
rect 2964 20742 3016 20748
rect 2870 19816 2926 19825
rect 2870 19751 2926 19760
rect 2320 19712 2372 19718
rect 2320 19654 2372 19660
rect 2872 19712 2924 19718
rect 2872 19654 2924 19660
rect 2332 19417 2360 19654
rect 2318 19408 2374 19417
rect 2318 19343 2374 19352
rect 2320 19236 2372 19242
rect 2320 19178 2372 19184
rect 2780 19236 2832 19242
rect 2780 19178 2832 19184
rect 2228 18828 2280 18834
rect 2228 18770 2280 18776
rect 2228 18624 2280 18630
rect 2228 18566 2280 18572
rect 2240 18465 2268 18566
rect 2226 18456 2282 18465
rect 2226 18391 2282 18400
rect 2226 18320 2282 18329
rect 2148 18278 2226 18306
rect 2226 18255 2228 18264
rect 2280 18255 2282 18264
rect 2228 18226 2280 18232
rect 2056 18142 2176 18170
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 1964 17678 1992 17709
rect 1768 17672 1820 17678
rect 1952 17672 2004 17678
rect 1768 17614 1820 17620
rect 1950 17640 1952 17649
rect 2004 17640 2006 17649
rect 1780 17134 1808 17614
rect 1950 17575 2006 17584
rect 1964 17270 1992 17575
rect 1952 17264 2004 17270
rect 1952 17206 2004 17212
rect 1768 17128 1820 17134
rect 1768 17070 1820 17076
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 1872 16794 1900 16934
rect 1860 16788 1912 16794
rect 1860 16730 1912 16736
rect 1964 14906 1992 17206
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 2056 16794 2084 17138
rect 2148 17066 2176 18142
rect 2332 17882 2360 19178
rect 2792 18766 2820 19178
rect 2688 18760 2740 18766
rect 2688 18702 2740 18708
rect 2780 18760 2832 18766
rect 2780 18702 2832 18708
rect 2596 18148 2648 18154
rect 2596 18090 2648 18096
rect 2320 17876 2372 17882
rect 2320 17818 2372 17824
rect 2332 17202 2360 17818
rect 2502 17640 2558 17649
rect 2608 17610 2636 18090
rect 2700 17882 2728 18702
rect 2780 18080 2832 18086
rect 2780 18022 2832 18028
rect 2688 17876 2740 17882
rect 2688 17818 2740 17824
rect 2792 17814 2820 18022
rect 2884 17921 2912 19654
rect 2976 19145 3004 20742
rect 3148 20256 3200 20262
rect 3148 20198 3200 20204
rect 3160 19786 3188 20198
rect 3148 19780 3200 19786
rect 3148 19722 3200 19728
rect 3160 19378 3188 19722
rect 3148 19372 3200 19378
rect 3148 19314 3200 19320
rect 2962 19136 3018 19145
rect 2962 19071 3018 19080
rect 2870 17912 2926 17921
rect 2870 17847 2926 17856
rect 2780 17808 2832 17814
rect 2780 17750 2832 17756
rect 2502 17575 2558 17584
rect 2596 17604 2648 17610
rect 2516 17338 2544 17575
rect 2596 17546 2648 17552
rect 2504 17332 2556 17338
rect 2504 17274 2556 17280
rect 2320 17196 2372 17202
rect 2320 17138 2372 17144
rect 2136 17060 2188 17066
rect 2136 17002 2188 17008
rect 2044 16788 2096 16794
rect 2044 16730 2096 16736
rect 2044 15904 2096 15910
rect 2044 15846 2096 15852
rect 2056 15570 2084 15846
rect 2044 15564 2096 15570
rect 2044 15506 2096 15512
rect 2056 15026 2084 15506
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 1964 14878 2084 14906
rect 2056 14822 2084 14878
rect 2044 14816 2096 14822
rect 2044 14758 2096 14764
rect 1858 14376 1914 14385
rect 1858 14311 1860 14320
rect 1912 14311 1914 14320
rect 1860 14282 1912 14288
rect 1872 14006 1900 14282
rect 1860 14000 1912 14006
rect 1860 13942 1912 13948
rect 2056 13569 2084 14758
rect 2042 13560 2098 13569
rect 1676 13524 1728 13530
rect 2042 13495 2098 13504
rect 1676 13466 1728 13472
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 1492 12776 1544 12782
rect 1492 12718 1544 12724
rect 1780 12481 1808 13330
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 2056 12782 2084 13262
rect 2044 12776 2096 12782
rect 2044 12718 2096 12724
rect 1766 12472 1822 12481
rect 2148 12442 2176 17002
rect 2792 16998 2820 17750
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 3252 17626 3280 22392
rect 3436 22114 3464 23462
rect 3516 22976 3568 22982
rect 3516 22918 3568 22924
rect 3528 22234 3556 22918
rect 3516 22228 3568 22234
rect 3516 22170 3568 22176
rect 3436 22086 3556 22114
rect 3332 22024 3384 22030
rect 3332 21966 3384 21972
rect 3344 21554 3372 21966
rect 3424 21616 3476 21622
rect 3424 21558 3476 21564
rect 3332 21548 3384 21554
rect 3332 21490 3384 21496
rect 3436 21146 3464 21558
rect 3424 21140 3476 21146
rect 3424 21082 3476 21088
rect 3332 20936 3384 20942
rect 3332 20878 3384 20884
rect 3344 20058 3372 20878
rect 3424 20460 3476 20466
rect 3424 20402 3476 20408
rect 3436 20369 3464 20402
rect 3422 20360 3478 20369
rect 3422 20295 3478 20304
rect 3528 20058 3556 22086
rect 3332 20052 3384 20058
rect 3332 19994 3384 20000
rect 3516 20052 3568 20058
rect 3516 19994 3568 20000
rect 3332 19916 3384 19922
rect 3332 19858 3384 19864
rect 3344 18737 3372 19858
rect 3422 19136 3478 19145
rect 3422 19071 3478 19080
rect 3330 18728 3386 18737
rect 3330 18663 3332 18672
rect 3384 18663 3386 18672
rect 3332 18634 3384 18640
rect 3436 18329 3464 19071
rect 3620 18850 3648 24806
rect 3804 21162 3832 25162
rect 4080 24834 4108 25191
rect 4172 24954 4200 25298
rect 4160 24948 4212 24954
rect 4160 24890 4212 24896
rect 4080 24806 4200 24834
rect 4172 24410 4200 24806
rect 4264 24732 4292 27520
rect 4712 25152 4764 25158
rect 4712 25094 4764 25100
rect 4724 24818 4752 25094
rect 4816 24834 4844 27520
rect 4896 26308 4948 26314
rect 4896 26250 4948 26256
rect 4908 25226 4936 26250
rect 5368 25430 5396 27520
rect 5540 26444 5592 26450
rect 5540 26386 5592 26392
rect 5356 25424 5408 25430
rect 5356 25366 5408 25372
rect 5264 25288 5316 25294
rect 5264 25230 5316 25236
rect 4896 25220 4948 25226
rect 4896 25162 4948 25168
rect 4712 24812 4764 24818
rect 4816 24806 5212 24834
rect 4712 24754 4764 24760
rect 4264 24704 4384 24732
rect 4160 24404 4212 24410
rect 4160 24346 4212 24352
rect 4068 24268 4120 24274
rect 4120 24228 4200 24256
rect 4068 24210 4120 24216
rect 4068 23588 4120 23594
rect 4068 23530 4120 23536
rect 4080 23202 4108 23530
rect 4172 23322 4200 24228
rect 4160 23316 4212 23322
rect 4160 23258 4212 23264
rect 3884 23180 3936 23186
rect 4080 23174 4200 23202
rect 3884 23122 3936 23128
rect 3896 22506 3924 23122
rect 3974 22536 4030 22545
rect 3884 22500 3936 22506
rect 3974 22471 4030 22480
rect 3884 22442 3936 22448
rect 3712 21134 3832 21162
rect 3712 20330 3740 21134
rect 3792 21072 3844 21078
rect 3792 21014 3844 21020
rect 3804 20602 3832 21014
rect 3896 21010 3924 22442
rect 3884 21004 3936 21010
rect 3884 20946 3936 20952
rect 3988 20942 4016 22471
rect 4172 21962 4200 23174
rect 4252 22432 4304 22438
rect 4252 22374 4304 22380
rect 4160 21956 4212 21962
rect 4160 21898 4212 21904
rect 4160 21548 4212 21554
rect 4160 21490 4212 21496
rect 4172 21146 4200 21490
rect 4160 21140 4212 21146
rect 4160 21082 4212 21088
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 4172 20602 4200 21082
rect 4264 21078 4292 22374
rect 4252 21072 4304 21078
rect 4252 21014 4304 21020
rect 3792 20596 3844 20602
rect 3792 20538 3844 20544
rect 4160 20596 4212 20602
rect 4160 20538 4212 20544
rect 3700 20324 3752 20330
rect 3700 20266 3752 20272
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 4080 18970 4108 19654
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 3528 18822 3648 18850
rect 3700 18828 3752 18834
rect 3422 18320 3478 18329
rect 3422 18255 3478 18264
rect 3332 17672 3384 17678
rect 3252 17620 3332 17626
rect 3252 17614 3384 17620
rect 3068 17338 3096 17614
rect 3252 17598 3372 17614
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 2780 16992 2832 16998
rect 2780 16934 2832 16940
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 2228 16720 2280 16726
rect 2228 16662 2280 16668
rect 2240 15162 2268 16662
rect 2412 16652 2464 16658
rect 2412 16594 2464 16600
rect 2228 15156 2280 15162
rect 2228 15098 2280 15104
rect 2240 14550 2268 15098
rect 2424 14618 2452 16594
rect 2412 14612 2464 14618
rect 2412 14554 2464 14560
rect 2228 14544 2280 14550
rect 2228 14486 2280 14492
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2424 14006 2452 14350
rect 2412 14000 2464 14006
rect 2412 13942 2464 13948
rect 2424 12594 2452 13942
rect 2516 13818 2544 16730
rect 2596 16584 2648 16590
rect 2596 16526 2648 16532
rect 2608 15910 2636 16526
rect 2596 15904 2648 15910
rect 2596 15846 2648 15852
rect 2608 15366 2636 15846
rect 2596 15360 2648 15366
rect 2596 15302 2648 15308
rect 2608 14278 2636 15302
rect 2792 14890 2820 16934
rect 3068 16794 3096 17274
rect 3252 17270 3280 17598
rect 3240 17264 3292 17270
rect 3240 17206 3292 17212
rect 3056 16788 3108 16794
rect 3056 16730 3108 16736
rect 3146 16280 3202 16289
rect 3146 16215 3202 16224
rect 2964 15020 3016 15026
rect 2964 14962 3016 14968
rect 2780 14884 2832 14890
rect 2780 14826 2832 14832
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 2884 14414 2912 14554
rect 2976 14414 3004 14962
rect 3056 14884 3108 14890
rect 3056 14826 3108 14832
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 3068 14346 3096 14826
rect 3056 14340 3108 14346
rect 3056 14282 3108 14288
rect 2596 14272 2648 14278
rect 2596 14214 2648 14220
rect 2608 13938 2636 14214
rect 2964 14000 3016 14006
rect 2962 13968 2964 13977
rect 3016 13968 3018 13977
rect 2596 13932 2648 13938
rect 2962 13903 3018 13912
rect 2596 13874 2648 13880
rect 2780 13864 2832 13870
rect 2516 13812 2780 13818
rect 2516 13806 2832 13812
rect 2516 13790 2820 13806
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 2872 13184 2924 13190
rect 2872 13126 2924 13132
rect 2424 12566 2544 12594
rect 2410 12472 2466 12481
rect 1766 12407 1822 12416
rect 2136 12436 2188 12442
rect 2410 12407 2412 12416
rect 2136 12378 2188 12384
rect 2464 12407 2466 12416
rect 2412 12378 2464 12384
rect 1584 12300 1636 12306
rect 1584 12242 1636 12248
rect 1398 11656 1454 11665
rect 1398 11591 1454 11600
rect 1412 11354 1440 11591
rect 1596 11558 1624 12242
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1596 11257 1624 11494
rect 1872 11354 1900 12038
rect 2148 11898 2176 12378
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1582 11248 1638 11257
rect 1582 11183 1638 11192
rect 2044 10804 2096 10810
rect 2044 10746 2096 10752
rect 2056 10198 2084 10746
rect 2134 10704 2190 10713
rect 2134 10639 2136 10648
rect 2188 10639 2190 10648
rect 2136 10610 2188 10616
rect 2516 10538 2544 12566
rect 2700 12458 2728 13126
rect 2884 12889 2912 13126
rect 2870 12880 2926 12889
rect 2926 12838 3004 12866
rect 2870 12815 2926 12824
rect 2872 12640 2924 12646
rect 2872 12582 2924 12588
rect 2700 12430 2820 12458
rect 2792 12374 2820 12430
rect 2780 12368 2832 12374
rect 2780 12310 2832 12316
rect 2884 12050 2912 12582
rect 2976 12442 3004 12838
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 2792 12022 2912 12050
rect 2792 11626 2820 12022
rect 2870 11928 2926 11937
rect 2870 11863 2926 11872
rect 2780 11620 2832 11626
rect 2780 11562 2832 11568
rect 2792 11286 2820 11562
rect 2780 11280 2832 11286
rect 2780 11222 2832 11228
rect 2504 10532 2556 10538
rect 2504 10474 2556 10480
rect 2688 10464 2740 10470
rect 2688 10406 2740 10412
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2044 10192 2096 10198
rect 2044 10134 2096 10140
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9586 1440 9998
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1412 8634 1440 9522
rect 1768 9444 1820 9450
rect 1768 9386 1820 9392
rect 1780 9178 1808 9386
rect 2056 9178 2084 10134
rect 2502 9616 2558 9625
rect 2502 9551 2558 9560
rect 2516 9382 2544 9551
rect 2608 9450 2636 10202
rect 2596 9444 2648 9450
rect 2596 9386 2648 9392
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2700 9194 2728 10406
rect 2700 9178 2820 9194
rect 1768 9172 1820 9178
rect 1768 9114 1820 9120
rect 2044 9172 2096 9178
rect 2700 9172 2832 9178
rect 2700 9166 2780 9172
rect 2044 9114 2096 9120
rect 2780 9114 2832 9120
rect 2884 9058 2912 11863
rect 3068 9110 3096 14282
rect 3160 14074 3188 16215
rect 3252 14618 3280 17206
rect 3436 17202 3464 18255
rect 3424 17196 3476 17202
rect 3424 17138 3476 17144
rect 3528 16454 3556 18822
rect 3700 18770 3752 18776
rect 4160 18828 4212 18834
rect 4160 18770 4212 18776
rect 3608 18760 3660 18766
rect 3608 18702 3660 18708
rect 3620 18426 3648 18702
rect 3712 18630 3740 18770
rect 3700 18624 3752 18630
rect 3700 18566 3752 18572
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 3712 17882 3740 18566
rect 4068 18352 4120 18358
rect 4068 18294 4120 18300
rect 4172 18306 4200 18770
rect 4252 18624 4304 18630
rect 4250 18592 4252 18601
rect 4304 18592 4306 18601
rect 4250 18527 4306 18536
rect 4250 18320 4306 18329
rect 3700 17876 3752 17882
rect 3700 17818 3752 17824
rect 3792 17536 3844 17542
rect 3792 17478 3844 17484
rect 3804 16658 3832 17478
rect 4080 17134 4108 18294
rect 4172 18278 4250 18306
rect 4250 18255 4252 18264
rect 4304 18255 4306 18264
rect 4252 18226 4304 18232
rect 4356 17746 4384 24704
rect 4724 24410 4752 24754
rect 4712 24404 4764 24410
rect 4712 24346 4764 24352
rect 4436 24336 4488 24342
rect 4436 24278 4488 24284
rect 4710 24304 4766 24313
rect 4448 24070 4476 24278
rect 4528 24268 4580 24274
rect 4710 24239 4766 24248
rect 4528 24210 4580 24216
rect 4436 24064 4488 24070
rect 4436 24006 4488 24012
rect 4448 23594 4476 24006
rect 4540 23662 4568 24210
rect 4528 23656 4580 23662
rect 4528 23598 4580 23604
rect 4436 23588 4488 23594
rect 4436 23530 4488 23536
rect 4448 23186 4476 23530
rect 4436 23180 4488 23186
rect 4436 23122 4488 23128
rect 4620 20324 4672 20330
rect 4620 20266 4672 20272
rect 4632 19854 4660 20266
rect 4620 19848 4672 19854
rect 4620 19790 4672 19796
rect 4632 19174 4660 19790
rect 4724 19310 4752 24239
rect 4988 23248 5040 23254
rect 4988 23190 5040 23196
rect 5078 23216 5134 23225
rect 5000 22778 5028 23190
rect 5078 23151 5134 23160
rect 4988 22772 5040 22778
rect 4988 22714 5040 22720
rect 5000 22030 5028 22714
rect 4804 22024 4856 22030
rect 4802 21992 4804 22001
rect 4988 22024 5040 22030
rect 4856 21992 4858 22001
rect 4988 21966 5040 21972
rect 4802 21927 4858 21936
rect 4816 21690 4844 21927
rect 4804 21684 4856 21690
rect 4804 21626 4856 21632
rect 4896 21548 4948 21554
rect 4896 21490 4948 21496
rect 4908 21078 4936 21490
rect 5092 21486 5120 23151
rect 5080 21480 5132 21486
rect 5080 21422 5132 21428
rect 4896 21072 4948 21078
rect 4896 21014 4948 21020
rect 4896 19712 4948 19718
rect 4896 19654 4948 19660
rect 4908 19310 4936 19654
rect 4712 19304 4764 19310
rect 4712 19246 4764 19252
rect 4896 19304 4948 19310
rect 4896 19246 4948 19252
rect 4988 19304 5040 19310
rect 4988 19246 5040 19252
rect 4528 19168 4580 19174
rect 4620 19168 4672 19174
rect 4528 19110 4580 19116
rect 4618 19136 4620 19145
rect 4672 19136 4674 19145
rect 4436 18624 4488 18630
rect 4436 18566 4488 18572
rect 4344 17740 4396 17746
rect 4344 17682 4396 17688
rect 4250 17368 4306 17377
rect 4250 17303 4306 17312
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 4080 16794 4108 17070
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 3792 16652 3844 16658
rect 3792 16594 3844 16600
rect 3884 16516 3936 16522
rect 3884 16458 3936 16464
rect 3516 16448 3568 16454
rect 3516 16390 3568 16396
rect 3790 16144 3846 16153
rect 3790 16079 3846 16088
rect 3804 15065 3832 16079
rect 3896 15706 3924 16458
rect 4160 16040 4212 16046
rect 3988 16000 4160 16028
rect 3884 15700 3936 15706
rect 3884 15642 3936 15648
rect 3884 15564 3936 15570
rect 3884 15506 3936 15512
rect 3896 15473 3924 15506
rect 3882 15464 3938 15473
rect 3882 15399 3938 15408
rect 3896 15162 3924 15399
rect 3884 15156 3936 15162
rect 3884 15098 3936 15104
rect 3790 15056 3846 15065
rect 3790 14991 3846 15000
rect 3988 14929 4016 16000
rect 4160 15982 4212 15988
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 4160 15904 4212 15910
rect 4160 15846 4212 15852
rect 4080 15162 4108 15846
rect 4172 15570 4200 15846
rect 4264 15706 4292 17303
rect 4356 16658 4384 17682
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 4252 15700 4304 15706
rect 4252 15642 4304 15648
rect 4160 15564 4212 15570
rect 4160 15506 4212 15512
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 3974 14920 4030 14929
rect 3974 14855 4030 14864
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3330 14512 3386 14521
rect 3240 14476 3292 14482
rect 3330 14447 3386 14456
rect 3240 14418 3292 14424
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 3252 13977 3280 14418
rect 3238 13968 3294 13977
rect 3238 13903 3294 13912
rect 3344 12084 3372 14447
rect 4080 13938 4108 15098
rect 4172 14958 4200 15506
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 4172 14482 4200 14894
rect 4252 14884 4304 14890
rect 4252 14826 4304 14832
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 3608 13932 3660 13938
rect 3608 13874 3660 13880
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 3424 13728 3476 13734
rect 3424 13670 3476 13676
rect 3436 12986 3464 13670
rect 3620 13530 3648 13874
rect 3792 13864 3844 13870
rect 3792 13806 3844 13812
rect 3804 13530 3832 13806
rect 4172 13682 4200 14418
rect 4264 14074 4292 14826
rect 4252 14068 4304 14074
rect 4252 14010 4304 14016
rect 4356 13977 4384 16594
rect 4342 13968 4398 13977
rect 4342 13903 4398 13912
rect 4080 13654 4200 13682
rect 3608 13524 3660 13530
rect 3608 13466 3660 13472
rect 3792 13524 3844 13530
rect 3792 13466 3844 13472
rect 3882 13152 3938 13161
rect 3882 13087 3938 13096
rect 3424 12980 3476 12986
rect 3424 12922 3476 12928
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3424 12164 3476 12170
rect 3424 12106 3476 12112
rect 3252 12056 3372 12084
rect 3148 10532 3200 10538
rect 3148 10474 3200 10480
rect 2792 9042 2912 9058
rect 3056 9104 3108 9110
rect 3056 9046 3108 9052
rect 2780 9036 2912 9042
rect 2832 9030 2912 9036
rect 2780 8978 2832 8984
rect 2412 8832 2464 8838
rect 2412 8774 2464 8780
rect 1400 8628 1452 8634
rect 1400 8570 1452 8576
rect 2424 8129 2452 8774
rect 2792 8634 2820 8978
rect 3068 8634 3096 9046
rect 3160 8974 3188 10474
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 3160 8566 3188 8910
rect 3148 8560 3200 8566
rect 3148 8502 3200 8508
rect 2410 8120 2466 8129
rect 2410 8055 2466 8064
rect 572 7744 624 7750
rect 572 7686 624 7692
rect 584 7585 612 7686
rect 570 7576 626 7585
rect 570 7511 626 7520
rect 572 7200 624 7206
rect 572 7142 624 7148
rect 584 7041 612 7142
rect 570 7032 626 7041
rect 570 6967 626 6976
rect 3252 2689 3280 12056
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 3344 10470 3372 10950
rect 3436 10810 3464 12106
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3528 11218 3556 11494
rect 3516 11212 3568 11218
rect 3516 11154 3568 11160
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3344 10266 3372 10406
rect 3436 10266 3464 10610
rect 3528 10538 3556 11154
rect 3516 10532 3568 10538
rect 3516 10474 3568 10480
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3436 9722 3464 10202
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 3332 9648 3384 9654
rect 3332 9590 3384 9596
rect 3344 3913 3372 9590
rect 3422 7440 3478 7449
rect 3422 7375 3478 7384
rect 3436 7206 3464 7375
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3330 3904 3386 3913
rect 3330 3839 3386 3848
rect 3620 3369 3648 12378
rect 3790 12336 3846 12345
rect 3790 12271 3846 12280
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3712 9654 3740 9862
rect 3700 9648 3752 9654
rect 3700 9590 3752 9596
rect 3804 9042 3832 12271
rect 3896 11830 3924 13087
rect 3976 12640 4028 12646
rect 3976 12582 4028 12588
rect 3884 11824 3936 11830
rect 3884 11766 3936 11772
rect 3884 10260 3936 10266
rect 3884 10202 3936 10208
rect 3896 9518 3924 10202
rect 3988 10146 4016 12582
rect 4080 12345 4108 13654
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 4066 12336 4122 12345
rect 4172 12306 4200 13262
rect 4448 12442 4476 18566
rect 4540 18426 4568 19110
rect 4724 19122 4752 19246
rect 5000 19122 5028 19246
rect 4724 19094 5028 19122
rect 4618 19071 4674 19080
rect 4632 18834 4660 19071
rect 4620 18828 4672 18834
rect 4620 18770 4672 18776
rect 5184 18578 5212 24806
rect 5276 24750 5304 25230
rect 5356 24812 5408 24818
rect 5356 24754 5408 24760
rect 5264 24744 5316 24750
rect 5264 24686 5316 24692
rect 5368 24585 5396 24754
rect 5354 24576 5410 24585
rect 5354 24511 5410 24520
rect 5368 24274 5396 24511
rect 5356 24268 5408 24274
rect 5356 24210 5408 24216
rect 5552 23848 5580 26386
rect 6012 25362 6040 27520
rect 6564 25514 6592 27520
rect 7116 26874 7144 27520
rect 6472 25486 6592 25514
rect 6932 26846 7144 26874
rect 6000 25356 6052 25362
rect 6000 25298 6052 25304
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6012 24818 6040 25298
rect 6000 24812 6052 24818
rect 6000 24754 6052 24760
rect 5998 24712 6054 24721
rect 5998 24647 6054 24656
rect 6012 24410 6040 24647
rect 6276 24608 6328 24614
rect 6276 24550 6328 24556
rect 6000 24404 6052 24410
rect 6000 24346 6052 24352
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 6012 23866 6040 24346
rect 6000 23860 6052 23866
rect 5552 23820 5672 23848
rect 5540 23520 5592 23526
rect 5354 23488 5410 23497
rect 5540 23462 5592 23468
rect 5354 23423 5410 23432
rect 5368 22953 5396 23423
rect 5448 23248 5500 23254
rect 5552 23236 5580 23462
rect 5500 23208 5580 23236
rect 5448 23190 5500 23196
rect 5644 23168 5672 23820
rect 6000 23802 6052 23808
rect 5814 23352 5870 23361
rect 5814 23287 5816 23296
rect 5868 23287 5870 23296
rect 5816 23258 5868 23264
rect 6288 23186 6316 24550
rect 6472 24313 6500 25486
rect 6552 25424 6604 25430
rect 6552 25366 6604 25372
rect 6564 24818 6592 25366
rect 6552 24812 6604 24818
rect 6552 24754 6604 24760
rect 6458 24304 6514 24313
rect 6458 24239 6514 24248
rect 6552 24268 6604 24274
rect 6552 24210 6604 24216
rect 6460 24200 6512 24206
rect 6460 24142 6512 24148
rect 6472 23594 6500 24142
rect 6564 24041 6592 24210
rect 6550 24032 6606 24041
rect 6550 23967 6606 23976
rect 6564 23866 6592 23967
rect 6552 23860 6604 23866
rect 6552 23802 6604 23808
rect 6460 23588 6512 23594
rect 6460 23530 6512 23536
rect 6472 23322 6500 23530
rect 6828 23520 6880 23526
rect 6828 23462 6880 23468
rect 6460 23316 6512 23322
rect 6460 23258 6512 23264
rect 5552 23140 5672 23168
rect 6276 23180 6328 23186
rect 5354 22944 5410 22953
rect 5354 22879 5410 22888
rect 5552 22778 5580 23140
rect 6276 23122 6328 23128
rect 6090 23080 6146 23089
rect 6090 23015 6146 23024
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5540 22772 5592 22778
rect 5540 22714 5592 22720
rect 5264 22432 5316 22438
rect 5262 22400 5264 22409
rect 5316 22400 5318 22409
rect 5262 22335 5318 22344
rect 5446 22400 5502 22409
rect 5446 22335 5502 22344
rect 5460 22166 5488 22335
rect 5448 22160 5500 22166
rect 5448 22102 5500 22108
rect 5264 22092 5316 22098
rect 5264 22034 5316 22040
rect 5276 21894 5304 22034
rect 5264 21888 5316 21894
rect 5264 21830 5316 21836
rect 5276 20330 5304 21830
rect 5460 21690 5488 22102
rect 6000 22092 6052 22098
rect 6000 22034 6052 22040
rect 5540 22024 5592 22030
rect 5540 21966 5592 21972
rect 5552 21690 5580 21966
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5448 21684 5500 21690
rect 5448 21626 5500 21632
rect 5540 21684 5592 21690
rect 5540 21626 5592 21632
rect 5816 21344 5868 21350
rect 5816 21286 5868 21292
rect 5828 20913 5856 21286
rect 6012 21185 6040 22034
rect 6104 21962 6132 23015
rect 6288 22778 6316 23122
rect 6840 22778 6868 23462
rect 6932 23225 6960 26846
rect 7104 26716 7156 26722
rect 7104 26658 7156 26664
rect 7116 25226 7144 26658
rect 7104 25220 7156 25226
rect 7104 25162 7156 25168
rect 7012 24676 7064 24682
rect 7012 24618 7064 24624
rect 7024 24410 7052 24618
rect 7104 24608 7156 24614
rect 7104 24550 7156 24556
rect 7012 24404 7064 24410
rect 7012 24346 7064 24352
rect 6918 23216 6974 23225
rect 6918 23151 6974 23160
rect 7012 23112 7064 23118
rect 7012 23054 7064 23060
rect 6276 22772 6328 22778
rect 6276 22714 6328 22720
rect 6828 22772 6880 22778
rect 6828 22714 6880 22720
rect 6840 22574 6868 22714
rect 6828 22568 6880 22574
rect 6828 22510 6880 22516
rect 7024 22522 7052 23054
rect 7116 22681 7144 24550
rect 7380 24268 7432 24274
rect 7380 24210 7432 24216
rect 7392 23526 7420 24210
rect 7380 23520 7432 23526
rect 7380 23462 7432 23468
rect 7288 22976 7340 22982
rect 7288 22918 7340 22924
rect 7102 22672 7158 22681
rect 7102 22607 7158 22616
rect 7300 22574 7328 22918
rect 7380 22636 7432 22642
rect 7380 22578 7432 22584
rect 7288 22568 7340 22574
rect 7024 22494 7144 22522
rect 7288 22510 7340 22516
rect 6828 22432 6880 22438
rect 6828 22374 6880 22380
rect 6840 22273 6868 22374
rect 6826 22264 6882 22273
rect 6826 22199 6882 22208
rect 7116 22030 7144 22494
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 6092 21956 6144 21962
rect 6092 21898 6144 21904
rect 6460 21480 6512 21486
rect 6460 21422 6512 21428
rect 5998 21176 6054 21185
rect 5998 21111 6000 21120
rect 6052 21111 6054 21120
rect 6000 21082 6052 21088
rect 5814 20904 5870 20913
rect 5540 20868 5592 20874
rect 6472 20874 6500 21422
rect 7116 21350 7144 21966
rect 7300 21690 7328 22510
rect 7392 22098 7420 22578
rect 7380 22092 7432 22098
rect 7380 22034 7432 22040
rect 7288 21684 7340 21690
rect 7288 21626 7340 21632
rect 7392 21418 7420 22034
rect 7668 22001 7696 27520
rect 8022 24848 8078 24857
rect 8022 24783 8078 24792
rect 7840 24744 7892 24750
rect 7840 24686 7892 24692
rect 7852 24342 7880 24686
rect 7840 24336 7892 24342
rect 7840 24278 7892 24284
rect 7852 23730 7880 24278
rect 7840 23724 7892 23730
rect 7840 23666 7892 23672
rect 7852 23322 7880 23666
rect 7840 23316 7892 23322
rect 7840 23258 7892 23264
rect 7654 21992 7710 22001
rect 7654 21927 7710 21936
rect 8036 21554 8064 24783
rect 8220 24721 8248 27520
rect 8206 24712 8262 24721
rect 8206 24647 8262 24656
rect 8208 24608 8260 24614
rect 8208 24550 8260 24556
rect 8482 24576 8538 24585
rect 8116 23588 8168 23594
rect 8116 23530 8168 23536
rect 8128 22250 8156 23530
rect 8220 22778 8248 24550
rect 8482 24511 8538 24520
rect 8496 24410 8524 24511
rect 8484 24404 8536 24410
rect 8484 24346 8536 24352
rect 8300 23520 8352 23526
rect 8300 23462 8352 23468
rect 8312 23322 8340 23462
rect 8300 23316 8352 23322
rect 8300 23258 8352 23264
rect 8208 22772 8260 22778
rect 8208 22714 8260 22720
rect 8864 22642 8892 27520
rect 9416 24857 9444 27520
rect 9968 25498 9996 27520
rect 10520 25786 10548 27520
rect 10060 25758 10548 25786
rect 9956 25492 10008 25498
rect 9956 25434 10008 25440
rect 9402 24848 9458 24857
rect 9220 24812 9272 24818
rect 9402 24783 9458 24792
rect 9772 24812 9824 24818
rect 9220 24754 9272 24760
rect 9772 24754 9824 24760
rect 9232 23866 9260 24754
rect 9220 23860 9272 23866
rect 9220 23802 9272 23808
rect 8852 22636 8904 22642
rect 8852 22578 8904 22584
rect 8944 22636 8996 22642
rect 8944 22578 8996 22584
rect 8760 22432 8812 22438
rect 8760 22374 8812 22380
rect 8128 22234 8340 22250
rect 8128 22228 8352 22234
rect 8128 22222 8300 22228
rect 8300 22170 8352 22176
rect 8772 22137 8800 22374
rect 8956 22234 8984 22578
rect 9680 22432 9732 22438
rect 9680 22374 9732 22380
rect 8944 22228 8996 22234
rect 8944 22170 8996 22176
rect 8758 22128 8814 22137
rect 9692 22114 9720 22374
rect 8758 22063 8814 22072
rect 9600 22086 9720 22114
rect 9784 22098 9812 24754
rect 10060 23610 10088 25758
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10784 25152 10836 25158
rect 10784 25094 10836 25100
rect 10796 24818 10824 25094
rect 10874 24848 10930 24857
rect 10784 24812 10836 24818
rect 10874 24783 10930 24792
rect 10968 24812 11020 24818
rect 10784 24754 10836 24760
rect 10140 24608 10192 24614
rect 10140 24550 10192 24556
rect 9968 23582 10088 23610
rect 9968 23361 9996 23582
rect 10048 23520 10100 23526
rect 10048 23462 10100 23468
rect 9954 23352 10010 23361
rect 9954 23287 10010 23296
rect 9956 22704 10008 22710
rect 9956 22646 10008 22652
rect 9772 22092 9824 22098
rect 9036 21888 9088 21894
rect 9036 21830 9088 21836
rect 9496 21888 9548 21894
rect 9496 21830 9548 21836
rect 8024 21548 8076 21554
rect 8024 21490 8076 21496
rect 7380 21412 7432 21418
rect 7380 21354 7432 21360
rect 7104 21344 7156 21350
rect 7104 21286 7156 21292
rect 8024 21344 8076 21350
rect 8024 21286 8076 21292
rect 8484 21344 8536 21350
rect 8484 21286 8536 21292
rect 7012 21004 7064 21010
rect 7012 20946 7064 20952
rect 5814 20839 5870 20848
rect 6460 20868 6512 20874
rect 5540 20810 5592 20816
rect 6460 20810 6512 20816
rect 5264 20324 5316 20330
rect 5264 20266 5316 20272
rect 5356 20256 5408 20262
rect 5356 20198 5408 20204
rect 5368 19922 5396 20198
rect 5356 19916 5408 19922
rect 5356 19858 5408 19864
rect 5368 19378 5396 19858
rect 5448 19712 5500 19718
rect 5552 19700 5580 20810
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 6274 20360 6330 20369
rect 6184 20324 6236 20330
rect 6274 20295 6330 20304
rect 6184 20266 6236 20272
rect 6196 20058 6224 20266
rect 6184 20052 6236 20058
rect 6184 19994 6236 20000
rect 6288 19718 6316 20295
rect 7024 20262 7052 20946
rect 7116 20942 7144 21286
rect 8036 21049 8064 21286
rect 8496 21146 8524 21286
rect 8484 21140 8536 21146
rect 8484 21082 8536 21088
rect 8022 21040 8078 21049
rect 7380 21004 7432 21010
rect 8022 20975 8078 20984
rect 7380 20946 7432 20952
rect 7104 20936 7156 20942
rect 7104 20878 7156 20884
rect 7392 20602 7420 20946
rect 9048 20806 9076 21830
rect 9128 21548 9180 21554
rect 9128 21490 9180 21496
rect 7748 20800 7800 20806
rect 7748 20742 7800 20748
rect 9036 20800 9088 20806
rect 9036 20742 9088 20748
rect 7380 20596 7432 20602
rect 7380 20538 7432 20544
rect 7760 20466 7788 20742
rect 9140 20602 9168 21490
rect 9128 20596 9180 20602
rect 9128 20538 9180 20544
rect 7748 20460 7800 20466
rect 7748 20402 7800 20408
rect 8482 20360 8538 20369
rect 8208 20324 8260 20330
rect 8482 20295 8538 20304
rect 8208 20266 8260 20272
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 7748 20256 7800 20262
rect 7748 20198 7800 20204
rect 7760 19718 7788 20198
rect 7932 19916 7984 19922
rect 7932 19858 7984 19864
rect 5500 19672 5580 19700
rect 6276 19712 6328 19718
rect 5448 19654 5500 19660
rect 7748 19712 7800 19718
rect 6276 19654 6328 19660
rect 7746 19680 7748 19689
rect 7800 19680 7802 19689
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5356 19372 5408 19378
rect 5356 19314 5408 19320
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 5276 18630 5304 19110
rect 5356 18964 5408 18970
rect 5356 18906 5408 18912
rect 4908 18550 5212 18578
rect 5264 18624 5316 18630
rect 5264 18566 5316 18572
rect 4528 18420 4580 18426
rect 4528 18362 4580 18368
rect 4710 18184 4766 18193
rect 4710 18119 4766 18128
rect 4724 18086 4752 18119
rect 4712 18080 4764 18086
rect 4712 18022 4764 18028
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4724 17338 4752 17614
rect 4712 17332 4764 17338
rect 4712 17274 4764 17280
rect 4724 17241 4752 17274
rect 4710 17232 4766 17241
rect 4710 17167 4766 17176
rect 4908 14793 4936 18550
rect 5170 18456 5226 18465
rect 5170 18391 5226 18400
rect 5184 18290 5212 18391
rect 5172 18284 5224 18290
rect 5172 18226 5224 18232
rect 5080 18080 5132 18086
rect 5080 18022 5132 18028
rect 5092 17649 5120 18022
rect 5184 17882 5212 18226
rect 5172 17876 5224 17882
rect 5172 17818 5224 17824
rect 5078 17640 5134 17649
rect 5078 17575 5134 17584
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 5080 16652 5132 16658
rect 5080 16594 5132 16600
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 5000 15366 5028 16526
rect 5092 16046 5120 16594
rect 5276 16590 5304 16934
rect 5264 16584 5316 16590
rect 5170 16552 5226 16561
rect 5264 16526 5316 16532
rect 5170 16487 5226 16496
rect 5184 16250 5212 16487
rect 5172 16244 5224 16250
rect 5172 16186 5224 16192
rect 5080 16040 5132 16046
rect 5080 15982 5132 15988
rect 5264 15972 5316 15978
rect 5264 15914 5316 15920
rect 5276 15706 5304 15914
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5368 15570 5396 18906
rect 5448 18896 5500 18902
rect 5448 18838 5500 18844
rect 5460 18034 5488 18838
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 6104 18086 6132 18770
rect 6092 18080 6144 18086
rect 5460 18006 5580 18034
rect 6092 18022 6144 18028
rect 5552 17814 5580 18006
rect 5540 17808 5592 17814
rect 5540 17750 5592 17756
rect 6000 17808 6052 17814
rect 6000 17750 6052 17756
rect 5540 17672 5592 17678
rect 5538 17640 5540 17649
rect 5592 17640 5594 17649
rect 5538 17575 5594 17584
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 6012 17338 6040 17750
rect 6000 17332 6052 17338
rect 6000 17274 6052 17280
rect 6012 16726 6040 17274
rect 6104 16726 6132 18022
rect 6288 17898 6316 19654
rect 7746 19615 7802 19624
rect 6918 19408 6974 19417
rect 6918 19343 6974 19352
rect 6368 19168 6420 19174
rect 6368 19110 6420 19116
rect 6380 18970 6408 19110
rect 6368 18964 6420 18970
rect 6368 18906 6420 18912
rect 6550 18864 6606 18873
rect 6550 18799 6606 18808
rect 6564 18426 6592 18799
rect 6932 18698 6960 19343
rect 7472 19236 7524 19242
rect 7472 19178 7524 19184
rect 7748 19236 7800 19242
rect 7748 19178 7800 19184
rect 7012 19168 7064 19174
rect 7484 19145 7512 19178
rect 7012 19110 7064 19116
rect 7470 19136 7526 19145
rect 7024 18902 7052 19110
rect 7470 19071 7526 19080
rect 7760 18970 7788 19178
rect 7748 18964 7800 18970
rect 7748 18906 7800 18912
rect 7012 18896 7064 18902
rect 7012 18838 7064 18844
rect 7840 18896 7892 18902
rect 7840 18838 7892 18844
rect 7380 18828 7432 18834
rect 7380 18770 7432 18776
rect 6920 18692 6972 18698
rect 6920 18634 6972 18640
rect 6644 18624 6696 18630
rect 6642 18592 6644 18601
rect 6696 18592 6698 18601
rect 6642 18527 6698 18536
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 6564 18086 6592 18362
rect 6552 18080 6604 18086
rect 6552 18022 6604 18028
rect 6196 17870 6316 17898
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 6092 16720 6144 16726
rect 6092 16662 6144 16668
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6012 16114 6040 16662
rect 6196 16572 6224 17870
rect 6656 17814 6684 18527
rect 7392 18290 7420 18770
rect 7852 18426 7880 18838
rect 7840 18420 7892 18426
rect 7840 18362 7892 18368
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7748 18148 7800 18154
rect 7748 18090 7800 18096
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 6644 17808 6696 17814
rect 6458 17776 6514 17785
rect 6644 17750 6696 17756
rect 6458 17711 6514 17720
rect 6276 16992 6328 16998
rect 6276 16934 6328 16940
rect 6288 16794 6316 16934
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 6104 16544 6224 16572
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 5356 15564 5408 15570
rect 5356 15506 5408 15512
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 4894 14784 4950 14793
rect 4894 14719 4950 14728
rect 4712 14544 4764 14550
rect 4712 14486 4764 14492
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 4526 14376 4582 14385
rect 4526 14311 4582 14320
rect 4540 14006 4568 14311
rect 4632 14074 4660 14418
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4528 14000 4580 14006
rect 4528 13942 4580 13948
rect 4724 13530 4752 14486
rect 4896 13864 4948 13870
rect 4896 13806 4948 13812
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4908 13258 4936 13806
rect 5368 13802 5396 15302
rect 5552 15144 5580 15302
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5460 15116 5580 15144
rect 5460 14890 5488 15116
rect 5448 14884 5500 14890
rect 5448 14826 5500 14832
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 5552 14550 5580 14758
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5552 13938 5580 14486
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5540 13932 5592 13938
rect 5460 13892 5540 13920
rect 5356 13796 5408 13802
rect 5356 13738 5408 13744
rect 5262 13696 5318 13705
rect 5262 13631 5318 13640
rect 5276 13530 5304 13631
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 5170 13424 5226 13433
rect 5170 13359 5226 13368
rect 4896 13252 4948 13258
rect 4896 13194 4948 13200
rect 5184 12866 5212 13359
rect 5276 12986 5304 13466
rect 5460 13326 5488 13892
rect 5540 13874 5592 13880
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 6012 13530 6040 13670
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 5184 12838 5304 12866
rect 5170 12744 5226 12753
rect 5080 12708 5132 12714
rect 5170 12679 5226 12688
rect 5080 12650 5132 12656
rect 4436 12436 4488 12442
rect 4436 12378 4488 12384
rect 4066 12271 4122 12280
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4066 12200 4122 12209
rect 4066 12135 4068 12144
rect 4120 12135 4122 12144
rect 4068 12106 4120 12112
rect 4448 11898 4476 12242
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 4172 11218 4200 11630
rect 4632 11354 4660 12174
rect 5092 11898 5120 12650
rect 5184 12646 5212 12679
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5276 12102 5304 12838
rect 5552 12832 5580 13398
rect 6000 13184 6052 13190
rect 6000 13126 6052 13132
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6012 12850 6040 13126
rect 6000 12844 6052 12850
rect 5552 12804 5672 12832
rect 5644 12442 5672 12804
rect 6000 12786 6052 12792
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5722 12336 5778 12345
rect 5722 12271 5724 12280
rect 5776 12271 5778 12280
rect 5724 12242 5776 12248
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 4896 11824 4948 11830
rect 4896 11766 4948 11772
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4908 11218 4936 11766
rect 5276 11558 5304 12038
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6104 11778 6132 16544
rect 6288 16046 6316 16730
rect 6472 16658 6500 17711
rect 6736 17060 6788 17066
rect 6736 17002 6788 17008
rect 6748 16794 6776 17002
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6460 16652 6512 16658
rect 6460 16594 6512 16600
rect 6748 16250 6776 16730
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6276 16040 6328 16046
rect 6276 15982 6328 15988
rect 6184 15632 6236 15638
rect 6184 15574 6236 15580
rect 6196 15162 6224 15574
rect 6184 15156 6236 15162
rect 6184 15098 6236 15104
rect 6748 14929 6776 16186
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 6920 15088 6972 15094
rect 6918 15056 6920 15065
rect 6972 15056 6974 15065
rect 6918 14991 6974 15000
rect 6734 14920 6790 14929
rect 6734 14855 6790 14864
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6184 14272 6236 14278
rect 6184 14214 6236 14220
rect 6196 13734 6224 14214
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6550 13696 6606 13705
rect 6196 12374 6224 13670
rect 6550 13631 6606 13640
rect 6564 13394 6592 13631
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 6184 12368 6236 12374
rect 6184 12310 6236 12316
rect 6196 11898 6224 12310
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6104 11750 6224 11778
rect 6092 11620 6144 11626
rect 6092 11562 6144 11568
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 4172 10674 4200 11154
rect 5644 11121 5672 11494
rect 6104 11354 6132 11562
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 5630 11112 5686 11121
rect 5630 11047 5686 11056
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4172 10266 4200 10610
rect 5460 10606 5488 10950
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 3988 10118 4200 10146
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 3792 9036 3844 9042
rect 3792 8978 3844 8984
rect 3896 8616 3924 9454
rect 4080 9110 4108 9998
rect 4068 9104 4120 9110
rect 4068 9046 4120 9052
rect 3974 8936 4030 8945
rect 3974 8871 3976 8880
rect 4028 8871 4030 8880
rect 3976 8842 4028 8848
rect 4080 8634 4108 9046
rect 4068 8628 4120 8634
rect 3896 8588 4016 8616
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3896 8090 3924 8434
rect 3988 8430 4016 8588
rect 4068 8570 4120 8576
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3988 8022 4016 8366
rect 4172 8022 4200 10118
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4724 8974 4752 9318
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4724 8430 4752 8910
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4526 8120 4582 8129
rect 4526 8055 4528 8064
rect 4580 8055 4582 8064
rect 4528 8026 4580 8032
rect 3976 8016 4028 8022
rect 3976 7958 4028 7964
rect 4160 8016 4212 8022
rect 4160 7958 4212 7964
rect 4066 7848 4122 7857
rect 4066 7783 4068 7792
rect 4120 7783 4122 7792
rect 4068 7754 4120 7760
rect 4172 7546 4200 7958
rect 4540 7546 4568 8026
rect 4816 7886 4844 10542
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5276 9110 5304 10066
rect 5368 9178 5396 10066
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5264 9104 5316 9110
rect 5264 9046 5316 9052
rect 5368 8634 5396 9114
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 4894 7984 4950 7993
rect 4894 7919 4950 7928
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4816 7410 4844 7822
rect 4908 7750 4936 7919
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6196 3505 6224 11750
rect 6380 11558 6408 13126
rect 6748 12073 6776 14758
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 6932 13841 6960 13942
rect 6918 13832 6974 13841
rect 6828 13796 6880 13802
rect 6918 13767 6974 13776
rect 6828 13738 6880 13744
rect 6840 13530 6868 13738
rect 7024 13530 7052 15642
rect 7116 14550 7144 18022
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7288 17536 7340 17542
rect 7288 17478 7340 17484
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7208 16250 7236 16390
rect 7196 16244 7248 16250
rect 7196 16186 7248 16192
rect 7104 14544 7156 14550
rect 7104 14486 7156 14492
rect 7116 14385 7144 14486
rect 7102 14376 7158 14385
rect 7208 14362 7236 16186
rect 7300 15638 7328 17478
rect 7392 17134 7420 17682
rect 7380 17128 7432 17134
rect 7656 17128 7708 17134
rect 7380 17070 7432 17076
rect 7654 17096 7656 17105
rect 7708 17096 7710 17105
rect 7654 17031 7710 17040
rect 7656 16652 7708 16658
rect 7656 16594 7708 16600
rect 7288 15632 7340 15638
rect 7288 15574 7340 15580
rect 7470 14920 7526 14929
rect 7470 14855 7526 14864
rect 7208 14334 7328 14362
rect 7102 14311 7158 14320
rect 7116 14006 7144 14311
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 7104 14000 7156 14006
rect 7104 13942 7156 13948
rect 7208 13870 7236 14214
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 7208 13326 7236 13806
rect 7300 13462 7328 14334
rect 7380 14340 7432 14346
rect 7380 14282 7432 14288
rect 7392 13938 7420 14282
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7484 13530 7512 14855
rect 7668 14618 7696 16594
rect 7760 14618 7788 18090
rect 7838 17912 7894 17921
rect 7838 17847 7894 17856
rect 7852 16658 7880 17847
rect 7840 16652 7892 16658
rect 7840 16594 7892 16600
rect 7944 16046 7972 19858
rect 8024 19712 8076 19718
rect 8024 19654 8076 19660
rect 8036 18970 8064 19654
rect 8116 19304 8168 19310
rect 8114 19272 8116 19281
rect 8168 19272 8170 19281
rect 8114 19207 8170 19216
rect 8220 19122 8248 20266
rect 8496 20058 8524 20295
rect 8484 20052 8536 20058
rect 8484 19994 8536 20000
rect 8392 19508 8444 19514
rect 8496 19496 8524 19994
rect 9404 19984 9456 19990
rect 9404 19926 9456 19932
rect 8576 19916 8628 19922
rect 8576 19858 8628 19864
rect 8444 19468 8524 19496
rect 8392 19450 8444 19456
rect 8392 19168 8444 19174
rect 8220 19116 8392 19122
rect 8588 19145 8616 19858
rect 8944 19780 8996 19786
rect 8944 19722 8996 19728
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 8220 19110 8444 19116
rect 8574 19136 8630 19145
rect 8220 19094 8432 19110
rect 8024 18964 8076 18970
rect 8024 18906 8076 18912
rect 8036 17882 8064 18906
rect 8220 18766 8248 19094
rect 8574 19071 8630 19080
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8220 18426 8248 18702
rect 8482 18592 8538 18601
rect 8482 18527 8538 18536
rect 8208 18420 8260 18426
rect 8208 18362 8260 18368
rect 8496 18290 8524 18527
rect 8588 18465 8616 19071
rect 8574 18456 8630 18465
rect 8574 18391 8630 18400
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 8392 18080 8444 18086
rect 8392 18022 8444 18028
rect 8024 17876 8076 17882
rect 8024 17818 8076 17824
rect 8404 16794 8432 18022
rect 8496 17882 8524 18226
rect 8772 18086 8800 19654
rect 8956 19242 8984 19722
rect 9416 19378 9444 19926
rect 9508 19836 9536 21830
rect 9600 21554 9628 22086
rect 9772 22034 9824 22040
rect 9680 21956 9732 21962
rect 9680 21898 9732 21904
rect 9588 21548 9640 21554
rect 9588 21490 9640 21496
rect 9692 21321 9720 21898
rect 9784 21690 9812 22034
rect 9772 21684 9824 21690
rect 9772 21626 9824 21632
rect 9862 21448 9918 21457
rect 9862 21383 9918 21392
rect 9678 21312 9734 21321
rect 9678 21247 9734 21256
rect 9876 20942 9904 21383
rect 9968 21010 9996 22646
rect 10060 22409 10088 23462
rect 10152 23322 10180 24550
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10692 24268 10744 24274
rect 10692 24210 10744 24216
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10140 23316 10192 23322
rect 10140 23258 10192 23264
rect 10704 23118 10732 24210
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 10046 22400 10102 22409
rect 10046 22335 10102 22344
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10704 22098 10732 23054
rect 10796 22642 10824 23462
rect 10784 22636 10836 22642
rect 10784 22578 10836 22584
rect 10692 22092 10744 22098
rect 10692 22034 10744 22040
rect 10888 21554 10916 24783
rect 10968 24754 11020 24760
rect 10980 24342 11008 24754
rect 10968 24336 11020 24342
rect 10968 24278 11020 24284
rect 10980 23866 11008 24278
rect 10968 23860 11020 23866
rect 10968 23802 11020 23808
rect 10980 23322 11008 23802
rect 10968 23316 11020 23322
rect 10968 23258 11020 23264
rect 10968 22976 11020 22982
rect 10968 22918 11020 22924
rect 10980 22642 11008 22918
rect 10968 22636 11020 22642
rect 10968 22578 11020 22584
rect 10980 22166 11008 22578
rect 10968 22160 11020 22166
rect 10968 22102 11020 22108
rect 10968 22024 11020 22030
rect 10968 21966 11020 21972
rect 10876 21548 10928 21554
rect 10876 21490 10928 21496
rect 10692 21344 10744 21350
rect 10692 21286 10744 21292
rect 10876 21344 10928 21350
rect 10876 21286 10928 21292
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 9956 21004 10008 21010
rect 9956 20946 10008 20952
rect 9864 20936 9916 20942
rect 9864 20878 9916 20884
rect 9588 20800 9640 20806
rect 9640 20748 9812 20754
rect 9588 20742 9812 20748
rect 9600 20726 9812 20742
rect 9680 20256 9732 20262
rect 9680 20198 9732 20204
rect 9692 19961 9720 20198
rect 9784 20058 9812 20726
rect 9968 20602 9996 20946
rect 10598 20904 10654 20913
rect 10598 20839 10654 20848
rect 10612 20806 10640 20839
rect 10600 20800 10652 20806
rect 10600 20742 10652 20748
rect 9956 20596 10008 20602
rect 9956 20538 10008 20544
rect 10612 20346 10640 20742
rect 10704 20466 10732 21286
rect 10888 20806 10916 21286
rect 10980 21010 11008 21966
rect 10968 21004 11020 21010
rect 10968 20946 11020 20952
rect 10876 20800 10928 20806
rect 10876 20742 10928 20748
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10980 20466 11008 20742
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10968 20460 11020 20466
rect 10968 20402 11020 20408
rect 10140 20324 10192 20330
rect 10612 20318 10732 20346
rect 10140 20266 10192 20272
rect 9772 20052 9824 20058
rect 9772 19994 9824 20000
rect 9678 19952 9734 19961
rect 9678 19887 9734 19896
rect 9680 19848 9732 19854
rect 9508 19808 9680 19836
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 9508 19281 9536 19808
rect 9680 19790 9732 19796
rect 10152 19378 10180 20266
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10140 19372 10192 19378
rect 10140 19314 10192 19320
rect 9494 19272 9550 19281
rect 8944 19236 8996 19242
rect 9494 19207 9550 19216
rect 9862 19272 9918 19281
rect 9862 19207 9918 19216
rect 8944 19178 8996 19184
rect 8956 18970 8984 19178
rect 9772 19168 9824 19174
rect 9772 19110 9824 19116
rect 8944 18964 8996 18970
rect 8944 18906 8996 18912
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 9232 18222 9260 18566
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9220 18216 9272 18222
rect 9220 18158 9272 18164
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 8484 17876 8536 17882
rect 8484 17818 8536 17824
rect 8772 17785 8800 18022
rect 8758 17776 8814 17785
rect 8758 17711 8814 17720
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 8758 17640 8814 17649
rect 8484 17264 8536 17270
rect 8482 17232 8484 17241
rect 8536 17232 8538 17241
rect 8482 17167 8538 17176
rect 8588 16794 8616 17614
rect 9692 17626 9720 18226
rect 9784 18222 9812 19110
rect 9772 18216 9824 18222
rect 9772 18158 9824 18164
rect 8758 17575 8814 17584
rect 9508 17598 9720 17626
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8772 16658 8800 17575
rect 9508 17105 9536 17598
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9494 17096 9550 17105
rect 9494 17031 9550 17040
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8760 16652 8812 16658
rect 8760 16594 8812 16600
rect 9036 16652 9088 16658
rect 9036 16594 9088 16600
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 7932 16040 7984 16046
rect 7932 15982 7984 15988
rect 8128 15910 8156 16526
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 8128 15570 8156 15846
rect 8220 15706 8248 16594
rect 9048 16561 9076 16594
rect 9220 16584 9272 16590
rect 9034 16552 9090 16561
rect 8956 16510 9034 16538
rect 8484 15972 8536 15978
rect 8484 15914 8536 15920
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 7932 15564 7984 15570
rect 8116 15564 8168 15570
rect 7984 15524 8064 15552
rect 7932 15506 7984 15512
rect 8036 15065 8064 15524
rect 8116 15506 8168 15512
rect 8022 15056 8078 15065
rect 8022 14991 8024 15000
rect 8076 14991 8078 15000
rect 8024 14962 8076 14968
rect 7932 14952 7984 14958
rect 7932 14894 7984 14900
rect 7944 14822 7972 14894
rect 8128 14890 8156 15506
rect 8116 14884 8168 14890
rect 8116 14826 8168 14832
rect 7932 14816 7984 14822
rect 7932 14758 7984 14764
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 7564 14272 7616 14278
rect 7564 14214 7616 14220
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7288 13456 7340 13462
rect 7288 13398 7340 13404
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 7300 12918 7328 13398
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 7288 12912 7340 12918
rect 7288 12854 7340 12860
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6840 12322 6868 12718
rect 6920 12368 6972 12374
rect 6840 12316 6920 12322
rect 6840 12310 6972 12316
rect 6840 12294 6960 12310
rect 6734 12064 6790 12073
rect 6734 11999 6790 12008
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6380 11354 6408 11494
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6472 10674 6500 10950
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 6472 9926 6500 10610
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6826 10568 6882 10577
rect 6564 10470 6592 10542
rect 6736 10532 6788 10538
rect 6826 10503 6882 10512
rect 6736 10474 6788 10480
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6472 9042 6500 9862
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 6472 8634 6500 8978
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6564 8090 6592 10406
rect 6748 9722 6776 10474
rect 6840 10470 6868 10503
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 7024 9450 7052 12854
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7300 12442 7328 12718
rect 7484 12646 7512 13466
rect 7576 13326 7604 14214
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7576 12986 7604 13262
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7116 11694 7144 12038
rect 7300 11914 7328 12378
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 7208 11898 7328 11914
rect 7196 11892 7328 11898
rect 7248 11886 7328 11892
rect 7196 11834 7248 11840
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7300 11354 7328 11886
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7576 11082 7604 12242
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7576 10266 7604 11018
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7300 9926 7328 10066
rect 7668 9994 7696 13670
rect 7760 13530 7788 14554
rect 7944 14414 7972 14758
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 8206 14104 8262 14113
rect 8206 14039 8262 14048
rect 7840 14000 7892 14006
rect 7840 13942 7892 13948
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7748 12708 7800 12714
rect 7748 12650 7800 12656
rect 7760 12102 7788 12650
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7760 11898 7788 12038
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7852 11830 7880 13942
rect 7840 11824 7892 11830
rect 7840 11766 7892 11772
rect 8024 11348 8076 11354
rect 8024 11290 8076 11296
rect 8036 11257 8064 11290
rect 8022 11248 8078 11257
rect 8022 11183 8078 11192
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8128 10810 8156 11086
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8220 10266 8248 14039
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8404 12986 8432 13670
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8404 10266 8432 10406
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 7656 9988 7708 9994
rect 7656 9930 7708 9936
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7300 9586 7328 9862
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7852 9518 7880 10066
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 7840 9512 7892 9518
rect 7838 9480 7840 9489
rect 7892 9480 7894 9489
rect 7012 9444 7064 9450
rect 7838 9415 7894 9424
rect 7012 9386 7064 9392
rect 8036 9178 8064 9998
rect 8220 9722 8248 10202
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 7012 9104 7064 9110
rect 7012 9046 7064 9052
rect 7024 8634 7052 9046
rect 8036 8634 8064 9114
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7668 8090 7696 8434
rect 8036 8362 8064 8570
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 8496 4049 8524 15914
rect 8850 14376 8906 14385
rect 8850 14311 8906 14320
rect 8864 14074 8892 14311
rect 8852 14068 8904 14074
rect 8852 14010 8904 14016
rect 8864 13938 8892 14010
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 8864 13530 8892 13874
rect 8956 13530 8984 16510
rect 9220 16526 9272 16532
rect 9034 16487 9090 16496
rect 9232 15638 9260 16526
rect 9312 15904 9364 15910
rect 9312 15846 9364 15852
rect 9220 15632 9272 15638
rect 9220 15574 9272 15580
rect 9324 15450 9352 15846
rect 9232 15422 9352 15450
rect 9508 15434 9536 17031
rect 9692 15570 9720 17478
rect 9680 15564 9732 15570
rect 9600 15524 9680 15552
rect 9496 15428 9548 15434
rect 9034 15328 9090 15337
rect 9034 15263 9090 15272
rect 9048 14618 9076 15263
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 9232 14482 9260 15422
rect 9496 15370 9548 15376
rect 9600 14498 9628 15524
rect 9680 15506 9732 15512
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 9416 14470 9628 14498
rect 9036 14408 9088 14414
rect 9036 14350 9088 14356
rect 9048 14249 9076 14350
rect 9128 14272 9180 14278
rect 9034 14240 9090 14249
rect 9128 14214 9180 14220
rect 9034 14175 9090 14184
rect 9048 13938 9076 14175
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 9140 13705 9168 14214
rect 9126 13696 9182 13705
rect 9126 13631 9182 13640
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8944 13524 8996 13530
rect 8944 13466 8996 13472
rect 8668 12912 8720 12918
rect 8666 12880 8668 12889
rect 8720 12880 8722 12889
rect 8666 12815 8722 12824
rect 8864 12306 8892 13466
rect 9232 12442 9260 14418
rect 9416 13530 9444 14470
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9586 13968 9642 13977
rect 9586 13903 9642 13912
rect 9600 13841 9628 13903
rect 9586 13832 9642 13841
rect 9586 13767 9642 13776
rect 9692 13530 9720 14350
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9324 12986 9352 13262
rect 9692 12986 9720 13466
rect 9784 13258 9812 18158
rect 9876 17814 9904 19207
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 9954 18864 10010 18873
rect 9954 18799 9956 18808
rect 10008 18799 10010 18808
rect 9956 18770 10008 18776
rect 9968 18426 9996 18770
rect 10140 18760 10192 18766
rect 10138 18728 10140 18737
rect 10192 18728 10194 18737
rect 10138 18663 10194 18672
rect 10140 18624 10192 18630
rect 10140 18566 10192 18572
rect 9956 18420 10008 18426
rect 9956 18362 10008 18368
rect 10152 18086 10180 18566
rect 9956 18080 10008 18086
rect 9956 18022 10008 18028
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 9864 17808 9916 17814
rect 9864 17750 9916 17756
rect 9876 17202 9904 17750
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9968 16697 9996 18022
rect 10152 17921 10180 18022
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10138 17912 10194 17921
rect 10289 17904 10585 17924
rect 10138 17847 10194 17856
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 10060 16794 10088 17682
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 10232 17672 10284 17678
rect 10232 17614 10284 17620
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 9954 16688 10010 16697
rect 9954 16623 10010 16632
rect 10152 16250 10180 17614
rect 10244 17338 10272 17614
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10704 16658 10732 20318
rect 10980 19990 11008 20402
rect 11072 20369 11100 27520
rect 11716 24857 11744 27520
rect 11702 24848 11758 24857
rect 11702 24783 11758 24792
rect 11980 24064 12032 24070
rect 11610 24032 11666 24041
rect 11980 24006 12032 24012
rect 11610 23967 11666 23976
rect 11428 23724 11480 23730
rect 11428 23666 11480 23672
rect 11440 23254 11468 23666
rect 11428 23248 11480 23254
rect 11428 23190 11480 23196
rect 11440 22778 11468 23190
rect 11428 22772 11480 22778
rect 11428 22714 11480 22720
rect 11520 22160 11572 22166
rect 11520 22102 11572 22108
rect 11152 21888 11204 21894
rect 11152 21830 11204 21836
rect 11164 21554 11192 21830
rect 11532 21690 11560 22102
rect 11520 21684 11572 21690
rect 11520 21626 11572 21632
rect 11152 21548 11204 21554
rect 11152 21490 11204 21496
rect 11164 21078 11192 21490
rect 11152 21072 11204 21078
rect 11152 21014 11204 21020
rect 11164 20602 11192 21014
rect 11152 20596 11204 20602
rect 11152 20538 11204 20544
rect 11058 20360 11114 20369
rect 11058 20295 11114 20304
rect 10968 19984 11020 19990
rect 10968 19926 11020 19932
rect 10980 19514 11008 19926
rect 11334 19680 11390 19689
rect 11334 19615 11390 19624
rect 10968 19508 11020 19514
rect 10968 19450 11020 19456
rect 11348 19310 11376 19615
rect 11336 19304 11388 19310
rect 11336 19246 11388 19252
rect 11348 18970 11376 19246
rect 11336 18964 11388 18970
rect 11336 18906 11388 18912
rect 11428 18828 11480 18834
rect 11428 18770 11480 18776
rect 11440 18465 11468 18770
rect 11426 18456 11482 18465
rect 11426 18391 11428 18400
rect 11480 18391 11482 18400
rect 11428 18362 11480 18368
rect 10876 17536 10928 17542
rect 10874 17504 10876 17513
rect 10928 17504 10930 17513
rect 10874 17439 10930 17448
rect 11242 17504 11298 17513
rect 11242 17439 11298 17448
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10692 16652 10744 16658
rect 10692 16594 10744 16600
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 9864 15496 9916 15502
rect 9862 15464 9864 15473
rect 9916 15464 9918 15473
rect 9862 15399 9918 15408
rect 10704 15366 10732 16594
rect 10796 16590 10824 17002
rect 10784 16584 10836 16590
rect 10784 16526 10836 16532
rect 11256 16114 11284 17439
rect 11440 16726 11468 18362
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 11532 17338 11560 17682
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11624 16946 11652 23967
rect 11992 23730 12020 24006
rect 12268 23798 12296 27520
rect 12820 24818 12848 27520
rect 12808 24812 12860 24818
rect 12808 24754 12860 24760
rect 13084 24812 13136 24818
rect 13084 24754 13136 24760
rect 12532 24608 12584 24614
rect 12532 24550 12584 24556
rect 12544 24070 12572 24550
rect 12532 24064 12584 24070
rect 12530 24032 12532 24041
rect 12584 24032 12586 24041
rect 12530 23967 12586 23976
rect 12256 23792 12308 23798
rect 12256 23734 12308 23740
rect 11980 23724 12032 23730
rect 11980 23666 12032 23672
rect 12440 23656 12492 23662
rect 12440 23598 12492 23604
rect 12452 23526 12480 23598
rect 13096 23594 13124 24754
rect 13268 24200 13320 24206
rect 13268 24142 13320 24148
rect 13084 23588 13136 23594
rect 13084 23530 13136 23536
rect 11980 23520 12032 23526
rect 11980 23462 12032 23468
rect 12440 23520 12492 23526
rect 12440 23462 12492 23468
rect 11992 19310 12020 23462
rect 12452 23186 12480 23462
rect 13280 23322 13308 24142
rect 13268 23316 13320 23322
rect 13268 23258 13320 23264
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12452 22114 12480 23122
rect 12900 22976 12952 22982
rect 12900 22918 12952 22924
rect 12716 22636 12768 22642
rect 12716 22578 12768 22584
rect 12728 22545 12756 22578
rect 12912 22574 12940 22918
rect 13280 22778 13308 23258
rect 13268 22772 13320 22778
rect 13268 22714 13320 22720
rect 12900 22568 12952 22574
rect 12714 22536 12770 22545
rect 12900 22510 12952 22516
rect 12714 22471 12770 22480
rect 12360 22098 12480 22114
rect 12348 22092 12480 22098
rect 12400 22086 12480 22092
rect 12348 22034 12400 22040
rect 12360 21690 12388 22034
rect 13372 22030 13400 27520
rect 13820 23656 13872 23662
rect 13542 23624 13598 23633
rect 13820 23598 13872 23604
rect 13542 23559 13598 23568
rect 13450 23488 13506 23497
rect 13450 23423 13506 23432
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13084 21888 13136 21894
rect 13084 21830 13136 21836
rect 12348 21684 12400 21690
rect 12348 21626 12400 21632
rect 13096 21486 13124 21830
rect 13084 21480 13136 21486
rect 13084 21422 13136 21428
rect 12808 21412 12860 21418
rect 12808 21354 12860 21360
rect 12164 21344 12216 21350
rect 12164 21286 12216 21292
rect 11980 19304 12032 19310
rect 11980 19246 12032 19252
rect 12176 19174 12204 21286
rect 12440 19916 12492 19922
rect 12440 19858 12492 19864
rect 12452 19802 12480 19858
rect 12360 19774 12480 19802
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12164 19168 12216 19174
rect 12164 19110 12216 19116
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 11808 18426 11836 18770
rect 11980 18760 12032 18766
rect 11980 18702 12032 18708
rect 11796 18420 11848 18426
rect 11796 18362 11848 18368
rect 11992 18358 12020 18702
rect 11980 18352 12032 18358
rect 11980 18294 12032 18300
rect 12176 18222 12204 19110
rect 12360 18970 12388 19774
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 12452 19378 12480 19654
rect 12544 19514 12572 19790
rect 12532 19508 12584 19514
rect 12532 19450 12584 19456
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12348 18964 12400 18970
rect 12348 18906 12400 18912
rect 12452 18766 12480 19314
rect 12544 19242 12572 19450
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 12532 19236 12584 19242
rect 12532 19178 12584 19184
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 12164 18216 12216 18222
rect 12164 18158 12216 18164
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11716 17814 11744 18022
rect 11704 17808 11756 17814
rect 11704 17750 11756 17756
rect 12176 17338 12204 18158
rect 12360 18068 12388 18362
rect 12360 18040 12480 18068
rect 12452 17882 12480 18040
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12636 17610 12664 18566
rect 12624 17604 12676 17610
rect 12624 17546 12676 17552
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 11532 16918 11652 16946
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 11428 16720 11480 16726
rect 11428 16662 11480 16668
rect 11336 16516 11388 16522
rect 11336 16458 11388 16464
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 10966 15872 11022 15881
rect 10966 15807 11022 15816
rect 10980 15706 11008 15807
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 11348 15570 11376 16458
rect 11440 16250 11468 16662
rect 11428 16244 11480 16250
rect 11428 16186 11480 16192
rect 11532 16046 11560 16918
rect 11610 16824 11666 16833
rect 11610 16759 11612 16768
rect 11664 16759 11666 16768
rect 12256 16788 12308 16794
rect 11612 16730 11664 16736
rect 12256 16730 12308 16736
rect 11624 16114 11652 16730
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 11520 16040 11572 16046
rect 11440 16000 11520 16028
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 10874 15464 10930 15473
rect 10874 15399 10876 15408
rect 10928 15399 10930 15408
rect 11150 15464 11206 15473
rect 11150 15399 11206 15408
rect 10876 15370 10928 15376
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10048 14884 10100 14890
rect 10048 14826 10100 14832
rect 10060 14793 10088 14826
rect 10140 14816 10192 14822
rect 10046 14784 10102 14793
rect 10140 14758 10192 14764
rect 10046 14719 10102 14728
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9968 14074 9996 14418
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 9772 13252 9824 13258
rect 9772 13194 9824 13200
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 8852 12300 8904 12306
rect 8852 12242 8904 12248
rect 8864 11898 8892 12242
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 8852 11892 8904 11898
rect 8852 11834 8904 11840
rect 9140 11830 9168 12174
rect 9588 12164 9640 12170
rect 9588 12106 9640 12112
rect 9128 11824 9180 11830
rect 9128 11766 9180 11772
rect 9404 11688 9456 11694
rect 9456 11648 9536 11676
rect 9404 11630 9456 11636
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 8772 10198 8800 11154
rect 8956 10810 8984 11290
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 9508 10554 9536 11648
rect 9600 11626 9628 12106
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9600 11082 9628 11562
rect 9692 11354 9720 12038
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9876 11218 9904 13942
rect 9968 12374 9996 14010
rect 10152 13512 10180 14758
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10704 14521 10732 15302
rect 11164 14958 11192 15399
rect 11348 15337 11376 15506
rect 11334 15328 11390 15337
rect 11334 15263 11390 15272
rect 11152 14952 11204 14958
rect 11152 14894 11204 14900
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 10690 14512 10746 14521
rect 10690 14447 10746 14456
rect 10968 14340 11020 14346
rect 10968 14282 11020 14288
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10244 14074 10272 14214
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10704 13870 10732 14214
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10152 13484 10272 13512
rect 10244 13326 10272 13484
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10244 12986 10272 13262
rect 10704 12986 10732 13670
rect 10784 13184 10836 13190
rect 10782 13152 10784 13161
rect 10836 13152 10838 13161
rect 10782 13087 10838 13096
rect 10888 12986 10916 14010
rect 10980 13938 11008 14282
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 10232 12980 10284 12986
rect 10232 12922 10284 12928
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 11072 12850 11100 14758
rect 11152 14544 11204 14550
rect 11152 14486 11204 14492
rect 11334 14512 11390 14521
rect 11164 13161 11192 14486
rect 11334 14447 11390 14456
rect 11244 14408 11296 14414
rect 11348 14396 11376 14447
rect 11296 14368 11376 14396
rect 11244 14350 11296 14356
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11256 13784 11284 14214
rect 11348 14074 11376 14368
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11336 13796 11388 13802
rect 11256 13756 11336 13784
rect 11336 13738 11388 13744
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11150 13152 11206 13161
rect 11150 13087 11206 13096
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 10784 12708 10836 12714
rect 10784 12650 10836 12656
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 9956 12368 10008 12374
rect 9956 12310 10008 12316
rect 9954 12064 10010 12073
rect 9954 11999 10010 12008
rect 9968 11286 9996 11999
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 9956 11280 10008 11286
rect 9956 11222 10008 11228
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9588 11076 9640 11082
rect 9588 11018 9640 11024
rect 9692 10826 9720 11154
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9600 10810 9720 10826
rect 9588 10804 9720 10810
rect 9640 10798 9720 10804
rect 9588 10746 9640 10752
rect 9784 10674 9812 11086
rect 10140 11076 10192 11082
rect 10140 11018 10192 11024
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 9680 10600 9732 10606
rect 9508 10548 9680 10554
rect 9508 10542 9732 10548
rect 9508 10526 9720 10542
rect 8760 10192 8812 10198
rect 8760 10134 8812 10140
rect 9508 9518 9536 10526
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9678 10024 9734 10033
rect 9678 9959 9680 9968
rect 9732 9959 9734 9968
rect 9772 9988 9824 9994
rect 9680 9930 9732 9936
rect 9772 9930 9824 9936
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 8680 9110 8708 9454
rect 8944 9444 8996 9450
rect 8944 9386 8996 9392
rect 8956 9178 8984 9386
rect 9784 9194 9812 9930
rect 9600 9178 9812 9194
rect 9876 9178 9904 10134
rect 10060 9722 10088 10202
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 10152 9382 10180 11018
rect 10704 10606 10732 11494
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10692 9648 10744 9654
rect 10692 9590 10744 9596
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 9588 9172 9812 9178
rect 9640 9166 9812 9172
rect 9864 9172 9916 9178
rect 9588 9114 9640 9120
rect 9864 9114 9916 9120
rect 8668 9104 8720 9110
rect 8668 9046 8720 9052
rect 8956 8634 8984 9114
rect 10152 9058 10180 9318
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10048 9036 10100 9042
rect 10152 9030 10272 9058
rect 10048 8978 10100 8984
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 9692 8566 9720 8910
rect 9680 8560 9732 8566
rect 9678 8528 9680 8537
rect 9732 8528 9734 8537
rect 10060 8498 10088 8978
rect 10244 8974 10272 9030
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10612 8634 10640 8910
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 9678 8463 9734 8472
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 10060 8090 10088 8434
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 7010 4040 7066 4049
rect 7010 3975 7066 3984
rect 8482 4040 8538 4049
rect 8482 3975 8538 3984
rect 6182 3496 6238 3505
rect 6182 3431 6238 3440
rect 3606 3360 3662 3369
rect 3606 3295 3662 3304
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 3238 2680 3294 2689
rect 3238 2615 3294 2624
rect 3422 2544 3478 2553
rect 3422 2479 3478 2488
rect 3436 1465 3464 2479
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 3422 1456 3478 1465
rect 3422 1391 3478 1400
rect 3514 1184 3570 1193
rect 3514 1119 3570 1128
rect 3528 377 3556 1119
rect 7024 480 7052 3975
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10704 1193 10732 9590
rect 10796 2553 10824 12650
rect 11072 12442 11100 12786
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10888 11354 10916 12242
rect 11256 12102 11284 13262
rect 11348 13190 11376 13738
rect 11336 13184 11388 13190
rect 11336 13126 11388 13132
rect 11348 12850 11376 13126
rect 11440 12918 11468 16000
rect 11520 15982 11572 15988
rect 11900 15706 11928 16390
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11900 15162 11928 15438
rect 12268 15366 12296 16730
rect 12452 16046 12480 16934
rect 12532 16108 12584 16114
rect 12532 16050 12584 16056
rect 12440 16040 12492 16046
rect 12544 16017 12572 16050
rect 12440 15982 12492 15988
rect 12530 16008 12586 16017
rect 12452 15881 12480 15982
rect 12530 15943 12586 15952
rect 12438 15872 12494 15881
rect 12438 15807 12494 15816
rect 12348 15700 12400 15706
rect 12348 15642 12400 15648
rect 12360 15450 12388 15642
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12360 15422 12480 15450
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 12452 15162 12480 15422
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12438 15056 12494 15065
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11796 15020 11848 15026
rect 12636 15042 12664 15506
rect 12494 15014 12664 15042
rect 12438 14991 12494 15000
rect 11796 14962 11848 14968
rect 11520 14952 11572 14958
rect 11520 14894 11572 14900
rect 11428 12912 11480 12918
rect 11428 12854 11480 12860
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 11348 12374 11376 12786
rect 11336 12368 11388 12374
rect 11336 12310 11388 12316
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 11072 11218 11100 12038
rect 11348 11898 11376 12174
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11348 11370 11376 11834
rect 11256 11342 11376 11370
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 11072 10538 11100 11154
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 11072 10266 11100 10474
rect 11256 10266 11284 11342
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11348 10470 11376 11154
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11256 9382 11284 10066
rect 11532 9654 11560 14894
rect 11716 13394 11744 14962
rect 11808 14618 11836 14962
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 11796 14612 11848 14618
rect 11796 14554 11848 14560
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11716 13002 11744 13330
rect 11716 12974 11836 13002
rect 11808 12646 11836 12974
rect 11796 12640 11848 12646
rect 11794 12608 11796 12617
rect 11848 12608 11850 12617
rect 11794 12543 11850 12552
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11624 12345 11652 12378
rect 11610 12336 11666 12345
rect 11610 12271 11666 12280
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 11992 11558 12020 12242
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11702 11112 11758 11121
rect 11702 11047 11758 11056
rect 11716 10062 11744 11047
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11992 10062 12020 10406
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11716 9722 11744 9998
rect 11992 9722 12020 9998
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11980 9716 12032 9722
rect 11980 9658 12032 9664
rect 11520 9648 11572 9654
rect 11520 9590 11572 9596
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11072 8401 11100 9318
rect 11058 8392 11114 8401
rect 11058 8327 11114 8336
rect 10782 2544 10838 2553
rect 10782 2479 10838 2488
rect 12176 2417 12204 14758
rect 12348 14544 12400 14550
rect 12348 14486 12400 14492
rect 12360 14074 12388 14486
rect 12452 14346 12480 14991
rect 12728 14890 12756 19246
rect 12820 18329 12848 21354
rect 13096 21146 13124 21422
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 13174 21040 13230 21049
rect 13174 20975 13230 20984
rect 13188 20806 13216 20975
rect 13176 20800 13228 20806
rect 13176 20742 13228 20748
rect 13188 20262 13216 20742
rect 13176 20256 13228 20262
rect 13176 20198 13228 20204
rect 12900 19712 12952 19718
rect 12900 19654 12952 19660
rect 12912 18873 12940 19654
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 13004 18970 13032 19110
rect 12992 18964 13044 18970
rect 12992 18906 13044 18912
rect 12898 18864 12954 18873
rect 12898 18799 12954 18808
rect 12806 18320 12862 18329
rect 12806 18255 12862 18264
rect 12808 18080 12860 18086
rect 12806 18048 12808 18057
rect 12860 18048 12862 18057
rect 12806 17983 12862 17992
rect 13188 16998 13216 20198
rect 13464 18970 13492 23423
rect 13556 19938 13584 23559
rect 13832 23474 13860 23598
rect 13648 23446 13860 23474
rect 13648 23050 13676 23446
rect 13728 23112 13780 23118
rect 13728 23054 13780 23060
rect 13636 23044 13688 23050
rect 13636 22986 13688 22992
rect 13648 22778 13676 22986
rect 13636 22772 13688 22778
rect 13636 22714 13688 22720
rect 13740 22234 13768 23054
rect 13728 22228 13780 22234
rect 13728 22170 13780 22176
rect 13924 22114 13952 27520
rect 14188 24268 14240 24274
rect 14188 24210 14240 24216
rect 14200 23526 14228 24210
rect 14188 23520 14240 23526
rect 14568 23497 14596 27520
rect 15120 25242 15148 27520
rect 14844 25214 15148 25242
rect 14648 24064 14700 24070
rect 14648 24006 14700 24012
rect 14660 23730 14688 24006
rect 14648 23724 14700 23730
rect 14648 23666 14700 23672
rect 14188 23462 14240 23468
rect 14554 23488 14610 23497
rect 14096 22976 14148 22982
rect 14096 22918 14148 22924
rect 14108 22438 14136 22918
rect 14096 22432 14148 22438
rect 14096 22374 14148 22380
rect 13648 22086 13952 22114
rect 14002 22128 14058 22137
rect 13648 20466 13676 22086
rect 14002 22063 14004 22072
rect 14056 22063 14058 22072
rect 14004 22034 14056 22040
rect 13912 22024 13964 22030
rect 13912 21966 13964 21972
rect 13924 21690 13952 21966
rect 13912 21684 13964 21690
rect 13912 21626 13964 21632
rect 14016 21570 14044 22034
rect 14108 22030 14136 22374
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 14108 21690 14136 21966
rect 14096 21684 14148 21690
rect 14096 21626 14148 21632
rect 13924 21542 14044 21570
rect 13924 21350 13952 21542
rect 13912 21344 13964 21350
rect 13912 21286 13964 21292
rect 13820 20936 13872 20942
rect 13820 20878 13872 20884
rect 13832 20618 13860 20878
rect 13740 20602 13860 20618
rect 13728 20596 13860 20602
rect 13780 20590 13860 20596
rect 13728 20538 13780 20544
rect 13636 20460 13688 20466
rect 13636 20402 13688 20408
rect 13556 19910 13768 19938
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 13556 19514 13584 19790
rect 13544 19508 13596 19514
rect 13544 19450 13596 19456
rect 13452 18964 13504 18970
rect 13452 18906 13504 18912
rect 13268 18828 13320 18834
rect 13268 18770 13320 18776
rect 13280 18057 13308 18770
rect 13360 18420 13412 18426
rect 13464 18408 13492 18906
rect 13636 18692 13688 18698
rect 13636 18634 13688 18640
rect 13412 18380 13492 18408
rect 13360 18362 13412 18368
rect 13648 18222 13676 18634
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 13636 18216 13688 18222
rect 13636 18158 13688 18164
rect 13266 18048 13322 18057
rect 13266 17983 13322 17992
rect 13372 17814 13400 18158
rect 13360 17808 13412 17814
rect 13360 17750 13412 17756
rect 13266 17504 13322 17513
rect 13266 17439 13322 17448
rect 13280 17338 13308 17439
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 13740 17134 13768 19910
rect 13924 18834 13952 21286
rect 13912 18828 13964 18834
rect 13912 18770 13964 18776
rect 13820 17536 13872 17542
rect 13820 17478 13872 17484
rect 13832 17202 13860 17478
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 13728 17128 13780 17134
rect 13728 17070 13780 17076
rect 13176 16992 13228 16998
rect 13176 16934 13228 16940
rect 13188 16726 13216 16934
rect 14200 16726 14228 23462
rect 14554 23423 14610 23432
rect 14660 23338 14688 23666
rect 14844 23633 14872 25214
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15568 24744 15620 24750
rect 15568 24686 15620 24692
rect 15580 24614 15608 24686
rect 15568 24608 15620 24614
rect 15568 24550 15620 24556
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 14830 23624 14886 23633
rect 14830 23559 14886 23568
rect 15476 23588 15528 23594
rect 15476 23530 15528 23536
rect 14568 23310 14688 23338
rect 14568 23186 14596 23310
rect 14556 23180 14608 23186
rect 14556 23122 14608 23128
rect 14568 22982 14596 23122
rect 14556 22976 14608 22982
rect 14556 22918 14608 22924
rect 14568 22506 14596 22918
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15488 22778 15516 23530
rect 15476 22772 15528 22778
rect 15476 22714 15528 22720
rect 14556 22500 14608 22506
rect 14556 22442 14608 22448
rect 14568 21486 14596 22442
rect 15580 22098 15608 24550
rect 15672 22114 15700 27520
rect 16224 24410 16252 27520
rect 16776 24800 16804 27520
rect 16500 24772 16804 24800
rect 16500 24682 16528 24772
rect 16488 24676 16540 24682
rect 16488 24618 16540 24624
rect 17420 24410 17448 27520
rect 16212 24404 16264 24410
rect 16212 24346 16264 24352
rect 17408 24404 17460 24410
rect 17408 24346 17460 24352
rect 16396 24268 16448 24274
rect 16396 24210 16448 24216
rect 17500 24268 17552 24274
rect 17500 24210 17552 24216
rect 16408 23526 16436 24210
rect 17512 23526 17540 24210
rect 17972 23746 18000 27520
rect 18524 24410 18552 27520
rect 19076 27418 19104 27520
rect 19076 27390 19196 27418
rect 19062 24712 19118 24721
rect 19062 24647 19118 24656
rect 19076 24410 19104 24647
rect 18512 24404 18564 24410
rect 18512 24346 18564 24352
rect 19064 24404 19116 24410
rect 19064 24346 19116 24352
rect 18880 24268 18932 24274
rect 18880 24210 18932 24216
rect 17880 23718 18000 23746
rect 18328 23724 18380 23730
rect 16396 23520 16448 23526
rect 16396 23462 16448 23468
rect 17500 23520 17552 23526
rect 17500 23462 17552 23468
rect 17774 23488 17830 23497
rect 16408 23254 16436 23462
rect 16396 23248 16448 23254
rect 16396 23190 16448 23196
rect 16028 23180 16080 23186
rect 16028 23122 16080 23128
rect 16580 23180 16632 23186
rect 16580 23122 16632 23128
rect 16040 22438 16068 23122
rect 16592 22438 16620 23122
rect 16028 22432 16080 22438
rect 16028 22374 16080 22380
rect 16580 22432 16632 22438
rect 16580 22374 16632 22380
rect 16856 22432 16908 22438
rect 16856 22374 16908 22380
rect 15568 22092 15620 22098
rect 15672 22086 15792 22114
rect 15568 22034 15620 22040
rect 15660 22024 15712 22030
rect 15660 21966 15712 21972
rect 14740 21888 14792 21894
rect 14740 21830 14792 21836
rect 14556 21480 14608 21486
rect 14556 21422 14608 21428
rect 14280 21004 14332 21010
rect 14280 20946 14332 20952
rect 14292 20602 14320 20946
rect 14568 20806 14596 21422
rect 14752 21418 14780 21830
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14740 21412 14792 21418
rect 14740 21354 14792 21360
rect 14752 20942 14780 21354
rect 14740 20936 14792 20942
rect 14740 20878 14792 20884
rect 14556 20800 14608 20806
rect 14556 20742 14608 20748
rect 14752 20602 14780 20878
rect 15672 20806 15700 21966
rect 14832 20800 14884 20806
rect 14832 20742 14884 20748
rect 15660 20800 15712 20806
rect 15660 20742 15712 20748
rect 14280 20596 14332 20602
rect 14280 20538 14332 20544
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14752 20058 14780 20538
rect 14844 20398 14872 20742
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14832 20392 14884 20398
rect 14832 20334 14884 20340
rect 15292 20392 15344 20398
rect 15292 20334 15344 20340
rect 15016 20324 15068 20330
rect 15016 20266 15068 20272
rect 15028 20233 15056 20266
rect 15014 20224 15070 20233
rect 15014 20159 15070 20168
rect 14740 20052 14792 20058
rect 14740 19994 14792 20000
rect 15304 19854 15332 20334
rect 15568 19916 15620 19922
rect 15568 19858 15620 19864
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14384 19378 14412 19654
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15304 19514 15332 19790
rect 15580 19514 15608 19858
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 15568 19508 15620 19514
rect 15568 19450 15620 19456
rect 14372 19372 14424 19378
rect 14372 19314 14424 19320
rect 14384 18630 14412 19314
rect 14740 19236 14792 19242
rect 14740 19178 14792 19184
rect 14372 18624 14424 18630
rect 14372 18566 14424 18572
rect 14384 17814 14412 18566
rect 14752 18426 14780 19178
rect 15580 18970 15608 19450
rect 15568 18964 15620 18970
rect 15568 18906 15620 18912
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14740 18420 14792 18426
rect 14740 18362 14792 18368
rect 15672 18193 15700 20742
rect 15658 18184 15714 18193
rect 15658 18119 15714 18128
rect 15658 18048 15714 18057
rect 15658 17983 15714 17992
rect 14372 17808 14424 17814
rect 14372 17750 14424 17756
rect 14384 17338 14412 17750
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14372 17332 14424 17338
rect 14372 17274 14424 17280
rect 14384 17134 14412 17274
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 15292 17060 15344 17066
rect 15292 17002 15344 17008
rect 13176 16720 13228 16726
rect 14188 16720 14240 16726
rect 13176 16662 13228 16668
rect 13910 16688 13966 16697
rect 13188 15473 13216 16662
rect 14188 16662 14240 16668
rect 13910 16623 13912 16632
rect 13964 16623 13966 16632
rect 13912 16594 13964 16600
rect 13268 16584 13320 16590
rect 13268 16526 13320 16532
rect 13280 15910 13308 16526
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13832 16114 13860 16390
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 13280 15570 13308 15846
rect 13648 15638 13676 15846
rect 13924 15706 13952 16594
rect 14740 16448 14792 16454
rect 14740 16390 14792 16396
rect 14752 15706 14780 16390
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 16250 15332 17002
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 14740 15700 14792 15706
rect 14740 15642 14792 15648
rect 13636 15632 13688 15638
rect 13636 15574 13688 15580
rect 14372 15632 14424 15638
rect 14372 15574 14424 15580
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 13174 15464 13230 15473
rect 13174 15399 13230 15408
rect 12990 15056 13046 15065
rect 13280 15026 13308 15506
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 12990 14991 12992 15000
rect 13044 14991 13046 15000
rect 13268 15020 13320 15026
rect 12992 14962 13044 14968
rect 13268 14962 13320 14968
rect 12716 14884 12768 14890
rect 12716 14826 12768 14832
rect 13280 14618 13308 14962
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 12348 14068 12400 14074
rect 12348 14010 12400 14016
rect 12452 13938 12480 14282
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12728 13530 12756 13806
rect 13372 13530 13400 14418
rect 13464 13530 13492 15302
rect 14384 15026 14412 15574
rect 15672 15570 15700 17983
rect 15764 15706 15792 22086
rect 16040 17649 16068 22374
rect 16302 21584 16358 21593
rect 16302 21519 16358 21528
rect 16316 21146 16344 21519
rect 16304 21140 16356 21146
rect 16304 21082 16356 21088
rect 16026 17640 16082 17649
rect 16026 17575 16082 17584
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 16224 16833 16252 16934
rect 16210 16824 16266 16833
rect 16210 16759 16266 16768
rect 16302 16144 16358 16153
rect 16592 16114 16620 22374
rect 16670 20224 16726 20233
rect 16670 20159 16726 20168
rect 16684 20058 16712 20159
rect 16672 20052 16724 20058
rect 16672 19994 16724 20000
rect 16302 16079 16358 16088
rect 16580 16108 16632 16114
rect 16316 16046 16344 16079
rect 16580 16050 16632 16056
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 15660 15564 15712 15570
rect 15660 15506 15712 15512
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15292 15360 15344 15366
rect 15292 15302 15344 15308
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15304 15065 15332 15302
rect 15290 15056 15346 15065
rect 14372 15020 14424 15026
rect 15290 14991 15346 15000
rect 14372 14962 14424 14968
rect 14096 14884 14148 14890
rect 14096 14826 14148 14832
rect 14108 14618 14136 14826
rect 14384 14618 14412 14962
rect 15396 14958 15424 15438
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 15672 14822 15700 15506
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14384 14278 14412 14554
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14462 14240 14518 14249
rect 14384 14074 14412 14214
rect 14462 14175 14518 14184
rect 14476 14074 14504 14175
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14384 13870 14412 14010
rect 15198 13968 15254 13977
rect 15198 13903 15254 13912
rect 15212 13870 15240 13903
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 14384 13462 14412 13806
rect 15198 13696 15254 13705
rect 15198 13631 15254 13640
rect 15212 13530 15240 13631
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 14372 13456 14424 13462
rect 14372 13398 14424 13404
rect 12438 13152 12494 13161
rect 12438 13087 12494 13096
rect 12452 12850 12480 13087
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 13818 12608 13874 12617
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 12268 11898 12296 12174
rect 13004 12102 13032 12582
rect 13818 12543 13874 12552
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 12808 11892 12860 11898
rect 13004 11880 13032 12038
rect 13832 11898 13860 12543
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 12860 11852 13032 11880
rect 12808 11834 12860 11840
rect 12268 11626 12296 11834
rect 12256 11620 12308 11626
rect 12256 11562 12308 11568
rect 12268 11354 12296 11562
rect 12348 11552 12400 11558
rect 12400 11500 12480 11506
rect 12348 11494 12480 11500
rect 12360 11478 12480 11494
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12452 10674 12480 11478
rect 13004 11354 13032 11852
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 13004 10810 13032 11290
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15304 9654 15332 14758
rect 15764 14618 15792 15642
rect 16488 15496 16540 15502
rect 16488 15438 16540 15444
rect 16500 15162 16528 15438
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16118 14648 16174 14657
rect 15752 14612 15804 14618
rect 16118 14583 16174 14592
rect 15752 14554 15804 14560
rect 16132 14550 16160 14583
rect 16120 14544 16172 14550
rect 16120 14486 16172 14492
rect 15844 14476 15896 14482
rect 15844 14418 15896 14424
rect 15856 13530 15884 14418
rect 15844 13524 15896 13530
rect 15844 13466 15896 13472
rect 16868 13462 16896 22374
rect 17512 14657 17540 23462
rect 17774 23423 17830 23432
rect 17684 23180 17736 23186
rect 17684 23122 17736 23128
rect 17696 22438 17724 23122
rect 17788 23050 17816 23423
rect 17880 23322 17908 23718
rect 18328 23666 18380 23672
rect 17960 23656 18012 23662
rect 17960 23598 18012 23604
rect 17868 23316 17920 23322
rect 17868 23258 17920 23264
rect 17776 23044 17828 23050
rect 17776 22986 17828 22992
rect 17684 22432 17736 22438
rect 17684 22374 17736 22380
rect 17498 14648 17554 14657
rect 17498 14583 17554 14592
rect 16856 13456 16908 13462
rect 16856 13398 16908 13404
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16684 12986 16712 13330
rect 16672 12980 16724 12986
rect 16672 12922 16724 12928
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 16210 12880 16266 12889
rect 16210 12815 16212 12824
rect 16264 12815 16266 12824
rect 16212 12786 16264 12792
rect 15936 12776 15988 12782
rect 15934 12744 15936 12753
rect 15988 12744 15990 12753
rect 15934 12679 15990 12688
rect 17052 12209 17080 12922
rect 17972 12889 18000 23598
rect 18144 23588 18196 23594
rect 18144 23530 18196 23536
rect 17958 12880 18014 12889
rect 17958 12815 18014 12824
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 17038 12200 17094 12209
rect 17038 12135 17094 12144
rect 17958 11656 18014 11665
rect 17958 11591 18014 11600
rect 17972 11218 18000 11591
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17972 10810 18000 11154
rect 17960 10804 18012 10810
rect 17960 10746 18012 10752
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 15292 9648 15344 9654
rect 15292 9590 15344 9596
rect 12162 2408 12218 2417
rect 12162 2343 12218 2352
rect 12452 1329 12480 9590
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 18064 7857 18092 12718
rect 18156 11286 18184 23530
rect 18340 12850 18368 23666
rect 18892 23594 18920 24210
rect 19168 23866 19196 27390
rect 19628 25786 19656 27520
rect 19444 25758 19656 25786
rect 19156 23860 19208 23866
rect 19156 23802 19208 23808
rect 18880 23588 18932 23594
rect 18880 23530 18932 23536
rect 19444 23497 19472 25758
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 20074 24576 20130 24585
rect 19622 24508 19918 24528
rect 20074 24511 20130 24520
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19984 23656 20036 23662
rect 19984 23598 20036 23604
rect 19430 23488 19486 23497
rect 19430 23423 19486 23432
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19432 23180 19484 23186
rect 19432 23122 19484 23128
rect 19444 22438 19472 23122
rect 19432 22432 19484 22438
rect 19432 22374 19484 22380
rect 18328 12844 18380 12850
rect 18328 12786 18380 12792
rect 18144 11280 18196 11286
rect 18144 11222 18196 11228
rect 19444 10674 19472 22374
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19996 10674 20024 23598
rect 20088 23322 20116 24511
rect 20272 23866 20300 27520
rect 20824 24721 20852 27520
rect 20810 24712 20866 24721
rect 20810 24647 20866 24656
rect 21376 24585 21404 27520
rect 21362 24576 21418 24585
rect 21362 24511 21418 24520
rect 21180 24268 21232 24274
rect 21180 24210 21232 24216
rect 20442 24032 20498 24041
rect 20442 23967 20498 23976
rect 20456 23866 20484 23967
rect 20260 23860 20312 23866
rect 20260 23802 20312 23808
rect 20444 23860 20496 23866
rect 20444 23802 20496 23808
rect 20996 23656 21048 23662
rect 20996 23598 21048 23604
rect 20076 23316 20128 23322
rect 20076 23258 20128 23264
rect 20812 23180 20864 23186
rect 20812 23122 20864 23128
rect 20824 22438 20852 23122
rect 20812 22432 20864 22438
rect 20812 22374 20864 22380
rect 20824 12345 20852 22374
rect 21008 12374 21036 23598
rect 21192 23526 21220 24210
rect 21928 24041 21956 27520
rect 22480 24410 22508 27520
rect 22468 24404 22520 24410
rect 22468 24346 22520 24352
rect 21914 24032 21970 24041
rect 21914 23967 21970 23976
rect 23124 23905 23152 27520
rect 23676 25106 23704 27520
rect 23400 25078 23704 25106
rect 21546 23896 21602 23905
rect 21546 23831 21548 23840
rect 21600 23831 21602 23840
rect 23110 23896 23166 23905
rect 23400 23866 23428 25078
rect 24228 24970 24256 27520
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 23492 24942 24256 24970
rect 23110 23831 23166 23840
rect 23388 23860 23440 23866
rect 21548 23802 21600 23808
rect 23388 23802 23440 23808
rect 22100 23656 22152 23662
rect 22020 23604 22100 23610
rect 22020 23598 22152 23604
rect 22020 23582 22140 23598
rect 21180 23520 21232 23526
rect 21180 23462 21232 23468
rect 20996 12368 21048 12374
rect 20810 12336 20866 12345
rect 20996 12310 21048 12316
rect 20810 12271 20866 12280
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20916 11558 20944 12242
rect 20904 11552 20956 11558
rect 20904 11494 20956 11500
rect 20916 11257 20944 11494
rect 20902 11248 20958 11257
rect 20902 11183 20958 11192
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 18420 10600 18472 10606
rect 19708 10600 19760 10606
rect 18420 10542 18472 10548
rect 19706 10568 19708 10577
rect 19760 10568 19762 10577
rect 18432 8945 18460 10542
rect 19706 10503 19762 10512
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 21192 10198 21220 23462
rect 22020 23254 22048 23582
rect 22008 23248 22060 23254
rect 22008 23190 22060 23196
rect 21180 10192 21232 10198
rect 21180 10134 21232 10140
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 19536 10033 19564 10066
rect 19522 10024 19578 10033
rect 19522 9959 19578 9968
rect 19536 9722 19564 9959
rect 19524 9716 19576 9722
rect 19524 9658 19576 9664
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 18418 8936 18474 8945
rect 18418 8871 18474 8880
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 23492 8106 23520 24942
rect 24780 24818 24808 27520
rect 23848 24812 23900 24818
rect 23848 24754 23900 24760
rect 24768 24812 24820 24818
rect 24768 24754 24820 24760
rect 23400 8090 23520 8106
rect 23388 8084 23520 8090
rect 23440 8078 23520 8084
rect 23388 8026 23440 8032
rect 22282 7984 22338 7993
rect 22282 7919 22284 7928
rect 22336 7919 22338 7928
rect 22284 7890 22336 7896
rect 18050 7848 18106 7857
rect 18050 7783 18106 7792
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 22296 7546 22324 7890
rect 23860 7546 23888 24754
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 25332 17218 25360 27520
rect 25976 24834 26004 27520
rect 24872 17190 25360 17218
rect 25424 24806 26004 24834
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 22284 7540 22336 7546
rect 22284 7482 22336 7488
rect 23848 7540 23900 7546
rect 23848 7482 23900 7488
rect 23662 7440 23718 7449
rect 23662 7375 23718 7384
rect 23676 7342 23704 7375
rect 23664 7336 23716 7342
rect 23664 7278 23716 7284
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24872 6474 24900 17190
rect 25424 17082 25452 24806
rect 26528 23746 26556 27520
rect 26344 23718 26556 23746
rect 26344 17218 26372 23718
rect 24780 6458 24900 6474
rect 24768 6452 24900 6458
rect 24820 6446 24900 6452
rect 24964 17054 25452 17082
rect 26252 17190 26372 17218
rect 24768 6394 24820 6400
rect 23662 6352 23718 6361
rect 23662 6287 23718 6296
rect 23676 6254 23704 6287
rect 23664 6248 23716 6254
rect 23664 6190 23716 6196
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 24964 5930 24992 17054
rect 24780 5914 24992 5930
rect 24768 5908 24992 5914
rect 24820 5902 24992 5908
rect 24768 5850 24820 5856
rect 24030 5808 24086 5817
rect 24030 5743 24032 5752
rect 24084 5743 24086 5752
rect 24032 5714 24084 5720
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 24044 5370 24072 5714
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 26252 5409 26280 17190
rect 27080 12866 27108 27520
rect 27632 14385 27660 27520
rect 27618 14376 27674 14385
rect 27618 14311 27674 14320
rect 26896 12838 27108 12866
rect 24674 5400 24730 5409
rect 24032 5364 24084 5370
rect 24674 5335 24676 5344
rect 24032 5306 24084 5312
rect 24728 5335 24730 5344
rect 26238 5400 26294 5409
rect 26238 5335 26294 5344
rect 24676 5306 24728 5312
rect 24490 5264 24546 5273
rect 24490 5199 24546 5208
rect 24504 5166 24532 5199
rect 24492 5160 24544 5166
rect 24492 5102 24544 5108
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 26896 4865 26924 12838
rect 24766 4856 24822 4865
rect 24766 4791 24768 4800
rect 24820 4791 24822 4800
rect 26882 4856 26938 4865
rect 26882 4791 26938 4800
rect 24768 4762 24820 4768
rect 24582 4720 24638 4729
rect 24582 4655 24584 4664
rect 24636 4655 24638 4664
rect 24584 4626 24636 4632
rect 24596 4570 24624 4626
rect 24596 4542 24716 4570
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24688 4282 24716 4542
rect 24676 4276 24728 4282
rect 24676 4218 24728 4224
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 20994 3496 21050 3505
rect 20994 3431 21050 3440
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 12438 1320 12494 1329
rect 12438 1255 12494 1264
rect 10690 1184 10746 1193
rect 10690 1119 10746 1128
rect 21008 480 21036 3431
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 3514 368 3570 377
rect 3514 303 3570 312
rect 7010 0 7066 480
rect 20994 0 21050 480
<< via2 >>
rect 3882 27648 3938 27704
rect 294 18808 350 18864
rect 1582 22208 1638 22264
rect 1398 20304 1454 20360
rect 1490 19916 1546 19952
rect 1490 19896 1492 19916
rect 1492 19896 1544 19916
rect 1544 19896 1546 19916
rect 1766 21120 1822 21176
rect 846 17584 902 17640
rect 1398 15988 1400 16008
rect 1400 15988 1452 16008
rect 1452 15988 1454 16008
rect 1398 15952 1454 15988
rect 1582 16632 1638 16688
rect 1490 15408 1546 15464
rect 2042 23588 2098 23624
rect 2042 23568 2044 23588
rect 2044 23568 2096 23588
rect 2096 23568 2098 23588
rect 2042 22208 2098 22264
rect 2318 22888 2374 22944
rect 2778 24656 2834 24712
rect 2686 22500 2742 22536
rect 2686 22480 2688 22500
rect 2688 22480 2740 22500
rect 2740 22480 2742 22500
rect 2594 22344 2650 22400
rect 2870 22752 2926 22808
rect 2686 21256 2742 21312
rect 3054 23976 3110 24032
rect 2962 21528 3018 21584
rect 3514 27104 3570 27160
rect 3330 25880 3386 25936
rect 4066 26444 4122 26480
rect 4066 26424 4068 26444
rect 4068 26424 4120 26444
rect 4120 26424 4122 26444
rect 4066 25200 4122 25256
rect 3238 23296 3294 23352
rect 3146 21528 3202 21584
rect 3054 20984 3110 21040
rect 2870 19760 2926 19816
rect 2318 19352 2374 19408
rect 2226 18400 2282 18456
rect 2226 18284 2282 18320
rect 2226 18264 2228 18284
rect 2228 18264 2280 18284
rect 2280 18264 2282 18284
rect 1950 17620 1952 17640
rect 1952 17620 2004 17640
rect 2004 17620 2006 17640
rect 1950 17584 2006 17620
rect 2502 17584 2558 17640
rect 2962 19080 3018 19136
rect 2870 17856 2926 17912
rect 1858 14340 1914 14376
rect 1858 14320 1860 14340
rect 1860 14320 1912 14340
rect 1912 14320 1914 14340
rect 2042 13504 2098 13560
rect 1766 12416 1822 12472
rect 3422 20304 3478 20360
rect 3422 19080 3478 19136
rect 3330 18692 3386 18728
rect 3330 18672 3332 18692
rect 3332 18672 3384 18692
rect 3384 18672 3386 18692
rect 3974 22480 4030 22536
rect 3422 18264 3478 18320
rect 3146 16224 3202 16280
rect 2962 13948 2964 13968
rect 2964 13948 3016 13968
rect 3016 13948 3018 13968
rect 2962 13912 3018 13948
rect 2410 12436 2466 12472
rect 2410 12416 2412 12436
rect 2412 12416 2464 12436
rect 2464 12416 2466 12436
rect 1398 11600 1454 11656
rect 1582 11192 1638 11248
rect 2134 10668 2190 10704
rect 2134 10648 2136 10668
rect 2136 10648 2188 10668
rect 2188 10648 2190 10668
rect 2870 12824 2926 12880
rect 2870 11872 2926 11928
rect 2502 9560 2558 9616
rect 4250 18572 4252 18592
rect 4252 18572 4304 18592
rect 4304 18572 4306 18592
rect 4250 18536 4306 18572
rect 4250 18284 4306 18320
rect 4250 18264 4252 18284
rect 4252 18264 4304 18284
rect 4304 18264 4306 18284
rect 4710 24248 4766 24304
rect 5078 23160 5134 23216
rect 4802 21972 4804 21992
rect 4804 21972 4856 21992
rect 4856 21972 4858 21992
rect 4802 21936 4858 21972
rect 4618 19116 4620 19136
rect 4620 19116 4672 19136
rect 4672 19116 4674 19136
rect 4250 17312 4306 17368
rect 3790 16088 3846 16144
rect 3882 15408 3938 15464
rect 3790 15000 3846 15056
rect 3974 14864 4030 14920
rect 3330 14456 3386 14512
rect 3238 13912 3294 13968
rect 4342 13912 4398 13968
rect 3882 13096 3938 13152
rect 2410 8064 2466 8120
rect 570 7520 626 7576
rect 570 6976 626 7032
rect 3422 7384 3478 7440
rect 3330 3848 3386 3904
rect 3790 12280 3846 12336
rect 4066 12280 4122 12336
rect 4618 19080 4674 19116
rect 5354 24520 5410 24576
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5998 24656 6054 24712
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5354 23432 5410 23488
rect 5814 23316 5870 23352
rect 5814 23296 5816 23316
rect 5816 23296 5868 23316
rect 5868 23296 5870 23316
rect 6458 24248 6514 24304
rect 6550 23976 6606 24032
rect 5354 22888 5410 22944
rect 6090 23024 6146 23080
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5262 22380 5264 22400
rect 5264 22380 5316 22400
rect 5316 22380 5318 22400
rect 5262 22344 5318 22380
rect 5446 22344 5502 22400
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 6918 23160 6974 23216
rect 7102 22616 7158 22672
rect 6826 22208 6882 22264
rect 5998 21140 6054 21176
rect 5998 21120 6000 21140
rect 6000 21120 6052 21140
rect 6052 21120 6054 21140
rect 5814 20848 5870 20904
rect 8022 24792 8078 24848
rect 7654 21936 7710 21992
rect 8206 24656 8262 24712
rect 8482 24520 8538 24576
rect 9402 24792 9458 24848
rect 8758 22072 8814 22128
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10874 24792 10930 24848
rect 9954 23296 10010 23352
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 6274 20304 6330 20360
rect 8022 20984 8078 21040
rect 8482 20304 8538 20360
rect 7746 19660 7748 19680
rect 7748 19660 7800 19680
rect 7800 19660 7802 19680
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 4710 18128 4766 18184
rect 4710 17176 4766 17232
rect 5170 18400 5226 18456
rect 5078 17584 5134 17640
rect 5170 16496 5226 16552
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5538 17620 5540 17640
rect 5540 17620 5592 17640
rect 5592 17620 5594 17640
rect 5538 17584 5594 17620
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 7746 19624 7802 19660
rect 6918 19352 6974 19408
rect 6550 18808 6606 18864
rect 7470 19080 7526 19136
rect 6642 18572 6644 18592
rect 6644 18572 6696 18592
rect 6696 18572 6698 18592
rect 6642 18536 6698 18572
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 6458 17720 6514 17776
rect 4894 14728 4950 14784
rect 4526 14320 4582 14376
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5262 13640 5318 13696
rect 5170 13368 5226 13424
rect 5170 12688 5226 12744
rect 4066 12164 4122 12200
rect 4066 12144 4068 12164
rect 4068 12144 4120 12164
rect 4120 12144 4122 12164
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5722 12300 5778 12336
rect 5722 12280 5724 12300
rect 5724 12280 5776 12300
rect 5776 12280 5778 12300
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 6918 15036 6920 15056
rect 6920 15036 6972 15056
rect 6972 15036 6974 15056
rect 6918 15000 6974 15036
rect 6734 14864 6790 14920
rect 6550 13640 6606 13696
rect 5630 11056 5686 11112
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 3974 8900 4030 8936
rect 3974 8880 3976 8900
rect 3976 8880 4028 8900
rect 4028 8880 4030 8900
rect 4526 8084 4582 8120
rect 4526 8064 4528 8084
rect 4528 8064 4580 8084
rect 4580 8064 4582 8084
rect 4066 7812 4122 7848
rect 4066 7792 4068 7812
rect 4068 7792 4120 7812
rect 4120 7792 4122 7812
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 4894 7928 4950 7984
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 6918 13776 6974 13832
rect 7102 14320 7158 14376
rect 7654 17076 7656 17096
rect 7656 17076 7708 17096
rect 7708 17076 7710 17096
rect 7654 17040 7710 17076
rect 7470 14864 7526 14920
rect 7838 17856 7894 17912
rect 8114 19252 8116 19272
rect 8116 19252 8168 19272
rect 8168 19252 8170 19272
rect 8114 19216 8170 19252
rect 8574 19080 8630 19136
rect 8482 18536 8538 18592
rect 8574 18400 8630 18456
rect 9862 21392 9918 21448
rect 9678 21256 9734 21312
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10046 22344 10102 22400
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10598 20848 10654 20904
rect 9678 19896 9734 19952
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 9494 19216 9550 19272
rect 9862 19216 9918 19272
rect 8758 17720 8814 17776
rect 8482 17212 8484 17232
rect 8484 17212 8536 17232
rect 8536 17212 8538 17232
rect 8482 17176 8538 17212
rect 8758 17584 8814 17640
rect 9494 17040 9550 17096
rect 8022 15020 8078 15056
rect 8022 15000 8024 15020
rect 8024 15000 8076 15020
rect 8076 15000 8078 15020
rect 6734 12008 6790 12064
rect 6826 10512 6882 10568
rect 8206 14048 8262 14104
rect 8022 11192 8078 11248
rect 7838 9460 7840 9480
rect 7840 9460 7892 9480
rect 7892 9460 7894 9480
rect 7838 9424 7894 9460
rect 8850 14320 8906 14376
rect 9034 16496 9090 16552
rect 9034 15272 9090 15328
rect 9034 14184 9090 14240
rect 9126 13640 9182 13696
rect 8666 12860 8668 12880
rect 8668 12860 8720 12880
rect 8720 12860 8722 12880
rect 8666 12824 8722 12860
rect 9586 13912 9642 13968
rect 9586 13776 9642 13832
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 9954 18828 10010 18864
rect 9954 18808 9956 18828
rect 9956 18808 10008 18828
rect 10008 18808 10010 18828
rect 10138 18708 10140 18728
rect 10140 18708 10192 18728
rect 10192 18708 10194 18728
rect 10138 18672 10194 18708
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10138 17856 10194 17912
rect 9954 16632 10010 16688
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 11702 24792 11758 24848
rect 11610 23976 11666 24032
rect 11058 20304 11114 20360
rect 11334 19624 11390 19680
rect 11426 18420 11482 18456
rect 11426 18400 11428 18420
rect 11428 18400 11480 18420
rect 11480 18400 11482 18420
rect 10874 17484 10876 17504
rect 10876 17484 10928 17504
rect 10928 17484 10930 17504
rect 10874 17448 10930 17484
rect 11242 17448 11298 17504
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 9862 15444 9864 15464
rect 9864 15444 9916 15464
rect 9916 15444 9918 15464
rect 9862 15408 9918 15444
rect 12530 24012 12532 24032
rect 12532 24012 12584 24032
rect 12584 24012 12586 24032
rect 12530 23976 12586 24012
rect 12714 22480 12770 22536
rect 13542 23568 13598 23624
rect 13450 23432 13506 23488
rect 10966 15816 11022 15872
rect 11610 16788 11666 16824
rect 11610 16768 11612 16788
rect 11612 16768 11664 16788
rect 11664 16768 11666 16788
rect 10874 15428 10930 15464
rect 10874 15408 10876 15428
rect 10876 15408 10928 15428
rect 10928 15408 10930 15428
rect 11150 15408 11206 15464
rect 10046 14728 10102 14784
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 11334 15272 11390 15328
rect 10690 14456 10746 14512
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10782 13132 10784 13152
rect 10784 13132 10836 13152
rect 10836 13132 10838 13152
rect 10782 13096 10838 13132
rect 11334 14456 11390 14512
rect 11150 13096 11206 13152
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 9954 12008 10010 12064
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 9678 9988 9734 10024
rect 9678 9968 9680 9988
rect 9680 9968 9732 9988
rect 9732 9968 9734 9988
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 9678 8508 9680 8528
rect 9680 8508 9732 8528
rect 9732 8508 9734 8528
rect 9678 8472 9734 8508
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 7010 3984 7066 4040
rect 8482 3984 8538 4040
rect 6182 3440 6238 3496
rect 3606 3304 3662 3360
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 3238 2624 3294 2680
rect 3422 2488 3478 2544
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 3422 1400 3478 1456
rect 3514 1128 3570 1184
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 12530 15952 12586 16008
rect 12438 15816 12494 15872
rect 12438 15000 12494 15056
rect 11794 12588 11796 12608
rect 11796 12588 11848 12608
rect 11848 12588 11850 12608
rect 11794 12552 11850 12588
rect 11610 12280 11666 12336
rect 11702 11056 11758 11112
rect 11058 8336 11114 8392
rect 10782 2488 10838 2544
rect 13174 20984 13230 21040
rect 12898 18808 12954 18864
rect 12806 18264 12862 18320
rect 12806 18028 12808 18048
rect 12808 18028 12860 18048
rect 12860 18028 12862 18048
rect 12806 17992 12862 18028
rect 14002 22092 14058 22128
rect 14002 22072 14004 22092
rect 14004 22072 14056 22092
rect 14056 22072 14058 22092
rect 13266 17992 13322 18048
rect 13266 17448 13322 17504
rect 14554 23432 14610 23488
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14830 23568 14886 23624
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 19062 24656 19118 24712
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 15014 20168 15070 20224
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 15658 18128 15714 18184
rect 15658 17992 15714 18048
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 13910 16652 13966 16688
rect 13910 16632 13912 16652
rect 13912 16632 13964 16652
rect 13964 16632 13966 16652
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 13174 15408 13230 15464
rect 12990 15020 13046 15056
rect 12990 15000 12992 15020
rect 12992 15000 13044 15020
rect 13044 15000 13046 15020
rect 16302 21528 16358 21584
rect 16026 17584 16082 17640
rect 16210 16768 16266 16824
rect 16302 16088 16358 16144
rect 16670 20168 16726 20224
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 15290 15000 15346 15056
rect 14462 14184 14518 14240
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 15198 13912 15254 13968
rect 15198 13640 15254 13696
rect 12438 13096 12494 13152
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 13818 12552 13874 12608
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 16118 14592 16174 14648
rect 17774 23432 17830 23488
rect 17498 14592 17554 14648
rect 16210 12844 16266 12880
rect 16210 12824 16212 12844
rect 16212 12824 16264 12844
rect 16264 12824 16266 12844
rect 15934 12724 15936 12744
rect 15936 12724 15988 12744
rect 15988 12724 15990 12744
rect 15934 12688 15990 12724
rect 17958 12824 18014 12880
rect 17038 12144 17094 12200
rect 17958 11600 18014 11656
rect 12162 2352 12218 2408
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 20074 24520 20130 24576
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19430 23432 19486 23488
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 20810 24656 20866 24712
rect 21362 24520 21418 24576
rect 20442 23976 20498 24032
rect 21914 23976 21970 24032
rect 21546 23860 21602 23896
rect 21546 23840 21548 23860
rect 21548 23840 21600 23860
rect 21600 23840 21602 23860
rect 23110 23840 23166 23896
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 20810 12280 20866 12336
rect 20902 11192 20958 11248
rect 19706 10548 19708 10568
rect 19708 10548 19760 10568
rect 19760 10548 19762 10568
rect 19706 10512 19762 10548
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19522 9968 19578 10024
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 18418 8880 18474 8936
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 22282 7948 22338 7984
rect 22282 7928 22284 7948
rect 22284 7928 22336 7948
rect 22336 7928 22338 7948
rect 18050 7792 18106 7848
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 23662 7384 23718 7440
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 23662 6296 23718 6352
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 24030 5772 24086 5808
rect 24030 5752 24032 5772
rect 24032 5752 24084 5772
rect 24084 5752 24086 5772
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 27618 14320 27674 14376
rect 24674 5364 24730 5400
rect 24674 5344 24676 5364
rect 24676 5344 24728 5364
rect 24728 5344 24730 5364
rect 26238 5344 26294 5400
rect 24490 5208 24546 5264
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 24766 4820 24822 4856
rect 24766 4800 24768 4820
rect 24768 4800 24820 4820
rect 24820 4800 24822 4820
rect 26882 4800 26938 4856
rect 24582 4684 24638 4720
rect 24582 4664 24584 4684
rect 24584 4664 24636 4684
rect 24636 4664 24638 4684
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 20994 3440 21050 3496
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 12438 1264 12494 1320
rect 10690 1128 10746 1184
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 3514 312 3570 368
<< metal3 >>
rect 0 27706 480 27736
rect 3877 27706 3943 27709
rect 0 27704 3943 27706
rect 0 27648 3882 27704
rect 3938 27648 3943 27704
rect 0 27646 3943 27648
rect 0 27616 480 27646
rect 3877 27643 3943 27646
rect 0 27162 480 27192
rect 3509 27162 3575 27165
rect 0 27160 3575 27162
rect 0 27104 3514 27160
rect 3570 27104 3575 27160
rect 0 27102 3575 27104
rect 0 27072 480 27102
rect 3509 27099 3575 27102
rect 0 26482 480 26512
rect 4061 26482 4127 26485
rect 0 26480 4127 26482
rect 0 26424 4066 26480
rect 4122 26424 4127 26480
rect 0 26422 4127 26424
rect 0 26392 480 26422
rect 4061 26419 4127 26422
rect 0 25938 480 25968
rect 3325 25938 3391 25941
rect 0 25936 3391 25938
rect 0 25880 3330 25936
rect 3386 25880 3391 25936
rect 0 25878 3391 25880
rect 0 25848 480 25878
rect 3325 25875 3391 25878
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25258 480 25288
rect 4061 25258 4127 25261
rect 0 25256 4127 25258
rect 0 25200 4066 25256
rect 4122 25200 4127 25256
rect 0 25198 4127 25200
rect 0 25168 480 25198
rect 4061 25195 4127 25198
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 8017 24850 8083 24853
rect 9397 24850 9463 24853
rect 8017 24848 9463 24850
rect 8017 24792 8022 24848
rect 8078 24792 9402 24848
rect 9458 24792 9463 24848
rect 8017 24790 9463 24792
rect 8017 24787 8083 24790
rect 9397 24787 9463 24790
rect 10869 24850 10935 24853
rect 11697 24850 11763 24853
rect 10869 24848 11763 24850
rect 10869 24792 10874 24848
rect 10930 24792 11702 24848
rect 11758 24792 11763 24848
rect 10869 24790 11763 24792
rect 10869 24787 10935 24790
rect 11697 24787 11763 24790
rect 0 24714 480 24744
rect 2773 24714 2839 24717
rect 0 24712 2839 24714
rect 0 24656 2778 24712
rect 2834 24656 2839 24712
rect 0 24654 2839 24656
rect 0 24624 480 24654
rect 2773 24651 2839 24654
rect 5993 24714 6059 24717
rect 8201 24714 8267 24717
rect 5993 24712 8267 24714
rect 5993 24656 5998 24712
rect 6054 24656 8206 24712
rect 8262 24656 8267 24712
rect 5993 24654 8267 24656
rect 5993 24651 6059 24654
rect 8201 24651 8267 24654
rect 19057 24714 19123 24717
rect 20805 24714 20871 24717
rect 19057 24712 20871 24714
rect 19057 24656 19062 24712
rect 19118 24656 20810 24712
rect 20866 24656 20871 24712
rect 19057 24654 20871 24656
rect 19057 24651 19123 24654
rect 20805 24651 20871 24654
rect 5349 24578 5415 24581
rect 8477 24578 8543 24581
rect 5349 24576 8543 24578
rect 5349 24520 5354 24576
rect 5410 24520 8482 24576
rect 8538 24520 8543 24576
rect 5349 24518 8543 24520
rect 5349 24515 5415 24518
rect 8477 24515 8543 24518
rect 20069 24578 20135 24581
rect 21357 24578 21423 24581
rect 20069 24576 21423 24578
rect 20069 24520 20074 24576
rect 20130 24520 21362 24576
rect 21418 24520 21423 24576
rect 20069 24518 21423 24520
rect 20069 24515 20135 24518
rect 21357 24515 21423 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 4705 24306 4771 24309
rect 6453 24306 6519 24309
rect 4705 24304 6519 24306
rect 4705 24248 4710 24304
rect 4766 24248 6458 24304
rect 6514 24248 6519 24304
rect 4705 24246 6519 24248
rect 4705 24243 4771 24246
rect 6453 24243 6519 24246
rect 0 24034 480 24064
rect 3049 24034 3115 24037
rect 0 24032 3115 24034
rect 0 23976 3054 24032
rect 3110 23976 3115 24032
rect 0 23974 3115 23976
rect 0 23944 480 23974
rect 3049 23971 3115 23974
rect 6545 24034 6611 24037
rect 11605 24034 11671 24037
rect 12525 24034 12591 24037
rect 6545 24032 12591 24034
rect 6545 23976 6550 24032
rect 6606 23976 11610 24032
rect 11666 23976 12530 24032
rect 12586 23976 12591 24032
rect 6545 23974 12591 23976
rect 6545 23971 6611 23974
rect 11605 23971 11671 23974
rect 12525 23971 12591 23974
rect 20437 24034 20503 24037
rect 21909 24034 21975 24037
rect 20437 24032 21975 24034
rect 20437 23976 20442 24032
rect 20498 23976 21914 24032
rect 21970 23976 21975 24032
rect 20437 23974 21975 23976
rect 20437 23971 20503 23974
rect 21909 23971 21975 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 21541 23898 21607 23901
rect 23105 23898 23171 23901
rect 21541 23896 23171 23898
rect 21541 23840 21546 23896
rect 21602 23840 23110 23896
rect 23166 23840 23171 23896
rect 21541 23838 23171 23840
rect 21541 23835 21607 23838
rect 23105 23835 23171 23838
rect 2037 23628 2103 23629
rect 2037 23626 2084 23628
rect 1992 23624 2084 23626
rect 1992 23568 2042 23624
rect 1992 23566 2084 23568
rect 2037 23564 2084 23566
rect 2148 23564 2154 23628
rect 13537 23626 13603 23629
rect 14825 23626 14891 23629
rect 13537 23624 14891 23626
rect 13537 23568 13542 23624
rect 13598 23568 14830 23624
rect 14886 23568 14891 23624
rect 13537 23566 14891 23568
rect 2037 23563 2103 23564
rect 13537 23563 13603 23566
rect 14825 23563 14891 23566
rect 0 23490 480 23520
rect 5349 23490 5415 23493
rect 13445 23490 13511 23493
rect 14549 23490 14615 23493
rect 0 23430 3066 23490
rect 0 23400 480 23430
rect 3006 23082 3066 23430
rect 5349 23488 6010 23490
rect 5349 23432 5354 23488
rect 5410 23432 6010 23488
rect 5349 23430 6010 23432
rect 5349 23427 5415 23430
rect 3233 23354 3299 23357
rect 5809 23354 5875 23357
rect 3233 23352 5875 23354
rect 3233 23296 3238 23352
rect 3294 23296 5814 23352
rect 5870 23296 5875 23352
rect 3233 23294 5875 23296
rect 5950 23354 6010 23430
rect 13445 23488 14615 23490
rect 13445 23432 13450 23488
rect 13506 23432 14554 23488
rect 14610 23432 14615 23488
rect 13445 23430 14615 23432
rect 13445 23427 13511 23430
rect 14549 23427 14615 23430
rect 17769 23490 17835 23493
rect 19425 23490 19491 23493
rect 17769 23488 19491 23490
rect 17769 23432 17774 23488
rect 17830 23432 19430 23488
rect 19486 23432 19491 23488
rect 17769 23430 19491 23432
rect 17769 23427 17835 23430
rect 19425 23427 19491 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 9949 23354 10015 23357
rect 5950 23352 10015 23354
rect 5950 23296 9954 23352
rect 10010 23296 10015 23352
rect 5950 23294 10015 23296
rect 3233 23291 3299 23294
rect 5809 23291 5875 23294
rect 9949 23291 10015 23294
rect 5073 23218 5139 23221
rect 6913 23218 6979 23221
rect 5073 23216 6979 23218
rect 5073 23160 5078 23216
rect 5134 23160 6918 23216
rect 6974 23160 6979 23216
rect 5073 23158 6979 23160
rect 5073 23155 5139 23158
rect 6913 23155 6979 23158
rect 6085 23082 6151 23085
rect 3006 23080 6151 23082
rect 3006 23024 6090 23080
rect 6146 23024 6151 23080
rect 3006 23022 6151 23024
rect 6085 23019 6151 23022
rect 2313 22946 2379 22949
rect 5349 22946 5415 22949
rect 2313 22944 5415 22946
rect 2313 22888 2318 22944
rect 2374 22888 5354 22944
rect 5410 22888 5415 22944
rect 2313 22886 5415 22888
rect 2313 22883 2379 22886
rect 5349 22883 5415 22886
rect 5610 22880 5930 22881
rect 0 22810 480 22840
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 2865 22810 2931 22813
rect 0 22808 2931 22810
rect 0 22752 2870 22808
rect 2926 22752 2931 22808
rect 0 22750 2931 22752
rect 0 22720 480 22750
rect 2865 22747 2931 22750
rect 7097 22674 7163 22677
rect 3742 22672 7163 22674
rect 3742 22616 7102 22672
rect 7158 22616 7163 22672
rect 3742 22614 7163 22616
rect 2681 22538 2747 22541
rect 3742 22538 3802 22614
rect 7097 22611 7163 22614
rect 2681 22536 3802 22538
rect 2681 22480 2686 22536
rect 2742 22480 3802 22536
rect 2681 22478 3802 22480
rect 3969 22538 4035 22541
rect 12709 22538 12775 22541
rect 3969 22536 12775 22538
rect 3969 22480 3974 22536
rect 4030 22480 12714 22536
rect 12770 22480 12775 22536
rect 3969 22478 12775 22480
rect 2681 22475 2747 22478
rect 3969 22475 4035 22478
rect 12709 22475 12775 22478
rect 2589 22402 2655 22405
rect 5257 22402 5323 22405
rect 2589 22400 5323 22402
rect 2589 22344 2594 22400
rect 2650 22344 5262 22400
rect 5318 22344 5323 22400
rect 2589 22342 5323 22344
rect 2589 22339 2655 22342
rect 5257 22339 5323 22342
rect 5441 22402 5507 22405
rect 10041 22402 10107 22405
rect 5441 22400 10107 22402
rect 5441 22344 5446 22400
rect 5502 22344 10046 22400
rect 10102 22344 10107 22400
rect 5441 22342 10107 22344
rect 5441 22339 5507 22342
rect 10041 22339 10107 22342
rect 10277 22336 10597 22337
rect 0 22266 480 22296
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 1577 22266 1643 22269
rect 0 22264 1643 22266
rect 0 22208 1582 22264
rect 1638 22208 1643 22264
rect 0 22206 1643 22208
rect 0 22176 480 22206
rect 1577 22203 1643 22206
rect 2037 22266 2103 22269
rect 6821 22266 6887 22269
rect 2037 22264 6887 22266
rect 2037 22208 2042 22264
rect 2098 22208 6826 22264
rect 6882 22208 6887 22264
rect 2037 22206 6887 22208
rect 2037 22203 2103 22206
rect 6821 22203 6887 22206
rect 8753 22130 8819 22133
rect 13997 22130 14063 22133
rect 8753 22128 14063 22130
rect 8753 22072 8758 22128
rect 8814 22072 14002 22128
rect 14058 22072 14063 22128
rect 8753 22070 14063 22072
rect 8753 22067 8819 22070
rect 13997 22067 14063 22070
rect 4797 21994 4863 21997
rect 7649 21994 7715 21997
rect 4797 21992 7715 21994
rect 4797 21936 4802 21992
rect 4858 21936 7654 21992
rect 7710 21936 7715 21992
rect 4797 21934 7715 21936
rect 4797 21931 4863 21934
rect 7649 21931 7715 21934
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 0 21586 480 21616
rect 2957 21586 3023 21589
rect 0 21584 3023 21586
rect 0 21528 2962 21584
rect 3018 21528 3023 21584
rect 0 21526 3023 21528
rect 0 21496 480 21526
rect 2957 21523 3023 21526
rect 3141 21586 3207 21589
rect 16297 21586 16363 21589
rect 3141 21584 16363 21586
rect 3141 21528 3146 21584
rect 3202 21528 16302 21584
rect 16358 21528 16363 21584
rect 3141 21526 16363 21528
rect 3141 21523 3207 21526
rect 16297 21523 16363 21526
rect 9622 21388 9628 21452
rect 9692 21450 9698 21452
rect 9857 21450 9923 21453
rect 9692 21448 9923 21450
rect 9692 21392 9862 21448
rect 9918 21392 9923 21448
rect 9692 21390 9923 21392
rect 9692 21388 9698 21390
rect 9857 21387 9923 21390
rect 2681 21314 2747 21317
rect 9673 21314 9739 21317
rect 2681 21312 9739 21314
rect 2681 21256 2686 21312
rect 2742 21256 9678 21312
rect 9734 21256 9739 21312
rect 2681 21254 9739 21256
rect 2681 21251 2747 21254
rect 9673 21251 9739 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 1761 21178 1827 21181
rect 5993 21178 6059 21181
rect 1761 21176 6059 21178
rect 1761 21120 1766 21176
rect 1822 21120 5998 21176
rect 6054 21120 6059 21176
rect 1761 21118 6059 21120
rect 1761 21115 1827 21118
rect 5993 21115 6059 21118
rect 0 21042 480 21072
rect 3049 21042 3115 21045
rect 0 21040 3115 21042
rect 0 20984 3054 21040
rect 3110 20984 3115 21040
rect 0 20982 3115 20984
rect 0 20952 480 20982
rect 3049 20979 3115 20982
rect 8017 21042 8083 21045
rect 13169 21042 13235 21045
rect 8017 21040 13235 21042
rect 8017 20984 8022 21040
rect 8078 20984 13174 21040
rect 13230 20984 13235 21040
rect 8017 20982 13235 20984
rect 8017 20979 8083 20982
rect 13169 20979 13235 20982
rect 5809 20906 5875 20909
rect 10593 20906 10659 20909
rect 5809 20904 10659 20906
rect 5809 20848 5814 20904
rect 5870 20848 10598 20904
rect 10654 20848 10659 20904
rect 5809 20846 10659 20848
rect 5809 20843 5875 20846
rect 10593 20843 10659 20846
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 0 20362 480 20392
rect 1393 20362 1459 20365
rect 0 20360 1459 20362
rect 0 20304 1398 20360
rect 1454 20304 1459 20360
rect 0 20302 1459 20304
rect 0 20272 480 20302
rect 1393 20299 1459 20302
rect 3417 20362 3483 20365
rect 6269 20362 6335 20365
rect 3417 20360 6335 20362
rect 3417 20304 3422 20360
rect 3478 20304 6274 20360
rect 6330 20304 6335 20360
rect 3417 20302 6335 20304
rect 3417 20299 3483 20302
rect 6269 20299 6335 20302
rect 8477 20362 8543 20365
rect 11053 20362 11119 20365
rect 8477 20360 11119 20362
rect 8477 20304 8482 20360
rect 8538 20304 11058 20360
rect 11114 20304 11119 20360
rect 8477 20302 11119 20304
rect 8477 20299 8543 20302
rect 11053 20299 11119 20302
rect 15009 20226 15075 20229
rect 16665 20226 16731 20229
rect 15009 20224 16731 20226
rect 15009 20168 15014 20224
rect 15070 20168 16670 20224
rect 16726 20168 16731 20224
rect 15009 20166 16731 20168
rect 15009 20163 15075 20166
rect 16665 20163 16731 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 1485 19954 1551 19957
rect 9673 19954 9739 19957
rect 1485 19952 9739 19954
rect 1485 19896 1490 19952
rect 1546 19896 9678 19952
rect 9734 19896 9739 19952
rect 1485 19894 9739 19896
rect 1485 19891 1551 19894
rect 9673 19891 9739 19894
rect 0 19818 480 19848
rect 2865 19818 2931 19821
rect 0 19816 2931 19818
rect 0 19760 2870 19816
rect 2926 19760 2931 19816
rect 0 19758 2931 19760
rect 0 19728 480 19758
rect 2865 19755 2931 19758
rect 7741 19682 7807 19685
rect 11329 19682 11395 19685
rect 7741 19680 11395 19682
rect 7741 19624 7746 19680
rect 7802 19624 11334 19680
rect 11390 19624 11395 19680
rect 7741 19622 11395 19624
rect 7741 19619 7807 19622
rect 11329 19619 11395 19622
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 2313 19410 2379 19413
rect 6913 19410 6979 19413
rect 2313 19408 6979 19410
rect 2313 19352 2318 19408
rect 2374 19352 6918 19408
rect 6974 19352 6979 19408
rect 2313 19350 6979 19352
rect 2313 19347 2379 19350
rect 6913 19347 6979 19350
rect 8109 19274 8175 19277
rect 9489 19274 9555 19277
rect 9857 19274 9923 19277
rect 8109 19272 9923 19274
rect 8109 19216 8114 19272
rect 8170 19216 9494 19272
rect 9550 19216 9862 19272
rect 9918 19216 9923 19272
rect 8109 19214 9923 19216
rect 8109 19211 8175 19214
rect 9489 19211 9555 19214
rect 9857 19211 9923 19214
rect 0 19138 480 19168
rect 2957 19138 3023 19141
rect 0 19136 3023 19138
rect 0 19080 2962 19136
rect 3018 19080 3023 19136
rect 0 19078 3023 19080
rect 0 19048 480 19078
rect 2957 19075 3023 19078
rect 3417 19138 3483 19141
rect 4613 19138 4679 19141
rect 3417 19136 4679 19138
rect 3417 19080 3422 19136
rect 3478 19080 4618 19136
rect 4674 19080 4679 19136
rect 3417 19078 4679 19080
rect 3417 19075 3483 19078
rect 4613 19075 4679 19078
rect 7465 19138 7531 19141
rect 8569 19138 8635 19141
rect 7465 19136 8635 19138
rect 7465 19080 7470 19136
rect 7526 19080 8574 19136
rect 8630 19080 8635 19136
rect 7465 19078 8635 19080
rect 7465 19075 7531 19078
rect 8569 19075 8635 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 289 18866 355 18869
rect 6545 18866 6611 18869
rect 289 18864 6611 18866
rect 289 18808 294 18864
rect 350 18808 6550 18864
rect 6606 18808 6611 18864
rect 289 18806 6611 18808
rect 289 18803 355 18806
rect 6545 18803 6611 18806
rect 9949 18866 10015 18869
rect 12893 18866 12959 18869
rect 9949 18864 12959 18866
rect 9949 18808 9954 18864
rect 10010 18808 12898 18864
rect 12954 18808 12959 18864
rect 9949 18806 12959 18808
rect 9949 18803 10015 18806
rect 12893 18803 12959 18806
rect 3325 18730 3391 18733
rect 10133 18730 10199 18733
rect 3325 18728 10199 18730
rect 3325 18672 3330 18728
rect 3386 18672 10138 18728
rect 10194 18672 10199 18728
rect 3325 18670 10199 18672
rect 3325 18667 3391 18670
rect 10133 18667 10199 18670
rect 0 18594 480 18624
rect 4245 18594 4311 18597
rect 0 18592 4311 18594
rect 0 18536 4250 18592
rect 4306 18536 4311 18592
rect 0 18534 4311 18536
rect 0 18504 480 18534
rect 4245 18531 4311 18534
rect 6637 18594 6703 18597
rect 8477 18594 8543 18597
rect 6637 18592 8543 18594
rect 6637 18536 6642 18592
rect 6698 18536 8482 18592
rect 8538 18536 8543 18592
rect 6637 18534 8543 18536
rect 6637 18531 6703 18534
rect 8477 18531 8543 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 2221 18458 2287 18461
rect 5165 18458 5231 18461
rect 2221 18456 5231 18458
rect 2221 18400 2226 18456
rect 2282 18400 5170 18456
rect 5226 18400 5231 18456
rect 2221 18398 5231 18400
rect 2221 18395 2287 18398
rect 5165 18395 5231 18398
rect 8569 18458 8635 18461
rect 11421 18458 11487 18461
rect 8569 18456 11487 18458
rect 8569 18400 8574 18456
rect 8630 18400 11426 18456
rect 11482 18400 11487 18456
rect 8569 18398 11487 18400
rect 8569 18395 8635 18398
rect 11421 18395 11487 18398
rect 2221 18322 2287 18325
rect 3417 18322 3483 18325
rect 2221 18320 3483 18322
rect 2221 18264 2226 18320
rect 2282 18264 3422 18320
rect 3478 18264 3483 18320
rect 2221 18262 3483 18264
rect 2221 18259 2287 18262
rect 3417 18259 3483 18262
rect 4245 18322 4311 18325
rect 12801 18322 12867 18325
rect 4245 18320 12867 18322
rect 4245 18264 4250 18320
rect 4306 18264 12806 18320
rect 12862 18264 12867 18320
rect 4245 18262 12867 18264
rect 4245 18259 4311 18262
rect 12801 18259 12867 18262
rect 4705 18186 4771 18189
rect 15653 18186 15719 18189
rect 4705 18184 15719 18186
rect 4705 18128 4710 18184
rect 4766 18128 15658 18184
rect 15714 18128 15719 18184
rect 4705 18126 15719 18128
rect 4705 18123 4771 18126
rect 15653 18123 15719 18126
rect 12801 18050 12867 18053
rect 13261 18050 13327 18053
rect 15653 18050 15719 18053
rect 12801 18048 15719 18050
rect 12801 17992 12806 18048
rect 12862 17992 13266 18048
rect 13322 17992 15658 18048
rect 15714 17992 15719 18048
rect 12801 17990 15719 17992
rect 12801 17987 12867 17990
rect 13261 17987 13327 17990
rect 15653 17987 15719 17990
rect 10277 17984 10597 17985
rect 0 17914 480 17944
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 2865 17914 2931 17917
rect 0 17912 2931 17914
rect 0 17856 2870 17912
rect 2926 17856 2931 17912
rect 0 17854 2931 17856
rect 0 17824 480 17854
rect 2865 17851 2931 17854
rect 7833 17914 7899 17917
rect 10133 17914 10199 17917
rect 7833 17912 10199 17914
rect 7833 17856 7838 17912
rect 7894 17856 10138 17912
rect 10194 17856 10199 17912
rect 7833 17854 10199 17856
rect 7833 17851 7899 17854
rect 10133 17851 10199 17854
rect 6453 17778 6519 17781
rect 8753 17778 8819 17781
rect 6453 17776 8819 17778
rect 6453 17720 6458 17776
rect 6514 17720 8758 17776
rect 8814 17720 8819 17776
rect 6453 17718 8819 17720
rect 6453 17715 6519 17718
rect 8753 17715 8819 17718
rect 841 17642 907 17645
rect 1945 17642 2011 17645
rect 841 17640 2011 17642
rect 841 17584 846 17640
rect 902 17584 1950 17640
rect 2006 17584 2011 17640
rect 841 17582 2011 17584
rect 841 17579 907 17582
rect 1945 17579 2011 17582
rect 2497 17642 2563 17645
rect 5073 17642 5139 17645
rect 5533 17642 5599 17645
rect 2497 17640 5599 17642
rect 2497 17584 2502 17640
rect 2558 17584 5078 17640
rect 5134 17584 5538 17640
rect 5594 17584 5599 17640
rect 2497 17582 5599 17584
rect 2497 17579 2563 17582
rect 5073 17579 5139 17582
rect 5533 17579 5599 17582
rect 8753 17642 8819 17645
rect 16021 17642 16087 17645
rect 8753 17640 16087 17642
rect 8753 17584 8758 17640
rect 8814 17584 16026 17640
rect 16082 17584 16087 17640
rect 8753 17582 16087 17584
rect 8753 17579 8819 17582
rect 16021 17579 16087 17582
rect 10869 17506 10935 17509
rect 11237 17506 11303 17509
rect 13261 17506 13327 17509
rect 10869 17504 13327 17506
rect 10869 17448 10874 17504
rect 10930 17448 11242 17504
rect 11298 17448 13266 17504
rect 13322 17448 13327 17504
rect 10869 17446 13327 17448
rect 10869 17443 10935 17446
rect 11237 17443 11303 17446
rect 13261 17443 13327 17446
rect 5610 17440 5930 17441
rect 0 17370 480 17400
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 4245 17370 4311 17373
rect 0 17368 4311 17370
rect 0 17312 4250 17368
rect 4306 17312 4311 17368
rect 0 17310 4311 17312
rect 0 17280 480 17310
rect 4245 17307 4311 17310
rect 4705 17234 4771 17237
rect 8477 17234 8543 17237
rect 4705 17232 8543 17234
rect 4705 17176 4710 17232
rect 4766 17176 8482 17232
rect 8538 17176 8543 17232
rect 4705 17174 8543 17176
rect 4705 17171 4771 17174
rect 8477 17171 8543 17174
rect 7649 17098 7715 17101
rect 9489 17098 9555 17101
rect 7649 17096 9555 17098
rect 7649 17040 7654 17096
rect 7710 17040 9494 17096
rect 9550 17040 9555 17096
rect 7649 17038 9555 17040
rect 7649 17035 7715 17038
rect 9489 17035 9555 17038
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 11605 16826 11671 16829
rect 16205 16826 16271 16829
rect 11605 16824 16271 16826
rect 11605 16768 11610 16824
rect 11666 16768 16210 16824
rect 16266 16768 16271 16824
rect 11605 16766 16271 16768
rect 11605 16763 11671 16766
rect 16205 16763 16271 16766
rect 0 16690 480 16720
rect 1577 16690 1643 16693
rect 0 16688 1643 16690
rect 0 16632 1582 16688
rect 1638 16632 1643 16688
rect 0 16630 1643 16632
rect 0 16600 480 16630
rect 1577 16627 1643 16630
rect 9949 16690 10015 16693
rect 13905 16690 13971 16693
rect 9949 16688 13971 16690
rect 9949 16632 9954 16688
rect 10010 16632 13910 16688
rect 13966 16632 13971 16688
rect 9949 16630 13971 16632
rect 9949 16627 10015 16630
rect 13905 16627 13971 16630
rect 5165 16554 5231 16557
rect 9029 16554 9095 16557
rect 5165 16552 9095 16554
rect 5165 16496 5170 16552
rect 5226 16496 9034 16552
rect 9090 16496 9095 16552
rect 5165 16494 9095 16496
rect 5165 16491 5231 16494
rect 9029 16491 9095 16494
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 3141 16282 3207 16285
rect 3141 16280 3986 16282
rect 3141 16224 3146 16280
rect 3202 16224 3986 16280
rect 3141 16222 3986 16224
rect 3141 16219 3207 16222
rect 0 16146 480 16176
rect 3785 16146 3851 16149
rect 0 16144 3851 16146
rect 0 16088 3790 16144
rect 3846 16088 3851 16144
rect 0 16086 3851 16088
rect 3926 16146 3986 16222
rect 16297 16146 16363 16149
rect 3926 16144 16363 16146
rect 3926 16088 16302 16144
rect 16358 16088 16363 16144
rect 3926 16086 16363 16088
rect 0 16056 480 16086
rect 3785 16083 3851 16086
rect 16297 16083 16363 16086
rect 1393 16010 1459 16013
rect 12525 16010 12591 16013
rect 1393 16008 12591 16010
rect 1393 15952 1398 16008
rect 1454 15952 12530 16008
rect 12586 15952 12591 16008
rect 1393 15950 12591 15952
rect 1393 15947 1459 15950
rect 12525 15947 12591 15950
rect 10961 15874 11027 15877
rect 12433 15874 12499 15877
rect 10961 15872 12499 15874
rect 10961 15816 10966 15872
rect 11022 15816 12438 15872
rect 12494 15816 12499 15872
rect 10961 15814 12499 15816
rect 10961 15811 11027 15814
rect 12433 15811 12499 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 0 15466 480 15496
rect 1485 15466 1551 15469
rect 0 15464 1551 15466
rect 0 15408 1490 15464
rect 1546 15408 1551 15464
rect 0 15406 1551 15408
rect 0 15376 480 15406
rect 1485 15403 1551 15406
rect 3877 15466 3943 15469
rect 9857 15466 9923 15469
rect 3877 15464 9923 15466
rect 3877 15408 3882 15464
rect 3938 15408 9862 15464
rect 9918 15408 9923 15464
rect 3877 15406 9923 15408
rect 3877 15403 3943 15406
rect 9857 15403 9923 15406
rect 10869 15466 10935 15469
rect 11145 15466 11211 15469
rect 13169 15466 13235 15469
rect 10869 15464 13235 15466
rect 10869 15408 10874 15464
rect 10930 15408 11150 15464
rect 11206 15408 13174 15464
rect 13230 15408 13235 15464
rect 10869 15406 13235 15408
rect 10869 15403 10935 15406
rect 11145 15403 11211 15406
rect 13169 15403 13235 15406
rect 9029 15330 9095 15333
rect 11329 15330 11395 15333
rect 9029 15328 11395 15330
rect 9029 15272 9034 15328
rect 9090 15272 11334 15328
rect 11390 15272 11395 15328
rect 9029 15270 11395 15272
rect 9029 15267 9095 15270
rect 11329 15267 11395 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 3785 15058 3851 15061
rect 6913 15058 6979 15061
rect 3785 15056 6979 15058
rect 3785 15000 3790 15056
rect 3846 15000 6918 15056
rect 6974 15000 6979 15056
rect 3785 14998 6979 15000
rect 3785 14995 3851 14998
rect 6913 14995 6979 14998
rect 8017 15058 8083 15061
rect 12433 15058 12499 15061
rect 8017 15056 12499 15058
rect 8017 15000 8022 15056
rect 8078 15000 12438 15056
rect 12494 15000 12499 15056
rect 8017 14998 12499 15000
rect 8017 14995 8083 14998
rect 12433 14995 12499 14998
rect 12985 15058 13051 15061
rect 15285 15058 15351 15061
rect 12985 15056 15351 15058
rect 12985 15000 12990 15056
rect 13046 15000 15290 15056
rect 15346 15000 15351 15056
rect 12985 14998 15351 15000
rect 12985 14995 13051 14998
rect 15285 14995 15351 14998
rect 0 14922 480 14952
rect 3969 14922 4035 14925
rect 0 14920 4035 14922
rect 0 14864 3974 14920
rect 4030 14864 4035 14920
rect 0 14862 4035 14864
rect 0 14832 480 14862
rect 3969 14859 4035 14862
rect 6729 14922 6795 14925
rect 7465 14922 7531 14925
rect 6729 14920 7531 14922
rect 6729 14864 6734 14920
rect 6790 14864 7470 14920
rect 7526 14864 7531 14920
rect 6729 14862 7531 14864
rect 6729 14859 6795 14862
rect 7465 14859 7531 14862
rect 4889 14786 4955 14789
rect 10041 14786 10107 14789
rect 4889 14784 10107 14786
rect 4889 14728 4894 14784
rect 4950 14728 10046 14784
rect 10102 14728 10107 14784
rect 4889 14726 10107 14728
rect 4889 14723 4955 14726
rect 10041 14723 10107 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 16113 14650 16179 14653
rect 17493 14650 17559 14653
rect 16113 14648 17559 14650
rect 16113 14592 16118 14648
rect 16174 14592 17498 14648
rect 17554 14592 17559 14648
rect 16113 14590 17559 14592
rect 16113 14587 16179 14590
rect 17493 14587 17559 14590
rect 3325 14514 3391 14517
rect 10685 14514 10751 14517
rect 11329 14514 11395 14517
rect 3325 14512 11395 14514
rect 3325 14456 3330 14512
rect 3386 14456 10690 14512
rect 10746 14456 11334 14512
rect 11390 14456 11395 14512
rect 3325 14454 11395 14456
rect 3325 14451 3391 14454
rect 10685 14451 10751 14454
rect 11329 14451 11395 14454
rect 0 14378 480 14408
rect 1853 14378 1919 14381
rect 0 14376 1919 14378
rect 0 14320 1858 14376
rect 1914 14320 1919 14376
rect 0 14318 1919 14320
rect 0 14288 480 14318
rect 1853 14315 1919 14318
rect 4521 14378 4587 14381
rect 7097 14378 7163 14381
rect 4521 14376 7163 14378
rect 4521 14320 4526 14376
rect 4582 14320 7102 14376
rect 7158 14320 7163 14376
rect 4521 14318 7163 14320
rect 4521 14315 4587 14318
rect 7097 14315 7163 14318
rect 8845 14378 8911 14381
rect 27613 14378 27679 14381
rect 8845 14376 27679 14378
rect 8845 14320 8850 14376
rect 8906 14320 27618 14376
rect 27674 14320 27679 14376
rect 8845 14318 27679 14320
rect 8845 14315 8911 14318
rect 27613 14315 27679 14318
rect 9029 14242 9095 14245
rect 14457 14242 14523 14245
rect 9029 14240 14523 14242
rect 9029 14184 9034 14240
rect 9090 14184 14462 14240
rect 14518 14184 14523 14240
rect 9029 14182 14523 14184
rect 9029 14179 9095 14182
rect 14457 14179 14523 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 8201 14106 8267 14109
rect 27520 14106 28000 14136
rect 6134 14104 8267 14106
rect 6134 14048 8206 14104
rect 8262 14048 8267 14104
rect 6134 14046 8267 14048
rect 2957 13970 3023 13973
rect 3233 13970 3299 13973
rect 4337 13970 4403 13973
rect 6134 13970 6194 14046
rect 8201 14043 8267 14046
rect 24902 14046 28000 14106
rect 9581 13970 9647 13973
rect 15193 13970 15259 13973
rect 24902 13970 24962 14046
rect 27520 14016 28000 14046
rect 2957 13968 6194 13970
rect 2957 13912 2962 13968
rect 3018 13912 3238 13968
rect 3294 13912 4342 13968
rect 4398 13912 6194 13968
rect 2957 13910 6194 13912
rect 9500 13968 9690 13970
rect 9500 13912 9586 13968
rect 9642 13912 9690 13968
rect 9500 13910 9690 13912
rect 2957 13907 3023 13910
rect 3233 13907 3299 13910
rect 4337 13907 4403 13910
rect 9581 13907 9690 13910
rect 15193 13968 24962 13970
rect 15193 13912 15198 13968
rect 15254 13912 24962 13968
rect 15193 13910 24962 13912
rect 15193 13907 15259 13910
rect 9630 13837 9690 13907
rect 6913 13834 6979 13837
rect 9581 13834 9690 13837
rect 6913 13832 14290 13834
rect 6913 13776 6918 13832
rect 6974 13776 9586 13832
rect 9642 13776 14290 13832
rect 6913 13774 14290 13776
rect 6913 13771 6979 13774
rect 9581 13771 9647 13774
rect 0 13698 480 13728
rect 5257 13698 5323 13701
rect 0 13696 5323 13698
rect 0 13640 5262 13696
rect 5318 13640 5323 13696
rect 0 13638 5323 13640
rect 0 13608 480 13638
rect 5257 13635 5323 13638
rect 6545 13698 6611 13701
rect 9121 13698 9187 13701
rect 6545 13696 9187 13698
rect 6545 13640 6550 13696
rect 6606 13640 9126 13696
rect 9182 13640 9187 13696
rect 6545 13638 9187 13640
rect 14230 13698 14290 13774
rect 15193 13698 15259 13701
rect 14230 13696 15259 13698
rect 14230 13640 15198 13696
rect 15254 13640 15259 13696
rect 14230 13638 15259 13640
rect 6545 13635 6611 13638
rect 9121 13635 9187 13638
rect 15193 13635 15259 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 2037 13562 2103 13565
rect 2037 13560 3986 13562
rect 2037 13504 2042 13560
rect 2098 13504 3986 13560
rect 2037 13502 3986 13504
rect 2037 13499 2103 13502
rect 3926 13426 3986 13502
rect 5165 13426 5231 13429
rect 3926 13424 5231 13426
rect 3926 13368 5170 13424
rect 5226 13368 5231 13424
rect 3926 13366 5231 13368
rect 5165 13363 5231 13366
rect 0 13154 480 13184
rect 3877 13154 3943 13157
rect 0 13152 3943 13154
rect 0 13096 3882 13152
rect 3938 13096 3943 13152
rect 0 13094 3943 13096
rect 0 13064 480 13094
rect 3877 13091 3943 13094
rect 10777 13154 10843 13157
rect 11145 13154 11211 13157
rect 12433 13154 12499 13157
rect 10777 13152 12499 13154
rect 10777 13096 10782 13152
rect 10838 13096 11150 13152
rect 11206 13096 12438 13152
rect 12494 13096 12499 13152
rect 10777 13094 12499 13096
rect 10777 13091 10843 13094
rect 11145 13091 11211 13094
rect 12433 13091 12499 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 2865 12882 2931 12885
rect 8661 12882 8727 12885
rect 2865 12880 8727 12882
rect 2865 12824 2870 12880
rect 2926 12824 8666 12880
rect 8722 12824 8727 12880
rect 2865 12822 8727 12824
rect 2865 12819 2931 12822
rect 8661 12819 8727 12822
rect 16205 12882 16271 12885
rect 17953 12882 18019 12885
rect 16205 12880 18019 12882
rect 16205 12824 16210 12880
rect 16266 12824 17958 12880
rect 18014 12824 18019 12880
rect 16205 12822 18019 12824
rect 16205 12819 16271 12822
rect 17953 12819 18019 12822
rect 5165 12746 5231 12749
rect 15929 12746 15995 12749
rect 5165 12744 15995 12746
rect 5165 12688 5170 12744
rect 5226 12688 15934 12744
rect 15990 12688 15995 12744
rect 5165 12686 15995 12688
rect 5165 12683 5231 12686
rect 15929 12683 15995 12686
rect 11789 12610 11855 12613
rect 13813 12610 13879 12613
rect 11789 12608 13879 12610
rect 11789 12552 11794 12608
rect 11850 12552 13818 12608
rect 13874 12552 13879 12608
rect 11789 12550 13879 12552
rect 11789 12547 11855 12550
rect 13813 12547 13879 12550
rect 10277 12544 10597 12545
rect 0 12474 480 12504
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 1761 12474 1827 12477
rect 2405 12474 2471 12477
rect 0 12472 2471 12474
rect 0 12416 1766 12472
rect 1822 12416 2410 12472
rect 2466 12416 2471 12472
rect 0 12414 2471 12416
rect 0 12384 480 12414
rect 1761 12411 1827 12414
rect 2405 12411 2471 12414
rect 3785 12338 3851 12341
rect 4061 12338 4127 12341
rect 5717 12338 5783 12341
rect 3785 12336 5783 12338
rect 3785 12280 3790 12336
rect 3846 12280 4066 12336
rect 4122 12280 5722 12336
rect 5778 12280 5783 12336
rect 3785 12278 5783 12280
rect 3785 12275 3851 12278
rect 4061 12275 4127 12278
rect 5717 12275 5783 12278
rect 11605 12338 11671 12341
rect 20805 12338 20871 12341
rect 11605 12336 20871 12338
rect 11605 12280 11610 12336
rect 11666 12280 20810 12336
rect 20866 12280 20871 12336
rect 11605 12278 20871 12280
rect 11605 12275 11671 12278
rect 20805 12275 20871 12278
rect 4061 12202 4127 12205
rect 17033 12202 17099 12205
rect 4061 12200 17099 12202
rect 4061 12144 4066 12200
rect 4122 12144 17038 12200
rect 17094 12144 17099 12200
rect 4061 12142 17099 12144
rect 4061 12139 4127 12142
rect 17033 12139 17099 12142
rect 6729 12066 6795 12069
rect 9949 12066 10015 12069
rect 6729 12064 10015 12066
rect 6729 12008 6734 12064
rect 6790 12008 9954 12064
rect 10010 12008 10015 12064
rect 6729 12006 10015 12008
rect 6729 12003 6795 12006
rect 9949 12003 10015 12006
rect 5610 12000 5930 12001
rect 0 11930 480 11960
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 2865 11930 2931 11933
rect 0 11928 2931 11930
rect 0 11872 2870 11928
rect 2926 11872 2931 11928
rect 0 11870 2931 11872
rect 0 11840 480 11870
rect 2865 11867 2931 11870
rect 1393 11658 1459 11661
rect 17953 11658 18019 11661
rect 1393 11656 18019 11658
rect 1393 11600 1398 11656
rect 1454 11600 17958 11656
rect 18014 11600 18019 11656
rect 1393 11598 18019 11600
rect 1393 11595 1459 11598
rect 17953 11595 18019 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 0 11250 480 11280
rect 1577 11250 1643 11253
rect 0 11248 1643 11250
rect 0 11192 1582 11248
rect 1638 11192 1643 11248
rect 0 11190 1643 11192
rect 0 11160 480 11190
rect 1577 11187 1643 11190
rect 8017 11250 8083 11253
rect 20897 11250 20963 11253
rect 8017 11248 20963 11250
rect 8017 11192 8022 11248
rect 8078 11192 20902 11248
rect 20958 11192 20963 11248
rect 8017 11190 20963 11192
rect 8017 11187 8083 11190
rect 20897 11187 20963 11190
rect 5625 11114 5691 11117
rect 11697 11114 11763 11117
rect 5625 11112 11763 11114
rect 5625 11056 5630 11112
rect 5686 11056 11702 11112
rect 11758 11056 11763 11112
rect 5625 11054 11763 11056
rect 5625 11051 5691 11054
rect 11697 11051 11763 11054
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 0 10706 480 10736
rect 2129 10706 2195 10709
rect 0 10704 2195 10706
rect 0 10648 2134 10704
rect 2190 10648 2195 10704
rect 0 10646 2195 10648
rect 0 10616 480 10646
rect 2129 10643 2195 10646
rect 6821 10570 6887 10573
rect 19701 10570 19767 10573
rect 6821 10568 19767 10570
rect 6821 10512 6826 10568
rect 6882 10512 19706 10568
rect 19762 10512 19767 10568
rect 6821 10510 19767 10512
rect 6821 10507 6887 10510
rect 19701 10507 19767 10510
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 0 10026 480 10056
rect 9673 10026 9739 10029
rect 19517 10026 19583 10029
rect 0 9966 2698 10026
rect 0 9936 480 9966
rect 2497 9618 2563 9621
rect 2638 9618 2698 9966
rect 9673 10024 19583 10026
rect 9673 9968 9678 10024
rect 9734 9968 19522 10024
rect 19578 9968 19583 10024
rect 9673 9966 19583 9968
rect 9673 9963 9739 9966
rect 19517 9963 19583 9966
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 2497 9616 2698 9618
rect 2497 9560 2502 9616
rect 2558 9560 2698 9616
rect 2497 9558 2698 9560
rect 2497 9555 2563 9558
rect 0 9482 480 9512
rect 7833 9482 7899 9485
rect 0 9480 7899 9482
rect 0 9424 7838 9480
rect 7894 9424 7899 9480
rect 0 9422 7899 9424
rect 0 9392 480 9422
rect 7833 9419 7899 9422
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 3969 8938 4035 8941
rect 18413 8938 18479 8941
rect 3969 8936 18479 8938
rect 3969 8880 3974 8936
rect 4030 8880 18418 8936
rect 18474 8880 18479 8936
rect 3969 8878 18479 8880
rect 3969 8875 4035 8878
rect 18413 8875 18479 8878
rect 0 8802 480 8832
rect 0 8742 2698 8802
rect 0 8712 480 8742
rect 2638 8666 2698 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 2638 8606 2882 8666
rect 2822 8530 2882 8606
rect 9673 8530 9739 8533
rect 2822 8528 9739 8530
rect 2822 8472 9678 8528
rect 9734 8472 9739 8528
rect 2822 8470 9739 8472
rect 9673 8467 9739 8470
rect 11053 8394 11119 8397
rect 9998 8392 11119 8394
rect 9998 8336 11058 8392
rect 11114 8336 11119 8392
rect 9998 8334 11119 8336
rect 0 8258 480 8288
rect 9998 8258 10058 8334
rect 11053 8331 11119 8334
rect 0 8198 10058 8258
rect 0 8168 480 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 2405 8122 2471 8125
rect 4521 8122 4587 8125
rect 2405 8120 4587 8122
rect 2405 8064 2410 8120
rect 2466 8064 4526 8120
rect 4582 8064 4587 8120
rect 2405 8062 4587 8064
rect 2405 8059 2471 8062
rect 4521 8059 4587 8062
rect 4889 7986 4955 7989
rect 22277 7986 22343 7989
rect 4889 7984 22343 7986
rect 4889 7928 4894 7984
rect 4950 7928 22282 7984
rect 22338 7928 22343 7984
rect 4889 7926 22343 7928
rect 4889 7923 4955 7926
rect 22277 7923 22343 7926
rect 4061 7850 4127 7853
rect 18045 7850 18111 7853
rect 4061 7848 18111 7850
rect 4061 7792 4066 7848
rect 4122 7792 18050 7848
rect 18106 7792 18111 7848
rect 4061 7790 18111 7792
rect 4061 7787 4127 7790
rect 18045 7787 18111 7790
rect 5610 7648 5930 7649
rect 0 7578 480 7608
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 565 7578 631 7581
rect 0 7576 631 7578
rect 0 7520 570 7576
rect 626 7520 631 7576
rect 0 7518 631 7520
rect 0 7488 480 7518
rect 565 7515 631 7518
rect 3417 7442 3483 7445
rect 23657 7442 23723 7445
rect 3417 7440 23723 7442
rect 3417 7384 3422 7440
rect 3478 7384 23662 7440
rect 23718 7384 23723 7440
rect 3417 7382 23723 7384
rect 3417 7379 3483 7382
rect 23657 7379 23723 7382
rect 10277 7104 10597 7105
rect 0 7034 480 7064
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 565 7034 631 7037
rect 0 7032 631 7034
rect 0 6976 570 7032
rect 626 6976 631 7032
rect 0 6974 631 6976
rect 0 6944 480 6974
rect 565 6971 631 6974
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 0 6354 480 6384
rect 23657 6354 23723 6357
rect 0 6352 23723 6354
rect 0 6296 23662 6352
rect 23718 6296 23723 6352
rect 0 6294 23723 6296
rect 0 6264 480 6294
rect 23657 6291 23723 6294
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 0 5810 480 5840
rect 24025 5810 24091 5813
rect 0 5808 24091 5810
rect 0 5752 24030 5808
rect 24086 5752 24091 5808
rect 0 5750 24091 5752
rect 0 5720 480 5750
rect 24025 5747 24091 5750
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 24669 5402 24735 5405
rect 26233 5402 26299 5405
rect 24669 5400 26299 5402
rect 24669 5344 24674 5400
rect 24730 5344 26238 5400
rect 26294 5344 26299 5400
rect 24669 5342 26299 5344
rect 24669 5339 24735 5342
rect 26233 5339 26299 5342
rect 24485 5266 24551 5269
rect 614 5264 24551 5266
rect 614 5208 24490 5264
rect 24546 5208 24551 5264
rect 614 5206 24551 5208
rect 0 5130 480 5160
rect 614 5130 674 5206
rect 24485 5203 24551 5206
rect 0 5070 674 5130
rect 0 5040 480 5070
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 24761 4858 24827 4861
rect 26877 4858 26943 4861
rect 24761 4856 26943 4858
rect 24761 4800 24766 4856
rect 24822 4800 26882 4856
rect 26938 4800 26943 4856
rect 24761 4798 26943 4800
rect 24761 4795 24827 4798
rect 26877 4795 26943 4798
rect 24577 4722 24643 4725
rect 614 4720 24643 4722
rect 614 4664 24582 4720
rect 24638 4664 24643 4720
rect 614 4662 24643 4664
rect 0 4586 480 4616
rect 614 4586 674 4662
rect 24577 4659 24643 4662
rect 0 4526 674 4586
rect 0 4496 480 4526
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 7005 4042 7071 4045
rect 8477 4042 8543 4045
rect 7005 4040 8543 4042
rect 7005 3984 7010 4040
rect 7066 3984 8482 4040
rect 8538 3984 8543 4040
rect 7005 3982 8543 3984
rect 7005 3979 7071 3982
rect 8477 3979 8543 3982
rect 0 3906 480 3936
rect 3325 3906 3391 3909
rect 0 3904 3391 3906
rect 0 3848 3330 3904
rect 3386 3848 3391 3904
rect 0 3846 3391 3848
rect 0 3816 480 3846
rect 3325 3843 3391 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 6177 3498 6243 3501
rect 20989 3498 21055 3501
rect 6177 3496 21055 3498
rect 6177 3440 6182 3496
rect 6238 3440 20994 3496
rect 21050 3440 21055 3496
rect 6177 3438 21055 3440
rect 6177 3435 6243 3438
rect 20989 3435 21055 3438
rect 0 3362 480 3392
rect 3601 3362 3667 3365
rect 0 3360 3667 3362
rect 0 3304 3606 3360
rect 3662 3304 3667 3360
rect 0 3302 3667 3304
rect 0 3272 480 3302
rect 3601 3299 3667 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 10277 2752 10597 2753
rect 0 2682 480 2712
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 3233 2682 3299 2685
rect 0 2680 3299 2682
rect 0 2624 3238 2680
rect 3294 2624 3299 2680
rect 0 2622 3299 2624
rect 0 2592 480 2622
rect 3233 2619 3299 2622
rect 3417 2546 3483 2549
rect 10777 2546 10843 2549
rect 3417 2544 10843 2546
rect 3417 2488 3422 2544
rect 3478 2488 10782 2544
rect 10838 2488 10843 2544
rect 3417 2486 10843 2488
rect 3417 2483 3483 2486
rect 10777 2483 10843 2486
rect 12157 2410 12223 2413
rect 1718 2408 12223 2410
rect 1718 2352 12162 2408
rect 12218 2352 12223 2408
rect 1718 2350 12223 2352
rect 0 2138 480 2168
rect 1718 2138 1778 2350
rect 12157 2347 12223 2350
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 0 2078 1778 2138
rect 0 2048 480 2078
rect 0 1458 480 1488
rect 3417 1458 3483 1461
rect 0 1456 3483 1458
rect 0 1400 3422 1456
rect 3478 1400 3483 1456
rect 0 1398 3483 1400
rect 0 1368 480 1398
rect 3417 1395 3483 1398
rect 12433 1322 12499 1325
rect 3374 1320 12499 1322
rect 3374 1264 12438 1320
rect 12494 1264 12499 1320
rect 3374 1262 12499 1264
rect 0 914 480 944
rect 3374 914 3434 1262
rect 12433 1259 12499 1262
rect 3509 1186 3575 1189
rect 10685 1186 10751 1189
rect 3509 1184 10751 1186
rect 3509 1128 3514 1184
rect 3570 1128 10690 1184
rect 10746 1128 10751 1184
rect 3509 1126 10751 1128
rect 3509 1123 3575 1126
rect 10685 1123 10751 1126
rect 0 854 3434 914
rect 0 824 480 854
rect 0 370 480 400
rect 3509 370 3575 373
rect 0 368 3575 370
rect 0 312 3514 368
rect 3570 312 3575 368
rect 0 310 3575 312
rect 0 280 480 310
rect 3509 307 3575 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 2084 23624 2148 23628
rect 2084 23568 2098 23624
rect 2098 23568 2148 23624
rect 2084 23564 2148 23568
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 9628 21388 9692 21452
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 2083 23628 2149 23629
rect 2083 23564 2084 23628
rect 2148 23564 2149 23628
rect 2083 23563 2149 23564
rect 2086 21538 2146 23563
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 1998 21302 2234 21538
rect 9542 21452 9778 21538
rect 9542 21388 9628 21452
rect 9628 21388 9692 21452
rect 9692 21388 9778 21452
rect 9542 21302 9778 21388
<< metal5 >>
rect 1956 21538 9820 21580
rect 1956 21302 1998 21538
rect 2234 21302 9542 21538
rect 9778 21302 9820 21538
rect 1956 21260 9820 21302
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1604681595
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1604681595
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604681595
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1604681595
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1604681595
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1604681595
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1604681595
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1604681595
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1604681595
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1604681595
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1604681595
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1604681595
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1604681595
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1604681595
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1604681595
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1604681595
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_220
timestamp 1604681595
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1604681595
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1604681595
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_249
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_232
timestamp 1604681595
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_261
timestamp 1604681595
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1604681595
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_269
timestamp 1604681595
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_273
timestamp 1604681595
transform 1 0 26220 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1604681595
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1604681595
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1604681595
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1604681595
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1604681595
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1604681595
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1604681595
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1604681595
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1604681595
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1604681595
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1604681595
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1604681595
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1604681595
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1604681595
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1604681595
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1604681595
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604681595
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1604681595
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1604681595
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1604681595
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1604681595
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1604681595
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1604681595
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1604681595
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1604681595
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1604681595
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1604681595
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 24564 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_253
timestamp 1604681595
transform 1 0 24380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1604681595
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_269
timestamp 1604681595
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1604681595
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1604681595
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1604681595
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1604681595
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1604681595
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1604681595
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1604681595
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1604681595
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1604681595
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1604681595
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1604681595
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1604681595
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _80_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 24564 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_251
timestamp 1604681595
transform 1 0 24196 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_259
timestamp 1604681595
transform 1 0 24932 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_271
timestamp 1604681595
transform 1 0 26036 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1604681595
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1604681595
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1604681595
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1604681595
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1604681595
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1604681595
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1604681595
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1604681595
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1604681595
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1604681595
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1604681595
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1604681595
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__82__A
timestamp 1604681595
transform 1 0 24012 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1604681595
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_245
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1604681595
transform 1 0 24472 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__81__A
timestamp 1604681595
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_251
timestamp 1604681595
transform 1 0 24196 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_258
timestamp 1604681595
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_262
timestamp 1604681595
transform 1 0 25208 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_274
timestamp 1604681595
transform 1 0 26312 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604681595
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1604681595
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1604681595
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1604681595
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1604681595
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1604681595
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1604681595
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1604681595
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1604681595
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1604681595
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1604681595
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1604681595
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1604681595
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1604681595
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1604681595
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1604681595
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1604681595
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1604681595
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1604681595
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1604681595
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1604681595
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1604681595
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1604681595
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1604681595
transform 1 0 24012 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_239
timestamp 1604681595
transform 1 0 23092 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_247
timestamp 1604681595
transform 1 0 23828 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_232
timestamp 1604681595
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_249
timestamp 1604681595
transform 1 0 24012 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__83__A
timestamp 1604681595
transform 1 0 24196 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1604681595
transform 1 0 24380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_265
timestamp 1604681595
transform 1 0 25484 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_253
timestamp 1604681595
transform 1 0 24380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_265
timestamp 1604681595
transform 1 0 25484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_273
timestamp 1604681595
transform 1 0 26220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1604681595
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1604681595
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1604681595
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1604681595
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1604681595
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1604681595
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1604681595
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1604681595
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1604681595
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1604681595
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1604681595
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1604681595
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_251
timestamp 1604681595
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1604681595
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_31
timestamp 1604681595
transform 1 0 3956 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_34
timestamp 1604681595
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_38
timestamp 1604681595
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_42
timestamp 1604681595
transform 1 0 4968 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_54
timestamp 1604681595
transform 1 0 6072 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1604681595
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1604681595
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1604681595
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_98
timestamp 1604681595
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_110
timestamp 1604681595
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1604681595
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1604681595
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1604681595
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1604681595
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1604681595
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1604681595
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_220
timestamp 1604681595
transform 1 0 21344 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_228
timestamp 1604681595
transform 1 0 22080 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__85__A
timestamp 1604681595
transform 1 0 22264 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_232
timestamp 1604681595
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_249
timestamp 1604681595
transform 1 0 24012 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__84__A
timestamp 1604681595
transform 1 0 24196 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_253
timestamp 1604681595
transform 1 0 24380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_265
timestamp 1604681595
transform 1 0 25484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_15
timestamp 1604681595
transform 1 0 2484 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_23
timestamp 1604681595
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_41
timestamp 1604681595
transform 1 0 4876 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _40_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5796 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_49
timestamp 1604681595
transform 1 0 5612 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_54
timestamp 1604681595
transform 1 0 6072 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_66
timestamp 1604681595
transform 1 0 7176 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_70
timestamp 1604681595
transform 1 0 7544 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_73
timestamp 1604681595
transform 1 0 7820 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_85
timestamp 1604681595
transform 1 0 8924 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1604681595
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1604681595
transform 1 0 10028 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1604681595
transform 1 0 11132 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1604681595
transform 1 0 12236 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_133
timestamp 1604681595
transform 1 0 13340 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_145
timestamp 1604681595
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1604681595
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1604681595
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1604681595
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1604681595
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_227
timestamp 1604681595
transform 1 0 21988 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1604681595
transform 1 0 22264 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_234
timestamp 1604681595
transform 1 0 22632 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_246
timestamp 1604681595
transform 1 0 23736 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_258
timestamp 1604681595
transform 1 0 24840 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_270
timestamp 1604681595
transform 1 0 25944 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_274
timestamp 1604681595
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_7
timestamp 1604681595
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_11
timestamp 1604681595
transform 1 0 2116 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_16
timestamp 1604681595
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_20
timestamp 1604681595
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4048 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3128 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3496 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_24
timestamp 1604681595
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_28
timestamp 1604681595
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_51
timestamp 1604681595
transform 1 0 5796 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7636 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7452 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6992 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_66
timestamp 1604681595
transform 1 0 7176 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1604681595
transform 1 0 10120 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_90
timestamp 1604681595
transform 1 0 9384 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_95
timestamp 1604681595
transform 1 0 9844 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1604681595
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_105
timestamp 1604681595
transform 1 0 10764 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_117
timestamp 1604681595
transform 1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1604681595
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1604681595
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1604681595
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1604681595
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1604681595
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1604681595
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_220
timestamp 1604681595
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_232
timestamp 1604681595
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1604681595
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_269
timestamp 1604681595
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_8
timestamp 1604681595
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_12
timestamp 1604681595
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_23
timestamp 1604681595
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_41
timestamp 1604681595
transform 1 0 4876 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6348 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_47
timestamp 1604681595
transform 1 0 5428 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_51
timestamp 1604681595
transform 1 0 5796 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 8648 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8280 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_76
timestamp 1604681595
transform 1 0 8096 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_80
timestamp 1604681595
transform 1 0 8464 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_84
timestamp 1604681595
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_88
timestamp 1604681595
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_102
timestamp 1604681595
transform 1 0 10488 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_114
timestamp 1604681595
transform 1 0 11592 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_126
timestamp 1604681595
transform 1 0 12696 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_138
timestamp 1604681595
transform 1 0 13800 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_150
timestamp 1604681595
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1604681595
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1604681595
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1604681595
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1604681595
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1604681595
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1604681595
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_251
timestamp 1604681595
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_263
timestamp 1604681595
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 1656 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_22
timestamp 1604681595
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3312 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_25
timestamp 1604681595
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1604681595
transform 1 0 3496 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3680 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_29
timestamp 1604681595
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1604681595
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_39
timestamp 1604681595
transform 1 0 4692 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_35
timestamp 1604681595
transform 1 0 4324 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 4508 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4140 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5244 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_52
timestamp 1604681595
transform 1 0 5888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1604681595
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_43
timestamp 1604681595
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_68
timestamp 1604681595
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_64
timestamp 1604681595
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_71
timestamp 1604681595
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 7544 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7728 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_81
timestamp 1604681595
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_79
timestamp 1604681595
transform 1 0 8372 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_75
timestamp 1604681595
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 8648 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_101
timestamp 1604681595
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp 1604681595
transform 1 0 8924 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_89
timestamp 1604681595
transform 1 0 9292 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_102
timestamp 1604681595
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_106
timestamp 1604681595
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_112
timestamp 1604681595
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_109
timestamp 1604681595
transform 1 0 11132 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_105
timestamp 1604681595
transform 1 0 10764 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11040 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11224 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1604681595
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_116
timestamp 1604681595
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_119
timestamp 1604681595
transform 1 0 12052 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1604681595
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_131
timestamp 1604681595
transform 1 0 13156 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_143
timestamp 1604681595
transform 1 0 14260 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_147
timestamp 1604681595
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_159
timestamp 1604681595
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1604681595
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1604681595
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_171
timestamp 1604681595
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1604681595
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 19504 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19504 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_196
timestamp 1604681595
transform 1 0 19136 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_202
timestamp 1604681595
transform 1 0 19688 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_190
timestamp 1604681595
transform 1 0 18584 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_198
timestamp 1604681595
transform 1 0 19320 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_206
timestamp 1604681595
transform 1 0 20056 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_214
timestamp 1604681595
transform 1 0 20792 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_226
timestamp 1604681595
transform 1 0 21896 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1604681595
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_238
timestamp 1604681595
transform 1 0 23000 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1604681595
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1604681595
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_269
timestamp 1604681595
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_251
timestamp 1604681595
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_263
timestamp 1604681595
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2300 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2116 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_9
timestamp 1604681595
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4232 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_22
timestamp 1604681595
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_26
timestamp 1604681595
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_30
timestamp 1604681595
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_53
timestamp 1604681595
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1604681595
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1604681595
transform 1 0 8372 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_71
timestamp 1604681595
transform 1 0 7636 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_77
timestamp 1604681595
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_82
timestamp 1604681595
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9844 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_86
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_91
timestamp 1604681595
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_114
timestamp 1604681595
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_118
timestamp 1604681595
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_126
timestamp 1604681595
transform 1 0 12696 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_138
timestamp 1604681595
transform 1 0 13800 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_150
timestamp 1604681595
transform 1 0 14904 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_162
timestamp 1604681595
transform 1 0 16008 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18216 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_174
timestamp 1604681595
transform 1 0 17112 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1604681595
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18400 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19688 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19136 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_194
timestamp 1604681595
transform 1 0 18952 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1604681595
transform 1 0 19320 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_208
timestamp 1604681595
transform 1 0 20240 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20424 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_212
timestamp 1604681595
transform 1 0 20608 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_224
timestamp 1604681595
transform 1 0 21712 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_236
timestamp 1604681595
transform 1 0 22816 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_257
timestamp 1604681595
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_269
timestamp 1604681595
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1604681595
transform 1 0 2944 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2392 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_12
timestamp 1604681595
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_16
timestamp 1604681595
transform 1 0 2576 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1604681595
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5980 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 6348 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_51
timestamp 1604681595
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_55
timestamp 1604681595
transform 1 0 6164 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_59
timestamp 1604681595
transform 1 0 6532 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_64
timestamp 1604681595
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_68
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_72
timestamp 1604681595
transform 1 0 7728 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10396 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9292 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_84
timestamp 1604681595
transform 1 0 8832 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_88
timestamp 1604681595
transform 1 0 9200 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1604681595
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_99
timestamp 1604681595
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_103
timestamp 1604681595
transform 1 0 10580 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11040 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 10856 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_127
timestamp 1604681595
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_131
timestamp 1604681595
transform 1 0 13156 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_143
timestamp 1604681595
transform 1 0 14260 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1604681595
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1604681595
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17940 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_178
timestamp 1604681595
transform 1 0 17480 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_182
timestamp 1604681595
transform 1 0 17848 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_189
timestamp 1604681595
transform 1 0 18492 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_201
timestamp 1604681595
transform 1 0 19596 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1604681595
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1604681595
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1604681595
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_251
timestamp 1604681595
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_263
timestamp 1604681595
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 2116 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4876 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_30
timestamp 1604681595
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_34
timestamp 1604681595
transform 1 0 4232 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_38
timestamp 1604681595
transform 1 0 4600 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_53
timestamp 1604681595
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1604681595
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_81
timestamp 1604681595
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9292 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_85
timestamp 1604681595
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_108
timestamp 1604681595
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_112
timestamp 1604681595
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_116
timestamp 1604681595
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_142
timestamp 1604681595
transform 1 0 14168 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_154
timestamp 1604681595
transform 1 0 15272 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_166
timestamp 1604681595
transform 1 0 16376 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_178
timestamp 1604681595
transform 1 0 17480 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_182
timestamp 1604681595
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1604681595
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_208
timestamp 1604681595
transform 1 0 20240 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_214
timestamp 1604681595
transform 1 0 20792 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_217
timestamp 1604681595
transform 1 0 21068 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_229
timestamp 1604681595
transform 1 0 22172 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_241
timestamp 1604681595
transform 1 0 23276 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1604681595
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1604681595
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2392 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_12
timestamp 1604681595
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_16
timestamp 1604681595
transform 1 0 2576 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_20
timestamp 1604681595
transform 1 0 2944 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3128 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1604681595
transform 1 0 3312 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_28
timestamp 1604681595
transform 1 0 3680 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_41
timestamp 1604681595
transform 1 0 4876 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 5704 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_46
timestamp 1604681595
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1604681595
transform 1 0 8188 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 7636 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8648 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_69
timestamp 1604681595
transform 1 0 7452 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_73
timestamp 1604681595
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_80
timestamp 1604681595
transform 1 0 8464 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_84
timestamp 1604681595
transform 1 0 8832 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_89
timestamp 1604681595
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1604681595
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11592 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 11224 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_106
timestamp 1604681595
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_113
timestamp 1604681595
transform 1 0 11500 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_123
timestamp 1604681595
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_127
timestamp 1604681595
transform 1 0 12788 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_139
timestamp 1604681595
transform 1 0 13892 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1604681595
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1604681595
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1604681595
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_190
timestamp 1604681595
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_202
timestamp 1604681595
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1604681595
transform 1 0 21436 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1604681595
transform 1 0 22540 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_245
timestamp 1604681595
transform 1 0 23644 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_257
timestamp 1604681595
transform 1 0 24748 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_269
timestamp 1604681595
transform 1 0 25852 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1604681595
transform 1 0 2944 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 2760 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_12
timestamp 1604681595
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_16
timestamp 1604681595
transform 1 0 2576 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_26
timestamp 1604681595
transform 1 0 3496 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_22
timestamp 1604681595
transform 1 0 3128 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3312 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1604681595
transform 1 0 3956 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 4232 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_34
timestamp 1604681595
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 4600 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_38
timestamp 1604681595
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_36
timestamp 1604681595
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4784 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_49
timestamp 1604681595
transform 1 0 5612 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_42
timestamp 1604681595
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_60
timestamp 1604681595
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_53
timestamp 1604681595
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1604681595
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1604681595
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 6164 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 6348 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1604681595
transform 1 0 8556 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7268 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6992 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8004 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6992 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_66
timestamp 1604681595
transform 1 0 7176 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_73
timestamp 1604681595
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_77
timestamp 1604681595
transform 1 0 8188 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_86
timestamp 1604681595
transform 1 0 9016 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1604681595
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_88
timestamp 1604681595
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9292 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_91
timestamp 1604681595
transform 1 0 9476 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_102
timestamp 1604681595
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_99
timestamp 1604681595
transform 1 0 10212 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_95
timestamp 1604681595
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10488 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10672 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_110
timestamp 1604681595
transform 1 0 11224 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_106
timestamp 1604681595
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1604681595
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1604681595
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_117
timestamp 1604681595
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 12052 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11408 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_20_135
timestamp 1604681595
transform 1 0 13524 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_131
timestamp 1604681595
transform 1 0 13156 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_126
timestamp 1604681595
transform 1 0 12696 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12880 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 13340 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_142
timestamp 1604681595
transform 1 0 14168 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 13708 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _56_
timestamp 1604681595
transform 1 0 13892 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_142
timestamp 1604681595
transform 1 0 14168 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_130
timestamp 1604681595
transform 1 0 13064 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15916 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15824 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14904 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_154
timestamp 1604681595
transform 1 0 15272 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_160
timestamp 1604681595
transform 1 0 15824 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1604681595
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_154
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_162
timestamp 1604681595
transform 1 0 16008 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_168
timestamp 1604681595
transform 1 0 16560 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_175
timestamp 1604681595
transform 1 0 17204 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_171
timestamp 1604681595
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_167
timestamp 1604681595
transform 1 0 16468 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16652 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_187
timestamp 1604681595
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_175
timestamp 1604681595
transform 1 0 17204 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18768 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_190
timestamp 1604681595
transform 1 0 18584 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_194
timestamp 1604681595
transform 1 0 18952 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_206
timestamp 1604681595
transform 1 0 20056 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_199
timestamp 1604681595
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_218
timestamp 1604681595
transform 1 0 21160 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_211
timestamp 1604681595
transform 1 0 20516 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_227
timestamp 1604681595
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_230
timestamp 1604681595
transform 1 0 22264 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_242
timestamp 1604681595
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_245
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_239
timestamp 1604681595
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_257
timestamp 1604681595
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_269
timestamp 1604681595
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_251
timestamp 1604681595
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_263
timestamp 1604681595
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 1472 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 2484 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_13
timestamp 1604681595
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_17
timestamp 1604681595
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 3036 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 4600 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_30
timestamp 1604681595
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_34
timestamp 1604681595
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_41
timestamp 1604681595
transform 1 0 4876 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1604681595
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1604681595
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 8372 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1604681595
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_75
timestamp 1604681595
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10396 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 9936 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9752 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_88
timestamp 1604681595
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_92
timestamp 1604681595
transform 1 0 9568 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_99
timestamp 1604681595
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1604681595
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1604681595
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_142
timestamp 1604681595
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14904 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14720 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_146
timestamp 1604681595
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1604681595
transform 1 0 16652 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1604681595
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1604681595
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1604681595
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_220
timestamp 1604681595
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_232
timestamp 1604681595
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_245
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_257
timestamp 1604681595
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_269
timestamp 1604681595
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_6
timestamp 1604681595
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_10
timestamp 1604681595
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4784 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 4416 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_38
timestamp 1604681595
transform 1 0 4600 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4968 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_22_61
timestamp 1604681595
transform 1 0 6716 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7544 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 8556 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6900 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_65
timestamp 1604681595
transform 1 0 7084 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_79
timestamp 1604681595
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_83
timestamp 1604681595
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1604681595
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8924 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 9108 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_103
timestamp 1604681595
transform 1 0 10580 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_100
timestamp 1604681595
transform 1 0 10304 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_96
timestamp 1604681595
transform 1 0 9936 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10396 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10672 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 12236 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11684 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_113
timestamp 1604681595
transform 1 0 11500 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_117
timestamp 1604681595
transform 1 0 11868 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_124
timestamp 1604681595
transform 1 0 12512 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12696 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1604681595
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15824 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15456 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1604681595
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_158
timestamp 1604681595
transform 1 0 15640 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1604681595
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1604681595
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1604681595
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1604681595
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_227
timestamp 1604681595
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_239
timestamp 1604681595
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_251
timestamp 1604681595
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_263
timestamp 1604681595
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2208 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_7
timestamp 1604681595
transform 1 0 1748 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4140 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1604681595
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_21
timestamp 1604681595
transform 1 0 3036 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_25
timestamp 1604681595
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_29
timestamp 1604681595
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6072 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_52
timestamp 1604681595
transform 1 0 5888 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_56
timestamp 1604681595
transform 1 0 6256 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 8004 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 7452 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_66
timestamp 1604681595
transform 1 0 7176 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_71
timestamp 1604681595
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_94
timestamp 1604681595
transform 1 0 9752 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_98
timestamp 1604681595
transform 1 0 10120 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_101
timestamp 1604681595
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12512 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_114
timestamp 1604681595
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1604681595
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 14352 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14168 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13524 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_133
timestamp 1604681595
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_137
timestamp 1604681595
transform 1 0 13708 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_141
timestamp 1604681595
transform 1 0 14076 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16284 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_163
timestamp 1604681595
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_167
timestamp 1604681595
transform 1 0 16468 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1604681595
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1604681595
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1604681595
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_220
timestamp 1604681595
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_232
timestamp 1604681595
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1604681595
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_269
timestamp 1604681595
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 1472 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4692 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_23
timestamp 1604681595
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_36
timestamp 1604681595
transform 1 0 4416 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_41
timestamp 1604681595
transform 1 0 4876 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 5336 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 7820 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7268 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_65
timestamp 1604681595
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_69
timestamp 1604681595
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10396 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_99
timestamp 1604681595
transform 1 0 10212 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_103
timestamp 1604681595
transform 1 0 10580 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 12512 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10948 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12052 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_116
timestamp 1604681595
transform 1 0 11776 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_121
timestamp 1604681595
transform 1 0 12236 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_143
timestamp 1604681595
transform 1 0 14260 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_147
timestamp 1604681595
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1604681595
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_163
timestamp 1604681595
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_175
timestamp 1604681595
transform 1 0 17204 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_187
timestamp 1604681595
transform 1 0 18308 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_199
timestamp 1604681595
transform 1 0 19412 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_211
timestamp 1604681595
transform 1 0 20516 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_227
timestamp 1604681595
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_239
timestamp 1604681595
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_251
timestamp 1604681595
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_263
timestamp 1604681595
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 2668 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_7
timestamp 1604681595
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_11
timestamp 1604681595
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_15
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 4692 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_36
timestamp 1604681595
transform 1 0 4416 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_41
timestamp 1604681595
transform 1 0 4876 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6256 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1604681595
transform 1 0 5980 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_58
timestamp 1604681595
transform 1 0 6440 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8372 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 7268 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_65
timestamp 1604681595
transform 1 0 7084 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 1604681595
transform 1 0 7452 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_75
timestamp 1604681595
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_99
timestamp 1604681595
transform 1 0 10212 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12052 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_114
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_118
timestamp 1604681595
transform 1 0 11960 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1604681595
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 13800 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 13156 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_129
timestamp 1604681595
transform 1 0 12972 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_133
timestamp 1604681595
transform 1 0 13340 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16284 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_157
timestamp 1604681595
transform 1 0 15548 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_171
timestamp 1604681595
transform 1 0 16836 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_175
timestamp 1604681595
transform 1 0 17204 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1604681595
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1604681595
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_220
timestamp 1604681595
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_232
timestamp 1604681595
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_245
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_257
timestamp 1604681595
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_269
timestamp 1604681595
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_7
timestamp 1604681595
transform 1 0 1748 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 1932 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 1564 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_16
timestamp 1604681595
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_12
timestamp 1604681595
transform 1 0 2208 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2116 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_27_20
timestamp 1604681595
transform 1 0 2944 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_20
timestamp 1604681595
transform 1 0 2944 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_25
timestamp 1604681595
transform 1 0 3404 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_28
timestamp 1604681595
transform 1 0 3680 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1604681595
transform 1 0 3312 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3128 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 3588 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_36
timestamp 1604681595
transform 1 0 4416 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4232 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4692 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 3772 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_27_48
timestamp 1604681595
transform 1 0 5520 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_48
timestamp 1604681595
transform 1 0 5520 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5704 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_58
timestamp 1604681595
transform 1 0 6440 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1604681595
transform 1 0 6072 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_52
timestamp 1604681595
transform 1 0 5888 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6256 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 5888 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 6072 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6256 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7360 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7820 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8648 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 7176 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7636 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_65
timestamp 1604681595
transform 1 0 7084 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_69
timestamp 1604681595
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_91
timestamp 1604681595
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_87
timestamp 1604681595
transform 1 0 9108 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1604681595
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 9292 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9660 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9936 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10120 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 9844 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_114
timestamp 1604681595
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_111
timestamp 1604681595
transform 1 0 11316 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_107
timestamp 1604681595
transform 1 0 10948 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11500 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11132 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_118
timestamp 1604681595
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_115
timestamp 1604681595
transform 1 0 11684 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11868 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12052 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12604 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_127
timestamp 1604681595
transform 1 0 12788 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_134
timestamp 1604681595
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_128
timestamp 1604681595
transform 1 0 12880 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13248 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13064 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13248 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_141
timestamp 1604681595
transform 1 0 14076 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_138
timestamp 1604681595
transform 1 0 13800 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 14260 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 13616 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_145
timestamp 1604681595
transform 1 0 14444 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_145
timestamp 1604681595
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 14812 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14628 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_149
timestamp 1604681595
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1604681595
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1604681595
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_168
timestamp 1604681595
transform 1 0 16560 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_180
timestamp 1604681595
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1604681595
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1604681595
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1604681595
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1604681595
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1604681595
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1604681595
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1604681595
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1604681595
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_251
timestamp 1604681595
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1604681595
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1604681595
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_269
timestamp 1604681595
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 1840 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_6
timestamp 1604681595
transform 1 0 1656 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_10
timestamp 1604681595
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_23
timestamp 1604681595
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_41
timestamp 1604681595
transform 1 0 4876 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 5888 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5060 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5428 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_45
timestamp 1604681595
transform 1 0 5244 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_49
timestamp 1604681595
transform 1 0 5612 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1604681595
transform 1 0 8556 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8372 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_71
timestamp 1604681595
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_75
timestamp 1604681595
transform 1 0 8004 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_84
timestamp 1604681595
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_88
timestamp 1604681595
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_102
timestamp 1604681595
transform 1 0 10488 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 11224 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10764 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_107
timestamp 1604681595
transform 1 0 10948 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604681595
transform 1 0 13708 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13248 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14168 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_129
timestamp 1604681595
transform 1 0 12972 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_134
timestamp 1604681595
transform 1 0 13432 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_140
timestamp 1604681595
transform 1 0 13984 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_144
timestamp 1604681595
transform 1 0 14352 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14812 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_148
timestamp 1604681595
transform 1 0 14720 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1604681595
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1604681595
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1604681595
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1604681595
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1604681595
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1604681595
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1604681595
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_251
timestamp 1604681595
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_263
timestamp 1604681595
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 2208 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 2024 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1604681595
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_7
timestamp 1604681595
transform 1 0 1748 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4692 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4508 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1604681595
transform 1 0 4140 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_31
timestamp 1604681595
transform 1 0 3956 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_35
timestamp 1604681595
transform 1 0 4324 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5704 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_48
timestamp 1604681595
transform 1 0 5520 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_52
timestamp 1604681595
transform 1 0 5888 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1604681595
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8372 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8188 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_71
timestamp 1604681595
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_75
timestamp 1604681595
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9936 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9752 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9384 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_88
timestamp 1604681595
transform 1 0 9200 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_92
timestamp 1604681595
transform 1 0 9568 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_105
timestamp 1604681595
transform 1 0 10764 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11040 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1604681595
transform 1 0 11224 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_114
timestamp 1604681595
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 11684 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604681595
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12604 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13340 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12972 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_127
timestamp 1604681595
transform 1 0 12788 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_131
timestamp 1604681595
transform 1 0 13156 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_152
timestamp 1604681595
transform 1 0 15088 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_164
timestamp 1604681595
transform 1 0 16192 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_176
timestamp 1604681595
transform 1 0 17296 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_182
timestamp 1604681595
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1604681595
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1604681595
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1604681595
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1604681595
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1604681595
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_269
timestamp 1604681595
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2208 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1932 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1604681595
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_11
timestamp 1604681595
transform 1 0 2116 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_25
timestamp 1604681595
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_21
timestamp 1604681595
transform 1 0 3036 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1604681595
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1604681595
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_40
timestamp 1604681595
transform 1 0 4784 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_36
timestamp 1604681595
transform 1 0 4416 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 4600 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5244 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_44
timestamp 1604681595
transform 1 0 5152 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7820 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7176 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_64
timestamp 1604681595
transform 1 0 6992 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_68
timestamp 1604681595
transform 1 0 7360 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1604681595
transform 1 0 8648 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9936 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_86
timestamp 1604681595
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1604681595
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_102
timestamp 1604681595
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 11408 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 11224 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_106
timestamp 1604681595
transform 1 0 10856 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_121
timestamp 1604681595
transform 1 0 12236 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_125
timestamp 1604681595
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12972 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12788 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13984 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14352 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1604681595
transform 1 0 13800 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_142
timestamp 1604681595
transform 1 0 14168 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15456 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14720 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_146
timestamp 1604681595
transform 1 0 14536 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_150
timestamp 1604681595
transform 1 0 14904 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_158
timestamp 1604681595
transform 1 0 15640 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_170
timestamp 1604681595
transform 1 0 16744 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_182
timestamp 1604681595
transform 1 0 17848 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_194
timestamp 1604681595
transform 1 0 18952 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_206
timestamp 1604681595
transform 1 0 20056 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1604681595
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1604681595
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1604681595
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1604681595
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 2024 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 1840 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_7
timestamp 1604681595
transform 1 0 1748 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 4692 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4508 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4140 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_29
timestamp 1604681595
transform 1 0 3772 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_35
timestamp 1604681595
transform 1 0 4324 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4968 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_51
timestamp 1604681595
transform 1 0 5796 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_55
timestamp 1604681595
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _52_
timestamp 1604681595
transform 1 0 6992 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 8004 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7452 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_67
timestamp 1604681595
transform 1 0 7268 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_71
timestamp 1604681595
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _51_
timestamp 1604681595
transform 1 0 10488 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9936 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 10304 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_94
timestamp 1604681595
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_98
timestamp 1604681595
transform 1 0 10120 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_109
timestamp 1604681595
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_105
timestamp 1604681595
transform 1 0 10764 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11316 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10948 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 11500 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_116
timestamp 1604681595
transform 1 0 11776 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12512 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 14352 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13524 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 14168 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_133
timestamp 1604681595
transform 1 0 13340 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_137
timestamp 1604681595
transform 1 0 13708 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_141
timestamp 1604681595
transform 1 0 14076 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 16284 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_163
timestamp 1604681595
transform 1 0 16100 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_167
timestamp 1604681595
transform 1 0 16468 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_179
timestamp 1604681595
transform 1 0 17572 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1604681595
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1604681595
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1604681595
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1604681595
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_269
timestamp 1604681595
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 2760 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 2576 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_10
timestamp 1604681595
transform 1 0 2024 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_14
timestamp 1604681595
transform 1 0 2392 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_22
timestamp 1604681595
transform 1 0 3128 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1604681595
transform 1 0 3312 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_30
timestamp 1604681595
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1604681595
transform 1 0 3496 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 3680 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_35
timestamp 1604681595
transform 1 0 4324 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _57_
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 4692 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_41
timestamp 1604681595
transform 1 0 4876 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5060 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_32_62
timestamp 1604681595
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 7728 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 7544 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6992 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_66
timestamp 1604681595
transform 1 0 7176 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_88
timestamp 1604681595
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_84
timestamp 1604681595
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_97
timestamp 1604681595
transform 1 0 10028 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9844 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10212 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10396 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12512 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_120
timestamp 1604681595
transform 1 0 12144 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12880 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13892 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14260 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_126
timestamp 1604681595
transform 1 0 12696 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_137
timestamp 1604681595
transform 1 0 13708 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1604681595
transform 1 0 14076 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_145
timestamp 1604681595
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_149
timestamp 1604681595
transform 1 0 14812 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_173
timestamp 1604681595
transform 1 0 17020 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_185
timestamp 1604681595
transform 1 0 18124 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1604681595
transform 1 0 19228 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_209
timestamp 1604681595
transform 1 0 20332 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1604681595
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1604681595
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1604681595
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_251
timestamp 1604681595
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_263
timestamp 1604681595
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_9
timestamp 1604681595
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_17
timestamp 1604681595
transform 1 0 2668 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_14
timestamp 1604681595
transform 1 0 2392 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_10
timestamp 1604681595
transform 1 0 2024 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_13
timestamp 1604681595
transform 1 0 2300 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2668 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 2760 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_26
timestamp 1604681595
transform 1 0 3496 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_22
timestamp 1604681595
transform 1 0 3128 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_30
timestamp 1604681595
transform 1 0 3864 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_26
timestamp 1604681595
transform 1 0 3496 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3312 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3680 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 4048 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4232 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_34_51
timestamp 1604681595
transform 1 0 5796 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_53
timestamp 1604681595
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604681595
transform 1 0 5980 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_55
timestamp 1604681595
transform 1 0 6164 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1604681595
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 6348 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_59
timestamp 1604681595
transform 1 0 6532 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 6808 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7728 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7084 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 7544 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7084 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_67
timestamp 1604681595
transform 1 0 7268 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_88
timestamp 1604681595
transform 1 0 9200 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_84
timestamp 1604681595
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_91
timestamp 1604681595
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_34_99
timestamp 1604681595
transform 1 0 10212 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_95
timestamp 1604681595
transform 1 0 9844 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10028 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10488 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10212 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_34_104
timestamp 1604681595
transform 1 0 10672 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_112
timestamp 1604681595
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_108
timestamp 1604681595
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_123
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_116
timestamp 1604681595
transform 1 0 11776 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12604 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10948 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_34_133
timestamp 1604681595
transform 1 0 13340 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_130
timestamp 1604681595
transform 1 0 13064 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_126
timestamp 1604681595
transform 1 0 12696 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_127
timestamp 1604681595
transform 1 0 12788 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13156 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12972 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13156 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_33_144
timestamp 1604681595
transform 1 0 14352 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_140
timestamp 1604681595
transform 1 0 13984 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14168 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_145
timestamp 1604681595
transform 1 0 14444 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_149
timestamp 1604681595
transform 1 0 14812 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14536 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_161
timestamp 1604681595
transform 1 0 15916 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_157
timestamp 1604681595
transform 1 0 15548 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15732 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _58_
timestamp 1604681595
transform 1 0 16284 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 14720 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_167
timestamp 1604681595
transform 1 0 16468 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_179
timestamp 1604681595
transform 1 0 17572 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_168
timestamp 1604681595
transform 1 0 16560 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_180
timestamp 1604681595
transform 1 0 17664 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1604681595
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1604681595
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_192
timestamp 1604681595
transform 1 0 18768 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_204
timestamp 1604681595
transform 1 0 19872 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_220
timestamp 1604681595
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_212
timestamp 1604681595
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604681595
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_232
timestamp 1604681595
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1604681595
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1604681595
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_269
timestamp 1604681595
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_251
timestamp 1604681595
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1604681595
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2760 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 2208 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2576 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_10
timestamp 1604681595
transform 1 0 2024 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_14
timestamp 1604681595
transform 1 0 2392 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4324 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4140 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_31
timestamp 1604681595
transform 1 0 3956 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_44
timestamp 1604681595
transform 1 0 5152 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_48
timestamp 1604681595
transform 1 0 5520 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 5336 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_52
timestamp 1604681595
transform 1 0 5888 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 5704 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6072 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 6256 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1604681595
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7636 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7452 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7084 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 8648 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_67
timestamp 1604681595
transform 1 0 7268 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_80
timestamp 1604681595
transform 1 0 8464 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _50_
timestamp 1604681595
transform 1 0 9476 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10488 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10304 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9016 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9936 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_84
timestamp 1604681595
transform 1 0 8832 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_88
timestamp 1604681595
transform 1 0 9200 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_94
timestamp 1604681595
transform 1 0 9752 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_98
timestamp 1604681595
transform 1 0 10120 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 12052 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11500 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 11868 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_111
timestamp 1604681595
transform 1 0 11316 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_115
timestamp 1604681595
transform 1 0 11684 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_123
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13064 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13800 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14168 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12880 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_127
timestamp 1604681595
transform 1 0 12788 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_136
timestamp 1604681595
transform 1 0 13616 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_140
timestamp 1604681595
transform 1 0 13984 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_144
timestamp 1604681595
transform 1 0 14352 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14536 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_35_165
timestamp 1604681595
transform 1 0 16284 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_177
timestamp 1604681595
transform 1 0 17388 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1604681595
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1604681595
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_220
timestamp 1604681595
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_232
timestamp 1604681595
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_245
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_257
timestamp 1604681595
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_269
timestamp 1604681595
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 2484 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1932 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2300 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_7
timestamp 1604681595
transform 1 0 1748 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_11
timestamp 1604681595
transform 1 0 2116 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_19
timestamp 1604681595
transform 1 0 2852 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4324 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3036 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_23
timestamp 1604681595
transform 1 0 3220 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_27
timestamp 1604681595
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_32
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 5888 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6808 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 5336 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 5704 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6440 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_44
timestamp 1604681595
transform 1 0 5152 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_48
timestamp 1604681595
transform 1 0 5520 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_56
timestamp 1604681595
transform 1 0 6256 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_60
timestamp 1604681595
transform 1 0 6624 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7084 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_36_64
timestamp 1604681595
transform 1 0 6992 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10488 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_84
timestamp 1604681595
transform 1 0 8832 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_88
timestamp 1604681595
transform 1 0 9200 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_99
timestamp 1604681595
transform 1 0 10212 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_104
timestamp 1604681595
transform 1 0 10672 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10948 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13432 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13248 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12880 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_126
timestamp 1604681595
transform 1 0 12696 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_130
timestamp 1604681595
transform 1 0 13064 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_143
timestamp 1604681595
transform 1 0 14260 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14536 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_148
timestamp 1604681595
transform 1 0 14720 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_152
timestamp 1604681595
transform 1 0 15088 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_160
timestamp 1604681595
transform 1 0 15824 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_172
timestamp 1604681595
transform 1 0 16928 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_184
timestamp 1604681595
transform 1 0 18032 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_196
timestamp 1604681595
transform 1 0 19136 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_208
timestamp 1604681595
transform 1 0 20240 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_227
timestamp 1604681595
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_239
timestamp 1604681595
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_251
timestamp 1604681595
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_263
timestamp 1604681595
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 2944 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 2760 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 2392 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_10
timestamp 1604681595
transform 1 0 2024 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_16
timestamp 1604681595
transform 1 0 2576 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 4876 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_39
timestamp 1604681595
transform 1 0 4692 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 5428 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604681595
transform 1 0 5244 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_43
timestamp 1604681595
transform 1 0 5060 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1604681595
transform 1 0 5796 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1604681595
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8372 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_71
timestamp 1604681595
transform 1 0 7636 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_75
timestamp 1604681595
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10304 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10120 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9752 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9384 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_88
timestamp 1604681595
transform 1 0 9200 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_92
timestamp 1604681595
transform 1 0 9568 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_96
timestamp 1604681595
transform 1 0 9936 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12512 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11316 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11684 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_109
timestamp 1604681595
transform 1 0 11132 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1604681595
transform 1 0 11500 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_117
timestamp 1604681595
transform 1 0 11868 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_123
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 14076 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13248 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13616 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_130
timestamp 1604681595
transform 1 0 13064 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_134
timestamp 1604681595
transform 1 0 13432 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_138
timestamp 1604681595
transform 1 0 13800 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16008 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_160
timestamp 1604681595
transform 1 0 15824 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1604681595
transform 1 0 16192 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__93__A
timestamp 1604681595
transform 1 0 17664 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__96__A
timestamp 1604681595
transform 1 0 16560 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_170
timestamp 1604681595
transform 1 0 16744 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_178
timestamp 1604681595
transform 1 0 17480 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_182
timestamp 1604681595
transform 1 0 17848 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__90__A
timestamp 1604681595
transform 1 0 19412 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_196
timestamp 1604681595
transform 1 0 19136 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_201
timestamp 1604681595
transform 1 0 19596 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20884 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_213
timestamp 1604681595
transform 1 0 20700 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_217
timestamp 1604681595
transform 1 0 21068 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_229
timestamp 1604681595
transform 1 0 22172 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_241
timestamp 1604681595
transform 1 0 23276 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_245
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_257
timestamp 1604681595
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_269
timestamp 1604681595
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 2852 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2576 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_11
timestamp 1604681595
transform 1 0 2116 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_15
timestamp 1604681595
transform 1 0 2484 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_18
timestamp 1604681595
transform 1 0 2760 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4416 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 4232 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_23
timestamp 1604681595
transform 1 0 3220 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_27
timestamp 1604681595
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_32
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6348 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6808 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_55
timestamp 1604681595
transform 1 0 6164 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_59
timestamp 1604681595
transform 1 0 6532 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7084 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_38_64
timestamp 1604681595
transform 1 0 6992 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _49_
timestamp 1604681595
transform 1 0 9752 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10580 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 10212 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_84
timestamp 1604681595
transform 1 0 8832 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_97
timestamp 1604681595
transform 1 0 10028 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_101
timestamp 1604681595
transform 1 0 10396 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10764 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_38_124
timestamp 1604681595
transform 1 0 12512 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13248 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14260 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12696 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_128
timestamp 1604681595
transform 1 0 12880 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1604681595
transform 1 0 14076 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_145
timestamp 1604681595
transform 1 0 14444 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_149
timestamp 1604681595
transform 1 0 14812 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_160
timestamp 1604681595
transform 1 0 15824 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _93_
timestamp 1604681595
transform 1 0 17664 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _96_
timestamp 1604681595
transform 1 0 16560 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_172
timestamp 1604681595
transform 1 0 16928 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_184
timestamp 1604681595
transform 1 0 18032 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _90_
timestamp 1604681595
transform 1 0 19412 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_196
timestamp 1604681595
transform 1 0 19136 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_203
timestamp 1604681595
transform 1 0 19780 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_211
timestamp 1604681595
transform 1 0 20516 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_221
timestamp 1604681595
transform 1 0 21436 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_233
timestamp 1604681595
transform 1 0 22540 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_245
timestamp 1604681595
transform 1 0 23644 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_257
timestamp 1604681595
transform 1 0 24748 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_269
timestamp 1604681595
transform 1 0 25852 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_7
timestamp 1604681595
transform 1 0 1748 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604681595
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_18
timestamp 1604681595
transform 1 0 2760 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_15
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_11
timestamp 1604681595
transform 1 0 2116 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_11
timestamp 1604681595
transform 1 0 2116 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 2576 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2392 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2576 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 2852 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1604681595
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_23
timestamp 1604681595
transform 1 0 3220 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_29
timestamp 1604681595
transform 1 0 3772 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_25
timestamp 1604681595
transform 1 0 3404 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 3588 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_40
timestamp 1604681595
transform 1 0 4784 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_36
timestamp 1604681595
transform 1 0 4416 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 4048 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4600 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4232 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_40_44
timestamp 1604681595
transform 1 0 5152 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 4968 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5520 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_61
timestamp 1604681595
transform 1 0 6716 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_57
timestamp 1604681595
transform 1 0 6348 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1604681595
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_53
timestamp 1604681595
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6532 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _53_
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7820 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7084 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6900 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7636 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7268 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_65
timestamp 1604681595
transform 1 0 7084 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_69
timestamp 1604681595
transform 1 0 7452 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_84
timestamp 1604681595
transform 1 0 8832 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_92
timestamp 1604681595
transform 1 0 9568 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_102
timestamp 1604681595
transform 1 0 10488 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_99
timestamp 1604681595
transform 1 0 10212 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_101
timestamp 1604681595
transform 1 0 10396 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_97
timestamp 1604681595
transform 1 0 10028 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9844 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10304 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10212 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10580 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12512 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_114
timestamp 1604681595
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 1604681595
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_122
timestamp 1604681595
transform 1 0 12328 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _48_
timestamp 1604681595
transform 1 0 13248 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__99__A
timestamp 1604681595
transform 1 0 14352 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_142
timestamp 1604681595
transform 1 0 14168 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_126
timestamp 1604681595
transform 1 0 12696 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_135
timestamp 1604681595
transform 1 0 13524 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_152
timestamp 1604681595
transform 1 0 15088 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_147
timestamp 1604681595
transform 1 0 14628 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_146
timestamp 1604681595
transform 1 0 14536 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14904 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14720 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _99_
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_158
timestamp 1604681595
transform 1 0 15640 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _97_
timestamp 1604681595
transform 1 0 16376 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14904 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_40_170
timestamp 1604681595
transform 1 0 16744 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_173
timestamp 1604681595
transform 1 0 17020 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1604681595
transform 1 0 16652 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__97__A
timestamp 1604681595
transform 1 0 16836 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_182
timestamp 1604681595
transform 1 0 17848 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_180
timestamp 1604681595
transform 1 0 17664 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_177
timestamp 1604681595
transform 1 0 17388 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__95__A
timestamp 1604681595
transform 1 0 17480 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _95_
timestamp 1604681595
transform 1 0 17480 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _94_
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_190
timestamp 1604681595
transform 1 0 18584 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_192
timestamp 1604681595
transform 1 0 18768 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_188
timestamp 1604681595
transform 1 0 18400 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__91__A
timestamp 1604681595
transform 1 0 18952 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__94__A
timestamp 1604681595
transform 1 0 18584 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _92_
timestamp 1604681595
transform 1 0 19136 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _91_
timestamp 1604681595
transform 1 0 18860 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_204
timestamp 1604681595
transform 1 0 19872 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_200
timestamp 1604681595
transform 1 0 19504 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__92__A
timestamp 1604681595
transform 1 0 19688 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _89_
timestamp 1604681595
transform 1 0 20240 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1604681595
transform 1 0 19228 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_213
timestamp 1604681595
transform 1 0 20700 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_209
timestamp 1604681595
transform 1 0 20332 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_216
timestamp 1604681595
transform 1 0 20976 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_212
timestamp 1604681595
transform 1 0 20608 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__88__A
timestamp 1604681595
transform 1 0 21160 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__89__A
timestamp 1604681595
transform 1 0 20792 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _88_
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_228
timestamp 1604681595
transform 1 0 22080 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_224
timestamp 1604681595
transform 1 0 21712 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__87__A
timestamp 1604681595
transform 1 0 21896 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _87_
timestamp 1604681595
transform 1 0 21344 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_219
timestamp 1604681595
transform 1 0 21252 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1604681595
transform 1 0 22448 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__86__A
timestamp 1604681595
transform 1 0 23000 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_236
timestamp 1604681595
transform 1 0 22816 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_240
timestamp 1604681595
transform 1 0 23184 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_245
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_231
timestamp 1604681595
transform 1 0 22356 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_243
timestamp 1604681595
transform 1 0 23460 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_257
timestamp 1604681595
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_269
timestamp 1604681595
transform 1 0 25852 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_255
timestamp 1604681595
transform 1 0 24564 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_267
timestamp 1604681595
transform 1 0 25668 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 2852 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 2300 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604681595
transform 1 0 2668 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_11
timestamp 1604681595
transform 1 0 2116 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_15
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4600 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4416 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604681595
transform 1 0 3404 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604681595
transform 1 0 4048 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_23
timestamp 1604681595
transform 1 0 3220 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_27
timestamp 1604681595
transform 1 0 3588 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_31
timestamp 1604681595
transform 1 0 3956 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_34
timestamp 1604681595
transform 1 0 4232 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604681595
transform 1 0 5612 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_47
timestamp 1604681595
transform 1 0 5428 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1604681595
transform 1 0 5796 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1604681595
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _54_
timestamp 1604681595
transform 1 0 8464 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6900 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7912 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8280 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_72
timestamp 1604681595
transform 1 0 7728 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_76
timestamp 1604681595
transform 1 0 8096 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_83
timestamp 1604681595
transform 1 0 8740 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10304 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10120 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_95
timestamp 1604681595
transform 1 0 9844 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_109
timestamp 1604681595
transform 1 0 11132 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_115
timestamp 1604681595
transform 1 0 11684 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_118
timestamp 1604681595
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_132
timestamp 1604681595
transform 1 0 13248 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_144
timestamp 1604681595
transform 1 0 14352 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _98_
timestamp 1604681595
transform 1 0 15180 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__98__A
timestamp 1604681595
transform 1 0 15732 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_152
timestamp 1604681595
transform 1 0 15088 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_157
timestamp 1604681595
transform 1 0 15548 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_161
timestamp 1604681595
transform 1 0 15916 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_173
timestamp 1604681595
transform 1 0 17020 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_181
timestamp 1604681595
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1604681595
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1604681595
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_220
timestamp 1604681595
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_232
timestamp 1604681595
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1604681595
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_269
timestamp 1604681595
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 2484 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1932 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2300 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_7
timestamp 1604681595
transform 1 0 1748 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_11
timestamp 1604681595
transform 1 0 2116 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_19
timestamp 1604681595
transform 1 0 2852 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4600 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_36
timestamp 1604681595
transform 1 0 4416 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_40
timestamp 1604681595
transform 1 0 4784 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 5152 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_48
timestamp 1604681595
transform 1 0 5520 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_60
timestamp 1604681595
transform 1 0 6624 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _55_
timestamp 1604681595
transform 1 0 8004 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_67
timestamp 1604681595
transform 1 0 7268 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_78
timestamp 1604681595
transform 1 0 8280 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _59_
timestamp 1604681595
transform 1 0 9752 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10304 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_90
timestamp 1604681595
transform 1 0 9384 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_97
timestamp 1604681595
transform 1 0 10028 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_102
timestamp 1604681595
transform 1 0 10488 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_114
timestamp 1604681595
transform 1 0 11592 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_122
timestamp 1604681595
transform 1 0 12328 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_125
timestamp 1604681595
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_137
timestamp 1604681595
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_149
timestamp 1604681595
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1604681595
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1604681595
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_180
timestamp 1604681595
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_187
timestamp 1604681595
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_199
timestamp 1604681595
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_211
timestamp 1604681595
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_218
timestamp 1604681595
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_230
timestamp 1604681595
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_242
timestamp 1604681595
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_249
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_261
timestamp 1604681595
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_273
timestamp 1604681595
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal3 s 27520 14016 28000 14136 6 ccff_head
port 0 nsew default input
rlabel metal2 s 20994 0 21050 480 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_in[0]
port 2 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[10]
port 3 nsew default input
rlabel metal3 s 0 10616 480 10736 6 chanx_left_in[11]
port 4 nsew default input
rlabel metal3 s 0 11160 480 11280 6 chanx_left_in[12]
port 5 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_in[13]
port 6 nsew default input
rlabel metal3 s 0 12384 480 12504 6 chanx_left_in[14]
port 7 nsew default input
rlabel metal3 s 0 13064 480 13184 6 chanx_left_in[15]
port 8 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chanx_left_in[16]
port 9 nsew default input
rlabel metal3 s 0 14288 480 14408 6 chanx_left_in[17]
port 10 nsew default input
rlabel metal3 s 0 14832 480 14952 6 chanx_left_in[18]
port 11 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chanx_left_in[19]
port 12 nsew default input
rlabel metal3 s 0 4496 480 4616 6 chanx_left_in[1]
port 13 nsew default input
rlabel metal3 s 0 5040 480 5160 6 chanx_left_in[2]
port 14 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[3]
port 15 nsew default input
rlabel metal3 s 0 6264 480 6384 6 chanx_left_in[4]
port 16 nsew default input
rlabel metal3 s 0 6944 480 7064 6 chanx_left_in[5]
port 17 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[6]
port 18 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[7]
port 19 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chanx_left_in[8]
port 20 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[9]
port 21 nsew default input
rlabel metal3 s 0 16056 480 16176 6 chanx_left_out[0]
port 22 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 chanx_left_out[10]
port 23 nsew default tristate
rlabel metal3 s 0 22720 480 22840 6 chanx_left_out[11]
port 24 nsew default tristate
rlabel metal3 s 0 23400 480 23520 6 chanx_left_out[12]
port 25 nsew default tristate
rlabel metal3 s 0 23944 480 24064 6 chanx_left_out[13]
port 26 nsew default tristate
rlabel metal3 s 0 24624 480 24744 6 chanx_left_out[14]
port 27 nsew default tristate
rlabel metal3 s 0 25168 480 25288 6 chanx_left_out[15]
port 28 nsew default tristate
rlabel metal3 s 0 25848 480 25968 6 chanx_left_out[16]
port 29 nsew default tristate
rlabel metal3 s 0 26392 480 26512 6 chanx_left_out[17]
port 30 nsew default tristate
rlabel metal3 s 0 27072 480 27192 6 chanx_left_out[18]
port 31 nsew default tristate
rlabel metal3 s 0 27616 480 27736 6 chanx_left_out[19]
port 32 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 chanx_left_out[1]
port 33 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[2]
port 34 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[3]
port 35 nsew default tristate
rlabel metal3 s 0 18504 480 18624 6 chanx_left_out[4]
port 36 nsew default tristate
rlabel metal3 s 0 19048 480 19168 6 chanx_left_out[5]
port 37 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_left_out[6]
port 38 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 chanx_left_out[7]
port 39 nsew default tristate
rlabel metal3 s 0 20952 480 21072 6 chanx_left_out[8]
port 40 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[9]
port 41 nsew default tristate
rlabel metal2 s 4802 27520 4858 28000 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 10506 27520 10562 28000 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 11058 27520 11114 28000 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 11702 27520 11758 28000 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 12254 27520 12310 28000 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 12806 27520 12862 28000 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 13358 27520 13414 28000 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 14554 27520 14610 28000 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 15106 27520 15162 28000 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 15658 27520 15714 28000 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 5354 27520 5410 28000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 5998 27520 6054 28000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 6550 27520 6606 28000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 7102 27520 7158 28000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 7654 27520 7710 28000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 8206 27520 8262 28000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 8850 27520 8906 28000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 9402 27520 9458 28000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 9954 27520 10010 28000 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 16210 27520 16266 28000 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 21914 27520 21970 28000 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 22466 27520 22522 28000 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 23110 27520 23166 28000 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 23662 27520 23718 28000 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 24214 27520 24270 28000 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 24766 27520 24822 28000 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 25318 27520 25374 28000 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 25962 27520 26018 28000 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 26514 27520 26570 28000 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 27066 27520 27122 28000 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 16762 27520 16818 28000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 17406 27520 17462 28000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 17958 27520 18014 28000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 18510 27520 18566 28000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 19062 27520 19118 28000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 19614 27520 19670 28000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 20258 27520 20314 28000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 20810 27520 20866 28000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 21362 27520 21418 28000 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 left_bottom_grid_pin_11_
port 82 nsew default input
rlabel metal3 s 0 280 480 400 6 left_bottom_grid_pin_1_
port 83 nsew default input
rlabel metal3 s 0 824 480 944 6 left_bottom_grid_pin_3_
port 84 nsew default input
rlabel metal3 s 0 1368 480 1488 6 left_bottom_grid_pin_5_
port 85 nsew default input
rlabel metal3 s 0 2048 480 2168 6 left_bottom_grid_pin_7_
port 86 nsew default input
rlabel metal3 s 0 2592 480 2712 6 left_bottom_grid_pin_9_
port 87 nsew default input
rlabel metal2 s 7010 0 7066 480 6 prog_clk
port 88 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_42_
port 89 nsew default input
rlabel metal2 s 846 27520 902 28000 6 top_left_grid_pin_43_
port 90 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 top_left_grid_pin_44_
port 91 nsew default input
rlabel metal2 s 1950 27520 2006 28000 6 top_left_grid_pin_45_
port 92 nsew default input
rlabel metal2 s 2502 27520 2558 28000 6 top_left_grid_pin_46_
port 93 nsew default input
rlabel metal2 s 3146 27520 3202 28000 6 top_left_grid_pin_47_
port 94 nsew default input
rlabel metal2 s 3698 27520 3754 28000 6 top_left_grid_pin_48_
port 95 nsew default input
rlabel metal2 s 4250 27520 4306 28000 6 top_left_grid_pin_49_
port 96 nsew default input
rlabel metal2 s 27618 27520 27674 28000 6 top_right_grid_pin_1_
port 97 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 98 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 99 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
