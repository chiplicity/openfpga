* NGSPICE file created from cbx_1__3_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

.subckt cbx_1__3_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_grid_pin_0_ bottom_grid_pin_4_ bottom_grid_pin_8_ chanx_left_in[0]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_out[0] chanx_left_out[1]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_right_in[0] chanx_right_in[1] chanx_right_in[2]
+ chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7]
+ chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ data_in enable top_grid_pin_0_ top_grid_pin_10_ top_grid_pin_12_ top_grid_pin_14_
+ top_grid_pin_2_ top_grid_pin_4_ top_grid_pin_6_ top_grid_pin_8_ vpwr vgnd
XFILLER_26_96 vgnd vpwr scs8hd_decap_6
XFILLER_3_56 vgnd vpwr scs8hd_decap_3
XANTENNA__113__B _114_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_67 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_1_.latch data_in mem_bottom_ipin_2.LATCH_1_.latch/Q _129_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_192 vpwr vgnd scs8hd_fill_2
XFILLER_27_214 vgnd vpwr scs8hd_fill_1
XFILLER_12_10 vpwr vgnd scs8hd_fill_2
XFILLER_12_32 vgnd vpwr scs8hd_decap_3
XFILLER_33_217 vgnd vpwr scs8hd_decap_12
XANTENNA__108__B _099_/D vgnd vpwr scs8hd_diode_2
XFILLER_5_173 vgnd vpwr scs8hd_decap_4
XANTENNA__124__A _124_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_195 vgnd vpwr scs8hd_decap_6
Xmem_bottom_ipin_4.LATCH_4_.latch data_in mem_bottom_ipin_4.LATCH_4_.latch/Q _070_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_062_ _056_/B _114_/A _062_/Y vgnd vpwr scs8hd_nor2_4
X_131_ _131_/HI _131_/LO vgnd vpwr scs8hd_conb_1
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_198 vgnd vpwr scs8hd_decap_12
XFILLER_2_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__110__C address[3] vgnd vpwr scs8hd_diode_2
XANTENNA__119__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_22 vpwr vgnd scs8hd_fill_2
XFILLER_9_33 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_231 vpwr vgnd scs8hd_fill_2
X_114_ _114_/A _114_/B _114_/Y vgnd vpwr scs8hd_nor2_4
X_045_ _045_/A _045_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__121__B _121_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_2_.latch/Q mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_7 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_5.LATCH_0_.latch_SLEEPB _082_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_4_227 vgnd vpwr scs8hd_decap_6
XFILLER_4_205 vgnd vpwr scs8hd_decap_8
XFILLER_20_32 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_0_.latch/Q mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_74 vgnd vpwr scs8hd_fill_1
XANTENNA__116__B _114_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_45 vpwr vgnd scs8hd_fill_2
XFILLER_6_89 vgnd vpwr scs8hd_decap_3
XFILLER_13_3 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _131_/HI mem_bottom_ipin_0.LATCH_5_.latch/Q
+ mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_1_208 vgnd vpwr scs8hd_decap_12
XANTENNA__042__A address[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_25_197 vpwr vgnd scs8hd_fill_2
XFILLER_15_98 vgnd vpwr scs8hd_decap_6
XFILLER_0_230 vgnd vpwr scs8hd_decap_3
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XANTENNA__127__A _127_/A vgnd vpwr scs8hd_diode_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_197 vgnd vpwr scs8hd_fill_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_10_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_145 vgnd vpwr scs8hd_decap_8
XFILLER_22_167 vgnd vpwr scs8hd_decap_12
XFILLER_26_64 vpwr vgnd scs8hd_fill_2
XFILLER_26_20 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_bottom_ipin_5.LATCH_0_.latch data_in mem_bottom_ipin_5.LATCH_0_.latch/Q _082_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_35 vpwr vgnd scs8hd_fill_2
XFILLER_3_24 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_171 vgnd vpwr scs8hd_decap_12
XFILLER_10_104 vpwr vgnd scs8hd_fill_2
XFILLER_12_77 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_7.LATCH_3_.latch data_in mem_bottom_ipin_7.LATCH_3_.latch/Q _094_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_3.LATCH_1_.latch_SLEEPB _064_/Y vgnd vpwr scs8hd_diode_2
XFILLER_33_229 vgnd vpwr scs8hd_decap_4
XANTENNA__108__C _059_/C vgnd vpwr scs8hd_diode_2
XFILLER_5_163 vgnd vpwr scs8hd_fill_1
XFILLER_5_152 vgnd vpwr scs8hd_decap_4
XANTENNA__124__B _124_/B vgnd vpwr scs8hd_diode_2
XFILLER_24_218 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_0_ vgnd vpwr scs8hd_inv_1
XANTENNA__050__A address[6] vgnd vpwr scs8hd_diode_2
X_130_ _074_/A _127_/B _130_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_87 vpwr vgnd scs8hd_fill_2
X_061_ _059_/A address[2] address[0] _114_/A vgnd vpwr scs8hd_or3_4
XFILLER_2_111 vgnd vpwr scs8hd_decap_4
XFILLER_2_166 vgnd vpwr scs8hd_decap_12
XANTENNA__110__D _124_/A vgnd vpwr scs8hd_diode_2
XANTENNA__119__B _121_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XFILLER_9_89 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_232 vgnd vpwr scs8hd_fill_1
XANTENNA__045__A _045_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_10 vpwr vgnd scs8hd_fill_2
XFILLER_11_210 vpwr vgnd scs8hd_fill_2
X_113_ _127_/A _114_/B _113_/Y vgnd vpwr scs8hd_nor2_4
X_044_ _044_/A _044_/Y vgnd vpwr scs8hd_inv_8
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XFILLER_29_107 vgnd vpwr scs8hd_decap_4
XFILLER_1_90 vpwr vgnd scs8hd_fill_2
XFILLER_20_44 vgnd vpwr scs8hd_decap_8
XFILLER_20_55 vpwr vgnd scs8hd_fill_2
XFILLER_29_86 vpwr vgnd scs8hd_fill_2
XFILLER_29_20 vpwr vgnd scs8hd_fill_2
XFILLER_28_173 vgnd vpwr scs8hd_fill_1
XFILLER_28_151 vpwr vgnd scs8hd_fill_2
XFILLER_6_24 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_ipin_1.LATCH_2_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_154 vpwr vgnd scs8hd_fill_2
XFILLER_15_55 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_31_87 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_121 vpwr vgnd scs8hd_fill_2
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_135 vgnd vpwr scs8hd_decap_12
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__B _127_/B vgnd vpwr scs8hd_diode_2
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_176 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__143__A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_22_179 vgnd vpwr scs8hd_decap_3
XANTENNA__053__A address[1] vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_0.LATCH_4_.latch data_in mem_top_ipin_0.LATCH_4_.latch/Q _101_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_43 vgnd vpwr scs8hd_decap_6
XFILLER_9_106 vpwr vgnd scs8hd_fill_2
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_14 vpwr vgnd scs8hd_fill_2
XANTENNA__048__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_12_23 vgnd vpwr scs8hd_decap_8
XFILLER_12_89 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_2_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _043_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_5.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_230 vgnd vpwr scs8hd_decap_3
XFILLER_23_66 vgnd vpwr scs8hd_fill_1
XFILLER_3_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_6.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_060_ _056_/B _127_/A _060_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_178 vgnd vpwr scs8hd_decap_6
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_230 vgnd vpwr scs8hd_decap_3
XFILLER_9_57 vgnd vpwr scs8hd_fill_1
XFILLER_9_79 vgnd vpwr scs8hd_decap_4
XANTENNA__151__A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__061__A _059_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_4_.latch data_in mem_bottom_ipin_0.LATCH_4_.latch/Q _112_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
X_043_ _043_/A _043_/Y vgnd vpwr scs8hd_inv_8
X_112_ _126_/A _114_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__146__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__056__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_185 vpwr vgnd scs8hd_fill_2
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_1.LATCH_0_.latch data_in _044_/A _107_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_130 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_15_45 vpwr vgnd scs8hd_fill_2
XFILLER_15_78 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_16_100 vgnd vpwr scs8hd_fill_1
XFILLER_16_133 vgnd vpwr scs8hd_decap_3
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_147 vgnd vpwr scs8hd_decap_12
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__053__B _053_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_9_129 vpwr vgnd scs8hd_fill_2
XFILLER_13_114 vgnd vpwr scs8hd_fill_1
XFILLER_13_158 vpwr vgnd scs8hd_fill_2
XFILLER_21_191 vpwr vgnd scs8hd_fill_2
XFILLER_3_48 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__154__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_8_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_2_.latch_SLEEPB _088_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_217 vgnd vpwr scs8hd_decap_12
XFILLER_10_139 vgnd vpwr scs8hd_decap_3
XFILLER_12_46 vgnd vpwr scs8hd_decap_12
XANTENNA__064__A _056_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_206 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_1.LATCH_0_.latch data_in mem_bottom_ipin_1.LATCH_0_.latch/Q _123_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__149__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__059__A _059_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_209 vgnd vpwr scs8hd_decap_8
XFILLER_23_78 vpwr vgnd scs8hd_fill_2
XFILLER_23_23 vpwr vgnd scs8hd_fill_2
XFILLER_2_135 vgnd vpwr scs8hd_decap_12
XFILLER_2_124 vpwr vgnd scs8hd_fill_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_3.LATCH_3_.latch data_in mem_bottom_ipin_3.LATCH_3_.latch/Q _060_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_3 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _045_/A mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__061__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_18_23 vgnd vpwr scs8hd_decap_6
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XFILLER_11_223 vpwr vgnd scs8hd_fill_2
X_042_ address[0] _059_/C vgnd vpwr scs8hd_inv_8
Xmux_top_ipin_1.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_111_ _125_/A _114_/B _111_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_bottom_ipin_4.LATCH_3_.latch_SLEEPB _071_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__056__B _056_/B vgnd vpwr scs8hd_diode_2
XANTENNA__072__A _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_33 vpwr vgnd scs8hd_fill_2
XFILLER_29_66 vpwr vgnd scs8hd_fill_2
XFILLER_28_120 vgnd vpwr scs8hd_decap_3
XFILLER_3_230 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XANTENNA__157__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_19_175 vpwr vgnd scs8hd_fill_2
XFILLER_19_197 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_2_.latch/Q mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_25_178 vgnd vpwr scs8hd_decap_3
XFILLER_25_134 vpwr vgnd scs8hd_fill_2
XANTENNA__067__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_0_211 vgnd vpwr scs8hd_decap_6
XFILLER_31_104 vgnd vpwr scs8hd_decap_12
XFILLER_16_145 vgnd vpwr scs8hd_decap_4
XFILLER_16_189 vgnd vpwr scs8hd_decap_8
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_159 vgnd vpwr scs8hd_decap_12
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__053__C _059_/C vgnd vpwr scs8hd_diode_2
XFILLER_3_27 vpwr vgnd scs8hd_fill_2
XFILLER_8_152 vgnd vpwr scs8hd_fill_1
XFILLER_8_196 vgnd vpwr scs8hd_decap_4
XFILLER_12_181 vgnd vpwr scs8hd_decap_4
XFILLER_27_229 vgnd vpwr scs8hd_decap_4
XANTENNA__064__B _073_/A vgnd vpwr scs8hd_diode_2
XANTENNA__080__A _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_58 vgnd vpwr scs8hd_decap_3
XFILLER_18_218 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB _126_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_111 vpwr vgnd scs8hd_fill_2
XFILLER_5_100 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_6.LATCH_2_.latch data_in mem_bottom_ipin_6.LATCH_2_.latch/Q _088_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__059__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__075__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XFILLER_2_147 vgnd vpwr scs8hd_decap_3
XFILLER_9_37 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_224 vgnd vpwr scs8hd_decap_8
XANTENNA__061__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_18_46 vgnd vpwr scs8hd_decap_4
XFILLER_18_57 vpwr vgnd scs8hd_fill_2
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
X_110_ _091_/A address[4] address[3] _124_/A _114_/B vgnd vpwr scs8hd_or4_4
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _131_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__072__B _073_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB _106_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_14 vpwr vgnd scs8hd_fill_2
XFILLER_29_12 vgnd vpwr scs8hd_decap_8
XFILLER_28_165 vgnd vpwr scs8hd_decap_8
XFILLER_28_143 vgnd vpwr scs8hd_decap_8
XFILLER_28_132 vgnd vpwr scs8hd_decap_8
XFILLER_6_16 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_6_49 vpwr vgnd scs8hd_fill_2
XFILLER_10_80 vgnd vpwr scs8hd_decap_8
XFILLER_19_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_146 vpwr vgnd scs8hd_fill_2
XFILLER_25_168 vgnd vpwr scs8hd_decap_4
XANTENNA__083__A _091_/A vgnd vpwr scs8hd_diode_2
XANTENNA__067__B _098_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_116 vgnd vpwr scs8hd_decap_6
Xmux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_157 vgnd vpwr scs8hd_decap_8
XFILLER_16_168 vgnd vpwr scs8hd_decap_8
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_68 vgnd vpwr scs8hd_decap_4
XFILLER_13_138 vgnd vpwr scs8hd_decap_4
XANTENNA__078__A _126_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _043_/A mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_160 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_230 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_119 vpwr vgnd scs8hd_fill_2
XANTENNA__080__B _082_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_156 vgnd vpwr scs8hd_fill_1
XFILLER_5_123 vgnd vpwr scs8hd_fill_1
XANTENNA__059__C _059_/C vgnd vpwr scs8hd_diode_2
XFILLER_23_222 vgnd vpwr scs8hd_decap_8
XFILLER_23_211 vgnd vpwr scs8hd_decap_4
XANTENNA__075__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_23_36 vgnd vpwr scs8hd_decap_3
XANTENNA__091__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_16 vgnd vpwr scs8hd_decap_4
XFILLER_13_80 vgnd vpwr scs8hd_fill_1
XFILLER_13_91 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_2_.latch/Q mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XANTENNA__086__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_7.LATCH_4_.latch_SLEEPB _093_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_94 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_26 vpwr vgnd scs8hd_fill_2
XFILLER_20_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_0_.latch/Q mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_90 vgnd vpwr scs8hd_decap_3
XFILLER_25_158 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_25_114 vpwr vgnd scs8hd_fill_2
XFILLER_15_15 vpwr vgnd scs8hd_fill_2
XFILLER_15_26 vpwr vgnd scs8hd_fill_2
XFILLER_33_180 vgnd vpwr scs8hd_decap_3
XANTENNA__083__B _091_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_59 vpwr vgnd scs8hd_fill_2
XFILLER_16_103 vgnd vpwr scs8hd_decap_6
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_125 vgnd vpwr scs8hd_decap_8
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_30_194 vgnd vpwr scs8hd_decap_4
XFILLER_30_161 vpwr vgnd scs8hd_fill_2
XFILLER_15_191 vpwr vgnd scs8hd_fill_2
XFILLER_22_128 vgnd vpwr scs8hd_decap_8
XANTENNA__078__B _082_/B vgnd vpwr scs8hd_diode_2
XANTENNA__094__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_106 vpwr vgnd scs8hd_fill_2
XFILLER_13_117 vpwr vgnd scs8hd_fill_2
XFILLER_21_161 vpwr vgnd scs8hd_fill_2
XFILLER_21_172 vgnd vpwr scs8hd_decap_4
XFILLER_3_18 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_154 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_7.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_12_194 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_5.LATCH_5_.latch_SLEEPB _077_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_231 vpwr vgnd scs8hd_fill_2
XANTENNA__089__A _073_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_179 vpwr vgnd scs8hd_fill_2
XFILLER_5_135 vpwr vgnd scs8hd_fill_2
XFILLER_17_231 vpwr vgnd scs8hd_fill_2
XFILLER_4_61 vgnd vpwr scs8hd_decap_4
XANTENNA__075__C _091_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__091__B _091_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__086__B _086_/B vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_2_.latch data_in mem_bottom_ipin_2.LATCH_2_.latch/Q _128_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_27_3 vgnd vpwr scs8hd_decap_4
X_099_ _091_/A address[4] address[3] _099_/D _100_/B vgnd vpwr scs8hd_or4_4
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _132_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_62 vgnd vpwr scs8hd_decap_3
XFILLER_1_84 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_29_58 vgnd vpwr scs8hd_decap_3
XFILLER_28_112 vgnd vpwr scs8hd_decap_8
Xmem_bottom_ipin_4.LATCH_5_.latch data_in mem_bottom_ipin_4.LATCH_5_.latch/Q _069_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_189 vgnd vpwr scs8hd_decap_4
XANTENNA__097__A _074_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_top_ipin_0.LATCH_3_.latch/Q mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_3_222 vgnd vpwr scs8hd_decap_8
XFILLER_19_134 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_126 vpwr vgnd scs8hd_fill_2
XFILLER_15_49 vgnd vpwr scs8hd_decap_4
XFILLER_31_59 vpwr vgnd scs8hd_fill_2
XFILLER_31_15 vgnd vpwr scs8hd_decap_12
XANTENNA__083__C address[3] vgnd vpwr scs8hd_diode_2
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_22_118 vgnd vpwr scs8hd_fill_1
XFILLER_30_151 vpwr vgnd scs8hd_fill_2
XFILLER_7_50 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_83 vpwr vgnd scs8hd_fill_2
XANTENNA__094__B _095_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_70 vpwr vgnd scs8hd_fill_2
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XFILLER_8_144 vgnd vpwr scs8hd_decap_8
XFILLER_16_81 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__089__B _086_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_202 vgnd vpwr scs8hd_decap_12
XFILLER_4_180 vgnd vpwr scs8hd_decap_4
XFILLER_4_40 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_0_.latch/Q mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_128 vgnd vpwr scs8hd_decap_4
XANTENNA__091__C _091_/C vgnd vpwr scs8hd_diode_2
XFILLER_14_202 vpwr vgnd scs8hd_fill_2
XFILLER_29_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_5.LATCH_1_.latch data_in mem_bottom_ipin_5.LATCH_1_.latch/Q _081_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_1_.latch/Q mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_227 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_4.LATCH_0_.latch_SLEEPB _074_/Y vgnd vpwr scs8hd_diode_2
X_098_ address[5] _098_/B _099_/D vgnd vpwr scs8hd_or2_4
Xmem_bottom_ipin_7.LATCH_4_.latch data_in mem_bottom_ipin_7.LATCH_4_.latch/Q _093_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_29_37 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_2_ vgnd vpwr scs8hd_inv_1
XANTENNA__097__B _095_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_201 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_113 vgnd vpwr scs8hd_decap_4
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XFILLER_19_179 vpwr vgnd scs8hd_fill_2
XFILLER_33_160 vgnd vpwr scs8hd_decap_12
XFILLER_25_138 vgnd vpwr scs8hd_decap_8
XFILLER_31_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_93 vpwr vgnd scs8hd_fill_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_182 vgnd vpwr scs8hd_fill_1
XFILLER_7_62 vpwr vgnd scs8hd_fill_2
XFILLER_26_16 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_112 vpwr vgnd scs8hd_fill_2
XFILLER_35_211 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ _046_/A mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_26_200 vpwr vgnd scs8hd_fill_2
XFILLER_5_115 vgnd vpwr scs8hd_decap_4
XFILLER_5_104 vpwr vgnd scs8hd_fill_2
XFILLER_5_159 vpwr vgnd scs8hd_fill_2
XFILLER_17_200 vpwr vgnd scs8hd_fill_2
XFILLER_17_211 vpwr vgnd scs8hd_fill_2
XFILLER_4_74 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_107 vpwr vgnd scs8hd_fill_2
XANTENNA__091__D _084_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_83 vgnd vpwr scs8hd_fill_1
Xmem_top_ipin_0.LATCH_5_.latch data_in mem_top_ipin_0.LATCH_5_.latch/Q _100_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XFILLER_20_206 vgnd vpwr scs8hd_decap_6
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XFILLER_11_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_93 vgnd vpwr scs8hd_decap_3
XFILLER_24_71 vpwr vgnd scs8hd_fill_2
X_097_ _074_/A _095_/B _097_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_31 vgnd vpwr scs8hd_fill_1
XFILLER_1_53 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _133_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_18 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_213 vpwr vgnd scs8hd_fill_2
XFILLER_10_73 vgnd vpwr scs8hd_decap_4
XFILLER_19_60 vgnd vpwr scs8hd_fill_1
XFILLER_19_71 vpwr vgnd scs8hd_fill_2
XFILLER_34_117 vgnd vpwr scs8hd_decap_12
XFILLER_27_180 vgnd vpwr scs8hd_fill_1
XFILLER_19_158 vpwr vgnd scs8hd_fill_2
X_149_ chanx_right_in[1] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_172 vgnd vpwr scs8hd_decap_8
XFILLER_31_39 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_150 vgnd vpwr scs8hd_decap_3
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_194 vgnd vpwr scs8hd_decap_6
Xmem_bottom_ipin_0.LATCH_5_.latch data_in mem_bottom_ipin_0.LATCH_5_.latch/Q _111_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_83 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_0_.latch/Q mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_15_172 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_96 vpwr vgnd scs8hd_fill_2
XFILLER_26_28 vgnd vpwr scs8hd_decap_3
XFILLER_21_142 vgnd vpwr scs8hd_decap_4
XFILLER_29_220 vpwr vgnd scs8hd_fill_2
XFILLER_12_164 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_212 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_1.LATCH_1_.latch data_in _043_/A _106_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_93 vpwr vgnd scs8hd_fill_2
XFILLER_27_82 vpwr vgnd scs8hd_fill_2
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_171 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_ipin_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_4.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_62 vpwr vgnd scs8hd_fill_2
XFILLER_1_196 vgnd vpwr scs8hd_decap_12
XANTENNA__100__A _125_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_7.LATCH_1_.latch_SLEEPB _096_/Y vgnd vpwr scs8hd_diode_2
X_096_ _073_/A _095_/B _096_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_98 vgnd vpwr scs8hd_decap_3
Xmem_bottom_ipin_1.LATCH_1_.latch data_in mem_bottom_ipin_1.LATCH_1_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ _044_/A mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_19_126 vpwr vgnd scs8hd_fill_2
XFILLER_34_129 vgnd vpwr scs8hd_decap_12
X_148_ chanx_right_in[2] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
X_079_ _127_/A _082_/B _079_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_118 vpwr vgnd scs8hd_fill_2
XFILLER_15_19 vpwr vgnd scs8hd_fill_2
XFILLER_18_192 vgnd vpwr scs8hd_decap_3
Xmem_bottom_ipin_3.LATCH_4_.latch data_in mem_bottom_ipin_3.LATCH_4_.latch/Q _058_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
XFILLER_33_151 vgnd vpwr scs8hd_fill_1
XFILLER_24_184 vgnd vpwr scs8hd_fill_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_73 vpwr vgnd scs8hd_fill_2
XFILLER_30_165 vgnd vpwr scs8hd_decap_3
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_195 vgnd vpwr scs8hd_decap_3
XFILLER_30_198 vgnd vpwr scs8hd_fill_1
XFILLER_7_42 vgnd vpwr scs8hd_decap_6
XFILLER_21_132 vgnd vpwr scs8hd_decap_4
XFILLER_21_176 vgnd vpwr scs8hd_fill_1
XFILLER_21_187 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_5.LATCH_2_.latch_SLEEPB _080_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_232 vgnd vpwr scs8hd_fill_1
XFILLER_8_136 vpwr vgnd scs8hd_fill_2
XFILLER_12_132 vgnd vpwr scs8hd_decap_4
XFILLER_12_143 vpwr vgnd scs8hd_fill_2
XFILLER_12_154 vgnd vpwr scs8hd_decap_3
XFILLER_16_84 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_198 vpwr vgnd scs8hd_fill_2
XANTENNA__103__A _114_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_139 vpwr vgnd scs8hd_fill_2
XFILLER_32_227 vgnd vpwr scs8hd_decap_6
XFILLER_4_32 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _141_/HI _045_/Y mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_19 vpwr vgnd scs8hd_fill_2
XFILLER_13_30 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__100__B _100_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_220 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_0_.latch/Q mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_ipin_4.LATCH_0_.latch data_in mem_bottom_ipin_4.LATCH_0_.latch/Q _074_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_24_84 vpwr vgnd scs8hd_fill_2
XFILLER_6_201 vgnd vpwr scs8hd_decap_12
X_095_ _114_/A _095_/B _095_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_bottom_ipin_3.LATCH_3_.latch_SLEEPB _060_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_7 vgnd vpwr scs8hd_fill_1
XANTENNA__111__A _125_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _134_/HI vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_ipin_6.LATCH_3_.latch data_in mem_bottom_ipin_6.LATCH_3_.latch/Q _087_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_171 vgnd vpwr scs8hd_decap_3
XFILLER_19_95 vgnd vpwr scs8hd_decap_3
XFILLER_19_138 vgnd vpwr scs8hd_decap_3
XFILLER_35_94 vgnd vpwr scs8hd_decap_12
XFILLER_27_193 vpwr vgnd scs8hd_fill_2
XANTENNA__106__A _076_/B vgnd vpwr scs8hd_diode_2
X_147_ chanx_right_in[3] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
X_078_ _126_/A _082_/B _078_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_18_171 vgnd vpwr scs8hd_decap_8
XFILLER_33_196 vgnd vpwr scs8hd_fill_1
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_41 vpwr vgnd scs8hd_fill_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_30_177 vgnd vpwr scs8hd_decap_12
XFILLER_7_21 vpwr vgnd scs8hd_fill_2
XFILLER_7_10 vpwr vgnd scs8hd_fill_2
XFILLER_7_54 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_104 vpwr vgnd scs8hd_fill_2
XFILLER_8_159 vgnd vpwr scs8hd_decap_3
XFILLER_12_177 vpwr vgnd scs8hd_fill_2
XFILLER_16_96 vgnd vpwr scs8hd_decap_4
XANTENNA__103__B _100_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_1.LATCH_4_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__114__A _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_217 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_14_206 vgnd vpwr scs8hd_decap_8
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_0_.latch/Q mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_110 vpwr vgnd scs8hd_fill_2
XFILLER_1_132 vpwr vgnd scs8hd_fill_2
XFILLER_1_143 vgnd vpwr scs8hd_decap_12
XANTENNA__109__A _124_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_232 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_24_30 vgnd vpwr scs8hd_fill_1
XFILLER_6_213 vgnd vpwr scs8hd_fill_1
X_094_ _127_/A _095_/B _094_/Y vgnd vpwr scs8hd_nor2_4
Xmux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_8_ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB _104_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__111__B _114_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_34 vgnd vpwr scs8hd_decap_3
XFILLER_1_67 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_43 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_7.LATCH_3_.latch/Q mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_150 vgnd vpwr scs8hd_decap_4
XFILLER_19_41 vpwr vgnd scs8hd_fill_2
XFILLER_19_52 vpwr vgnd scs8hd_fill_2
XANTENNA__106__B _099_/D vgnd vpwr scs8hd_diode_2
XANTENNA__122__A _073_/A vgnd vpwr scs8hd_diode_2
X_077_ _125_/A _082_/B _077_/Y vgnd vpwr scs8hd_nor2_4
X_146_ chanx_right_in[4] chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_33_120 vpwr vgnd scs8hd_fill_2
XFILLER_24_120 vgnd vpwr scs8hd_decap_3
XFILLER_16_109 vgnd vpwr scs8hd_fill_1
XFILLER_24_142 vgnd vpwr scs8hd_decap_8
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XFILLER_21_97 vpwr vgnd scs8hd_fill_2
XPHY_6 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _140_/HI _043_/Y mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_142 vpwr vgnd scs8hd_fill_2
XFILLER_30_189 vgnd vpwr scs8hd_decap_3
XFILLER_30_123 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _124_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_66 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_129_ _073_/A _127_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_21_112 vgnd vpwr scs8hd_decap_4
XFILLER_32_96 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_193 vgnd vpwr scs8hd_decap_6
Xmux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_0_.latch/Q mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_204 vgnd vpwr scs8hd_decap_8
XFILLER_5_119 vgnd vpwr scs8hd_fill_1
XFILLER_27_52 vgnd vpwr scs8hd_fill_1
XFILLER_17_204 vpwr vgnd scs8hd_fill_2
XFILLER_17_215 vpwr vgnd scs8hd_fill_2
XFILLER_4_141 vpwr vgnd scs8hd_fill_2
XFILLER_4_130 vgnd vpwr scs8hd_fill_1
XANTENNA__114__B _114_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_78 vgnd vpwr scs8hd_decap_12
XFILLER_4_23 vgnd vpwr scs8hd_decap_8
XFILLER_4_12 vpwr vgnd scs8hd_fill_2
XANTENNA__130__A _074_/A vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_0.LATCH_0_.latch data_in mem_top_ipin_0.LATCH_0_.latch/Q _105_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_218 vgnd vpwr scs8hd_decap_12
XFILLER_13_76 vgnd vpwr scs8hd_decap_4
XFILLER_13_87 vpwr vgnd scs8hd_fill_2
XFILLER_1_155 vgnd vpwr scs8hd_decap_12
XFILLER_8_3 vgnd vpwr scs8hd_decap_3
XANTENNA__109__B _099_/D vgnd vpwr scs8hd_diode_2
XANTENNA__125__A _125_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_4_.latch_SLEEPB _086_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_1_.latch/Q mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_42 vpwr vgnd scs8hd_fill_2
XFILLER_10_232 vgnd vpwr scs8hd_fill_1
X_093_ _126_/A _095_/B _093_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _135_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_55 vgnd vpwr scs8hd_fill_1
XFILLER_10_88 vpwr vgnd scs8hd_fill_2
XFILLER_19_20 vgnd vpwr scs8hd_fill_1
XFILLER_35_63 vgnd vpwr scs8hd_decap_12
XFILLER_19_75 vgnd vpwr scs8hd_decap_4
XANTENNA__106__C _059_/C vgnd vpwr scs8hd_diode_2
X_145_ chanx_right_in[5] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA__122__B _121_/B vgnd vpwr scs8hd_diode_2
X_076_ _084_/A _076_/B _082_/B vgnd vpwr scs8hd_or2_4
Xmem_bottom_ipin_0.LATCH_0_.latch data_in mem_bottom_ipin_0.LATCH_0_.latch/Q _116_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_176 vgnd vpwr scs8hd_decap_8
XFILLER_24_165 vpwr vgnd scs8hd_fill_2
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_21 vgnd vpwr scs8hd_decap_4
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_132 vgnd vpwr scs8hd_decap_4
XFILLER_15_176 vgnd vpwr scs8hd_decap_4
XFILLER_15_187 vpwr vgnd scs8hd_fill_2
XFILLER_30_157 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_2.LATCH_3_.latch data_in mem_bottom_ipin_2.LATCH_3_.latch/Q _127_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_128_ _114_/A _127_/B _128_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__117__B _076_/B vgnd vpwr scs8hd_diode_2
X_059_ _059_/A address[2] _059_/C _127_/A vgnd vpwr scs8hd_or3_4
XFILLER_23_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_157 vpwr vgnd scs8hd_fill_2
XFILLER_21_168 vpwr vgnd scs8hd_fill_2
XFILLER_21_179 vpwr vgnd scs8hd_fill_2
XANTENNA__043__A _043_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_224 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_4.LATCH_5_.latch_SLEEPB _069_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_102 vpwr vgnd scs8hd_fill_2
XFILLER_16_10 vpwr vgnd scs8hd_fill_2
XFILLER_16_32 vpwr vgnd scs8hd_fill_2
XFILLER_8_117 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_5.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__128__A _114_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_150 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_86 vgnd vpwr scs8hd_decap_4
XFILLER_27_31 vpwr vgnd scs8hd_fill_2
XFILLER_27_97 vpwr vgnd scs8hd_fill_2
XFILLER_4_186 vgnd vpwr scs8hd_decap_4
XFILLER_4_57 vpwr vgnd scs8hd_fill_2
XFILLER_4_46 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__130__B _127_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_230 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_6.LATCH_3_.latch/Q mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_22 vpwr vgnd scs8hd_fill_2
XFILLER_13_44 vpwr vgnd scs8hd_fill_2
XFILLER_13_66 vgnd vpwr scs8hd_fill_1
XFILLER_1_167 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__125__B _127_/B vgnd vpwr scs8hd_diode_2
XANTENNA__109__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__051__A address[4] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_ipin_0.LATCH_4_.latch/Q mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_24_32 vgnd vpwr scs8hd_decap_6
XFILLER_24_10 vpwr vgnd scs8hd_fill_2
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
X_092_ _125_/A _095_/B _092_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _046_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__046__A _046_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_218 vpwr vgnd scs8hd_fill_2
XFILLER_10_12 vpwr vgnd scs8hd_fill_2
XFILLER_10_23 vpwr vgnd scs8hd_fill_2
XFILLER_19_119 vgnd vpwr scs8hd_decap_3
XFILLER_35_75 vgnd vpwr scs8hd_decap_12
X_144_ chanx_right_in[6] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
X_075_ _091_/A address[4] _091_/C _076_/B vgnd vpwr scs8hd_or3_4
XFILLER_25_7 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_0_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_6 vpwr vgnd scs8hd_fill_2
XFILLER_24_133 vgnd vpwr scs8hd_fill_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_ipin_5.LATCH_2_.latch data_in mem_bottom_ipin_5.LATCH_2_.latch/Q _080_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_77 vgnd vpwr scs8hd_decap_4
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_155 vpwr vgnd scs8hd_fill_2
X_127_ _127_/A _127_/B _127_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_79 vpwr vgnd scs8hd_fill_2
X_058_ _056_/B _126_/A _058_/Y vgnd vpwr scs8hd_nor2_4
Xmem_bottom_ipin_7.LATCH_5_.latch data_in mem_bottom_ipin_7.LATCH_5_.latch/Q _092_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_203 vgnd vpwr scs8hd_decap_6
XFILLER_12_114 vgnd vpwr scs8hd_decap_3
XFILLER_12_147 vgnd vpwr scs8hd_decap_6
XFILLER_16_66 vpwr vgnd scs8hd_fill_2
XFILLER_16_77 vgnd vpwr scs8hd_decap_4
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_191 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__144__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__128__B _127_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_180 vgnd vpwr scs8hd_fill_1
XFILLER_11_191 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_1_.latch/Q mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__054__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_27_65 vpwr vgnd scs8hd_fill_2
XFILLER_27_21 vpwr vgnd scs8hd_fill_2
XFILLER_27_10 vpwr vgnd scs8hd_fill_2
XFILLER_4_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__049__A enable vgnd vpwr scs8hd_diode_2
XFILLER_13_34 vgnd vpwr scs8hd_fill_1
XFILLER_13_56 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_2_.latch/Q mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_1_179 vgnd vpwr scs8hd_decap_4
XFILLER_9_213 vpwr vgnd scs8hd_fill_2
XFILLER_9_224 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_3.LATCH_0_.latch_SLEEPB _066_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_88 vgnd vpwr scs8hd_decap_4
XFILLER_6_227 vgnd vpwr scs8hd_decap_6
X_091_ _091_/A _091_/B _091_/C _084_/A _095_/B vgnd vpwr scs8hd_or4_4
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_48 vgnd vpwr scs8hd_decap_3
XANTENNA__152__A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _136_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__062__A _056_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_109 vpwr vgnd scs8hd_fill_2
XFILLER_35_87 vgnd vpwr scs8hd_decap_6
XFILLER_35_32 vgnd vpwr scs8hd_decap_12
XFILLER_27_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_143_ chanx_right_in[7] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
X_074_ _074_/A _073_/B _074_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
XFILLER_33_112 vgnd vpwr scs8hd_decap_8
XFILLER_18_142 vgnd vpwr scs8hd_fill_1
XFILLER_33_156 vpwr vgnd scs8hd_fill_2
XANTENNA__147__A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__057__A address[1] vgnd vpwr scs8hd_diode_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_45 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_30_104 vgnd vpwr scs8hd_decap_8
XFILLER_7_14 vgnd vpwr scs8hd_decap_4
X_126_ _126_/A _127_/B _126_/Y vgnd vpwr scs8hd_nor2_4
X_057_ address[1] _053_/B address[0] _126_/A vgnd vpwr scs8hd_or3_4
XFILLER_7_58 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_5.LATCH_3_.latch/Q mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_6 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ _046_/Y mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_23 vpwr vgnd scs8hd_fill_2
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_8_108 vpwr vgnd scs8hd_fill_2
XFILLER_35_218 vgnd vpwr scs8hd_decap_12
XFILLER_11_170 vpwr vgnd scs8hd_fill_2
X_109_ _124_/B _099_/D address[0] _109_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__054__B address[6] vgnd vpwr scs8hd_diode_2
XANTENNA__070__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_55 vgnd vpwr scs8hd_decap_6
XFILLER_27_44 vpwr vgnd scs8hd_fill_2
XFILLER_4_177 vgnd vpwr scs8hd_fill_1
XFILLER_4_133 vgnd vpwr scs8hd_fill_1
XANTENNA__155__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__065__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_22_232 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_114 vpwr vgnd scs8hd_fill_2
XFILLER_1_136 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_0_.latch/Q mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_210 vgnd vpwr scs8hd_decap_4
XFILLER_13_232 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_14_ vgnd vpwr scs8hd_inv_1
XFILLER_24_67 vpwr vgnd scs8hd_fill_2
XFILLER_10_213 vgnd vpwr scs8hd_fill_1
XFILLER_10_224 vgnd vpwr scs8hd_decap_8
X_090_ _074_/A _086_/B _090_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_3 vpwr vgnd scs8hd_fill_2
XFILLER_1_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_47 vgnd vpwr scs8hd_decap_8
XFILLER_10_69 vpwr vgnd scs8hd_fill_2
XANTENNA__062__B _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_12 vpwr vgnd scs8hd_fill_2
XFILLER_27_176 vgnd vpwr scs8hd_decap_4
XFILLER_27_132 vgnd vpwr scs8hd_decap_3
XFILLER_27_110 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_45 vpwr vgnd scs8hd_fill_2
XFILLER_19_56 vpwr vgnd scs8hd_fill_2
XFILLER_35_44 vgnd vpwr scs8hd_decap_12
X_142_ chanx_right_in[8] chanx_left_out[8] vgnd vpwr scs8hd_buf_2
X_073_ _073_/A _073_/B _073_/Y vgnd vpwr scs8hd_nor2_4
Xmux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_1_.latch/Q mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_33_135 vgnd vpwr scs8hd_decap_12
XFILLER_33_102 vpwr vgnd scs8hd_fill_2
XFILLER_18_121 vpwr vgnd scs8hd_fill_2
XFILLER_18_154 vgnd vpwr scs8hd_decap_6
XFILLER_2_81 vgnd vpwr scs8hd_decap_8
XFILLER_32_190 vgnd vpwr scs8hd_decap_12
XANTENNA__057__B _053_/B vgnd vpwr scs8hd_diode_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__073__A _073_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_13 vpwr vgnd scs8hd_fill_2
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_8_ vgnd vpwr scs8hd_inv_1
XFILLER_15_168 vpwr vgnd scs8hd_fill_2
XFILLER_30_127 vgnd vpwr scs8hd_decap_12
X_125_ _125_/A _127_/B _125_/Y vgnd vpwr scs8hd_nor2_4
X_056_ _125_/A _056_/B _056_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__158__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_21_138 vpwr vgnd scs8hd_fill_2
XANTENNA__068__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_1.LATCH_2_.latch data_in mem_bottom_ipin_1.LATCH_2_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_108_ _124_/B _099_/D _059_/C _108_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_7_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_3 vgnd vpwr scs8hd_fill_1
XFILLER_26_219 vgnd vpwr scs8hd_decap_12
XANTENNA__070__B _073_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_219 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_3.LATCH_5_.latch data_in mem_bottom_ipin_3.LATCH_5_.latch/Q _056_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_167 vpwr vgnd scs8hd_fill_2
XFILLER_4_145 vgnd vpwr scs8hd_decap_8
XFILLER_4_16 vgnd vpwr scs8hd_decap_4
XFILLER_31_222 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__065__B address[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_0_.latch/Q mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_14 vpwr vgnd scs8hd_fill_2
XANTENNA__081__A _073_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_1_.latch_SLEEPB _089_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_222 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_24_46 vgnd vpwr scs8hd_decap_4
XANTENNA__076__A _084_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_4.LATCH_3_.latch/Q mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ _044_/Y mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _137_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_24 vpwr vgnd scs8hd_fill_2
XFILLER_35_56 vgnd vpwr scs8hd_decap_6
X_141_ _141_/HI _141_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_210 vgnd vpwr scs8hd_decap_4
X_072_ _114_/A _073_/B _072_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_147 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _140_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_188 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_6.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_24_125 vpwr vgnd scs8hd_fill_2
XFILLER_2_93 vgnd vpwr scs8hd_decap_3
XFILLER_2_60 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_7.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_169 vgnd vpwr scs8hd_decap_4
XANTENNA__057__C address[0] vgnd vpwr scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__073__B _073_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_25 vgnd vpwr scs8hd_fill_1
XFILLER_15_114 vpwr vgnd scs8hd_fill_2
XFILLER_30_139 vgnd vpwr scs8hd_decap_12
XFILLER_7_38 vpwr vgnd scs8hd_fill_2
X_055_ _091_/A _091_/B _091_/C _124_/A _056_/B vgnd vpwr scs8hd_or4_4
X_124_ _124_/A _124_/B _127_/B vgnd vpwr scs8hd_or2_4
XANTENNA_mem_bottom_ipin_4.LATCH_2_.latch_SLEEPB _072_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_7 vgnd vpwr scs8hd_fill_1
XFILLER_16_6 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_4.LATCH_1_.latch data_in mem_bottom_ipin_4.LATCH_1_.latch/Q _073_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_0_.latch/Q mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__068__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_12_106 vgnd vpwr scs8hd_decap_8
XFILLER_16_36 vpwr vgnd scs8hd_fill_2
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XANTENNA__084__A _084_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_128 vpwr vgnd scs8hd_fill_2
XFILLER_12_139 vpwr vgnd scs8hd_fill_2
XFILLER_20_150 vgnd vpwr scs8hd_decap_3
X_107_ _076_/B _099_/D address[0] _107_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_7_132 vpwr vgnd scs8hd_fill_2
XFILLER_7_165 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_3 vgnd vpwr scs8hd_fill_1
Xmem_bottom_ipin_6.LATCH_4_.latch data_in mem_bottom_ipin_6.LATCH_4_.latch/Q _086_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__079__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_102 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _045_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__065__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__081__B _082_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_26 vpwr vgnd scs8hd_fill_2
XFILLER_13_48 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_1_.latch/Q mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_0_182 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_5_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_14 vpwr vgnd scs8hd_fill_2
XANTENNA__076__B _076_/B vgnd vpwr scs8hd_diode_2
XANTENNA__092__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_80 vgnd vpwr scs8hd_fill_1
XFILLER_14_91 vgnd vpwr scs8hd_fill_1
XFILLER_10_16 vpwr vgnd scs8hd_fill_2
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XFILLER_27_167 vpwr vgnd scs8hd_fill_2
XFILLER_27_156 vpwr vgnd scs8hd_fill_2
XANTENNA__087__A _127_/A vgnd vpwr scs8hd_diode_2
X_071_ _127_/A _073_/B _071_/Y vgnd vpwr scs8hd_nor2_4
X_140_ _140_/HI _140_/LO vgnd vpwr scs8hd_conb_1
XFILLER_18_145 vgnd vpwr scs8hd_decap_8
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_50 vgnd vpwr scs8hd_fill_1
XFILLER_24_137 vgnd vpwr scs8hd_decap_3
XFILLER_21_37 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_7.LATCH_0_.latch data_in mem_bottom_ipin_7.LATCH_0_.latch/Q _097_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_192 vgnd vpwr scs8hd_decap_6
XFILLER_15_104 vgnd vpwr scs8hd_fill_1
XFILLER_15_159 vgnd vpwr scs8hd_decap_6
X_054_ address[5] address[6] _124_/A vgnd vpwr scs8hd_or2_4
X_123_ _074_/A _121_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_0_.latch/Q mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XANTENNA__068__C address[3] vgnd vpwr scs8hd_diode_2
XANTENNA__084__B _124_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_173 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_100 vpwr vgnd scs8hd_fill_2
XFILLER_11_151 vgnd vpwr scs8hd_fill_1
X_106_ _076_/B _099_/D _059_/C _106_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_93 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_1_.latch/Q mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_3.LATCH_3_.latch/Q mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_69 vpwr vgnd scs8hd_fill_2
XFILLER_27_25 vgnd vpwr scs8hd_decap_4
XANTENNA__079__B _082_/B vgnd vpwr scs8hd_diode_2
XANTENNA__095__A _114_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[7] mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_17_80 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_22_202 vgnd vpwr scs8hd_decap_12
XFILLER_22_224 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_0_ vgnd vpwr scs8hd_inv_1
Xmux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_150 vgnd vpwr scs8hd_decap_4
XFILLER_5_83 vpwr vgnd scs8hd_fill_2
XFILLER_24_59 vgnd vpwr scs8hd_decap_6
XANTENNA__092__B _095_/B vgnd vpwr scs8hd_diode_2
XFILLER_10_205 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_7.LATCH_4_.latch/Q mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _138_/HI vgnd vpwr
+ scs8hd_diode_2
Xmem_top_ipin_0.LATCH_1_.latch data_in mem_top_ipin_0.LATCH_1_.latch/Q _104_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__087__B _086_/B vgnd vpwr scs8hd_diode_2
X_070_ _126_/A _073_/B _070_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_18_102 vpwr vgnd scs8hd_fill_2
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_80 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _141_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_7.LATCH_3_.latch_SLEEPB _094_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_49 vgnd vpwr scs8hd_fill_1
XANTENNA__098__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_7_18 vgnd vpwr scs8hd_fill_1
XFILLER_15_138 vpwr vgnd scs8hd_fill_2
X_122_ _073_/A _121_/B _122_/Y vgnd vpwr scs8hd_nor2_4
X_053_ address[1] _053_/B _059_/C _125_/A vgnd vpwr scs8hd_or3_4
XFILLER_11_93 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_1_.latch/Q mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__068__D _084_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_27 vgnd vpwr scs8hd_decap_4
XFILLER_16_49 vgnd vpwr scs8hd_decap_6
XFILLER_7_123 vpwr vgnd scs8hd_fill_2
XFILLER_7_145 vgnd vpwr scs8hd_decap_3
XFILLER_11_174 vgnd vpwr scs8hd_decap_6
X_105_ _074_/A _100_/B _105_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_61 vgnd vpwr scs8hd_fill_1
XFILLER_8_83 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_0.LATCH_1_.latch data_in mem_bottom_ipin_0.LATCH_1_.latch/Q _115_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_48 vgnd vpwr scs8hd_decap_4
XANTENNA__095__B _095_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_126 vgnd vpwr scs8hd_decap_4
XFILLER_31_214 vgnd vpwr scs8hd_fill_1
Xmem_bottom_ipin_2.LATCH_4_.latch data_in mem_bottom_ipin_2.LATCH_4_.latch/Q _126_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_2_.latch/Q mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_5.LATCH_4_.latch_SLEEPB _078_/Y vgnd vpwr scs8hd_diode_2
XFILLER_13_214 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_38 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_0_.latch/Q mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_232 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_114 vpwr vgnd scs8hd_fill_2
XFILLER_19_16 vpwr vgnd scs8hd_fill_2
XFILLER_35_180 vgnd vpwr scs8hd_decap_6
XFILLER_18_125 vgnd vpwr scs8hd_decap_4
XPHY_70 vgnd vpwr scs8hd_decap_3
XFILLER_25_92 vgnd vpwr scs8hd_fill_1
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_81 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_2.LATCH_3_.latch/Q mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_41 vpwr vgnd scs8hd_fill_2
XFILLER_21_17 vpwr vgnd scs8hd_fill_2
XANTENNA__098__B _098_/B vgnd vpwr scs8hd_diode_2
X_121_ _114_/A _121_/B _121_/Y vgnd vpwr scs8hd_nor2_4
X_052_ address[3] _091_/C vgnd vpwr scs8hd_inv_8
XANTENNA_mem_bottom_ipin_3.LATCH_5_.latch_SLEEPB _056_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_183 vpwr vgnd scs8hd_fill_2
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_120 vgnd vpwr scs8hd_decap_3
XFILLER_28_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _046_/Y vgnd vpwr
+ scs8hd_diode_2
X_104_ _073_/A _100_/B _104_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_bottom_ipin_4.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_113 vpwr vgnd scs8hd_fill_2
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_3.LATCH_0_.latch data_in mem_bottom_ipin_3.LATCH_0_.latch/Q _066_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_71 vpwr vgnd scs8hd_fill_2
XFILLER_22_93 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_6.LATCH_4_.latch/Q mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_201 vgnd vpwr scs8hd_decap_12
XFILLER_4_116 vgnd vpwr scs8hd_fill_1
Xmem_bottom_ipin_5.LATCH_3_.latch data_in mem_bottom_ipin_5.LATCH_3_.latch/Q _079_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_201 vpwr vgnd scs8hd_fill_2
XFILLER_17_93 vpwr vgnd scs8hd_fill_2
XFILLER_3_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_13_18 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _139_/HI mem_top_ipin_0.LATCH_5_.latch/Q
+ mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_13_226 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_5_30 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_72 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_1_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_28 vpwr vgnd scs8hd_fill_2
XFILLER_35_27 vgnd vpwr scs8hd_decap_4
XFILLER_27_137 vpwr vgnd scs8hd_fill_2
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_26_181 vpwr vgnd scs8hd_fill_2
XFILLER_25_71 vpwr vgnd scs8hd_fill_2
XPHY_82 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_64 vgnd vpwr scs8hd_fill_1
XFILLER_24_129 vgnd vpwr scs8hd_decap_4
XFILLER_17_181 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_107 vpwr vgnd scs8hd_fill_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
XFILLER_23_184 vpwr vgnd scs8hd_fill_2
XFILLER_23_173 vpwr vgnd scs8hd_fill_2
X_051_ address[4] _091_/B vgnd vpwr scs8hd_inv_8
X_120_ _127_/A _121_/B _120_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_62 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB _102_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_2_.latch/Q mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_154 vgnd vpwr scs8hd_decap_6
XFILLER_20_187 vpwr vgnd scs8hd_fill_2
XFILLER_28_210 vgnd vpwr scs8hd_fill_1
XFILLER_11_132 vgnd vpwr scs8hd_decap_4
X_103_ _114_/A _100_/B _103_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_169 vgnd vpwr scs8hd_decap_4
XFILLER_11_143 vpwr vgnd scs8hd_fill_2
XFILLER_11_165 vgnd vpwr scs8hd_decap_3
XFILLER_11_187 vpwr vgnd scs8hd_fill_2
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
XFILLER_8_30 vgnd vpwr scs8hd_fill_1
XFILLER_8_41 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_191 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_0_.latch/Q mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_213 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_16_213 vgnd vpwr scs8hd_fill_1
XFILLER_33_82 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_209 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_1.LATCH_3_.latch/Q mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XFILLER_28_93 vpwr vgnd scs8hd_fill_2
XFILLER_5_75 vpwr vgnd scs8hd_fill_2
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_5_20 vpwr vgnd scs8hd_fill_2
XFILLER_24_18 vgnd vpwr scs8hd_decap_12
XFILLER_5_212 vgnd vpwr scs8hd_decap_12
XFILLER_14_84 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__101__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_138 vgnd vpwr scs8hd_decap_4
XFILLER_33_108 vpwr vgnd scs8hd_fill_2
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_26_171 vgnd vpwr scs8hd_fill_1
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_83 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_72 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_5.LATCH_4_.latch/Q mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_160 vpwr vgnd scs8hd_fill_2
XFILLER_17_171 vpwr vgnd scs8hd_fill_2
XFILLER_32_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_050_ address[6] _098_/B vgnd vpwr scs8hd_inv_8
XFILLER_2_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB _115_/Y vgnd vpwr scs8hd_diode_2
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_20_177 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_102_ _127_/A _100_/B _102_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_84 vgnd vpwr scs8hd_decap_8
Xmux_top_ipin_0.INVTX1_0_.scs8hd_inv_1 chanx_left_in[3] mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_211 vgnd vpwr scs8hd_decap_4
XFILLER_8_64 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_6_170 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_1_.latch/Q mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_73 vgnd vpwr scs8hd_decap_4
XFILLER_33_94 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_6_ vgnd vpwr scs8hd_inv_1
XANTENNA__104__A _073_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_140 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_217 vgnd vpwr scs8hd_fill_1
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
XFILLER_0_154 vgnd vpwr scs8hd_fill_1
Xmem_bottom_ipin_1.LATCH_3_.latch data_in mem_bottom_ipin_1.LATCH_3_.latch/Q _120_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_87 vpwr vgnd scs8hd_fill_2
XFILLER_10_209 vgnd vpwr scs8hd_decap_4
XFILLER_30_40 vgnd vpwr scs8hd_fill_1
XFILLER_5_224 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_2_.latch/Q mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__101__B _100_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_227 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_ipin_7.LATCH_0_.latch_SLEEPB _097_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_106 vgnd vpwr scs8hd_decap_4
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_95 vpwr vgnd scs8hd_fill_2
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_84 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_73 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_2_77 vpwr vgnd scs8hd_fill_2
XFILLER_2_11 vgnd vpwr scs8hd_decap_12
XANTENNA__112__A _126_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_0_.latch/Q mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_153 vgnd vpwr scs8hd_fill_1
XFILLER_11_20 vpwr vgnd scs8hd_fill_2
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__107__A _076_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_3 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_0.LATCH_3_.latch/Q mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_145 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_101_ _126_/A _100_/B _101_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_112 vgnd vpwr scs8hd_decap_4
XFILLER_19_223 vpwr vgnd scs8hd_fill_2
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_21 vgnd vpwr scs8hd_decap_3
XFILLER_8_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_1_.latch/Q mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_31_218 vpwr vgnd scs8hd_fill_2
XFILLER_16_215 vgnd vpwr scs8hd_decap_12
XFILLER_17_41 vgnd vpwr scs8hd_fill_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XANTENNA__104__B _100_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_163 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_5.LATCH_1_.latch_SLEEPB _081_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_4.LATCH_2_.latch data_in mem_bottom_ipin_4.LATCH_2_.latch/Q _072_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_4.LATCH_4_.latch/Q mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_199 vgnd vpwr scs8hd_decap_12
XFILLER_8_200 vgnd vpwr scs8hd_fill_1
XANTENNA__115__A _073_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_bottom_ipin_6.LATCH_5_.latch data_in mem_bottom_ipin_6.LATCH_5_.latch/Q _085_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_30 vgnd vpwr scs8hd_fill_1
XFILLER_29_170 vpwr vgnd scs8hd_fill_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _045_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_140 vpwr vgnd scs8hd_fill_2
XFILLER_25_30 vpwr vgnd scs8hd_fill_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_85 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_74 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_4.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_89 vgnd vpwr scs8hd_decap_3
XFILLER_2_67 vgnd vpwr scs8hd_fill_1
XFILLER_2_45 vgnd vpwr scs8hd_decap_3
XFILLER_2_23 vgnd vpwr scs8hd_decap_8
XANTENNA__112__B _114_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_5.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_140 vgnd vpwr scs8hd_decap_6
XFILLER_17_184 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_1_.latch/Q mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_3.LATCH_2_.latch_SLEEPB _062_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_132 vpwr vgnd scs8hd_fill_2
XFILLER_11_32 vpwr vgnd scs8hd_fill_2
XFILLER_14_154 vgnd vpwr scs8hd_fill_1
XANTENNA__107__B _099_/D vgnd vpwr scs8hd_diode_2
XFILLER_14_187 vgnd vpwr scs8hd_decap_4
XANTENNA__123__A _074_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_102 vpwr vgnd scs8hd_fill_2
XFILLER_20_135 vgnd vpwr scs8hd_fill_1
XFILLER_9_191 vgnd vpwr scs8hd_decap_4
XFILLER_28_213 vgnd vpwr scs8hd_fill_1
XFILLER_28_202 vpwr vgnd scs8hd_fill_2
X_100_ _125_/A _100_/B _100_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_117 vgnd vpwr scs8hd_decap_3
XFILLER_7_128 vpwr vgnd scs8hd_fill_2
XFILLER_22_75 vgnd vpwr scs8hd_decap_6
XFILLER_34_227 vgnd vpwr scs8hd_decap_6
XANTENNA__118__A _125_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_2_.latch/Q mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_205 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_6
XFILLER_16_227 vgnd vpwr scs8hd_decap_6
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XFILLER_17_97 vpwr vgnd scs8hd_fill_2
XFILLER_3_197 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_7.LATCH_1_.latch data_in mem_bottom_ipin_7.LATCH_1_.latch/Q _096_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__120__B _121_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_1.LATCH_3_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_134 vpwr vgnd scs8hd_fill_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_12
XFILLER_0_178 vpwr vgnd scs8hd_fill_2
XFILLER_28_30 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_0_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_34 vpwr vgnd scs8hd_fill_2
XANTENNA__115__B _114_/B vgnd vpwr scs8hd_diode_2
XFILLER_14_43 vpwr vgnd scs8hd_fill_2
XFILLER_14_76 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_182 vgnd vpwr scs8hd_fill_1
XANTENNA__126__A _126_/A vgnd vpwr scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_185 vpwr vgnd scs8hd_fill_2
XFILLER_26_163 vpwr vgnd scs8hd_fill_2
XFILLER_26_152 vgnd vpwr scs8hd_fill_1
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_25_75 vpwr vgnd scs8hd_fill_2
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_75 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_32_166 vgnd vpwr scs8hd_decap_8
XFILLER_32_100 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_1_.latch/Q mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_100 vpwr vgnd scs8hd_fill_2
XFILLER_23_188 vpwr vgnd scs8hd_fill_2
XFILLER_23_177 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_66 vgnd vpwr scs8hd_fill_1
XFILLER_14_166 vgnd vpwr scs8hd_decap_8
XANTENNA__107__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__123__B _121_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_170 vpwr vgnd scs8hd_fill_2
XFILLER_20_114 vgnd vpwr scs8hd_decap_3
XFILLER_20_125 vpwr vgnd scs8hd_fill_2
XFILLER_20_169 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_3.LATCH_4_.latch/Q mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_2_.latch/Q mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_147 vgnd vpwr scs8hd_decap_4
XFILLER_22_43 vpwr vgnd scs8hd_fill_2
XFILLER_22_98 vgnd vpwr scs8hd_fill_1
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_0.LATCH_2_.latch data_in mem_top_ipin_0.LATCH_2_.latch/Q _103_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__118__B _121_/B vgnd vpwr scs8hd_diode_2
X_159_ chanx_left_in[0] chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_6_140 vpwr vgnd scs8hd_fill_2
XFILLER_8_89 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_25_217 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__044__A _044_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_53 vpwr vgnd scs8hd_fill_2
XFILLER_3_132 vpwr vgnd scs8hd_fill_2
XANTENNA__129__A _073_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_231 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _138_/HI mem_bottom_ipin_7.LATCH_5_.latch/Q
+ mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_0_146 vpwr vgnd scs8hd_fill_2
XFILLER_0_168 vgnd vpwr scs8hd_decap_6
XFILLER_28_97 vgnd vpwr scs8hd_decap_4
XFILLER_28_64 vpwr vgnd scs8hd_fill_2
XFILLER_8_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_79 vpwr vgnd scs8hd_fill_2
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XFILLER_5_24 vgnd vpwr scs8hd_decap_4
XFILLER_14_88 vgnd vpwr scs8hd_fill_1
XFILLER_30_43 vgnd vpwr scs8hd_decap_12
XFILLER_30_32 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_2_.latch data_in mem_bottom_ipin_0.LATCH_2_.latch/Q _114_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__126__B _127_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__142__A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__052__A address[3] vgnd vpwr scs8hd_diode_2
XPHY_65 vgnd vpwr scs8hd_decap_3
Xmem_bottom_ipin_2.LATCH_5_.latch data_in mem_bottom_ipin_2.LATCH_5_.latch/Q _125_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_76 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_6.LATCH_3_.latch_SLEEPB _087_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_164 vpwr vgnd scs8hd_fill_2
XFILLER_32_178 vgnd vpwr scs8hd_decap_12
XFILLER_32_112 vgnd vpwr scs8hd_decap_12
XFILLER_17_175 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_2_.latch/Q mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_156 vgnd vpwr scs8hd_decap_4
XANTENNA__047__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_11_12 vpwr vgnd scs8hd_fill_2
XFILLER_2_7 vpwr vgnd scs8hd_fill_2
XFILLER_11_45 vpwr vgnd scs8hd_fill_2
XFILLER_11_78 vgnd vpwr scs8hd_decap_6
XFILLER_11_89 vpwr vgnd scs8hd_fill_2
XFILLER_14_145 vgnd vpwr scs8hd_decap_8
XFILLER_9_182 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_0_.latch/Q mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_46 vpwr vgnd scs8hd_fill_2
XFILLER_8_57 vgnd vpwr scs8hd_decap_4
XFILLER_8_68 vpwr vgnd scs8hd_fill_2
XFILLER_8_79 vpwr vgnd scs8hd_fill_2
X_158_ chanx_left_in[1] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_6_152 vgnd vpwr scs8hd_fill_1
XFILLER_6_174 vgnd vpwr scs8hd_decap_4
X_089_ _073_/A _086_/B _089_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__150__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_12_ vgnd vpwr scs8hd_inv_1
XFILLER_25_229 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__060__A _056_/B vgnd vpwr scs8hd_diode_2
XFILLER_17_11 vgnd vpwr scs8hd_decap_3
XFILLER_17_33 vpwr vgnd scs8hd_fill_2
XFILLER_17_77 vgnd vpwr scs8hd_fill_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_10 vgnd vpwr scs8hd_decap_12
XANTENNA__129__B _127_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_4.LATCH_4_.latch_SLEEPB _070_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__145__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_0_80 vgnd vpwr scs8hd_fill_1
XANTENNA__055__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_210 vpwr vgnd scs8hd_fill_2
XFILLER_28_32 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_1_.latch/Q mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_210 vgnd vpwr scs8hd_decap_4
XFILLER_8_203 vpwr vgnd scs8hd_fill_2
XFILLER_12_232 vgnd vpwr scs8hd_fill_1
Xmem_bottom_ipin_3.LATCH_1_.latch data_in mem_bottom_ipin_3.LATCH_1_.latch/Q _064_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_4_ vgnd vpwr scs8hd_inv_1
XFILLER_30_55 vgnd vpwr scs8hd_decap_4
XFILLER_29_184 vgnd vpwr scs8hd_decap_6
XFILLER_29_140 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_2.LATCH_4_.latch/Q mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_5.LATCH_4_.latch data_in mem_bottom_ipin_5.LATCH_4_.latch/Q _078_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_187 vgnd vpwr scs8hd_decap_12
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_154 vpwr vgnd scs8hd_fill_2
XFILLER_25_99 vpwr vgnd scs8hd_fill_2
XFILLER_25_88 vgnd vpwr scs8hd_decap_4
XFILLER_25_11 vgnd vpwr scs8hd_decap_3
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_77 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_1_220 vgnd vpwr scs8hd_decap_12
XFILLER_17_110 vpwr vgnd scs8hd_fill_2
XFILLER_17_132 vpwr vgnd scs8hd_fill_2
XFILLER_32_124 vgnd vpwr scs8hd_decap_12
XANTENNA__153__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__063__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_11_24 vgnd vpwr scs8hd_fill_1
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__148__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_150 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _137_/HI mem_bottom_ipin_6.LATCH_5_.latch/Q
+ mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_3_91 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_138 vpwr vgnd scs8hd_fill_2
XANTENNA__058__A _056_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_23 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_227 vgnd vpwr scs8hd_decap_6
X_157_ chanx_left_in[2] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_10_193 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_ipin_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_197 vgnd vpwr scs8hd_fill_1
X_088_ _114_/A _086_/B _088_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__060__B _127_/A vgnd vpwr scs8hd_diode_2
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_230 vgnd vpwr scs8hd_decap_3
XFILLER_33_22 vgnd vpwr scs8hd_decap_12
XFILLER_3_167 vgnd vpwr scs8hd_decap_12
XFILLER_3_112 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__055__B _091_/B vgnd vpwr scs8hd_diode_2
XANTENNA__071__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_77 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_6.LATCH_0_.latch data_in mem_bottom_ipin_6.LATCH_0_.latch/Q _090_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_2_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XANTENNA__156__A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_6.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__066__A _056_/B vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_7.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_174 vgnd vpwr scs8hd_decap_8
XFILLER_29_163 vgnd vpwr scs8hd_decap_4
XFILLER_35_199 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_0_.latch/Q mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_144 vgnd vpwr scs8hd_decap_8
XFILLER_26_111 vgnd vpwr scs8hd_fill_1
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_25_34 vpwr vgnd scs8hd_fill_2
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_78 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_232 vgnd vpwr scs8hd_fill_1
XFILLER_32_136 vgnd vpwr scs8hd_decap_12
XFILLER_23_136 vpwr vgnd scs8hd_fill_2
XFILLER_23_114 vgnd vpwr scs8hd_decap_3
XANTENNA__063__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_22_191 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_106 vgnd vpwr scs8hd_decap_8
XFILLER_9_195 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_1_.latch/Q mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_206 vgnd vpwr scs8hd_decap_4
XANTENNA__058__B _126_/A vgnd vpwr scs8hd_diode_2
XANTENNA__074__A _074_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _044_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_19_217 vpwr vgnd scs8hd_fill_2
X_156_ chanx_left_in[3] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_6_110 vpwr vgnd scs8hd_fill_2
XFILLER_6_154 vgnd vpwr scs8hd_decap_4
XFILLER_8_26 vgnd vpwr scs8hd_decap_4
XFILLER_8_37 vpwr vgnd scs8hd_fill_2
XFILLER_10_161 vpwr vgnd scs8hd_fill_2
X_087_ _127_/A _086_/B _087_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_6 vpwr vgnd scs8hd_fill_2
XFILLER_6_187 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__159__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__069__A _125_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_7.LATCH_5_.latch_SLEEPB _092_/Y vgnd vpwr scs8hd_diode_2
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_34 vgnd vpwr scs8hd_decap_12
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
XFILLER_33_78 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_1.LATCH_4_.latch/Q mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
X_139_ _139_/HI _139_/LO vgnd vpwr scs8hd_conb_1
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XANTENNA__055__C _091_/C vgnd vpwr scs8hd_diode_2
XFILLER_21_223 vpwr vgnd scs8hd_fill_2
XANTENNA__071__B _073_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_105 vpwr vgnd scs8hd_fill_2
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_0_138 vgnd vpwr scs8hd_decap_4
XFILLER_28_89 vgnd vpwr scs8hd_decap_3
XFILLER_28_56 vgnd vpwr scs8hd_decap_8
XFILLER_28_45 vgnd vpwr scs8hd_decap_8
XFILLER_28_23 vgnd vpwr scs8hd_fill_1
XFILLER_8_227 vgnd vpwr scs8hd_decap_6
XFILLER_5_38 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _139_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_47 vgnd vpwr scs8hd_decap_12
XANTENNA__066__B _074_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_79 vgnd vpwr scs8hd_decap_12
XANTENNA__082__A _074_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _136_/HI mem_bottom_ipin_5.LATCH_5_.latch/Q
+ mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_156 vgnd vpwr scs8hd_decap_12
XFILLER_6_81 vgnd vpwr scs8hd_decap_6
XFILLER_26_167 vgnd vpwr scs8hd_decap_4
XFILLER_26_123 vpwr vgnd scs8hd_fill_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A _125_/A vgnd vpwr scs8hd_diode_2
XPHY_35 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XPHY_79 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_3 vpwr vgnd scs8hd_fill_2
XFILLER_32_148 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_104 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_1.LATCH_4_.latch data_in mem_bottom_ipin_1.LATCH_4_.latch/Q _119_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__063__C _059_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_129 vgnd vpwr scs8hd_decap_6
XFILLER_9_174 vgnd vpwr scs8hd_decap_8
XFILLER_3_71 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_2_.latch/Q mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
XFILLER_22_47 vgnd vpwr scs8hd_decap_12
XANTENNA__074__B _073_/B vgnd vpwr scs8hd_diode_2
XANTENNA__090__A _074_/A vgnd vpwr scs8hd_diode_2
X_155_ chanx_left_in[4] chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_6_144 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_086_ _126_/A _086_/B _086_/Y vgnd vpwr scs8hd_nor2_4
Xmem_top_ipin_2.LATCH_0_.latch data_in _046_/A _109_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__069__B _073_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_57 vgnd vpwr scs8hd_decap_4
XFILLER_33_46 vgnd vpwr scs8hd_decap_3
XANTENNA__085__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_136 vpwr vgnd scs8hd_fill_2
XFILLER_15_221 vpwr vgnd scs8hd_fill_2
XFILLER_30_202 vgnd vpwr scs8hd_decap_12
X_069_ _125_/A _073_/B _069_/Y vgnd vpwr scs8hd_nor2_4
X_138_ _138_/HI _138_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_72 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__055__D _124_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_202 vgnd vpwr scs8hd_fill_1
XFILLER_12_224 vgnd vpwr scs8hd_decap_8
XFILLER_14_15 vpwr vgnd scs8hd_fill_2
XFILLER_14_59 vpwr vgnd scs8hd_fill_2
XFILLER_30_69 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__082__B _082_/B vgnd vpwr scs8hd_diode_2
XFILLER_29_132 vgnd vpwr scs8hd_decap_8
Xmem_bottom_ipin_2.LATCH_0_.latch data_in mem_bottom_ipin_2.LATCH_0_.latch/Q _130_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_80 vgnd vpwr scs8hd_fill_1
XFILLER_20_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_ipin_6.LATCH_0_.latch_SLEEPB _090_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_1_.latch/Q mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_168 vgnd vpwr scs8hd_decap_12
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_102 vgnd vpwr scs8hd_fill_1
XFILLER_25_25 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XANTENNA__077__B _082_/B vgnd vpwr scs8hd_diode_2
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__093__A _126_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_4.LATCH_3_.latch data_in mem_bottom_ipin_4.LATCH_3_.latch/Q _071_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_146 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_182 vgnd vpwr scs8hd_fill_1
XFILLER_31_171 vgnd vpwr scs8hd_decap_3
XFILLER_23_149 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_0.LATCH_4_.latch/Q mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_16 vpwr vgnd scs8hd_fill_2
XFILLER_11_49 vpwr vgnd scs8hd_fill_2
XANTENNA__088__A _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_116 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_193 vpwr vgnd scs8hd_fill_2
XFILLER_28_219 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_108 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_2_.latch/Q mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_59 vgnd vpwr scs8hd_fill_1
XANTENNA__090__B _086_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_154_ chanx_left_in[5] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_6_123 vpwr vgnd scs8hd_fill_2
X_085_ _125_/A _086_/B _085_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_18_230 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_4.LATCH_1_.latch_SLEEPB _073_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_37 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _135_/HI mem_bottom_ipin_4.LATCH_5_.latch/Q
+ mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__085__B _086_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_159 vpwr vgnd scs8hd_fill_2
XFILLER_3_115 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_137_ _137_/HI _137_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB _100_/Y vgnd vpwr scs8hd_diode_2
X_068_ _091_/A address[4] address[3] _084_/A _073_/B vgnd vpwr scs8hd_or4_4
XFILLER_9_60 vgnd vpwr scs8hd_fill_1
XANTENNA__096__A _073_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_207 vgnd vpwr scs8hd_decap_6
XFILLER_18_91 vgnd vpwr scs8hd_fill_1
XFILLER_30_59 vgnd vpwr scs8hd_fill_1
XFILLER_29_111 vgnd vpwr scs8hd_fill_1
XFILLER_35_125 vgnd vpwr scs8hd_decap_12
XFILLER_29_90 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_2_.latch/Q mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_ipin_7.LATCH_2_.latch data_in mem_bottom_ipin_7.LATCH_2_.latch/Q _095_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_59 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA__093__B _095_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_136 vpwr vgnd scs8hd_fill_2
XFILLER_31_91 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_28 vpwr vgnd scs8hd_fill_2
XANTENNA__088__B _086_/B vgnd vpwr scs8hd_diode_2
XFILLER_14_128 vgnd vpwr scs8hd_decap_6
XFILLER_9_110 vgnd vpwr scs8hd_fill_1
XFILLER_9_187 vpwr vgnd scs8hd_fill_2
XFILLER_3_95 vpwr vgnd scs8hd_fill_2
XFILLER_3_62 vgnd vpwr scs8hd_decap_3
XANTENNA__099__A _091_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
X_153_ chanx_left_in[6] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_6_102 vpwr vgnd scs8hd_fill_2
X_084_ _084_/A _124_/B _086_/B vgnd vpwr scs8hd_or2_4
XFILLER_33_201 vpwr vgnd scs8hd_fill_2
XFILLER_17_16 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_7.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_1_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_136_ _136_/HI _136_/LO vgnd vpwr scs8hd_conb_1
X_067_ address[5] _098_/B _084_/A vgnd vpwr scs8hd_nand2_4
XANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB _113_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_26 vgnd vpwr scs8hd_decap_4
XANTENNA__096__B _095_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_70 vpwr vgnd scs8hd_fill_2
XFILLER_18_81 vpwr vgnd scs8hd_fill_2
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_0.INVTX1_2_.scs8hd_inv_1 chanx_left_in[7] mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_119_ _126_/A _121_/B _119_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_230 vgnd vpwr scs8hd_decap_3
Xmem_top_ipin_0.LATCH_3_.latch data_in mem_top_ipin_0.LATCH_3_.latch/Q _102_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_167 vgnd vpwr scs8hd_fill_1
XFILLER_29_145 vpwr vgnd scs8hd_fill_2
XFILLER_35_137 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_2_.latch/Q mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _043_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_159 vpwr vgnd scs8hd_fill_2
XFILLER_25_38 vpwr vgnd scs8hd_fill_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _134_/HI mem_bottom_ipin_3.LATCH_5_.latch/Q
+ mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_31_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_9_133 vpwr vgnd scs8hd_fill_2
XFILLER_9_166 vpwr vgnd scs8hd_fill_2
XFILLER_13_162 vpwr vgnd scs8hd_fill_2
XFILLER_3_52 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_0.LATCH_3_.latch data_in mem_bottom_ipin_0.LATCH_3_.latch/Q _113_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_210 vgnd vpwr scs8hd_decap_4
XANTENNA__099__B address[4] vgnd vpwr scs8hd_diode_2
X_152_ chanx_left_in[7] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
X_083_ _091_/A _091_/B address[3] _124_/B vgnd vpwr scs8hd_or3_4
XFILLER_6_158 vgnd vpwr scs8hd_fill_1
XFILLER_10_165 vgnd vpwr scs8hd_decap_3
XFILLER_10_187 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_ipin_7.LATCH_2_.latch_SLEEPB _095_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_210 vgnd vpwr scs8hd_decap_4
XFILLER_24_202 vgnd vpwr scs8hd_decap_12
XFILLER_3_106 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_135_ _135_/HI _135_/LO vgnd vpwr scs8hd_conb_1
XFILLER_23_82 vgnd vpwr scs8hd_decap_3
X_066_ _056_/B _074_/A _066_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_6 vpwr vgnd scs8hd_fill_2
XFILLER_9_62 vpwr vgnd scs8hd_fill_2
XFILLER_9_73 vgnd vpwr scs8hd_decap_4
XFILLER_21_227 vpwr vgnd scs8hd_fill_2
XFILLER_0_109 vgnd vpwr scs8hd_decap_4
X_118_ _125_/A _121_/B _118_/Y vgnd vpwr scs8hd_nor2_4
X_049_ enable _091_/A vgnd vpwr scs8hd_inv_8
XFILLER_22_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_201 vpwr vgnd scs8hd_fill_2
XFILLER_20_72 vgnd vpwr scs8hd_decap_8
XFILLER_20_83 vgnd vpwr scs8hd_decap_8
XFILLER_29_70 vgnd vpwr scs8hd_decap_4
XFILLER_35_149 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.LATCH_3_.latch_SLEEPB _079_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_127 vpwr vgnd scs8hd_fill_2
XFILLER_26_105 vgnd vpwr scs8hd_decap_6
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_25_193 vpwr vgnd scs8hd_fill_2
XFILLER_31_82 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_23_119 vgnd vpwr scs8hd_decap_3
XFILLER_23_108 vgnd vpwr scs8hd_fill_1
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_1_.latch/Q mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_108 vgnd vpwr scs8hd_decap_8
Xmem_bottom_ipin_3.LATCH_2_.latch data_in mem_bottom_ipin_3.LATCH_2_.latch/Q _062_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_4_ vgnd vpwr scs8hd_inv_1
XFILLER_26_60 vpwr vgnd scs8hd_fill_2
XFILLER_9_123 vgnd vpwr scs8hd_decap_3
XFILLER_9_156 vgnd vpwr scs8hd_fill_1
XFILLER_3_31 vpwr vgnd scs8hd_fill_2
XFILLER_22_29 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__099__C address[3] vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_5.LATCH_5_.latch data_in mem_bottom_ipin_5.LATCH_5_.latch/Q _077_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_100 vpwr vgnd scs8hd_fill_2
X_151_ chanx_left_in[8] chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_10_177 vgnd vpwr scs8hd_decap_8
XFILLER_12_73 vpwr vgnd scs8hd_fill_2
X_082_ _074_/A _082_/B _082_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_18_222 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_3.LATCH_4_.latch_SLEEPB _058_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_2_.latch/Q mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_225 vgnd vpwr scs8hd_decap_8
X_134_ _134_/HI _134_/LO vgnd vpwr scs8hd_conb_1
X_065_ address[1] address[2] address[0] _074_/A vgnd vpwr scs8hd_or3_4
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XFILLER_0_76 vpwr vgnd scs8hd_fill_2
XFILLER_21_206 vpwr vgnd scs8hd_fill_2
XFILLER_9_41 vgnd vpwr scs8hd_fill_1
XFILLER_9_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _133_/HI mem_bottom_ipin_2.LATCH_5_.latch/Q
+ mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
X_117_ _124_/A _076_/B _121_/B vgnd vpwr scs8hd_or2_4
XFILLER_7_210 vgnd vpwr scs8hd_decap_12
X_048_ address[2] _053_/B vgnd vpwr scs8hd_inv_8
XFILLER_15_3 vgnd vpwr scs8hd_decap_3
XFILLER_14_19 vgnd vpwr scs8hd_decap_12
XFILLER_30_18 vgnd vpwr scs8hd_decap_12
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XFILLER_29_103 vpwr vgnd scs8hd_fill_2
XFILLER_4_213 vgnd vpwr scs8hd_fill_1
XFILLER_35_106 vgnd vpwr scs8hd_decap_12
XFILLER_6_20 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB _108_/Y vgnd vpwr scs8hd_diode_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_25_150 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_5_.latch_SLEEPB _118_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_62 vgnd vpwr scs8hd_decap_3
XANTENNA__102__A _127_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_6.LATCH_1_.latch data_in mem_bottom_ipin_6.LATCH_1_.latch/Q _089_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_197 vpwr vgnd scs8hd_fill_2
XFILLER_26_72 vgnd vpwr scs8hd_fill_1
XFILLER_9_102 vpwr vgnd scs8hd_fill_2
XFILLER_9_146 vpwr vgnd scs8hd_fill_2
XFILLER_13_142 vgnd vpwr scs8hd_fill_1
XFILLER_13_175 vpwr vgnd scs8hd_fill_2
XFILLER_13_197 vpwr vgnd scs8hd_fill_2
XFILLER_3_87 vpwr vgnd scs8hd_fill_2
XANTENNA__099__D _099_/D vgnd vpwr scs8hd_diode_2
X_150_ chanx_right_in[0] chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_10_123 vpwr vgnd scs8hd_fill_2
XFILLER_10_134 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_127 vgnd vpwr scs8hd_decap_4
X_081_ _073_/A _082_/B _081_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_145 vgnd vpwr scs8hd_decap_8
XFILLER_12_63 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_119 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB _103_/Y vgnd vpwr scs8hd_diode_2
X_133_ _133_/HI _133_/LO vgnd vpwr scs8hd_conb_1
Xmux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_62 vgnd vpwr scs8hd_decap_4
XFILLER_2_152 vgnd vpwr scs8hd_fill_1
X_064_ _056_/B _073_/A _064_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_44 vgnd vpwr scs8hd_decap_6
XANTENNA__110__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_7 vpwr vgnd scs8hd_fill_2
XFILLER_9_53 vgnd vpwr scs8hd_decap_4
XFILLER_7_222 vgnd vpwr scs8hd_decap_8
X_116_ _074_/A _114_/B _116_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__105__A _074_/A vgnd vpwr scs8hd_diode_2
X_047_ address[1] _059_/A vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _044_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_1_.latch/Q mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_4.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_30 vgnd vpwr scs8hd_fill_1
XFILLER_35_118 vgnd vpwr scs8hd_decap_6
XFILLER_29_50 vgnd vpwr scs8hd_decap_8
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_15_30 vpwr vgnd scs8hd_fill_2
XFILLER_15_74 vpwr vgnd scs8hd_fill_2
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XFILLER_31_51 vgnd vpwr scs8hd_decap_8
XANTENNA__102__B _100_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_151 vpwr vgnd scs8hd_fill_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_176 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_2_.latch/Q mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_22_110 vgnd vpwr scs8hd_decap_8
XFILLER_22_154 vpwr vgnd scs8hd_fill_2
XFILLER_7_6 vpwr vgnd scs8hd_fill_2
XFILLER_26_84 vgnd vpwr scs8hd_decap_8
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_110 vgnd vpwr scs8hd_decap_4
XFILLER_13_121 vgnd vpwr scs8hd_fill_1
XFILLER_13_132 vgnd vpwr scs8hd_decap_4
XFILLER_13_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__113__A _127_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _132_/HI mem_bottom_ipin_1.LATCH_5_.latch/Q
+ mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_6_106 vpwr vgnd scs8hd_fill_2
X_080_ _114_/A _082_/B _080_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_157 vpwr vgnd scs8hd_fill_2
XFILLER_5_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_6.LATCH_5_.latch_SLEEPB _085_/Y vgnd vpwr scs8hd_diode_2
XFILLER_33_205 vgnd vpwr scs8hd_decap_12
XANTENNA__108__A _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_219 vgnd vpwr scs8hd_decap_12
X_063_ address[1] address[2] _059_/C _073_/A vgnd vpwr scs8hd_or3_4
Xmem_bottom_ipin_1.LATCH_5_.latch data_in mem_bottom_ipin_1.LATCH_5_.latch/Q _118_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_132_ _132_/HI _132_/LO vgnd vpwr scs8hd_conb_1
XFILLER_23_41 vgnd vpwr scs8hd_decap_3
XFILLER_2_186 vgnd vpwr scs8hd_decap_12
XANTENNA__110__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_19 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_41 vgnd vpwr scs8hd_decap_3
XFILLER_18_74 vgnd vpwr scs8hd_decap_4
XFILLER_18_85 vgnd vpwr scs8hd_decap_6
X_046_ _046_/A _046_/Y vgnd vpwr scs8hd_inv_8
X_115_ _073_/A _114_/B _115_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__105__B _100_/B vgnd vpwr scs8hd_diode_2
XANTENNA__121__A _114_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_149 vgnd vpwr scs8hd_decap_3
Xmem_top_ipin_2.LATCH_1_.latch data_in _045_/A _108_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XFILLER_29_62 vpwr vgnd scs8hd_fill_2
XANTENNA__116__A _074_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_66 vpwr vgnd scs8hd_fill_2
XFILLER_6_77 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_34_141 vgnd vpwr scs8hd_decap_12
XFILLER_19_171 vpwr vgnd scs8hd_fill_2
XFILLER_19_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_25_130 vpwr vgnd scs8hd_fill_2
XFILLER_25_174 vpwr vgnd scs8hd_fill_2
XFILLER_15_86 vgnd vpwr scs8hd_fill_1
XFILLER_31_74 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

