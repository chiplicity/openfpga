VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cby_3__1_
  CLASS BLOCK ;
  FOREIGN cby_3__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 200.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.070 197.600 29.350 200.000 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.830 197.600 32.110 200.000 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.050 197.600 35.330 200.000 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 197.600 38.550 200.000 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.490 197.600 41.770 200.000 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 197.600 44.530 200.000 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.470 197.600 47.750 200.000 ;
    END
  END address[6]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 197.600 1.750 200.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.230 197.600 4.510 200.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 197.600 7.730 200.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.670 197.600 10.950 200.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.430 197.600 13.710 200.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 197.600 16.930 200.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.870 197.600 20.150 200.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.630 197.600 22.910 200.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.850 197.600 26.130 200.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 53.450 197.600 53.730 200.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.670 197.600 56.950 200.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.890 197.600 60.170 200.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 62.650 197.600 62.930 200.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.870 197.600 66.150 200.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.090 197.600 69.370 200.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.850 197.600 72.130 200.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.070 197.600 75.350 200.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.290 197.600 78.570 200.000 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 197.600 50.970 200.000 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 2.400 ;
    END
  END enable
  PIN left_grid_pin_1_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.400 33.960 ;
    END
  END left_grid_pin_1_
  PIN left_grid_pin_5_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END left_grid_pin_5_
  PIN left_grid_pin_9_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 2.400 167.240 ;
    END
  END left_grid_pin_9_
  PIN right_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 12.280 80.000 12.880 ;
    END
  END right_grid_pin_0_
  PIN right_grid_pin_10_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 136.720 80.000 137.320 ;
    END
  END right_grid_pin_10_
  PIN right_grid_pin_12_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 161.880 80.000 162.480 ;
    END
  END right_grid_pin_12_
  PIN right_grid_pin_14_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 187.040 80.000 187.640 ;
    END
  END right_grid_pin_14_
  PIN right_grid_pin_2_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 36.760 80.000 37.360 ;
    END
  END right_grid_pin_2_
  PIN right_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 61.920 80.000 62.520 ;
    END
  END right_grid_pin_4_
  PIN right_grid_pin_6_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 87.080 80.000 87.680 ;
    END
  END right_grid_pin_6_
  PIN right_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 112.240 80.000 112.840 ;
    END
  END right_grid_pin_8_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 18.055 10.640 19.655 187.920 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 31.385 10.640 32.985 187.920 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 74.060 187.765 ;
      LAYER met1 ;
        RECT 0.530 0.380 79.050 198.180 ;
      LAYER met2 ;
        RECT 0.550 197.320 1.190 198.290 ;
        RECT 2.030 197.320 3.950 198.290 ;
        RECT 4.790 197.320 7.170 198.290 ;
        RECT 8.010 197.320 10.390 198.290 ;
        RECT 11.230 197.320 13.150 198.290 ;
        RECT 13.990 197.320 16.370 198.290 ;
        RECT 17.210 197.320 19.590 198.290 ;
        RECT 20.430 197.320 22.350 198.290 ;
        RECT 23.190 197.320 25.570 198.290 ;
        RECT 26.410 197.320 28.790 198.290 ;
        RECT 29.630 197.320 31.550 198.290 ;
        RECT 32.390 197.320 34.770 198.290 ;
        RECT 35.610 197.320 37.990 198.290 ;
        RECT 38.830 197.320 41.210 198.290 ;
        RECT 42.050 197.320 43.970 198.290 ;
        RECT 44.810 197.320 47.190 198.290 ;
        RECT 48.030 197.320 50.410 198.290 ;
        RECT 51.250 197.320 53.170 198.290 ;
        RECT 54.010 197.320 56.390 198.290 ;
        RECT 57.230 197.320 59.610 198.290 ;
        RECT 60.450 197.320 62.370 198.290 ;
        RECT 63.210 197.320 65.590 198.290 ;
        RECT 66.430 197.320 68.810 198.290 ;
        RECT 69.650 197.320 71.570 198.290 ;
        RECT 72.410 197.320 74.790 198.290 ;
        RECT 75.630 197.320 78.010 198.290 ;
        RECT 78.850 197.320 79.020 198.290 ;
        RECT 0.550 2.680 79.020 197.320 ;
        RECT 0.550 0.270 1.650 2.680 ;
        RECT 2.490 0.270 5.790 2.680 ;
        RECT 6.630 0.270 9.930 2.680 ;
        RECT 10.770 0.270 14.070 2.680 ;
        RECT 14.910 0.270 18.210 2.680 ;
        RECT 19.050 0.270 22.350 2.680 ;
        RECT 23.190 0.270 26.490 2.680 ;
        RECT 27.330 0.270 31.090 2.680 ;
        RECT 31.930 0.270 35.230 2.680 ;
        RECT 36.070 0.270 39.370 2.680 ;
        RECT 40.210 0.270 43.510 2.680 ;
        RECT 44.350 0.270 47.650 2.680 ;
        RECT 48.490 0.270 51.790 2.680 ;
        RECT 52.630 0.270 56.390 2.680 ;
        RECT 57.230 0.270 60.530 2.680 ;
        RECT 61.370 0.270 64.670 2.680 ;
        RECT 65.510 0.270 68.810 2.680 ;
        RECT 69.650 0.270 72.950 2.680 ;
        RECT 73.790 0.270 77.090 2.680 ;
        RECT 77.930 0.270 79.020 2.680 ;
      LAYER met3 ;
        RECT 0.310 186.640 77.200 187.845 ;
        RECT 0.310 167.640 77.890 186.640 ;
        RECT 2.800 166.240 77.890 167.640 ;
        RECT 0.310 162.880 77.890 166.240 ;
        RECT 0.310 161.480 77.200 162.880 ;
        RECT 0.310 137.720 77.890 161.480 ;
        RECT 0.310 136.320 77.200 137.720 ;
        RECT 0.310 113.240 77.890 136.320 ;
        RECT 0.310 111.840 77.200 113.240 ;
        RECT 0.310 101.000 77.890 111.840 ;
        RECT 2.800 99.600 77.890 101.000 ;
        RECT 0.310 88.080 77.890 99.600 ;
        RECT 0.310 86.680 77.200 88.080 ;
        RECT 0.310 62.920 77.890 86.680 ;
        RECT 0.310 61.520 77.200 62.920 ;
        RECT 0.310 37.760 77.890 61.520 ;
        RECT 0.310 36.360 77.200 37.760 ;
        RECT 0.310 34.360 77.890 36.360 ;
        RECT 2.800 32.960 77.890 34.360 ;
        RECT 0.310 13.280 77.890 32.960 ;
        RECT 0.310 11.880 77.200 13.280 ;
        RECT 0.310 0.175 77.890 11.880 ;
      LAYER met4 ;
        RECT 20.055 10.240 30.985 187.920 ;
        RECT 33.385 10.240 72.985 187.920 ;
        RECT 18.050 0.175 72.985 10.240 ;
  END
END cby_3__1_
END LIBRARY

