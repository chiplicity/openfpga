magic
tech sky130A
magscale 1 2
timestamp 1608763569
<< checkpaint >>
rect -1260 -1260 21260 18260
<< locali >>
rect 12357 10999 12391 11101
rect 12357 10965 12449 10999
rect 3525 8347 3559 8585
rect 7389 8347 7423 8585
rect 3249 6647 3283 6817
rect 3893 5627 3927 5729
rect 4445 5695 4479 5865
rect 2145 4471 2179 4641
rect 6193 4471 6227 4777
rect 6837 3587 6871 3689
rect 12265 3383 12299 3621
rect 14013 3383 14047 3485
rect 14473 3451 14507 3553
rect 8861 2499 8895 2601
rect 14749 2295 14783 2533
<< viali >>
rect 1961 14569 1995 14603
rect 1777 14433 1811 14467
rect 1869 14025 1903 14059
rect 2421 14025 2455 14059
rect 3525 14025 3559 14059
rect 7021 14025 7055 14059
rect 2973 13957 3007 13991
rect 6193 13957 6227 13991
rect 14657 13957 14691 13991
rect 1685 13821 1719 13855
rect 2237 13821 2271 13855
rect 2789 13821 2823 13855
rect 3341 13821 3375 13855
rect 6009 13821 6043 13855
rect 6837 13821 6871 13855
rect 13645 13821 13679 13855
rect 14473 13821 14507 13855
rect 15117 13821 15151 13855
rect 15669 13821 15703 13855
rect 13829 13685 13863 13719
rect 15301 13685 15335 13719
rect 15853 13685 15887 13719
rect 2237 13345 2271 13379
rect 2329 13277 2363 13311
rect 2513 13277 2547 13311
rect 1869 13141 1903 13175
rect 2237 12937 2271 12971
rect 4537 12937 4571 12971
rect 2789 12801 2823 12835
rect 3893 12801 3927 12835
rect 4997 12801 5031 12835
rect 5181 12801 5215 12835
rect 3617 12733 3651 12767
rect 4905 12733 4939 12767
rect 2605 12665 2639 12699
rect 2697 12597 2731 12631
rect 3249 12597 3283 12631
rect 3709 12597 3743 12631
rect 3709 12393 3743 12427
rect 5825 12393 5859 12427
rect 2596 12325 2630 12359
rect 4690 12325 4724 12359
rect 6346 12325 6380 12359
rect 4445 12257 4479 12291
rect 6101 12257 6135 12291
rect 1869 12189 1903 12223
rect 2329 12189 2363 12223
rect 7481 12053 7515 12087
rect 2237 11849 2271 11883
rect 4905 11849 4939 11883
rect 5365 11849 5399 11883
rect 2789 11713 2823 11747
rect 3525 11713 3559 11747
rect 6009 11713 6043 11747
rect 10425 11713 10459 11747
rect 2605 11645 2639 11679
rect 7849 11645 7883 11679
rect 10241 11645 10275 11679
rect 3770 11577 3804 11611
rect 5825 11577 5859 11611
rect 8585 11577 8619 11611
rect 10149 11577 10183 11611
rect 2697 11509 2731 11543
rect 5733 11509 5767 11543
rect 9781 11509 9815 11543
rect 1685 11305 1719 11339
rect 4629 11305 4663 11339
rect 6101 11305 6135 11339
rect 11897 11305 11931 11339
rect 2053 11169 2087 11203
rect 3065 11169 3099 11203
rect 4997 11169 5031 11203
rect 5089 11169 5123 11203
rect 6009 11169 6043 11203
rect 7012 11169 7046 11203
rect 9689 11169 9723 11203
rect 9956 11169 9990 11203
rect 11989 11169 12023 11203
rect 12808 11169 12842 11203
rect 2145 11101 2179 11135
rect 2329 11101 2363 11135
rect 3157 11101 3191 11135
rect 3341 11101 3375 11135
rect 5273 11101 5307 11135
rect 6193 11101 6227 11135
rect 6745 11101 6779 11135
rect 12173 11101 12207 11135
rect 12357 11101 12391 11135
rect 12541 11101 12575 11135
rect 11069 11033 11103 11067
rect 13921 11033 13955 11067
rect 2697 10965 2731 10999
rect 5641 10965 5675 10999
rect 8125 10965 8159 10999
rect 11529 10965 11563 10999
rect 12449 10965 12483 10999
rect 1409 10761 1443 10795
rect 5365 10761 5399 10795
rect 8861 10761 8895 10795
rect 9413 10761 9447 10795
rect 11805 10761 11839 10795
rect 12633 10761 12667 10795
rect 15393 10761 15427 10795
rect 4353 10693 4387 10727
rect 1869 10625 1903 10659
rect 2053 10625 2087 10659
rect 4997 10625 5031 10659
rect 5825 10625 5859 10659
rect 6009 10625 6043 10659
rect 10057 10625 10091 10659
rect 13093 10625 13127 10659
rect 13277 10625 13311 10659
rect 16497 10625 16531 10659
rect 17417 10625 17451 10659
rect 17601 10625 17635 10659
rect 2421 10557 2455 10591
rect 7481 10557 7515 10591
rect 7748 10557 7782 10591
rect 10425 10557 10459 10591
rect 13001 10557 13035 10591
rect 14013 10557 14047 10591
rect 1777 10489 1811 10523
rect 2688 10489 2722 10523
rect 5733 10489 5767 10523
rect 10692 10489 10726 10523
rect 14280 10489 14314 10523
rect 16313 10489 16347 10523
rect 17325 10489 17359 10523
rect 18061 10489 18095 10523
rect 3801 10421 3835 10455
rect 4721 10421 4755 10455
rect 4813 10421 4847 10455
rect 9781 10421 9815 10455
rect 9873 10421 9907 10455
rect 15945 10421 15979 10455
rect 16405 10421 16439 10455
rect 16957 10421 16991 10455
rect 1961 10217 1995 10251
rect 2421 10217 2455 10251
rect 2973 10217 3007 10251
rect 3433 10217 3467 10251
rect 4077 10217 4111 10251
rect 9689 10217 9723 10251
rect 10057 10217 10091 10251
rect 10149 10217 10183 10251
rect 12357 10217 12391 10251
rect 14933 10217 14967 10251
rect 17049 10217 17083 10251
rect 17509 10217 17543 10251
rect 2329 10149 2363 10183
rect 6101 10149 6135 10183
rect 7818 10149 7852 10183
rect 1409 10081 1443 10115
rect 3341 10081 3375 10115
rect 4445 10081 4479 10115
rect 5273 10081 5307 10115
rect 7573 10081 7607 10115
rect 11069 10081 11103 10115
rect 12725 10081 12759 10115
rect 13553 10081 13587 10115
rect 13820 10081 13854 10115
rect 15393 10081 15427 10115
rect 15660 10081 15694 10115
rect 17417 10081 17451 10115
rect 18061 10081 18095 10115
rect 2605 10013 2639 10047
rect 3617 10013 3651 10047
rect 4537 10013 4571 10047
rect 4629 10013 4663 10047
rect 6193 10013 6227 10047
rect 6285 10013 6319 10047
rect 6745 10013 6779 10047
rect 10333 10013 10367 10047
rect 11161 10013 11195 10047
rect 11345 10013 11379 10047
rect 12817 10013 12851 10047
rect 12909 10013 12943 10047
rect 17601 10013 17635 10047
rect 10701 9945 10735 9979
rect 1593 9877 1627 9911
rect 5089 9877 5123 9911
rect 5733 9877 5767 9911
rect 8953 9877 8987 9911
rect 16773 9877 16807 9911
rect 18245 9877 18279 9911
rect 3341 9673 3375 9707
rect 10609 9673 10643 9707
rect 12909 9673 12943 9707
rect 6837 9605 6871 9639
rect 7849 9605 7883 9639
rect 4445 9537 4479 9571
rect 6285 9537 6319 9571
rect 7389 9537 7423 9571
rect 8401 9537 8435 9571
rect 9413 9537 9447 9571
rect 11069 9537 11103 9571
rect 11253 9537 11287 9571
rect 11621 9537 11655 9571
rect 13553 9537 13587 9571
rect 14933 9537 14967 9571
rect 15853 9537 15887 9571
rect 16865 9537 16899 9571
rect 1409 9469 1443 9503
rect 1961 9469 1995 9503
rect 4905 9469 4939 9503
rect 7205 9469 7239 9503
rect 8217 9469 8251 9503
rect 9229 9469 9263 9503
rect 10977 9469 11011 9503
rect 14657 9469 14691 9503
rect 17417 9469 17451 9503
rect 18061 9469 18095 9503
rect 2228 9401 2262 9435
rect 5181 9401 5215 9435
rect 7297 9401 7331 9435
rect 1593 9333 1627 9367
rect 3893 9333 3927 9367
rect 4261 9333 4295 9367
rect 4353 9333 4387 9367
rect 5733 9333 5767 9367
rect 6101 9333 6135 9367
rect 6193 9333 6227 9367
rect 8309 9333 8343 9367
rect 8861 9333 8895 9367
rect 9321 9333 9355 9367
rect 13277 9333 13311 9367
rect 13369 9333 13403 9367
rect 14289 9333 14323 9367
rect 14749 9333 14783 9367
rect 15301 9333 15335 9367
rect 15669 9333 15703 9367
rect 15761 9333 15795 9367
rect 16313 9333 16347 9367
rect 16681 9333 16715 9367
rect 16773 9333 16807 9367
rect 17601 9333 17635 9367
rect 18245 9333 18279 9367
rect 4905 9129 4939 9163
rect 8585 9129 8619 9163
rect 10149 9129 10183 9163
rect 12909 9129 12943 9163
rect 15761 9129 15795 9163
rect 16129 9129 16163 9163
rect 16773 9129 16807 9163
rect 17141 9129 17175 9163
rect 8953 9061 8987 9095
rect 10057 9061 10091 9095
rect 13277 9061 13311 9095
rect 1593 8993 1627 9027
rect 1860 8993 1894 9027
rect 5273 8993 5307 9027
rect 6837 8993 6871 9027
rect 7104 8993 7138 9027
rect 11244 8993 11278 9027
rect 12817 8993 12851 9027
rect 13369 8993 13403 9027
rect 16221 8993 16255 9027
rect 17877 8993 17911 9027
rect 5365 8925 5399 8959
rect 5457 8925 5491 8959
rect 9045 8925 9079 8959
rect 9229 8925 9263 8959
rect 10241 8925 10275 8959
rect 10977 8925 11011 8959
rect 13553 8925 13587 8959
rect 16405 8925 16439 8959
rect 17233 8925 17267 8959
rect 17325 8925 17359 8959
rect 8217 8857 8251 8891
rect 2973 8789 3007 8823
rect 9689 8789 9723 8823
rect 12357 8789 12391 8823
rect 12633 8789 12667 8823
rect 18061 8789 18095 8823
rect 3525 8585 3559 8619
rect 4997 8585 5031 8619
rect 5457 8585 5491 8619
rect 7389 8585 7423 8619
rect 11713 8585 11747 8619
rect 15853 8585 15887 8619
rect 16773 8585 16807 8619
rect 3249 8449 3283 8483
rect 1685 8381 1719 8415
rect 6469 8517 6503 8551
rect 6009 8449 6043 8483
rect 3617 8381 3651 8415
rect 5825 8381 5859 8415
rect 6653 8381 6687 8415
rect 9781 8517 9815 8551
rect 8125 8449 8159 8483
rect 13461 8449 13495 8483
rect 17325 8449 17359 8483
rect 8493 8381 8527 8415
rect 10333 8381 10367 8415
rect 13277 8381 13311 8415
rect 14473 8381 14507 8415
rect 14740 8381 14774 8415
rect 16164 8381 16198 8415
rect 17141 8381 17175 8415
rect 18061 8381 18095 8415
rect 3525 8313 3559 8347
rect 3884 8313 3918 8347
rect 5917 8313 5951 8347
rect 7389 8313 7423 8347
rect 7849 8313 7883 8347
rect 7941 8313 7975 8347
rect 10578 8313 10612 8347
rect 16267 8313 16301 8347
rect 1869 8245 1903 8279
rect 2605 8245 2639 8279
rect 2973 8245 3007 8279
rect 3065 8245 3099 8279
rect 7481 8245 7515 8279
rect 12909 8245 12943 8279
rect 13369 8245 13403 8279
rect 17233 8245 17267 8279
rect 18245 8245 18279 8279
rect 2053 8041 2087 8075
rect 4537 8041 4571 8075
rect 6929 8041 6963 8075
rect 8033 8041 8067 8075
rect 8125 8041 8159 8075
rect 12357 8041 12391 8075
rect 12909 8041 12943 8075
rect 13277 8041 13311 8075
rect 16681 8041 16715 8075
rect 16957 8041 16991 8075
rect 17325 8041 17359 8075
rect 3065 7973 3099 8007
rect 5816 7973 5850 8007
rect 9934 7973 9968 8007
rect 12265 7973 12299 8007
rect 13369 7973 13403 8007
rect 1961 7905 1995 7939
rect 2973 7905 3007 7939
rect 4905 7905 4939 7939
rect 5549 7905 5583 7939
rect 8953 7905 8987 7939
rect 11529 7905 11563 7939
rect 14289 7905 14323 7939
rect 14381 7905 14415 7939
rect 15557 7905 15591 7939
rect 17417 7905 17451 7939
rect 17969 7905 18003 7939
rect 2237 7837 2271 7871
rect 3249 7837 3283 7871
rect 4997 7837 5031 7871
rect 5181 7837 5215 7871
rect 8217 7837 8251 7871
rect 9045 7837 9079 7871
rect 9229 7837 9263 7871
rect 9689 7837 9723 7871
rect 12541 7837 12575 7871
rect 13461 7837 13495 7871
rect 14473 7837 14507 7871
rect 15301 7837 15335 7871
rect 17509 7837 17543 7871
rect 8585 7769 8619 7803
rect 11345 7769 11379 7803
rect 1593 7701 1627 7735
rect 2605 7701 2639 7735
rect 7665 7701 7699 7735
rect 11069 7701 11103 7735
rect 11897 7701 11931 7735
rect 13921 7701 13955 7735
rect 18153 7701 18187 7735
rect 1777 7497 1811 7531
rect 2145 7497 2179 7531
rect 3617 7497 3651 7531
rect 9689 7497 9723 7531
rect 2697 7361 2731 7395
rect 3157 7361 3191 7395
rect 4261 7361 4295 7395
rect 5181 7361 5215 7395
rect 6193 7361 6227 7395
rect 7757 7361 7791 7395
rect 7941 7361 7975 7395
rect 10977 7361 11011 7395
rect 11805 7361 11839 7395
rect 11897 7361 11931 7395
rect 12909 7361 12943 7395
rect 13001 7361 13035 7395
rect 13737 7361 13771 7395
rect 16129 7361 16163 7395
rect 17141 7361 17175 7395
rect 1593 7293 1627 7327
rect 5089 7293 5123 7327
rect 8309 7293 8343 7327
rect 8565 7293 8599 7327
rect 12817 7293 12851 7327
rect 14004 7293 14038 7327
rect 18061 7293 18095 7327
rect 2513 7225 2547 7259
rect 2605 7225 2639 7259
rect 3985 7225 4019 7259
rect 7665 7225 7699 7259
rect 10701 7225 10735 7259
rect 11713 7225 11747 7259
rect 16865 7225 16899 7259
rect 17509 7225 17543 7259
rect 4077 7157 4111 7191
rect 4629 7157 4663 7191
rect 4997 7157 5031 7191
rect 5641 7157 5675 7191
rect 6009 7157 6043 7191
rect 6101 7157 6135 7191
rect 7297 7157 7331 7191
rect 10333 7157 10367 7191
rect 10793 7157 10827 7191
rect 11345 7157 11379 7191
rect 12449 7157 12483 7191
rect 15117 7157 15151 7191
rect 15485 7157 15519 7191
rect 15853 7157 15887 7191
rect 15945 7157 15979 7191
rect 16497 7157 16531 7191
rect 16957 7157 16991 7191
rect 18245 7157 18279 7191
rect 3525 6953 3559 6987
rect 5457 6953 5491 6987
rect 6285 6953 6319 6987
rect 8033 6953 8067 6987
rect 8401 6953 8435 6987
rect 11621 6953 11655 6987
rect 12449 6953 12483 6987
rect 14565 6953 14599 6987
rect 16681 6953 16715 6987
rect 17325 6953 17359 6987
rect 6653 6885 6687 6919
rect 1685 6817 1719 6851
rect 2237 6817 2271 6851
rect 2789 6817 2823 6851
rect 3249 6817 3283 6851
rect 3341 6817 3375 6851
rect 4333 6817 4367 6851
rect 6745 6817 6779 6851
rect 7297 6817 7331 6851
rect 10508 6817 10542 6851
rect 13461 6817 13495 6851
rect 13553 6817 13587 6851
rect 15568 6817 15602 6851
rect 17969 6817 18003 6851
rect 2973 6681 3007 6715
rect 4077 6749 4111 6783
rect 6837 6749 6871 6783
rect 8493 6749 8527 6783
rect 8585 6749 8619 6783
rect 9045 6749 9079 6783
rect 10241 6749 10275 6783
rect 12541 6749 12575 6783
rect 12633 6749 12667 6783
rect 13645 6749 13679 6783
rect 14657 6749 14691 6783
rect 14841 6749 14875 6783
rect 15301 6749 15335 6783
rect 17417 6749 17451 6783
rect 17509 6749 17543 6783
rect 14197 6681 14231 6715
rect 16957 6681 16991 6715
rect 1869 6613 1903 6647
rect 2421 6613 2455 6647
rect 3249 6613 3283 6647
rect 12081 6613 12115 6647
rect 13093 6613 13127 6647
rect 18153 6613 18187 6647
rect 6837 6409 6871 6443
rect 8033 6409 8067 6443
rect 11345 6409 11379 6443
rect 16129 6409 16163 6443
rect 17601 6409 17635 6443
rect 15485 6341 15519 6375
rect 7389 6273 7423 6307
rect 8493 6273 8527 6307
rect 8585 6273 8619 6307
rect 10885 6273 10919 6307
rect 11805 6273 11839 6307
rect 11897 6273 11931 6307
rect 12541 6273 12575 6307
rect 13185 6273 13219 6307
rect 14105 6273 14139 6307
rect 16773 6273 16807 6307
rect 1685 6205 1719 6239
rect 2421 6205 2455 6239
rect 4077 6205 4111 6239
rect 4721 6205 4755 6239
rect 8401 6205 8435 6239
rect 9137 6205 9171 6239
rect 11713 6205 11747 6239
rect 17417 6205 17451 6239
rect 18061 6205 18095 6239
rect 2688 6137 2722 6171
rect 4966 6137 5000 6171
rect 7205 6137 7239 6171
rect 9404 6137 9438 6171
rect 12633 6137 12667 6171
rect 14350 6137 14384 6171
rect 1869 6069 1903 6103
rect 3801 6069 3835 6103
rect 4261 6069 4295 6103
rect 6101 6069 6135 6103
rect 7297 6069 7331 6103
rect 10517 6069 10551 6103
rect 16497 6069 16531 6103
rect 16589 6069 16623 6103
rect 18245 6069 18279 6103
rect 2421 5865 2455 5899
rect 2973 5865 3007 5899
rect 4445 5865 4479 5899
rect 4537 5865 4571 5899
rect 6009 5865 6043 5899
rect 6561 5865 6595 5899
rect 7481 5865 7515 5899
rect 7573 5865 7607 5899
rect 12541 5865 12575 5899
rect 14289 5865 14323 5899
rect 15669 5865 15703 5899
rect 16681 5865 16715 5899
rect 17049 5865 17083 5899
rect 1409 5729 1443 5763
rect 2329 5729 2363 5763
rect 3341 5729 3375 5763
rect 3893 5729 3927 5763
rect 2605 5661 2639 5695
rect 3433 5661 3467 5695
rect 3617 5661 3651 5695
rect 11428 5797 11462 5831
rect 13154 5797 13188 5831
rect 16037 5797 16071 5831
rect 4905 5729 4939 5763
rect 5917 5729 5951 5763
rect 6745 5729 6779 5763
rect 9689 5729 9723 5763
rect 10057 5729 10091 5763
rect 10425 5729 10459 5763
rect 10768 5729 10802 5763
rect 11161 5729 11195 5763
rect 14657 5729 14691 5763
rect 16129 5729 16163 5763
rect 17141 5729 17175 5763
rect 17877 5729 17911 5763
rect 4445 5661 4479 5695
rect 4997 5661 5031 5695
rect 5181 5661 5215 5695
rect 6101 5661 6135 5695
rect 7757 5661 7791 5695
rect 12909 5661 12943 5695
rect 16313 5661 16347 5695
rect 17233 5661 17267 5695
rect 3893 5593 3927 5627
rect 5549 5593 5583 5627
rect 1593 5525 1627 5559
rect 1961 5525 1995 5559
rect 7113 5525 7147 5559
rect 10839 5525 10873 5559
rect 14841 5525 14875 5559
rect 18061 5525 18095 5559
rect 3065 5321 3099 5355
rect 6469 5321 6503 5355
rect 16681 5321 16715 5355
rect 6929 5253 6963 5287
rect 3709 5185 3743 5219
rect 4721 5185 4755 5219
rect 5089 5185 5123 5219
rect 14841 5185 14875 5219
rect 15669 5185 15703 5219
rect 15761 5185 15795 5219
rect 17233 5185 17267 5219
rect 1869 5117 1903 5151
rect 7297 5117 7331 5151
rect 8309 5117 8343 5151
rect 9965 5117 9999 5151
rect 11805 5117 11839 5151
rect 16256 5117 16290 5151
rect 17049 5117 17083 5151
rect 18061 5117 18095 5151
rect 2145 5049 2179 5083
rect 3433 5049 3467 5083
rect 4537 5049 4571 5083
rect 5356 5049 5390 5083
rect 7665 5049 7699 5083
rect 8576 5049 8610 5083
rect 10210 5049 10244 5083
rect 12541 5049 12575 5083
rect 12633 5049 12667 5083
rect 13553 5049 13587 5083
rect 13921 5049 13955 5083
rect 14013 5049 14047 5083
rect 16359 5049 16393 5083
rect 3525 4981 3559 5015
rect 4077 4981 4111 5015
rect 4445 4981 4479 5015
rect 9689 4981 9723 5015
rect 11345 4981 11379 5015
rect 11989 4981 12023 5015
rect 15209 4981 15243 5015
rect 15577 4981 15611 5015
rect 17141 4981 17175 5015
rect 18245 4981 18279 5015
rect 2421 4777 2455 4811
rect 4537 4777 4571 4811
rect 4997 4777 5031 4811
rect 6193 4777 6227 4811
rect 16681 4777 16715 4811
rect 17049 4777 17083 4811
rect 1685 4641 1719 4675
rect 2145 4641 2179 4675
rect 2237 4641 2271 4675
rect 3065 4641 3099 4675
rect 4905 4641 4939 4675
rect 3249 4573 3283 4607
rect 5181 4573 5215 4607
rect 1869 4437 1903 4471
rect 2145 4437 2179 4471
rect 9321 4709 9355 4743
rect 10324 4709 10358 4743
rect 13093 4709 13127 4743
rect 14013 4709 14047 4743
rect 15485 4709 15519 4743
rect 6285 4641 6319 4675
rect 6552 4641 6586 4675
rect 8953 4641 8987 4675
rect 11713 4641 11747 4675
rect 12357 4641 12391 4675
rect 14657 4641 14691 4675
rect 17877 4641 17911 4675
rect 10057 4573 10091 4607
rect 13001 4573 13035 4607
rect 15393 4573 15427 4607
rect 16221 4573 16255 4607
rect 17141 4573 17175 4607
rect 17233 4573 17267 4607
rect 8585 4505 8619 4539
rect 6193 4437 6227 4471
rect 7665 4437 7699 4471
rect 11437 4437 11471 4471
rect 11897 4437 11931 4471
rect 12541 4437 12575 4471
rect 14841 4437 14875 4471
rect 18061 4437 18095 4471
rect 5457 4233 5491 4267
rect 9137 4233 9171 4267
rect 12633 4165 12667 4199
rect 4077 4097 4111 4131
rect 7757 4097 7791 4131
rect 10057 4097 10091 4131
rect 10793 4097 10827 4131
rect 15117 4097 15151 4131
rect 15669 4097 15703 4131
rect 16589 4097 16623 4131
rect 1593 4029 1627 4063
rect 2329 4029 2363 4063
rect 9413 4029 9447 4063
rect 10425 4029 10459 4063
rect 11069 4029 11103 4063
rect 11437 4029 11471 4063
rect 11805 4029 11839 4063
rect 12265 4029 12299 4063
rect 12449 4029 12483 4063
rect 13093 4029 13127 4063
rect 13645 4029 13679 4063
rect 16992 4029 17026 4063
rect 17417 4029 17451 4063
rect 18061 4029 18095 4063
rect 1869 3961 1903 3995
rect 4344 3961 4378 3995
rect 8024 3961 8058 3995
rect 14289 3961 14323 3995
rect 14381 3961 14415 3995
rect 15761 3961 15795 3995
rect 2513 3893 2547 3927
rect 9597 3893 9631 3927
rect 12081 3893 12115 3927
rect 13277 3893 13311 3927
rect 13829 3893 13863 3927
rect 17095 3893 17129 3927
rect 17601 3893 17635 3927
rect 18245 3893 18279 3927
rect 6653 3689 6687 3723
rect 6837 3689 6871 3723
rect 8309 3689 8343 3723
rect 5540 3621 5574 3655
rect 11060 3621 11094 3655
rect 12265 3621 12299 3655
rect 12633 3621 12667 3655
rect 13553 3621 13587 3655
rect 15439 3621 15473 3655
rect 15853 3621 15887 3655
rect 15945 3621 15979 3655
rect 16865 3621 16899 3655
rect 1685 3553 1719 3587
rect 2237 3553 2271 3587
rect 2789 3553 2823 3587
rect 5273 3553 5307 3587
rect 6837 3553 6871 3587
rect 7185 3553 7219 3587
rect 8953 3553 8987 3587
rect 9781 3553 9815 3587
rect 10149 3553 10183 3587
rect 6929 3485 6963 3519
rect 8585 3485 8619 3519
rect 10793 3485 10827 3519
rect 1869 3417 1903 3451
rect 10333 3417 10367 3451
rect 14105 3553 14139 3587
rect 14473 3553 14507 3587
rect 14657 3553 14691 3587
rect 15336 3553 15370 3587
rect 17141 3553 17175 3587
rect 17877 3553 17911 3587
rect 12541 3485 12575 3519
rect 14013 3485 14047 3519
rect 2421 3349 2455 3383
rect 2973 3349 3007 3383
rect 9045 3349 9079 3383
rect 12173 3349 12207 3383
rect 12265 3349 12299 3383
rect 14473 3417 14507 3451
rect 14841 3417 14875 3451
rect 14013 3349 14047 3383
rect 14289 3349 14323 3383
rect 17325 3349 17359 3383
rect 18061 3349 18095 3383
rect 2421 3077 2455 3111
rect 8125 3077 8159 3111
rect 7573 3009 7607 3043
rect 8677 3009 8711 3043
rect 9689 3009 9723 3043
rect 11713 3009 11747 3043
rect 13001 3009 13035 3043
rect 14013 3009 14047 3043
rect 14381 3009 14415 3043
rect 15853 3009 15887 3043
rect 1685 2941 1719 2975
rect 2237 2941 2271 2975
rect 2973 2941 3007 2975
rect 3709 2941 3743 2975
rect 6320 2941 6354 2975
rect 6929 2941 6963 2975
rect 7297 2941 7331 2975
rect 7941 2941 7975 2975
rect 9965 2941 9999 2975
rect 12484 2941 12518 2975
rect 17417 2941 17451 2975
rect 18061 2941 18095 2975
rect 3249 2873 3283 2907
rect 6423 2873 6457 2907
rect 8769 2873 8803 2907
rect 10701 2873 10735 2907
rect 10793 2873 10827 2907
rect 13093 2873 13127 2907
rect 14473 2873 14507 2907
rect 15393 2873 15427 2907
rect 15945 2873 15979 2907
rect 16865 2873 16899 2907
rect 1869 2805 1903 2839
rect 3893 2805 3927 2839
rect 10149 2805 10183 2839
rect 12587 2805 12621 2839
rect 17601 2805 17635 2839
rect 18245 2805 18279 2839
rect 8125 2601 8159 2635
rect 8861 2601 8895 2635
rect 15071 2601 15105 2635
rect 3341 2533 3375 2567
rect 6285 2533 6319 2567
rect 7665 2533 7699 2567
rect 9965 2533 9999 2567
rect 10885 2533 10919 2567
rect 11345 2533 11379 2567
rect 13185 2533 13219 2567
rect 14105 2533 14139 2567
rect 14749 2533 14783 2567
rect 15669 2533 15703 2567
rect 1593 2465 1627 2499
rect 2329 2465 2363 2499
rect 3065 2465 3099 2499
rect 4077 2465 4111 2499
rect 5616 2465 5650 2499
rect 6009 2465 6043 2499
rect 7297 2465 7331 2499
rect 7941 2465 7975 2499
rect 8493 2465 8527 2499
rect 8861 2465 8895 2499
rect 9045 2465 9079 2499
rect 14381 2465 14415 2499
rect 1777 2397 1811 2431
rect 2513 2397 2547 2431
rect 4261 2397 4295 2431
rect 6929 2397 6963 2431
rect 9873 2397 9907 2431
rect 11253 2397 11287 2431
rect 12081 2397 12115 2431
rect 13093 2397 13127 2431
rect 8677 2329 8711 2363
rect 14968 2465 15002 2499
rect 17141 2465 17175 2499
rect 17693 2465 17727 2499
rect 15577 2397 15611 2431
rect 15853 2397 15887 2431
rect 5687 2261 5721 2295
rect 9229 2261 9263 2295
rect 14565 2261 14599 2295
rect 14749 2261 14783 2295
rect 17325 2261 17359 2295
rect 17877 2261 17911 2295
<< metal1 >>
rect 3602 15240 3608 15292
rect 3660 15280 3666 15292
rect 4338 15280 4344 15292
rect 3660 15252 4344 15280
rect 3660 15240 3666 15252
rect 4338 15240 4344 15252
rect 4396 15240 4402 15292
rect 4062 15172 4068 15224
rect 4120 15212 4126 15224
rect 7282 15212 7288 15224
rect 4120 15184 7288 15212
rect 4120 15172 4126 15184
rect 7282 15172 7288 15184
rect 7340 15172 7346 15224
rect 1104 14714 18860 14736
rect 1104 14662 6912 14714
rect 6964 14662 6976 14714
rect 7028 14662 7040 14714
rect 7092 14662 7104 14714
rect 7156 14662 12843 14714
rect 12895 14662 12907 14714
rect 12959 14662 12971 14714
rect 13023 14662 13035 14714
rect 13087 14662 18860 14714
rect 1104 14640 18860 14662
rect 1578 14560 1584 14612
rect 1636 14600 1642 14612
rect 1949 14603 2007 14609
rect 1949 14600 1961 14603
rect 1636 14572 1961 14600
rect 1636 14560 1642 14572
rect 1949 14569 1961 14572
rect 1995 14569 2007 14603
rect 1949 14563 2007 14569
rect 13906 14532 13912 14544
rect 1780 14504 13912 14532
rect 1780 14473 1808 14504
rect 13906 14492 13912 14504
rect 13964 14532 13970 14544
rect 18322 14532 18328 14544
rect 13964 14504 18328 14532
rect 13964 14492 13970 14504
rect 18322 14492 18328 14504
rect 18380 14492 18386 14544
rect 1765 14467 1823 14473
rect 1765 14433 1777 14467
rect 1811 14433 1823 14467
rect 11054 14464 11060 14476
rect 1765 14427 1823 14433
rect 3620 14436 11060 14464
rect 2590 14356 2596 14408
rect 2648 14396 2654 14408
rect 3620 14396 3648 14436
rect 11054 14424 11060 14436
rect 11112 14424 11118 14476
rect 2648 14368 3648 14396
rect 2648 14356 2654 14368
rect 9950 14356 9956 14408
rect 10008 14396 10014 14408
rect 12434 14396 12440 14408
rect 10008 14368 12440 14396
rect 10008 14356 10014 14368
rect 12434 14356 12440 14368
rect 12492 14356 12498 14408
rect 3326 14288 3332 14340
rect 3384 14328 3390 14340
rect 13998 14328 14004 14340
rect 3384 14300 14004 14328
rect 3384 14288 3390 14300
rect 13998 14288 14004 14300
rect 14056 14288 14062 14340
rect 2774 14220 2780 14272
rect 2832 14260 2838 14272
rect 14182 14260 14188 14272
rect 2832 14232 14188 14260
rect 2832 14220 2838 14232
rect 14182 14220 14188 14232
rect 14240 14220 14246 14272
rect 1104 14170 18860 14192
rect 1104 14118 3947 14170
rect 3999 14118 4011 14170
rect 4063 14118 4075 14170
rect 4127 14118 4139 14170
rect 4191 14118 9878 14170
rect 9930 14118 9942 14170
rect 9994 14118 10006 14170
rect 10058 14118 10070 14170
rect 10122 14118 15808 14170
rect 15860 14118 15872 14170
rect 15924 14118 15936 14170
rect 15988 14118 16000 14170
rect 16052 14118 18860 14170
rect 1104 14096 18860 14118
rect 290 14016 296 14068
rect 348 14056 354 14068
rect 1857 14059 1915 14065
rect 1857 14056 1869 14059
rect 348 14028 1869 14056
rect 348 14016 354 14028
rect 1857 14025 1869 14028
rect 1903 14025 1915 14059
rect 2409 14059 2467 14065
rect 2409 14056 2421 14059
rect 1857 14019 1915 14025
rect 1964 14028 2421 14056
rect 934 13948 940 14000
rect 992 13988 998 14000
rect 1964 13988 1992 14028
rect 2409 14025 2421 14028
rect 2455 14025 2467 14059
rect 2409 14019 2467 14025
rect 2866 14016 2872 14068
rect 2924 14056 2930 14068
rect 3513 14059 3571 14065
rect 3513 14056 3525 14059
rect 2924 14028 3525 14056
rect 2924 14016 2930 14028
rect 3513 14025 3525 14028
rect 3559 14025 3571 14059
rect 3513 14019 3571 14025
rect 6914 14016 6920 14068
rect 6972 14056 6978 14068
rect 7009 14059 7067 14065
rect 7009 14056 7021 14059
rect 6972 14028 7021 14056
rect 6972 14016 6978 14028
rect 7009 14025 7021 14028
rect 7055 14025 7067 14059
rect 7009 14019 7067 14025
rect 992 13960 1992 13988
rect 992 13948 998 13960
rect 2222 13948 2228 14000
rect 2280 13988 2286 14000
rect 2961 13991 3019 13997
rect 2961 13988 2973 13991
rect 2280 13960 2973 13988
rect 2280 13948 2286 13960
rect 2961 13957 2973 13960
rect 3007 13957 3019 13991
rect 2961 13951 3019 13957
rect 6181 13991 6239 13997
rect 6181 13957 6193 13991
rect 6227 13988 6239 13991
rect 6270 13988 6276 14000
rect 6227 13960 6276 13988
rect 6227 13957 6239 13960
rect 6181 13951 6239 13957
rect 6270 13948 6276 13960
rect 6328 13948 6334 14000
rect 13538 13948 13544 14000
rect 13596 13988 13602 14000
rect 14645 13991 14703 13997
rect 14645 13988 14657 13991
rect 13596 13960 14657 13988
rect 13596 13948 13602 13960
rect 14645 13957 14657 13960
rect 14691 13957 14703 13991
rect 14645 13951 14703 13957
rect 15654 13948 15660 14000
rect 15712 13948 15718 14000
rect 10686 13920 10692 13932
rect 1688 13892 10692 13920
rect 1688 13861 1716 13892
rect 10686 13880 10692 13892
rect 10744 13880 10750 13932
rect 15672 13920 15700 13948
rect 16206 13920 16212 13932
rect 15120 13892 16212 13920
rect 1673 13855 1731 13861
rect 1673 13821 1685 13855
rect 1719 13821 1731 13855
rect 1673 13815 1731 13821
rect 2225 13855 2283 13861
rect 2225 13821 2237 13855
rect 2271 13852 2283 13855
rect 2590 13852 2596 13864
rect 2271 13824 2596 13852
rect 2271 13821 2283 13824
rect 2225 13815 2283 13821
rect 2590 13812 2596 13824
rect 2648 13812 2654 13864
rect 2774 13812 2780 13864
rect 2832 13852 2838 13864
rect 3326 13852 3332 13864
rect 2832 13824 2877 13852
rect 3287 13824 3332 13852
rect 2832 13812 2838 13824
rect 3326 13812 3332 13824
rect 3384 13812 3390 13864
rect 5997 13855 6055 13861
rect 5997 13821 6009 13855
rect 6043 13852 6055 13855
rect 6086 13852 6092 13864
rect 6043 13824 6092 13852
rect 6043 13821 6055 13824
rect 5997 13815 6055 13821
rect 6086 13812 6092 13824
rect 6144 13812 6150 13864
rect 6546 13812 6552 13864
rect 6604 13852 6610 13864
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6604 13824 6837 13852
rect 6604 13812 6610 13824
rect 6825 13821 6837 13824
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 13633 13855 13691 13861
rect 13633 13821 13645 13855
rect 13679 13852 13691 13855
rect 14366 13852 14372 13864
rect 13679 13824 14372 13852
rect 13679 13821 13691 13824
rect 13633 13815 13691 13821
rect 14366 13812 14372 13824
rect 14424 13812 14430 13864
rect 14461 13855 14519 13861
rect 14461 13821 14473 13855
rect 14507 13852 14519 13855
rect 15010 13852 15016 13864
rect 14507 13824 15016 13852
rect 14507 13821 14519 13824
rect 14461 13815 14519 13821
rect 15010 13812 15016 13824
rect 15068 13812 15074 13864
rect 15120 13861 15148 13892
rect 16206 13880 16212 13892
rect 16264 13880 16270 13932
rect 15105 13855 15163 13861
rect 15105 13821 15117 13855
rect 15151 13821 15163 13855
rect 15105 13815 15163 13821
rect 15378 13812 15384 13864
rect 15436 13852 15442 13864
rect 15657 13855 15715 13861
rect 15657 13852 15669 13855
rect 15436 13824 15669 13852
rect 15436 13812 15442 13824
rect 15657 13821 15669 13824
rect 15703 13852 15715 13855
rect 16390 13852 16396 13864
rect 15703 13824 16396 13852
rect 15703 13821 15715 13824
rect 15657 13815 15715 13821
rect 16390 13812 16396 13824
rect 16448 13812 16454 13864
rect 7374 13744 7380 13796
rect 7432 13784 7438 13796
rect 9214 13784 9220 13796
rect 7432 13756 9220 13784
rect 7432 13744 7438 13756
rect 9214 13744 9220 13756
rect 9272 13744 9278 13796
rect 14384 13784 14412 13812
rect 14826 13784 14832 13796
rect 14384 13756 14832 13784
rect 14826 13744 14832 13756
rect 14884 13744 14890 13796
rect 3510 13676 3516 13728
rect 3568 13716 3574 13728
rect 13817 13719 13875 13725
rect 13817 13716 13829 13719
rect 3568 13688 13829 13716
rect 3568 13676 3574 13688
rect 13817 13685 13829 13688
rect 13863 13685 13875 13719
rect 15286 13716 15292 13728
rect 15247 13688 15292 13716
rect 13817 13679 13875 13685
rect 15286 13676 15292 13688
rect 15344 13676 15350 13728
rect 15838 13716 15844 13728
rect 15799 13688 15844 13716
rect 15838 13676 15844 13688
rect 15896 13676 15902 13728
rect 1104 13626 18860 13648
rect 1104 13574 6912 13626
rect 6964 13574 6976 13626
rect 7028 13574 7040 13626
rect 7092 13574 7104 13626
rect 7156 13574 12843 13626
rect 12895 13574 12907 13626
rect 12959 13574 12971 13626
rect 13023 13574 13035 13626
rect 13087 13574 18860 13626
rect 1104 13552 18860 13574
rect 4798 13472 4804 13524
rect 4856 13512 4862 13524
rect 15286 13512 15292 13524
rect 4856 13484 15292 13512
rect 4856 13472 4862 13484
rect 15286 13472 15292 13484
rect 15344 13472 15350 13524
rect 4246 13404 4252 13456
rect 4304 13444 4310 13456
rect 13538 13444 13544 13456
rect 4304 13416 13544 13444
rect 4304 13404 4310 13416
rect 13538 13404 13544 13416
rect 13596 13404 13602 13456
rect 14182 13404 14188 13456
rect 14240 13444 14246 13456
rect 18966 13444 18972 13456
rect 14240 13416 18972 13444
rect 14240 13404 14246 13416
rect 18966 13404 18972 13416
rect 19024 13404 19030 13456
rect 2222 13376 2228 13388
rect 2183 13348 2228 13376
rect 2222 13336 2228 13348
rect 2280 13336 2286 13388
rect 5442 13336 5448 13388
rect 5500 13376 5506 13388
rect 15838 13376 15844 13388
rect 5500 13348 15844 13376
rect 5500 13336 5506 13348
rect 15838 13336 15844 13348
rect 15896 13336 15902 13388
rect 2314 13308 2320 13320
rect 2275 13280 2320 13308
rect 2314 13268 2320 13280
rect 2372 13268 2378 13320
rect 2498 13308 2504 13320
rect 2459 13280 2504 13308
rect 2498 13268 2504 13280
rect 2556 13268 2562 13320
rect 10686 13268 10692 13320
rect 10744 13308 10750 13320
rect 17034 13308 17040 13320
rect 10744 13280 17040 13308
rect 10744 13268 10750 13280
rect 17034 13268 17040 13280
rect 17092 13268 17098 13320
rect 3418 13200 3424 13252
rect 3476 13240 3482 13252
rect 10870 13240 10876 13252
rect 3476 13212 10876 13240
rect 3476 13200 3482 13212
rect 10870 13200 10876 13212
rect 10928 13200 10934 13252
rect 11054 13200 11060 13252
rect 11112 13240 11118 13252
rect 12066 13240 12072 13252
rect 11112 13212 12072 13240
rect 11112 13200 11118 13212
rect 12066 13200 12072 13212
rect 12124 13240 12130 13252
rect 12124 13212 13768 13240
rect 12124 13200 12130 13212
rect 1857 13175 1915 13181
rect 1857 13141 1869 13175
rect 1903 13172 1915 13175
rect 3602 13172 3608 13184
rect 1903 13144 3608 13172
rect 1903 13141 1915 13144
rect 1857 13135 1915 13141
rect 3602 13132 3608 13144
rect 3660 13132 3666 13184
rect 13740 13172 13768 13212
rect 13814 13200 13820 13252
rect 13872 13240 13878 13252
rect 15010 13240 15016 13252
rect 13872 13212 15016 13240
rect 13872 13200 13878 13212
rect 15010 13200 15016 13212
rect 15068 13200 15074 13252
rect 17678 13172 17684 13184
rect 13740 13144 17684 13172
rect 17678 13132 17684 13144
rect 17736 13132 17742 13184
rect 1104 13082 18860 13104
rect 1104 13030 3947 13082
rect 3999 13030 4011 13082
rect 4063 13030 4075 13082
rect 4127 13030 4139 13082
rect 4191 13030 9878 13082
rect 9930 13030 9942 13082
rect 9994 13030 10006 13082
rect 10058 13030 10070 13082
rect 10122 13030 15808 13082
rect 15860 13030 15872 13082
rect 15924 13030 15936 13082
rect 15988 13030 16000 13082
rect 16052 13030 18860 13082
rect 1104 13008 18860 13030
rect 2225 12971 2283 12977
rect 2225 12937 2237 12971
rect 2271 12968 2283 12971
rect 2314 12968 2320 12980
rect 2271 12940 2320 12968
rect 2271 12937 2283 12940
rect 2225 12931 2283 12937
rect 2314 12928 2320 12940
rect 2372 12928 2378 12980
rect 4525 12971 4583 12977
rect 4525 12937 4537 12971
rect 4571 12968 4583 12971
rect 5258 12968 5264 12980
rect 4571 12940 5264 12968
rect 4571 12937 4583 12940
rect 4525 12931 4583 12937
rect 5258 12928 5264 12940
rect 5316 12928 5322 12980
rect 13998 12928 14004 12980
rect 14056 12968 14062 12980
rect 19610 12968 19616 12980
rect 14056 12940 19616 12968
rect 14056 12928 14062 12940
rect 19610 12928 19616 12940
rect 19668 12928 19674 12980
rect 3510 12860 3516 12912
rect 3568 12900 3574 12912
rect 6362 12900 6368 12912
rect 3568 12872 6368 12900
rect 3568 12860 3574 12872
rect 6362 12860 6368 12872
rect 6420 12860 6426 12912
rect 2590 12792 2596 12844
rect 2648 12832 2654 12844
rect 2777 12835 2835 12841
rect 2777 12832 2789 12835
rect 2648 12804 2789 12832
rect 2648 12792 2654 12804
rect 2777 12801 2789 12804
rect 2823 12801 2835 12835
rect 2777 12795 2835 12801
rect 3881 12835 3939 12841
rect 3881 12801 3893 12835
rect 3927 12832 3939 12835
rect 4614 12832 4620 12844
rect 3927 12804 4620 12832
rect 3927 12801 3939 12804
rect 3881 12795 3939 12801
rect 4614 12792 4620 12804
rect 4672 12792 4678 12844
rect 4706 12792 4712 12844
rect 4764 12832 4770 12844
rect 4985 12835 5043 12841
rect 4985 12832 4997 12835
rect 4764 12804 4997 12832
rect 4764 12792 4770 12804
rect 4985 12801 4997 12804
rect 5031 12801 5043 12835
rect 4985 12795 5043 12801
rect 5169 12835 5227 12841
rect 5169 12801 5181 12835
rect 5215 12832 5227 12835
rect 7650 12832 7656 12844
rect 5215 12804 7656 12832
rect 5215 12801 5227 12804
rect 5169 12795 5227 12801
rect 7650 12792 7656 12804
rect 7708 12792 7714 12844
rect 13722 12832 13728 12844
rect 7760 12804 13728 12832
rect 3602 12764 3608 12776
rect 3563 12736 3608 12764
rect 3602 12724 3608 12736
rect 3660 12724 3666 12776
rect 4890 12764 4896 12776
rect 4851 12736 4896 12764
rect 4890 12724 4896 12736
rect 4948 12724 4954 12776
rect 2593 12699 2651 12705
rect 2593 12665 2605 12699
rect 2639 12696 2651 12699
rect 3418 12696 3424 12708
rect 2639 12668 3424 12696
rect 2639 12665 2651 12668
rect 2593 12659 2651 12665
rect 3418 12656 3424 12668
rect 3476 12656 3482 12708
rect 7760 12696 7788 12804
rect 13722 12792 13728 12804
rect 13780 12792 13786 12844
rect 15194 12724 15200 12776
rect 15252 12764 15258 12776
rect 15562 12764 15568 12776
rect 15252 12736 15568 12764
rect 15252 12724 15258 12736
rect 15562 12724 15568 12736
rect 15620 12724 15626 12776
rect 4908 12668 7788 12696
rect 2685 12631 2743 12637
rect 2685 12597 2697 12631
rect 2731 12628 2743 12631
rect 2774 12628 2780 12640
rect 2731 12600 2780 12628
rect 2731 12597 2743 12600
rect 2685 12591 2743 12597
rect 2774 12588 2780 12600
rect 2832 12588 2838 12640
rect 3142 12588 3148 12640
rect 3200 12628 3206 12640
rect 3237 12631 3295 12637
rect 3237 12628 3249 12631
rect 3200 12600 3249 12628
rect 3200 12588 3206 12600
rect 3237 12597 3249 12600
rect 3283 12597 3295 12631
rect 3694 12628 3700 12640
rect 3655 12600 3700 12628
rect 3237 12591 3295 12597
rect 3694 12588 3700 12600
rect 3752 12588 3758 12640
rect 4062 12588 4068 12640
rect 4120 12628 4126 12640
rect 4908 12628 4936 12668
rect 10594 12656 10600 12708
rect 10652 12696 10658 12708
rect 14366 12696 14372 12708
rect 10652 12668 14372 12696
rect 10652 12656 10658 12668
rect 14366 12656 14372 12668
rect 14424 12656 14430 12708
rect 4120 12600 4936 12628
rect 4120 12588 4126 12600
rect 1104 12538 18860 12560
rect 1104 12486 6912 12538
rect 6964 12486 6976 12538
rect 7028 12486 7040 12538
rect 7092 12486 7104 12538
rect 7156 12486 12843 12538
rect 12895 12486 12907 12538
rect 12959 12486 12971 12538
rect 13023 12486 13035 12538
rect 13087 12486 18860 12538
rect 1104 12464 18860 12486
rect 2314 12384 2320 12436
rect 2372 12424 2378 12436
rect 2498 12424 2504 12436
rect 2372 12396 2504 12424
rect 2372 12384 2378 12396
rect 2498 12384 2504 12396
rect 2556 12424 2562 12436
rect 3697 12427 3755 12433
rect 3697 12424 3709 12427
rect 2556 12396 3709 12424
rect 2556 12384 2562 12396
rect 3697 12393 3709 12396
rect 3743 12393 3755 12427
rect 3697 12387 3755 12393
rect 5813 12427 5871 12433
rect 5813 12393 5825 12427
rect 5859 12393 5871 12427
rect 5813 12387 5871 12393
rect 2590 12365 2596 12368
rect 2584 12356 2596 12365
rect 2551 12328 2596 12356
rect 2584 12319 2596 12328
rect 2590 12316 2596 12319
rect 2648 12316 2654 12368
rect 2682 12316 2688 12368
rect 2740 12356 2746 12368
rect 2740 12328 4476 12356
rect 2740 12316 2746 12328
rect 3602 12248 3608 12300
rect 3660 12288 3666 12300
rect 3786 12288 3792 12300
rect 3660 12260 3792 12288
rect 3660 12248 3666 12260
rect 3786 12248 3792 12260
rect 3844 12248 3850 12300
rect 4448 12297 4476 12328
rect 4614 12316 4620 12368
rect 4672 12365 4678 12368
rect 4672 12359 4736 12365
rect 4672 12325 4690 12359
rect 4724 12325 4736 12359
rect 5828 12356 5856 12387
rect 15562 12384 15568 12436
rect 15620 12384 15626 12436
rect 6178 12356 6184 12368
rect 5828 12328 6184 12356
rect 4672 12319 4736 12325
rect 4672 12316 4678 12319
rect 6178 12316 6184 12328
rect 6236 12356 6242 12368
rect 6334 12359 6392 12365
rect 6334 12356 6346 12359
rect 6236 12328 6346 12356
rect 6236 12316 6242 12328
rect 6334 12325 6346 12328
rect 6380 12325 6392 12359
rect 6334 12319 6392 12325
rect 15378 12316 15384 12368
rect 15436 12356 15442 12368
rect 15580 12356 15608 12384
rect 15436 12328 15608 12356
rect 15436 12316 15442 12328
rect 4433 12291 4491 12297
rect 4433 12257 4445 12291
rect 4479 12288 4491 12291
rect 6089 12291 6147 12297
rect 6089 12288 6101 12291
rect 4479 12260 6101 12288
rect 4479 12257 4491 12260
rect 4433 12251 4491 12257
rect 6089 12257 6101 12260
rect 6135 12257 6147 12291
rect 6089 12251 6147 12257
rect 6196 12260 7880 12288
rect 1854 12220 1860 12232
rect 1815 12192 1860 12220
rect 1854 12180 1860 12192
rect 1912 12180 1918 12232
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12189 2375 12223
rect 2317 12183 2375 12189
rect 2332 12084 2360 12183
rect 5442 12180 5448 12232
rect 5500 12220 5506 12232
rect 6196 12220 6224 12260
rect 5500 12192 6224 12220
rect 5500 12180 5506 12192
rect 7742 12152 7748 12164
rect 7300 12124 7748 12152
rect 2682 12084 2688 12096
rect 2332 12056 2688 12084
rect 2682 12044 2688 12056
rect 2740 12044 2746 12096
rect 3786 12044 3792 12096
rect 3844 12084 3850 12096
rect 7300 12084 7328 12124
rect 7742 12112 7748 12124
rect 7800 12112 7806 12164
rect 7852 12152 7880 12260
rect 13170 12248 13176 12300
rect 13228 12288 13234 12300
rect 14550 12288 14556 12300
rect 13228 12260 14556 12288
rect 13228 12248 13234 12260
rect 14550 12248 14556 12260
rect 14608 12248 14614 12300
rect 12158 12180 12164 12232
rect 12216 12220 12222 12232
rect 16390 12220 16396 12232
rect 12216 12192 16396 12220
rect 12216 12180 12222 12192
rect 16390 12180 16396 12192
rect 16448 12180 16454 12232
rect 16574 12152 16580 12164
rect 7852 12124 16580 12152
rect 16574 12112 16580 12124
rect 16632 12112 16638 12164
rect 3844 12056 7328 12084
rect 3844 12044 3850 12056
rect 7374 12044 7380 12096
rect 7432 12084 7438 12096
rect 7469 12087 7527 12093
rect 7469 12084 7481 12087
rect 7432 12056 7481 12084
rect 7432 12044 7438 12056
rect 7469 12053 7481 12056
rect 7515 12053 7527 12087
rect 7469 12047 7527 12053
rect 10594 12044 10600 12096
rect 10652 12084 10658 12096
rect 16482 12084 16488 12096
rect 10652 12056 16488 12084
rect 10652 12044 10658 12056
rect 16482 12044 16488 12056
rect 16540 12044 16546 12096
rect 1104 11994 18860 12016
rect 1104 11942 3947 11994
rect 3999 11942 4011 11994
rect 4063 11942 4075 11994
rect 4127 11942 4139 11994
rect 4191 11942 9878 11994
rect 9930 11942 9942 11994
rect 9994 11942 10006 11994
rect 10058 11942 10070 11994
rect 10122 11942 15808 11994
rect 15860 11942 15872 11994
rect 15924 11942 15936 11994
rect 15988 11942 16000 11994
rect 16052 11942 18860 11994
rect 1104 11920 18860 11942
rect 2222 11880 2228 11892
rect 2183 11852 2228 11880
rect 2222 11840 2228 11852
rect 2280 11840 2286 11892
rect 3786 11840 3792 11892
rect 3844 11880 3850 11892
rect 3844 11852 4476 11880
rect 3844 11840 3850 11852
rect 2590 11772 2596 11824
rect 2648 11772 2654 11824
rect 2682 11772 2688 11824
rect 2740 11812 2746 11824
rect 4448 11812 4476 11852
rect 4614 11840 4620 11892
rect 4672 11880 4678 11892
rect 4893 11883 4951 11889
rect 4893 11880 4905 11883
rect 4672 11852 4905 11880
rect 4672 11840 4678 11852
rect 4893 11849 4905 11852
rect 4939 11849 4951 11883
rect 4893 11843 4951 11849
rect 4982 11840 4988 11892
rect 5040 11880 5046 11892
rect 5353 11883 5411 11889
rect 5353 11880 5365 11883
rect 5040 11852 5365 11880
rect 5040 11840 5046 11852
rect 5353 11849 5365 11852
rect 5399 11849 5411 11883
rect 5353 11843 5411 11849
rect 5810 11840 5816 11892
rect 5868 11880 5874 11892
rect 17770 11880 17776 11892
rect 5868 11852 17776 11880
rect 5868 11840 5874 11852
rect 17770 11840 17776 11852
rect 17828 11840 17834 11892
rect 6086 11812 6092 11824
rect 2740 11784 3556 11812
rect 4448 11784 6092 11812
rect 2740 11772 2746 11784
rect 2608 11744 2636 11772
rect 3528 11753 3556 11784
rect 6086 11772 6092 11784
rect 6144 11812 6150 11824
rect 17310 11812 17316 11824
rect 6144 11784 17316 11812
rect 6144 11772 6150 11784
rect 17310 11772 17316 11784
rect 17368 11772 17374 11824
rect 2777 11747 2835 11753
rect 2777 11744 2789 11747
rect 2608 11716 2789 11744
rect 2777 11713 2789 11716
rect 2823 11713 2835 11747
rect 2777 11707 2835 11713
rect 3513 11747 3571 11753
rect 3513 11713 3525 11747
rect 3559 11713 3571 11747
rect 3513 11707 3571 11713
rect 5258 11704 5264 11756
rect 5316 11744 5322 11756
rect 5997 11747 6055 11753
rect 5997 11744 6009 11747
rect 5316 11716 6009 11744
rect 5316 11704 5322 11716
rect 5997 11713 6009 11716
rect 6043 11744 6055 11747
rect 8110 11744 8116 11756
rect 6043 11716 8116 11744
rect 6043 11713 6055 11716
rect 5997 11707 6055 11713
rect 8110 11704 8116 11716
rect 8168 11704 8174 11756
rect 10318 11744 10324 11756
rect 8404 11716 10324 11744
rect 1854 11636 1860 11688
rect 1912 11676 1918 11688
rect 2593 11679 2651 11685
rect 2593 11676 2605 11679
rect 1912 11648 2605 11676
rect 1912 11636 1918 11648
rect 2593 11645 2605 11648
rect 2639 11645 2651 11679
rect 2593 11639 2651 11645
rect 3050 11636 3056 11688
rect 3108 11676 3114 11688
rect 5350 11676 5356 11688
rect 3108 11648 5356 11676
rect 3108 11636 3114 11648
rect 5350 11636 5356 11648
rect 5408 11636 5414 11688
rect 5460 11648 7788 11676
rect 2314 11568 2320 11620
rect 2372 11608 2378 11620
rect 3758 11611 3816 11617
rect 3758 11608 3770 11611
rect 2372 11580 3770 11608
rect 2372 11568 2378 11580
rect 3758 11577 3770 11580
rect 3804 11577 3816 11611
rect 3758 11571 3816 11577
rect 1762 11500 1768 11552
rect 1820 11540 1826 11552
rect 2685 11543 2743 11549
rect 2685 11540 2697 11543
rect 1820 11512 2697 11540
rect 1820 11500 1826 11512
rect 2685 11509 2697 11512
rect 2731 11540 2743 11543
rect 5460 11540 5488 11648
rect 5534 11568 5540 11620
rect 5592 11608 5598 11620
rect 5813 11611 5871 11617
rect 5813 11608 5825 11611
rect 5592 11580 5825 11608
rect 5592 11568 5598 11580
rect 5813 11577 5825 11580
rect 5859 11577 5871 11611
rect 7760 11608 7788 11648
rect 7834 11636 7840 11688
rect 7892 11676 7898 11688
rect 7892 11648 7937 11676
rect 7892 11636 7898 11648
rect 8404 11608 8432 11716
rect 10318 11704 10324 11716
rect 10376 11704 10382 11756
rect 10413 11747 10471 11753
rect 10413 11713 10425 11747
rect 10459 11744 10471 11747
rect 10962 11744 10968 11756
rect 10459 11716 10968 11744
rect 10459 11713 10471 11716
rect 10413 11707 10471 11713
rect 10962 11704 10968 11716
rect 11020 11704 11026 11756
rect 9674 11636 9680 11688
rect 9732 11676 9738 11688
rect 10229 11679 10287 11685
rect 10229 11676 10241 11679
rect 9732 11648 10241 11676
rect 9732 11636 9738 11648
rect 10229 11645 10241 11648
rect 10275 11645 10287 11679
rect 10336 11676 10364 11704
rect 11146 11676 11152 11688
rect 10336 11648 11152 11676
rect 10229 11639 10287 11645
rect 11146 11636 11152 11648
rect 11204 11636 11210 11688
rect 7760 11580 8432 11608
rect 8573 11611 8631 11617
rect 5813 11571 5871 11577
rect 8573 11577 8585 11611
rect 8619 11608 8631 11611
rect 9030 11608 9036 11620
rect 8619 11580 9036 11608
rect 8619 11577 8631 11580
rect 8573 11571 8631 11577
rect 9030 11568 9036 11580
rect 9088 11568 9094 11620
rect 9398 11568 9404 11620
rect 9456 11608 9462 11620
rect 10137 11611 10195 11617
rect 10137 11608 10149 11611
rect 9456 11580 10149 11608
rect 9456 11568 9462 11580
rect 10137 11577 10149 11580
rect 10183 11577 10195 11611
rect 10137 11571 10195 11577
rect 10778 11568 10784 11620
rect 10836 11608 10842 11620
rect 15470 11608 15476 11620
rect 10836 11580 15476 11608
rect 10836 11568 10842 11580
rect 15470 11568 15476 11580
rect 15528 11568 15534 11620
rect 2731 11512 5488 11540
rect 5721 11543 5779 11549
rect 2731 11509 2743 11512
rect 2685 11503 2743 11509
rect 5721 11509 5733 11543
rect 5767 11540 5779 11543
rect 7834 11540 7840 11552
rect 5767 11512 7840 11540
rect 5767 11509 5779 11512
rect 5721 11503 5779 11509
rect 7834 11500 7840 11512
rect 7892 11500 7898 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 9769 11543 9827 11549
rect 9769 11540 9781 11543
rect 8352 11512 9781 11540
rect 8352 11500 8358 11512
rect 9769 11509 9781 11512
rect 9815 11509 9827 11543
rect 9769 11503 9827 11509
rect 12526 11500 12532 11552
rect 12584 11540 12590 11552
rect 13170 11540 13176 11552
rect 12584 11512 13176 11540
rect 12584 11500 12590 11512
rect 13170 11500 13176 11512
rect 13228 11500 13234 11552
rect 1104 11450 18860 11472
rect 1104 11398 6912 11450
rect 6964 11398 6976 11450
rect 7028 11398 7040 11450
rect 7092 11398 7104 11450
rect 7156 11398 12843 11450
rect 12895 11398 12907 11450
rect 12959 11398 12971 11450
rect 13023 11398 13035 11450
rect 13087 11398 18860 11450
rect 1104 11376 18860 11398
rect 1673 11339 1731 11345
rect 1673 11305 1685 11339
rect 1719 11336 1731 11339
rect 3694 11336 3700 11348
rect 1719 11308 3700 11336
rect 1719 11305 1731 11308
rect 1673 11299 1731 11305
rect 3694 11296 3700 11308
rect 3752 11296 3758 11348
rect 4617 11339 4675 11345
rect 4617 11305 4629 11339
rect 4663 11336 4675 11339
rect 5074 11336 5080 11348
rect 4663 11308 5080 11336
rect 4663 11305 4675 11308
rect 4617 11299 4675 11305
rect 5074 11296 5080 11308
rect 5132 11296 5138 11348
rect 6086 11336 6092 11348
rect 6047 11308 6092 11336
rect 6086 11296 6092 11308
rect 6144 11296 6150 11348
rect 10778 11336 10784 11348
rect 6196 11308 10784 11336
rect 2406 11228 2412 11280
rect 2464 11268 2470 11280
rect 2682 11268 2688 11280
rect 2464 11240 2688 11268
rect 2464 11228 2470 11240
rect 2682 11228 2688 11240
rect 2740 11228 2746 11280
rect 2774 11228 2780 11280
rect 2832 11268 2838 11280
rect 6196 11268 6224 11308
rect 10778 11296 10784 11308
rect 10836 11296 10842 11348
rect 11885 11339 11943 11345
rect 11885 11305 11897 11339
rect 11931 11336 11943 11339
rect 11931 11308 13400 11336
rect 11931 11305 11943 11308
rect 11885 11299 11943 11305
rect 2832 11240 6224 11268
rect 2832 11228 2838 11240
rect 6730 11228 6736 11280
rect 6788 11268 6794 11280
rect 11900 11268 11928 11299
rect 6788 11240 11928 11268
rect 6788 11228 6794 11240
rect 2038 11200 2044 11212
rect 1999 11172 2044 11200
rect 2038 11160 2044 11172
rect 2096 11160 2102 11212
rect 3050 11200 3056 11212
rect 3011 11172 3056 11200
rect 3050 11160 3056 11172
rect 3108 11160 3114 11212
rect 4982 11200 4988 11212
rect 4943 11172 4988 11200
rect 4982 11160 4988 11172
rect 5040 11160 5046 11212
rect 5077 11203 5135 11209
rect 5077 11169 5089 11203
rect 5123 11200 5135 11203
rect 5902 11200 5908 11212
rect 5123 11172 5908 11200
rect 5123 11169 5135 11172
rect 5077 11163 5135 11169
rect 5902 11160 5908 11172
rect 5960 11160 5966 11212
rect 5997 11203 6055 11209
rect 5997 11169 6009 11203
rect 6043 11169 6055 11203
rect 5997 11163 6055 11169
rect 7000 11203 7058 11209
rect 7000 11169 7012 11203
rect 7046 11200 7058 11203
rect 7374 11200 7380 11212
rect 7046 11172 7380 11200
rect 7046 11169 7058 11172
rect 7000 11163 7058 11169
rect 2130 11132 2136 11144
rect 2091 11104 2136 11132
rect 2130 11092 2136 11104
rect 2188 11092 2194 11144
rect 2314 11132 2320 11144
rect 2275 11104 2320 11132
rect 2314 11092 2320 11104
rect 2372 11092 2378 11144
rect 2498 11092 2504 11144
rect 2556 11132 2562 11144
rect 2556 11104 2912 11132
rect 2556 11092 2562 11104
rect 1670 11024 1676 11076
rect 1728 11064 1734 11076
rect 2774 11064 2780 11076
rect 1728 11036 2780 11064
rect 1728 11024 1734 11036
rect 2774 11024 2780 11036
rect 2832 11024 2838 11076
rect 2884 11064 2912 11104
rect 2958 11092 2964 11144
rect 3016 11132 3022 11144
rect 3145 11135 3203 11141
rect 3145 11132 3157 11135
rect 3016 11104 3157 11132
rect 3016 11092 3022 11104
rect 3145 11101 3157 11104
rect 3191 11101 3203 11135
rect 3145 11095 3203 11101
rect 3329 11135 3387 11141
rect 3329 11101 3341 11135
rect 3375 11132 3387 11135
rect 3418 11132 3424 11144
rect 3375 11104 3424 11132
rect 3375 11101 3387 11104
rect 3329 11095 3387 11101
rect 3418 11092 3424 11104
rect 3476 11092 3482 11144
rect 5258 11132 5264 11144
rect 5219 11104 5264 11132
rect 5258 11092 5264 11104
rect 5316 11092 5322 11144
rect 5810 11092 5816 11144
rect 5868 11132 5874 11144
rect 6012 11132 6040 11163
rect 7374 11160 7380 11172
rect 7432 11160 7438 11212
rect 9677 11203 9735 11209
rect 9677 11169 9689 11203
rect 9723 11200 9735 11203
rect 9766 11200 9772 11212
rect 9723 11172 9772 11200
rect 9723 11169 9735 11172
rect 9677 11163 9735 11169
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 9944 11203 10002 11209
rect 9944 11169 9956 11203
rect 9990 11200 10002 11203
rect 10318 11200 10324 11212
rect 9990 11172 10324 11200
rect 9990 11169 10002 11172
rect 9944 11163 10002 11169
rect 10318 11160 10324 11172
rect 10376 11160 10382 11212
rect 11977 11203 12035 11209
rect 11977 11169 11989 11203
rect 12023 11200 12035 11203
rect 12618 11200 12624 11212
rect 12023 11172 12624 11200
rect 12023 11169 12035 11172
rect 11977 11163 12035 11169
rect 12618 11160 12624 11172
rect 12676 11160 12682 11212
rect 12796 11203 12854 11209
rect 12796 11169 12808 11203
rect 12842 11200 12854 11203
rect 13262 11200 13268 11212
rect 12842 11172 13268 11200
rect 12842 11169 12854 11172
rect 12796 11163 12854 11169
rect 13262 11160 13268 11172
rect 13320 11160 13326 11212
rect 13372 11200 13400 11308
rect 18046 11200 18052 11212
rect 13372 11172 18052 11200
rect 18046 11160 18052 11172
rect 18104 11160 18110 11212
rect 5868 11104 6040 11132
rect 5868 11092 5874 11104
rect 6178 11092 6184 11144
rect 6236 11132 6242 11144
rect 6236 11104 6281 11132
rect 6236 11092 6242 11104
rect 6638 11092 6644 11144
rect 6696 11132 6702 11144
rect 6733 11135 6791 11141
rect 6733 11132 6745 11135
rect 6696 11104 6745 11132
rect 6696 11092 6702 11104
rect 6733 11101 6745 11104
rect 6779 11101 6791 11135
rect 6733 11095 6791 11101
rect 12161 11135 12219 11141
rect 12161 11101 12173 11135
rect 12207 11132 12219 11135
rect 12342 11132 12348 11144
rect 12207 11104 12348 11132
rect 12207 11101 12219 11104
rect 12161 11095 12219 11101
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 12434 11092 12440 11144
rect 12492 11132 12498 11144
rect 12529 11135 12587 11141
rect 12529 11132 12541 11135
rect 12492 11104 12541 11132
rect 12492 11092 12498 11104
rect 12529 11101 12541 11104
rect 12575 11101 12587 11135
rect 12529 11095 12587 11101
rect 15194 11092 15200 11144
rect 15252 11132 15258 11144
rect 15470 11132 15476 11144
rect 15252 11104 15476 11132
rect 15252 11092 15258 11104
rect 15470 11092 15476 11104
rect 15528 11092 15534 11144
rect 5442 11064 5448 11076
rect 2884 11036 5448 11064
rect 5442 11024 5448 11036
rect 5500 11024 5506 11076
rect 10962 11024 10968 11076
rect 11020 11064 11026 11076
rect 11057 11067 11115 11073
rect 11057 11064 11069 11067
rect 11020 11036 11069 11064
rect 11020 11024 11026 11036
rect 11057 11033 11069 11036
rect 11103 11033 11115 11067
rect 13909 11067 13967 11073
rect 13909 11064 13921 11067
rect 11057 11027 11115 11033
rect 11348 11036 11652 11064
rect 1854 10956 1860 11008
rect 1912 10996 1918 11008
rect 2685 10999 2743 11005
rect 2685 10996 2697 10999
rect 1912 10968 2697 10996
rect 1912 10956 1918 10968
rect 2685 10965 2697 10968
rect 2731 10965 2743 10999
rect 5626 10996 5632 11008
rect 5587 10968 5632 10996
rect 2685 10959 2743 10965
rect 5626 10956 5632 10968
rect 5684 10956 5690 11008
rect 8110 10996 8116 11008
rect 8071 10968 8116 10996
rect 8110 10956 8116 10968
rect 8168 10956 8174 11008
rect 8202 10956 8208 11008
rect 8260 10996 8266 11008
rect 11348 10996 11376 11036
rect 11514 10996 11520 11008
rect 8260 10968 11376 10996
rect 11475 10968 11520 10996
rect 8260 10956 8266 10968
rect 11514 10956 11520 10968
rect 11572 10956 11578 11008
rect 11624 10996 11652 11036
rect 13464 11036 13921 11064
rect 12158 10996 12164 11008
rect 11624 10968 12164 10996
rect 12158 10956 12164 10968
rect 12216 10956 12222 11008
rect 12437 10999 12495 11005
rect 12437 10965 12449 10999
rect 12483 10996 12495 10999
rect 13464 10996 13492 11036
rect 13909 11033 13921 11036
rect 13955 11033 13967 11067
rect 13909 11027 13967 11033
rect 14200 11036 15700 11064
rect 12483 10968 13492 10996
rect 12483 10965 12495 10968
rect 12437 10959 12495 10965
rect 13630 10956 13636 11008
rect 13688 10996 13694 11008
rect 14200 10996 14228 11036
rect 13688 10968 14228 10996
rect 13688 10956 13694 10968
rect 14274 10956 14280 11008
rect 14332 10996 14338 11008
rect 15562 10996 15568 11008
rect 14332 10968 15568 10996
rect 14332 10956 14338 10968
rect 15562 10956 15568 10968
rect 15620 10956 15626 11008
rect 15672 10996 15700 11036
rect 17862 10996 17868 11008
rect 15672 10968 17868 10996
rect 17862 10956 17868 10968
rect 17920 10956 17926 11008
rect 1104 10906 18860 10928
rect 1104 10854 3947 10906
rect 3999 10854 4011 10906
rect 4063 10854 4075 10906
rect 4127 10854 4139 10906
rect 4191 10854 9878 10906
rect 9930 10854 9942 10906
rect 9994 10854 10006 10906
rect 10058 10854 10070 10906
rect 10122 10854 15808 10906
rect 15860 10854 15872 10906
rect 15924 10854 15936 10906
rect 15988 10854 16000 10906
rect 16052 10854 18860 10906
rect 1104 10832 18860 10854
rect 1397 10795 1455 10801
rect 1397 10761 1409 10795
rect 1443 10792 1455 10795
rect 2038 10792 2044 10804
rect 1443 10764 2044 10792
rect 1443 10761 1455 10764
rect 1397 10755 1455 10761
rect 2038 10752 2044 10764
rect 2096 10752 2102 10804
rect 4982 10752 4988 10804
rect 5040 10792 5046 10804
rect 5353 10795 5411 10801
rect 5353 10792 5365 10795
rect 5040 10764 5365 10792
rect 5040 10752 5046 10764
rect 5353 10761 5365 10764
rect 5399 10761 5411 10795
rect 5353 10755 5411 10761
rect 7650 10752 7656 10804
rect 7708 10792 7714 10804
rect 8849 10795 8907 10801
rect 8849 10792 8861 10795
rect 7708 10764 8861 10792
rect 7708 10752 7714 10764
rect 8849 10761 8861 10764
rect 8895 10761 8907 10795
rect 9398 10792 9404 10804
rect 9359 10764 9404 10792
rect 8849 10755 8907 10761
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 11793 10795 11851 10801
rect 11793 10792 11805 10795
rect 10428 10764 11805 10792
rect 4341 10727 4399 10733
rect 4341 10693 4353 10727
rect 4387 10724 4399 10727
rect 5534 10724 5540 10736
rect 4387 10696 5540 10724
rect 4387 10693 4399 10696
rect 4341 10687 4399 10693
rect 5534 10684 5540 10696
rect 5592 10684 5598 10736
rect 1854 10656 1860 10668
rect 1815 10628 1860 10656
rect 1854 10616 1860 10628
rect 1912 10616 1918 10668
rect 2038 10656 2044 10668
rect 1999 10628 2044 10656
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 4985 10659 5043 10665
rect 4985 10625 4997 10659
rect 5031 10625 5043 10659
rect 4985 10619 5043 10625
rect 2406 10588 2412 10600
rect 2367 10560 2412 10588
rect 2406 10548 2412 10560
rect 2464 10548 2470 10600
rect 2608 10560 3556 10588
rect 1578 10480 1584 10532
rect 1636 10520 1642 10532
rect 1765 10523 1823 10529
rect 1765 10520 1777 10523
rect 1636 10492 1777 10520
rect 1636 10480 1642 10492
rect 1765 10489 1777 10492
rect 1811 10520 1823 10523
rect 2608 10520 2636 10560
rect 2682 10529 2688 10532
rect 1811 10492 2636 10520
rect 1811 10489 1823 10492
rect 1765 10483 1823 10489
rect 2676 10483 2688 10529
rect 2740 10520 2746 10532
rect 3418 10520 3424 10532
rect 2740 10492 3424 10520
rect 2682 10480 2688 10483
rect 2740 10480 2746 10492
rect 3418 10480 3424 10492
rect 3476 10480 3482 10532
rect 3528 10520 3556 10560
rect 3602 10548 3608 10600
rect 3660 10588 3666 10600
rect 4798 10588 4804 10600
rect 3660 10560 4804 10588
rect 3660 10548 3666 10560
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 5000 10588 5028 10619
rect 5626 10616 5632 10668
rect 5684 10656 5690 10668
rect 5813 10659 5871 10665
rect 5813 10656 5825 10659
rect 5684 10628 5825 10656
rect 5684 10616 5690 10628
rect 5813 10625 5825 10628
rect 5859 10625 5871 10659
rect 5813 10619 5871 10625
rect 5997 10659 6055 10665
rect 5997 10625 6009 10659
rect 6043 10656 6055 10659
rect 7374 10656 7380 10668
rect 6043 10628 7380 10656
rect 6043 10625 6055 10628
rect 5997 10619 6055 10625
rect 6012 10588 6040 10619
rect 7374 10616 7380 10628
rect 7432 10616 7438 10668
rect 10045 10659 10103 10665
rect 10045 10625 10057 10659
rect 10091 10656 10103 10659
rect 10318 10656 10324 10668
rect 10091 10628 10324 10656
rect 10091 10625 10103 10628
rect 10045 10619 10103 10625
rect 10318 10616 10324 10628
rect 10376 10656 10382 10668
rect 10428 10656 10456 10764
rect 11793 10761 11805 10764
rect 11839 10761 11851 10795
rect 12618 10792 12624 10804
rect 12579 10764 12624 10792
rect 11793 10755 11851 10761
rect 12618 10752 12624 10764
rect 12676 10752 12682 10804
rect 15381 10795 15439 10801
rect 15381 10792 15393 10795
rect 13740 10764 15393 10792
rect 11422 10684 11428 10736
rect 11480 10724 11486 10736
rect 13630 10724 13636 10736
rect 11480 10696 13636 10724
rect 11480 10684 11486 10696
rect 13096 10665 13124 10696
rect 13630 10684 13636 10696
rect 13688 10684 13694 10736
rect 10376 10628 10456 10656
rect 13081 10659 13139 10665
rect 10376 10616 10382 10628
rect 13081 10625 13093 10659
rect 13127 10625 13139 10659
rect 13262 10656 13268 10668
rect 13175 10628 13268 10656
rect 13081 10619 13139 10625
rect 13262 10616 13268 10628
rect 13320 10656 13326 10668
rect 13538 10656 13544 10668
rect 13320 10628 13544 10656
rect 13320 10616 13326 10628
rect 13538 10616 13544 10628
rect 13596 10656 13602 10668
rect 13740 10656 13768 10764
rect 15381 10761 15393 10764
rect 15427 10761 15439 10795
rect 15381 10755 15439 10761
rect 15654 10684 15660 10736
rect 15712 10724 15718 10736
rect 15712 10696 17448 10724
rect 15712 10684 15718 10696
rect 16482 10656 16488 10668
rect 13596 10628 13768 10656
rect 16443 10628 16488 10656
rect 13596 10616 13602 10628
rect 16482 10616 16488 10628
rect 16540 10616 16546 10668
rect 17420 10665 17448 10696
rect 17405 10659 17463 10665
rect 17405 10625 17417 10659
rect 17451 10625 17463 10659
rect 17586 10656 17592 10668
rect 17547 10628 17592 10656
rect 17405 10619 17463 10625
rect 17586 10616 17592 10628
rect 17644 10616 17650 10668
rect 5000 10560 6040 10588
rect 6638 10548 6644 10600
rect 6696 10588 6702 10600
rect 7469 10591 7527 10597
rect 7469 10588 7481 10591
rect 6696 10560 7481 10588
rect 6696 10548 6702 10560
rect 7469 10557 7481 10560
rect 7515 10557 7527 10591
rect 7469 10551 7527 10557
rect 7736 10591 7794 10597
rect 7736 10557 7748 10591
rect 7782 10588 7794 10591
rect 8110 10588 8116 10600
rect 7782 10560 8116 10588
rect 7782 10557 7794 10560
rect 7736 10551 7794 10557
rect 8110 10548 8116 10560
rect 8168 10548 8174 10600
rect 9766 10548 9772 10600
rect 9824 10588 9830 10600
rect 10410 10588 10416 10600
rect 9824 10560 10416 10588
rect 9824 10548 9830 10560
rect 10410 10548 10416 10560
rect 10468 10588 10474 10600
rect 12434 10588 12440 10600
rect 10468 10560 12440 10588
rect 10468 10548 10474 10560
rect 12434 10548 12440 10560
rect 12492 10548 12498 10600
rect 12989 10591 13047 10597
rect 12989 10557 13001 10591
rect 13035 10588 13047 10591
rect 13446 10588 13452 10600
rect 13035 10560 13452 10588
rect 13035 10557 13047 10560
rect 12989 10551 13047 10557
rect 13446 10548 13452 10560
rect 13504 10548 13510 10600
rect 13630 10548 13636 10600
rect 13688 10588 13694 10600
rect 14001 10591 14059 10597
rect 14001 10588 14013 10591
rect 13688 10560 14013 10588
rect 13688 10548 13694 10560
rect 14001 10557 14013 10560
rect 14047 10557 14059 10591
rect 18506 10588 18512 10600
rect 14001 10551 14059 10557
rect 14108 10560 18512 10588
rect 3528 10492 5028 10520
rect 2038 10412 2044 10464
rect 2096 10452 2102 10464
rect 2590 10452 2596 10464
rect 2096 10424 2596 10452
rect 2096 10412 2102 10424
rect 2590 10412 2596 10424
rect 2648 10452 2654 10464
rect 3789 10455 3847 10461
rect 3789 10452 3801 10455
rect 2648 10424 3801 10452
rect 2648 10412 2654 10424
rect 3789 10421 3801 10424
rect 3835 10421 3847 10455
rect 3789 10415 3847 10421
rect 4338 10412 4344 10464
rect 4396 10452 4402 10464
rect 4706 10452 4712 10464
rect 4396 10424 4712 10452
rect 4396 10412 4402 10424
rect 4706 10412 4712 10424
rect 4764 10412 4770 10464
rect 4801 10455 4859 10461
rect 4801 10421 4813 10455
rect 4847 10452 4859 10455
rect 4890 10452 4896 10464
rect 4847 10424 4896 10452
rect 4847 10421 4859 10424
rect 4801 10415 4859 10421
rect 4890 10412 4896 10424
rect 4948 10412 4954 10464
rect 5000 10452 5028 10492
rect 5442 10480 5448 10532
rect 5500 10520 5506 10532
rect 5721 10523 5779 10529
rect 5721 10520 5733 10523
rect 5500 10492 5733 10520
rect 5500 10480 5506 10492
rect 5721 10489 5733 10492
rect 5767 10520 5779 10523
rect 10680 10523 10738 10529
rect 5767 10492 10640 10520
rect 5767 10489 5779 10492
rect 5721 10483 5779 10489
rect 6730 10452 6736 10464
rect 5000 10424 6736 10452
rect 6730 10412 6736 10424
rect 6788 10412 6794 10464
rect 7742 10412 7748 10464
rect 7800 10452 7806 10464
rect 9582 10452 9588 10464
rect 7800 10424 9588 10452
rect 7800 10412 7806 10424
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 9766 10452 9772 10464
rect 9727 10424 9772 10452
rect 9766 10412 9772 10424
rect 9824 10412 9830 10464
rect 9861 10455 9919 10461
rect 9861 10421 9873 10455
rect 9907 10452 9919 10455
rect 10502 10452 10508 10464
rect 9907 10424 10508 10452
rect 9907 10421 9919 10424
rect 9861 10415 9919 10421
rect 10502 10412 10508 10424
rect 10560 10412 10566 10464
rect 10612 10452 10640 10492
rect 10680 10489 10692 10523
rect 10726 10520 10738 10523
rect 11330 10520 11336 10532
rect 10726 10492 11336 10520
rect 10726 10489 10738 10492
rect 10680 10483 10738 10489
rect 11330 10480 11336 10492
rect 11388 10480 11394 10532
rect 14108 10452 14136 10560
rect 18506 10548 18512 10560
rect 18564 10548 18570 10600
rect 14268 10523 14326 10529
rect 14268 10489 14280 10523
rect 14314 10520 14326 10523
rect 14918 10520 14924 10532
rect 14314 10492 14924 10520
rect 14314 10489 14326 10492
rect 14268 10483 14326 10489
rect 14918 10480 14924 10492
rect 14976 10480 14982 10532
rect 16301 10523 16359 10529
rect 16301 10489 16313 10523
rect 16347 10520 16359 10523
rect 17313 10523 17371 10529
rect 16347 10492 16988 10520
rect 16347 10489 16359 10492
rect 16301 10483 16359 10489
rect 10612 10424 14136 10452
rect 15470 10412 15476 10464
rect 15528 10452 15534 10464
rect 15933 10455 15991 10461
rect 15933 10452 15945 10455
rect 15528 10424 15945 10452
rect 15528 10412 15534 10424
rect 15933 10421 15945 10424
rect 15979 10421 15991 10455
rect 16390 10452 16396 10464
rect 16351 10424 16396 10452
rect 15933 10415 15991 10421
rect 16390 10412 16396 10424
rect 16448 10412 16454 10464
rect 16960 10461 16988 10492
rect 17313 10489 17325 10523
rect 17359 10520 17371 10523
rect 18049 10523 18107 10529
rect 18049 10520 18061 10523
rect 17359 10492 18061 10520
rect 17359 10489 17371 10492
rect 17313 10483 17371 10489
rect 18049 10489 18061 10492
rect 18095 10489 18107 10523
rect 18049 10483 18107 10489
rect 16945 10455 17003 10461
rect 16945 10421 16957 10455
rect 16991 10421 17003 10455
rect 16945 10415 17003 10421
rect 1104 10362 18860 10384
rect 1104 10310 6912 10362
rect 6964 10310 6976 10362
rect 7028 10310 7040 10362
rect 7092 10310 7104 10362
rect 7156 10310 12843 10362
rect 12895 10310 12907 10362
rect 12959 10310 12971 10362
rect 13023 10310 13035 10362
rect 13087 10310 18860 10362
rect 1104 10288 18860 10310
rect 1949 10251 2007 10257
rect 1949 10217 1961 10251
rect 1995 10248 2007 10251
rect 2130 10248 2136 10260
rect 1995 10220 2136 10248
rect 1995 10217 2007 10220
rect 1949 10211 2007 10217
rect 2130 10208 2136 10220
rect 2188 10208 2194 10260
rect 2409 10251 2467 10257
rect 2409 10217 2421 10251
rect 2455 10248 2467 10251
rect 2961 10251 3019 10257
rect 2961 10248 2973 10251
rect 2455 10220 2973 10248
rect 2455 10217 2467 10220
rect 2409 10211 2467 10217
rect 2961 10217 2973 10220
rect 3007 10217 3019 10251
rect 2961 10211 3019 10217
rect 3421 10251 3479 10257
rect 3421 10217 3433 10251
rect 3467 10248 3479 10251
rect 3602 10248 3608 10260
rect 3467 10220 3608 10248
rect 3467 10217 3479 10220
rect 3421 10211 3479 10217
rect 3602 10208 3608 10220
rect 3660 10208 3666 10260
rect 4065 10251 4123 10257
rect 4065 10217 4077 10251
rect 4111 10217 4123 10251
rect 4065 10211 4123 10217
rect 2317 10183 2375 10189
rect 2317 10149 2329 10183
rect 2363 10180 2375 10183
rect 4080 10180 4108 10211
rect 4614 10208 4620 10260
rect 4672 10248 4678 10260
rect 4890 10248 4896 10260
rect 4672 10220 4896 10248
rect 4672 10208 4678 10220
rect 4890 10208 4896 10220
rect 4948 10248 4954 10260
rect 9674 10248 9680 10260
rect 4948 10220 7972 10248
rect 9635 10220 9680 10248
rect 4948 10208 4954 10220
rect 2363 10152 4108 10180
rect 4172 10152 4752 10180
rect 2363 10149 2375 10152
rect 2317 10143 2375 10149
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10072 1458 10124
rect 3050 10072 3056 10124
rect 3108 10112 3114 10124
rect 3329 10115 3387 10121
rect 3329 10112 3341 10115
rect 3108 10084 3341 10112
rect 3108 10072 3114 10084
rect 3329 10081 3341 10084
rect 3375 10081 3387 10115
rect 3329 10075 3387 10081
rect 3510 10072 3516 10124
rect 3568 10112 3574 10124
rect 3568 10084 3740 10112
rect 3568 10072 3574 10084
rect 2590 10044 2596 10056
rect 2551 10016 2596 10044
rect 2590 10004 2596 10016
rect 2648 10004 2654 10056
rect 3418 10004 3424 10056
rect 3476 10044 3482 10056
rect 3605 10047 3663 10053
rect 3605 10044 3617 10047
rect 3476 10016 3617 10044
rect 3476 10004 3482 10016
rect 3605 10013 3617 10016
rect 3651 10013 3663 10047
rect 3712 10044 3740 10084
rect 4062 10072 4068 10124
rect 4120 10112 4126 10124
rect 4172 10112 4200 10152
rect 4430 10112 4436 10124
rect 4120 10084 4200 10112
rect 4391 10084 4436 10112
rect 4120 10072 4126 10084
rect 4430 10072 4436 10084
rect 4488 10072 4494 10124
rect 4522 10044 4528 10056
rect 3712 10016 4528 10044
rect 3605 10007 3663 10013
rect 3620 9976 3648 10007
rect 4522 10004 4528 10016
rect 4580 10004 4586 10056
rect 4617 10047 4675 10053
rect 4617 10013 4629 10047
rect 4663 10013 4675 10047
rect 4724 10044 4752 10152
rect 5810 10140 5816 10192
rect 5868 10180 5874 10192
rect 6089 10183 6147 10189
rect 6089 10180 6101 10183
rect 5868 10152 6101 10180
rect 5868 10140 5874 10152
rect 6089 10149 6101 10152
rect 6135 10149 6147 10183
rect 6089 10143 6147 10149
rect 6178 10140 6184 10192
rect 6236 10140 6242 10192
rect 7650 10140 7656 10192
rect 7708 10180 7714 10192
rect 7806 10183 7864 10189
rect 7806 10180 7818 10183
rect 7708 10152 7818 10180
rect 7708 10140 7714 10152
rect 7806 10149 7818 10152
rect 7852 10149 7864 10183
rect 7806 10143 7864 10149
rect 5261 10115 5319 10121
rect 5261 10081 5273 10115
rect 5307 10112 5319 10115
rect 5994 10112 6000 10124
rect 5307 10084 6000 10112
rect 5307 10081 5319 10084
rect 5261 10075 5319 10081
rect 5994 10072 6000 10084
rect 6052 10072 6058 10124
rect 6196 10112 6224 10140
rect 6196 10084 6316 10112
rect 5626 10044 5632 10056
rect 4724 10016 5632 10044
rect 4617 10007 4675 10013
rect 4632 9976 4660 10007
rect 5626 10004 5632 10016
rect 5684 10044 5690 10056
rect 6288 10053 6316 10084
rect 6638 10072 6644 10124
rect 6696 10112 6702 10124
rect 7561 10115 7619 10121
rect 7561 10112 7573 10115
rect 6696 10084 7573 10112
rect 6696 10072 6702 10084
rect 7561 10081 7573 10084
rect 7607 10081 7619 10115
rect 7944 10112 7972 10220
rect 9674 10208 9680 10220
rect 9732 10208 9738 10260
rect 10042 10248 10048 10260
rect 10003 10220 10048 10248
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 10137 10251 10195 10257
rect 10137 10217 10149 10251
rect 10183 10248 10195 10251
rect 12345 10251 12403 10257
rect 12345 10248 12357 10251
rect 10183 10220 12357 10248
rect 10183 10217 10195 10220
rect 10137 10211 10195 10217
rect 12345 10217 12357 10220
rect 12391 10217 12403 10251
rect 12345 10211 12403 10217
rect 12434 10208 12440 10260
rect 12492 10248 12498 10260
rect 14918 10248 14924 10260
rect 12492 10220 13584 10248
rect 14879 10220 14924 10248
rect 12492 10208 12498 10220
rect 12618 10140 12624 10192
rect 12676 10180 12682 10192
rect 13446 10180 13452 10192
rect 12676 10152 13452 10180
rect 12676 10140 12682 10152
rect 13446 10140 13452 10152
rect 13504 10140 13510 10192
rect 13556 10180 13584 10220
rect 14918 10208 14924 10220
rect 14976 10208 14982 10260
rect 16390 10208 16396 10260
rect 16448 10248 16454 10260
rect 17037 10251 17095 10257
rect 17037 10248 17049 10251
rect 16448 10220 17049 10248
rect 16448 10208 16454 10220
rect 17037 10217 17049 10220
rect 17083 10217 17095 10251
rect 17494 10248 17500 10260
rect 17455 10220 17500 10248
rect 17037 10211 17095 10217
rect 17494 10208 17500 10220
rect 17552 10208 17558 10260
rect 17586 10180 17592 10192
rect 13556 10152 15424 10180
rect 10594 10112 10600 10124
rect 7944 10084 10600 10112
rect 7561 10075 7619 10081
rect 10594 10072 10600 10084
rect 10652 10072 10658 10124
rect 11054 10112 11060 10124
rect 11015 10084 11060 10112
rect 11054 10072 11060 10084
rect 11112 10072 11118 10124
rect 12710 10112 12716 10124
rect 12671 10084 12716 10112
rect 12710 10072 12716 10084
rect 12768 10072 12774 10124
rect 13556 10121 13584 10152
rect 13541 10115 13599 10121
rect 13541 10081 13553 10115
rect 13587 10112 13599 10115
rect 13630 10112 13636 10124
rect 13587 10084 13636 10112
rect 13587 10081 13599 10084
rect 13541 10075 13599 10081
rect 13630 10072 13636 10084
rect 13688 10072 13694 10124
rect 13808 10115 13866 10121
rect 13808 10081 13820 10115
rect 13854 10112 13866 10115
rect 15194 10112 15200 10124
rect 13854 10084 15200 10112
rect 13854 10081 13866 10084
rect 13808 10075 13866 10081
rect 15194 10072 15200 10084
rect 15252 10072 15258 10124
rect 15396 10121 15424 10152
rect 17144 10152 17592 10180
rect 15381 10115 15439 10121
rect 15381 10081 15393 10115
rect 15427 10081 15439 10115
rect 15381 10075 15439 10081
rect 15648 10115 15706 10121
rect 15648 10081 15660 10115
rect 15694 10112 15706 10115
rect 16114 10112 16120 10124
rect 15694 10084 16120 10112
rect 15694 10081 15706 10084
rect 15648 10075 15706 10081
rect 16114 10072 16120 10084
rect 16172 10112 16178 10124
rect 17144 10112 17172 10152
rect 17586 10140 17592 10152
rect 17644 10140 17650 10192
rect 16172 10084 17172 10112
rect 16172 10072 16178 10084
rect 17218 10072 17224 10124
rect 17276 10112 17282 10124
rect 17405 10115 17463 10121
rect 17405 10112 17417 10115
rect 17276 10084 17417 10112
rect 17276 10072 17282 10084
rect 17405 10081 17417 10084
rect 17451 10081 17463 10115
rect 17405 10075 17463 10081
rect 6181 10047 6239 10053
rect 6181 10044 6193 10047
rect 5684 10016 6193 10044
rect 5684 10004 5690 10016
rect 6181 10013 6193 10016
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 6273 10047 6331 10053
rect 6273 10013 6285 10047
rect 6319 10013 6331 10047
rect 6273 10007 6331 10013
rect 6733 10047 6791 10053
rect 6733 10013 6745 10047
rect 6779 10044 6791 10047
rect 7466 10044 7472 10056
rect 6779 10016 7472 10044
rect 6779 10013 6791 10016
rect 6733 10007 6791 10013
rect 7466 10004 7472 10016
rect 7524 10004 7530 10056
rect 10318 10044 10324 10056
rect 10279 10016 10324 10044
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 11146 10004 11152 10056
rect 11204 10044 11210 10056
rect 11204 10016 11249 10044
rect 11204 10004 11210 10016
rect 11330 10004 11336 10056
rect 11388 10044 11394 10056
rect 12802 10044 12808 10056
rect 11388 10016 11433 10044
rect 12763 10016 12808 10044
rect 11388 10004 11394 10016
rect 12802 10004 12808 10016
rect 12860 10004 12866 10056
rect 17604 10053 17632 10140
rect 18046 10112 18052 10124
rect 18007 10084 18052 10112
rect 18046 10072 18052 10084
rect 18104 10072 18110 10124
rect 12897 10047 12955 10053
rect 12897 10013 12909 10047
rect 12943 10013 12955 10047
rect 12897 10007 12955 10013
rect 17589 10047 17647 10053
rect 17589 10013 17601 10047
rect 17635 10013 17647 10047
rect 17589 10007 17647 10013
rect 3620 9948 4660 9976
rect 4706 9936 4712 9988
rect 4764 9976 4770 9988
rect 4764 9948 7328 9976
rect 4764 9936 4770 9948
rect 1394 9868 1400 9920
rect 1452 9908 1458 9920
rect 1581 9911 1639 9917
rect 1581 9908 1593 9911
rect 1452 9880 1593 9908
rect 1452 9868 1458 9880
rect 1581 9877 1593 9880
rect 1627 9877 1639 9911
rect 1581 9871 1639 9877
rect 4246 9868 4252 9920
rect 4304 9908 4310 9920
rect 5077 9911 5135 9917
rect 5077 9908 5089 9911
rect 4304 9880 5089 9908
rect 4304 9868 4310 9880
rect 5077 9877 5089 9880
rect 5123 9908 5135 9911
rect 5534 9908 5540 9920
rect 5123 9880 5540 9908
rect 5123 9877 5135 9880
rect 5077 9871 5135 9877
rect 5534 9868 5540 9880
rect 5592 9868 5598 9920
rect 5721 9911 5779 9917
rect 5721 9877 5733 9911
rect 5767 9908 5779 9911
rect 7190 9908 7196 9920
rect 5767 9880 7196 9908
rect 5767 9877 5779 9880
rect 5721 9871 5779 9877
rect 7190 9868 7196 9880
rect 7248 9868 7254 9920
rect 7300 9908 7328 9948
rect 8496 9948 9076 9976
rect 8496 9908 8524 9948
rect 7300 9880 8524 9908
rect 8846 9868 8852 9920
rect 8904 9908 8910 9920
rect 8941 9911 8999 9917
rect 8941 9908 8953 9911
rect 8904 9880 8953 9908
rect 8904 9868 8910 9880
rect 8941 9877 8953 9880
rect 8987 9877 8999 9911
rect 9048 9908 9076 9948
rect 9766 9936 9772 9988
rect 9824 9976 9830 9988
rect 10689 9979 10747 9985
rect 10689 9976 10701 9979
rect 9824 9948 10701 9976
rect 9824 9936 9830 9948
rect 10689 9945 10701 9948
rect 10735 9945 10747 9979
rect 10689 9939 10747 9945
rect 11882 9936 11888 9988
rect 11940 9976 11946 9988
rect 12250 9976 12256 9988
rect 11940 9948 12256 9976
rect 11940 9936 11946 9948
rect 12250 9936 12256 9948
rect 12308 9936 12314 9988
rect 12342 9936 12348 9988
rect 12400 9976 12406 9988
rect 12912 9976 12940 10007
rect 12400 9948 12940 9976
rect 12400 9936 12406 9948
rect 10594 9908 10600 9920
rect 9048 9880 10600 9908
rect 8941 9871 8999 9877
rect 10594 9868 10600 9880
rect 10652 9868 10658 9920
rect 15194 9868 15200 9920
rect 15252 9908 15258 9920
rect 16482 9908 16488 9920
rect 15252 9880 16488 9908
rect 15252 9868 15258 9880
rect 16482 9868 16488 9880
rect 16540 9908 16546 9920
rect 16761 9911 16819 9917
rect 16761 9908 16773 9911
rect 16540 9880 16773 9908
rect 16540 9868 16546 9880
rect 16761 9877 16773 9880
rect 16807 9877 16819 9911
rect 16761 9871 16819 9877
rect 18233 9911 18291 9917
rect 18233 9877 18245 9911
rect 18279 9908 18291 9911
rect 18414 9908 18420 9920
rect 18279 9880 18420 9908
rect 18279 9877 18291 9880
rect 18233 9871 18291 9877
rect 18414 9868 18420 9880
rect 18472 9868 18478 9920
rect 1104 9818 18860 9840
rect 1104 9766 3947 9818
rect 3999 9766 4011 9818
rect 4063 9766 4075 9818
rect 4127 9766 4139 9818
rect 4191 9766 9878 9818
rect 9930 9766 9942 9818
rect 9994 9766 10006 9818
rect 10058 9766 10070 9818
rect 10122 9766 15808 9818
rect 15860 9766 15872 9818
rect 15924 9766 15936 9818
rect 15988 9766 16000 9818
rect 16052 9766 18860 9818
rect 1104 9744 18860 9766
rect 2682 9664 2688 9716
rect 2740 9704 2746 9716
rect 3329 9707 3387 9713
rect 3329 9704 3341 9707
rect 2740 9676 3341 9704
rect 2740 9664 2746 9676
rect 3329 9673 3341 9676
rect 3375 9673 3387 9707
rect 3329 9667 3387 9673
rect 3418 9664 3424 9716
rect 3476 9664 3482 9716
rect 7668 9676 7972 9704
rect 3436 9568 3464 9664
rect 5902 9596 5908 9648
rect 5960 9636 5966 9648
rect 6825 9639 6883 9645
rect 6825 9636 6837 9639
rect 5960 9608 6837 9636
rect 5960 9596 5966 9608
rect 6825 9605 6837 9608
rect 6871 9605 6883 9639
rect 7668 9636 7696 9676
rect 7834 9636 7840 9648
rect 6825 9599 6883 9605
rect 7024 9608 7696 9636
rect 7795 9608 7840 9636
rect 3786 9568 3792 9580
rect 3436 9540 3792 9568
rect 3786 9528 3792 9540
rect 3844 9528 3850 9580
rect 4062 9528 4068 9580
rect 4120 9568 4126 9580
rect 4433 9571 4491 9577
rect 4433 9568 4445 9571
rect 4120 9540 4445 9568
rect 4120 9528 4126 9540
rect 4433 9537 4445 9540
rect 4479 9537 4491 9571
rect 4433 9531 4491 9537
rect 6178 9528 6184 9580
rect 6236 9568 6242 9580
rect 6273 9571 6331 9577
rect 6273 9568 6285 9571
rect 6236 9540 6285 9568
rect 6236 9528 6242 9540
rect 6273 9537 6285 9540
rect 6319 9537 6331 9571
rect 6273 9531 6331 9537
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 1762 9500 1768 9512
rect 1443 9472 1768 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1762 9460 1768 9472
rect 1820 9460 1826 9512
rect 1946 9460 1952 9512
rect 2004 9500 2010 9512
rect 4893 9503 4951 9509
rect 2004 9472 2452 9500
rect 2004 9460 2010 9472
rect 2424 9444 2452 9472
rect 4893 9469 4905 9503
rect 4939 9500 4951 9503
rect 7024 9500 7052 9608
rect 7834 9596 7840 9608
rect 7892 9596 7898 9648
rect 7944 9636 7972 9676
rect 8478 9664 8484 9716
rect 8536 9704 8542 9716
rect 9030 9704 9036 9716
rect 8536 9676 9036 9704
rect 8536 9664 8542 9676
rect 9030 9664 9036 9676
rect 9088 9664 9094 9716
rect 10502 9664 10508 9716
rect 10560 9704 10566 9716
rect 10597 9707 10655 9713
rect 10597 9704 10609 9707
rect 10560 9676 10609 9704
rect 10560 9664 10566 9676
rect 10597 9673 10609 9676
rect 10643 9673 10655 9707
rect 11330 9704 11336 9716
rect 11243 9676 11336 9704
rect 10597 9667 10655 9673
rect 8294 9636 8300 9648
rect 7944 9608 8300 9636
rect 8294 9596 8300 9608
rect 8352 9596 8358 9648
rect 8570 9596 8576 9648
rect 8628 9596 8634 9648
rect 9490 9596 9496 9648
rect 9548 9636 9554 9648
rect 9548 9608 11192 9636
rect 9548 9596 9554 9608
rect 7374 9568 7380 9580
rect 7287 9540 7380 9568
rect 7374 9528 7380 9540
rect 7432 9568 7438 9580
rect 8389 9571 8447 9577
rect 8389 9568 8401 9571
rect 7432 9540 8401 9568
rect 7432 9528 7438 9540
rect 8389 9537 8401 9540
rect 8435 9537 8447 9571
rect 8579 9568 8607 9596
rect 9398 9568 9404 9580
rect 8579 9540 8708 9568
rect 9359 9540 9404 9568
rect 8389 9531 8447 9537
rect 7190 9500 7196 9512
rect 4939 9472 7052 9500
rect 7151 9472 7196 9500
rect 4939 9469 4951 9472
rect 4893 9463 4951 9469
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 7466 9460 7472 9512
rect 7524 9500 7530 9512
rect 8205 9503 8263 9509
rect 8205 9500 8217 9503
rect 7524 9472 8217 9500
rect 7524 9460 7530 9472
rect 8205 9469 8217 9472
rect 8251 9469 8263 9503
rect 8680 9500 8708 9540
rect 9398 9528 9404 9540
rect 9456 9528 9462 9580
rect 10778 9528 10784 9580
rect 10836 9568 10842 9580
rect 11057 9571 11115 9577
rect 11057 9568 11069 9571
rect 10836 9540 11069 9568
rect 10836 9528 10842 9540
rect 11057 9537 11069 9540
rect 11103 9537 11115 9571
rect 11057 9531 11115 9537
rect 9217 9503 9275 9509
rect 9217 9500 9229 9503
rect 8680 9472 9229 9500
rect 8205 9463 8263 9469
rect 9217 9469 9229 9472
rect 9263 9500 9275 9503
rect 10594 9500 10600 9512
rect 9263 9472 10600 9500
rect 9263 9469 9275 9472
rect 9217 9463 9275 9469
rect 10594 9460 10600 9472
rect 10652 9460 10658 9512
rect 10870 9460 10876 9512
rect 10928 9500 10934 9512
rect 10965 9503 11023 9509
rect 10965 9500 10977 9503
rect 10928 9472 10977 9500
rect 10928 9460 10934 9472
rect 10965 9469 10977 9472
rect 11011 9469 11023 9503
rect 11164 9500 11192 9608
rect 11256 9577 11284 9676
rect 11330 9664 11336 9676
rect 11388 9704 11394 9716
rect 12342 9704 12348 9716
rect 11388 9676 12348 9704
rect 11388 9664 11394 9676
rect 12342 9664 12348 9676
rect 12400 9664 12406 9716
rect 12434 9664 12440 9716
rect 12492 9704 12498 9716
rect 12492 9676 12756 9704
rect 12492 9664 12498 9676
rect 12728 9636 12756 9676
rect 12802 9664 12808 9716
rect 12860 9704 12866 9716
rect 12897 9707 12955 9713
rect 12897 9704 12909 9707
rect 12860 9676 12909 9704
rect 12860 9664 12866 9676
rect 12897 9673 12909 9676
rect 12943 9673 12955 9707
rect 15378 9704 15384 9716
rect 12897 9667 12955 9673
rect 13004 9676 15384 9704
rect 13004 9636 13032 9676
rect 15378 9664 15384 9676
rect 15436 9664 15442 9716
rect 17494 9704 17500 9716
rect 16500 9676 17500 9704
rect 16500 9636 16528 9676
rect 17494 9664 17500 9676
rect 17552 9664 17558 9716
rect 12728 9608 13032 9636
rect 13096 9608 16528 9636
rect 11241 9571 11299 9577
rect 11241 9537 11253 9571
rect 11287 9537 11299 9571
rect 11606 9568 11612 9580
rect 11567 9540 11612 9568
rect 11241 9531 11299 9537
rect 11606 9528 11612 9540
rect 11664 9528 11670 9580
rect 13096 9500 13124 9608
rect 13538 9528 13544 9580
rect 13596 9568 13602 9580
rect 14918 9568 14924 9580
rect 13596 9540 13641 9568
rect 14879 9540 14924 9568
rect 13596 9528 13602 9540
rect 14918 9528 14924 9540
rect 14976 9528 14982 9580
rect 15194 9528 15200 9580
rect 15252 9568 15258 9580
rect 15841 9571 15899 9577
rect 15841 9568 15853 9571
rect 15252 9540 15853 9568
rect 15252 9528 15258 9540
rect 15841 9537 15853 9540
rect 15887 9537 15899 9571
rect 15841 9531 15899 9537
rect 16114 9528 16120 9580
rect 16172 9568 16178 9580
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16172 9540 16865 9568
rect 16172 9528 16178 9540
rect 16853 9537 16865 9540
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 17218 9528 17224 9580
rect 17276 9568 17282 9580
rect 17954 9568 17960 9580
rect 17276 9540 17960 9568
rect 17276 9528 17282 9540
rect 17954 9528 17960 9540
rect 18012 9528 18018 9580
rect 11164 9472 13124 9500
rect 14645 9503 14703 9509
rect 10965 9463 11023 9469
rect 14645 9469 14657 9503
rect 14691 9500 14703 9503
rect 15470 9500 15476 9512
rect 14691 9472 15476 9500
rect 14691 9469 14703 9472
rect 14645 9463 14703 9469
rect 15470 9460 15476 9472
rect 15528 9460 15534 9512
rect 16574 9460 16580 9512
rect 16632 9500 16638 9512
rect 17405 9503 17463 9509
rect 17405 9500 17417 9503
rect 16632 9472 17417 9500
rect 16632 9460 16638 9472
rect 17405 9469 17417 9472
rect 17451 9469 17463 9503
rect 17405 9463 17463 9469
rect 18049 9503 18107 9509
rect 18049 9469 18061 9503
rect 18095 9469 18107 9503
rect 18049 9463 18107 9469
rect 2222 9441 2228 9444
rect 2216 9432 2228 9441
rect 2183 9404 2228 9432
rect 2216 9395 2228 9404
rect 2222 9392 2228 9395
rect 2280 9392 2286 9444
rect 2406 9392 2412 9444
rect 2464 9432 2470 9444
rect 3326 9432 3332 9444
rect 2464 9404 3332 9432
rect 2464 9392 2470 9404
rect 3326 9392 3332 9404
rect 3384 9432 3390 9444
rect 4154 9432 4160 9444
rect 3384 9404 4160 9432
rect 3384 9392 3390 9404
rect 4154 9392 4160 9404
rect 4212 9392 4218 9444
rect 4430 9392 4436 9444
rect 4488 9432 4494 9444
rect 5169 9435 5227 9441
rect 5169 9432 5181 9435
rect 4488 9404 5181 9432
rect 4488 9392 4494 9404
rect 5169 9401 5181 9404
rect 5215 9401 5227 9435
rect 7285 9435 7343 9441
rect 7285 9432 7297 9435
rect 5169 9395 5227 9401
rect 5736 9404 7297 9432
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 3418 9324 3424 9376
rect 3476 9364 3482 9376
rect 3881 9367 3939 9373
rect 3881 9364 3893 9367
rect 3476 9336 3893 9364
rect 3476 9324 3482 9336
rect 3881 9333 3893 9336
rect 3927 9333 3939 9367
rect 4246 9364 4252 9376
rect 4207 9336 4252 9364
rect 3881 9327 3939 9333
rect 4246 9324 4252 9336
rect 4304 9324 4310 9376
rect 4338 9324 4344 9376
rect 4396 9364 4402 9376
rect 4396 9336 4441 9364
rect 4396 9324 4402 9336
rect 4522 9324 4528 9376
rect 4580 9364 4586 9376
rect 5074 9364 5080 9376
rect 4580 9336 5080 9364
rect 4580 9324 4586 9336
rect 5074 9324 5080 9336
rect 5132 9324 5138 9376
rect 5736 9373 5764 9404
rect 7285 9401 7297 9404
rect 7331 9401 7343 9435
rect 12158 9432 12164 9444
rect 7285 9395 7343 9401
rect 7392 9404 12164 9432
rect 5721 9367 5779 9373
rect 5721 9333 5733 9367
rect 5767 9333 5779 9367
rect 6086 9364 6092 9376
rect 6047 9336 6092 9364
rect 5721 9327 5779 9333
rect 6086 9324 6092 9336
rect 6144 9324 6150 9376
rect 6178 9324 6184 9376
rect 6236 9364 6242 9376
rect 6236 9336 6281 9364
rect 6236 9324 6242 9336
rect 6454 9324 6460 9376
rect 6512 9364 6518 9376
rect 7392 9364 7420 9404
rect 12158 9392 12164 9404
rect 12216 9392 12222 9444
rect 12802 9392 12808 9444
rect 12860 9432 12866 9444
rect 18064 9432 18092 9463
rect 12860 9404 18092 9432
rect 12860 9392 12866 9404
rect 6512 9336 7420 9364
rect 6512 9324 6518 9336
rect 7558 9324 7564 9376
rect 7616 9364 7622 9376
rect 8202 9364 8208 9376
rect 7616 9336 8208 9364
rect 7616 9324 7622 9336
rect 8202 9324 8208 9336
rect 8260 9364 8266 9376
rect 8297 9367 8355 9373
rect 8297 9364 8309 9367
rect 8260 9336 8309 9364
rect 8260 9324 8266 9336
rect 8297 9333 8309 9336
rect 8343 9333 8355 9367
rect 8297 9327 8355 9333
rect 8386 9324 8392 9376
rect 8444 9364 8450 9376
rect 8662 9364 8668 9376
rect 8444 9336 8668 9364
rect 8444 9324 8450 9336
rect 8662 9324 8668 9336
rect 8720 9324 8726 9376
rect 8849 9367 8907 9373
rect 8849 9333 8861 9367
rect 8895 9364 8907 9367
rect 9030 9364 9036 9376
rect 8895 9336 9036 9364
rect 8895 9333 8907 9336
rect 8849 9327 8907 9333
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 9122 9324 9128 9376
rect 9180 9364 9186 9376
rect 9309 9367 9367 9373
rect 9309 9364 9321 9367
rect 9180 9336 9321 9364
rect 9180 9324 9186 9336
rect 9309 9333 9321 9336
rect 9355 9364 9367 9367
rect 11974 9364 11980 9376
rect 9355 9336 11980 9364
rect 9355 9333 9367 9336
rect 9309 9327 9367 9333
rect 11974 9324 11980 9336
rect 12032 9324 12038 9376
rect 12342 9324 12348 9376
rect 12400 9364 12406 9376
rect 13265 9367 13323 9373
rect 13265 9364 13277 9367
rect 12400 9336 13277 9364
rect 12400 9324 12406 9336
rect 13265 9333 13277 9336
rect 13311 9333 13323 9367
rect 13265 9327 13323 9333
rect 13357 9367 13415 9373
rect 13357 9333 13369 9367
rect 13403 9364 13415 9367
rect 14090 9364 14096 9376
rect 13403 9336 14096 9364
rect 13403 9333 13415 9336
rect 13357 9327 13415 9333
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 14277 9367 14335 9373
rect 14277 9333 14289 9367
rect 14323 9364 14335 9367
rect 14458 9364 14464 9376
rect 14323 9336 14464 9364
rect 14323 9333 14335 9336
rect 14277 9327 14335 9333
rect 14458 9324 14464 9336
rect 14516 9324 14522 9376
rect 14737 9367 14795 9373
rect 14737 9333 14749 9367
rect 14783 9364 14795 9367
rect 15289 9367 15347 9373
rect 15289 9364 15301 9367
rect 14783 9336 15301 9364
rect 14783 9333 14795 9336
rect 14737 9327 14795 9333
rect 15289 9333 15301 9336
rect 15335 9333 15347 9367
rect 15654 9364 15660 9376
rect 15615 9336 15660 9364
rect 15289 9327 15347 9333
rect 15654 9324 15660 9336
rect 15712 9324 15718 9376
rect 15749 9367 15807 9373
rect 15749 9333 15761 9367
rect 15795 9364 15807 9367
rect 16301 9367 16359 9373
rect 16301 9364 16313 9367
rect 15795 9336 16313 9364
rect 15795 9333 15807 9336
rect 15749 9327 15807 9333
rect 16301 9333 16313 9336
rect 16347 9333 16359 9367
rect 16666 9364 16672 9376
rect 16627 9336 16672 9364
rect 16301 9327 16359 9333
rect 16666 9324 16672 9336
rect 16724 9324 16730 9376
rect 16758 9324 16764 9376
rect 16816 9364 16822 9376
rect 17586 9364 17592 9376
rect 16816 9336 16861 9364
rect 17547 9336 17592 9364
rect 16816 9324 16822 9336
rect 17586 9324 17592 9336
rect 17644 9324 17650 9376
rect 18233 9367 18291 9373
rect 18233 9333 18245 9367
rect 18279 9364 18291 9367
rect 18322 9364 18328 9376
rect 18279 9336 18328 9364
rect 18279 9333 18291 9336
rect 18233 9327 18291 9333
rect 18322 9324 18328 9336
rect 18380 9324 18386 9376
rect 1104 9274 18860 9296
rect 1104 9222 6912 9274
rect 6964 9222 6976 9274
rect 7028 9222 7040 9274
rect 7092 9222 7104 9274
rect 7156 9222 12843 9274
rect 12895 9222 12907 9274
rect 12959 9222 12971 9274
rect 13023 9222 13035 9274
rect 13087 9222 18860 9274
rect 1104 9200 18860 9222
rect 4338 9120 4344 9172
rect 4396 9160 4402 9172
rect 4893 9163 4951 9169
rect 4893 9160 4905 9163
rect 4396 9132 4905 9160
rect 4396 9120 4402 9132
rect 4893 9129 4905 9132
rect 4939 9129 4951 9163
rect 4893 9123 4951 9129
rect 8573 9163 8631 9169
rect 8573 9129 8585 9163
rect 8619 9160 8631 9163
rect 10137 9163 10195 9169
rect 10137 9160 10149 9163
rect 8619 9132 10149 9160
rect 8619 9129 8631 9132
rect 8573 9123 8631 9129
rect 10137 9129 10149 9132
rect 10183 9129 10195 9163
rect 10137 9123 10195 9129
rect 11882 9120 11888 9172
rect 11940 9160 11946 9172
rect 12250 9160 12256 9172
rect 11940 9132 12256 9160
rect 11940 9120 11946 9132
rect 12250 9120 12256 9132
rect 12308 9120 12314 9172
rect 12710 9120 12716 9172
rect 12768 9160 12774 9172
rect 12897 9163 12955 9169
rect 12897 9160 12909 9163
rect 12768 9132 12909 9160
rect 12768 9120 12774 9132
rect 12897 9129 12909 9132
rect 12943 9129 12955 9163
rect 12897 9123 12955 9129
rect 13170 9120 13176 9172
rect 13228 9160 13234 9172
rect 15286 9160 15292 9172
rect 13228 9132 15292 9160
rect 13228 9120 13234 9132
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 15654 9120 15660 9172
rect 15712 9160 15718 9172
rect 15749 9163 15807 9169
rect 15749 9160 15761 9163
rect 15712 9132 15761 9160
rect 15712 9120 15718 9132
rect 15749 9129 15761 9132
rect 15795 9129 15807 9163
rect 15749 9123 15807 9129
rect 16117 9163 16175 9169
rect 16117 9129 16129 9163
rect 16163 9160 16175 9163
rect 16390 9160 16396 9172
rect 16163 9132 16396 9160
rect 16163 9129 16175 9132
rect 16117 9123 16175 9129
rect 16390 9120 16396 9132
rect 16448 9120 16454 9172
rect 16666 9120 16672 9172
rect 16724 9160 16730 9172
rect 16761 9163 16819 9169
rect 16761 9160 16773 9163
rect 16724 9132 16773 9160
rect 16724 9120 16730 9132
rect 16761 9129 16773 9132
rect 16807 9129 16819 9163
rect 17126 9160 17132 9172
rect 17087 9132 17132 9160
rect 16761 9123 16819 9129
rect 17126 9120 17132 9132
rect 17184 9120 17190 9172
rect 1946 9092 1952 9104
rect 1596 9064 1952 9092
rect 1596 9033 1624 9064
rect 1946 9052 1952 9064
rect 2004 9052 2010 9104
rect 8941 9095 8999 9101
rect 8941 9092 8953 9095
rect 5092 9064 8953 9092
rect 1854 9033 1860 9036
rect 1581 9027 1639 9033
rect 1581 8993 1593 9027
rect 1627 8993 1639 9027
rect 1581 8987 1639 8993
rect 1848 8987 1860 9033
rect 1912 9024 1918 9036
rect 4062 9024 4068 9036
rect 1912 8996 4068 9024
rect 1854 8984 1860 8987
rect 1912 8984 1918 8996
rect 4062 8984 4068 8996
rect 4120 9024 4126 9036
rect 4890 9024 4896 9036
rect 4120 8996 4896 9024
rect 4120 8984 4126 8996
rect 4890 8984 4896 8996
rect 4948 8984 4954 9036
rect 3050 8916 3056 8968
rect 3108 8956 3114 8968
rect 5092 8956 5120 9064
rect 8941 9061 8953 9064
rect 8987 9092 8999 9095
rect 9030 9092 9036 9104
rect 8987 9064 9036 9092
rect 8987 9061 8999 9064
rect 8941 9055 8999 9061
rect 9030 9052 9036 9064
rect 9088 9052 9094 9104
rect 9122 9052 9128 9104
rect 9180 9092 9186 9104
rect 10045 9095 10103 9101
rect 10045 9092 10057 9095
rect 9180 9064 10057 9092
rect 9180 9052 9186 9064
rect 10045 9061 10057 9064
rect 10091 9061 10103 9095
rect 10045 9055 10103 9061
rect 13078 9052 13084 9104
rect 13136 9092 13142 9104
rect 13265 9095 13323 9101
rect 13265 9092 13277 9095
rect 13136 9064 13277 9092
rect 13136 9052 13142 9064
rect 13265 9061 13277 9064
rect 13311 9092 13323 9095
rect 18598 9092 18604 9104
rect 13311 9064 18604 9092
rect 13311 9061 13323 9064
rect 13265 9055 13323 9061
rect 18598 9052 18604 9064
rect 18656 9052 18662 9104
rect 5258 9024 5264 9036
rect 5219 8996 5264 9024
rect 5258 8984 5264 8996
rect 5316 8984 5322 9036
rect 5534 8984 5540 9036
rect 5592 9024 5598 9036
rect 6638 9024 6644 9036
rect 5592 8996 6644 9024
rect 5592 8984 5598 8996
rect 6638 8984 6644 8996
rect 6696 9024 6702 9036
rect 6825 9027 6883 9033
rect 6825 9024 6837 9027
rect 6696 8996 6837 9024
rect 6696 8984 6702 8996
rect 6825 8993 6837 8996
rect 6871 8993 6883 9027
rect 6825 8987 6883 8993
rect 7092 9027 7150 9033
rect 7092 8993 7104 9027
rect 7138 9024 7150 9027
rect 9398 9024 9404 9036
rect 7138 8996 9404 9024
rect 7138 8993 7150 8996
rect 7092 8987 7150 8993
rect 8956 8968 8984 8996
rect 5350 8956 5356 8968
rect 3108 8928 5120 8956
rect 5311 8928 5356 8956
rect 3108 8916 3114 8928
rect 5350 8916 5356 8928
rect 5408 8916 5414 8968
rect 5442 8916 5448 8968
rect 5500 8956 5506 8968
rect 5500 8928 5545 8956
rect 5500 8916 5506 8928
rect 8938 8916 8944 8968
rect 8996 8916 9002 8968
rect 9030 8916 9036 8968
rect 9088 8956 9094 8968
rect 9232 8965 9260 8996
rect 9398 8984 9404 8996
rect 9456 8984 9462 9036
rect 9582 8984 9588 9036
rect 9640 9024 9646 9036
rect 11054 9024 11060 9036
rect 9640 8996 11060 9024
rect 9640 8984 9646 8996
rect 11054 8984 11060 8996
rect 11112 8984 11118 9036
rect 11232 9027 11290 9033
rect 11232 8993 11244 9027
rect 11278 9024 11290 9027
rect 11698 9024 11704 9036
rect 11278 8996 11704 9024
rect 11278 8993 11290 8996
rect 11232 8987 11290 8993
rect 11698 8984 11704 8996
rect 11756 8984 11762 9036
rect 12158 8984 12164 9036
rect 12216 9024 12222 9036
rect 12805 9027 12863 9033
rect 12805 9024 12817 9027
rect 12216 8996 12817 9024
rect 12216 8984 12222 8996
rect 12805 8993 12817 8996
rect 12851 8993 12863 9027
rect 12805 8987 12863 8993
rect 12986 8984 12992 9036
rect 13044 9024 13050 9036
rect 13357 9027 13415 9033
rect 13357 9024 13369 9027
rect 13044 8996 13369 9024
rect 13044 8984 13050 8996
rect 13357 8993 13369 8996
rect 13403 9024 13415 9027
rect 14734 9024 14740 9036
rect 13403 8996 14740 9024
rect 13403 8993 13415 8996
rect 13357 8987 13415 8993
rect 14734 8984 14740 8996
rect 14792 8984 14798 9036
rect 16209 9027 16267 9033
rect 16209 8993 16221 9027
rect 16255 9024 16267 9027
rect 16942 9024 16948 9036
rect 16255 8996 16948 9024
rect 16255 8993 16267 8996
rect 16209 8987 16267 8993
rect 16942 8984 16948 8996
rect 17000 8984 17006 9036
rect 17865 9027 17923 9033
rect 17865 8993 17877 9027
rect 17911 9024 17923 9027
rect 17954 9024 17960 9036
rect 17911 8996 17960 9024
rect 17911 8993 17923 8996
rect 17865 8987 17923 8993
rect 17954 8984 17960 8996
rect 18012 8984 18018 9036
rect 9217 8959 9275 8965
rect 9088 8928 9133 8956
rect 9088 8916 9094 8928
rect 9217 8925 9229 8959
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 9490 8916 9496 8968
rect 9548 8956 9554 8968
rect 10229 8959 10287 8965
rect 10229 8956 10241 8959
rect 9548 8928 10241 8956
rect 9548 8916 9554 8928
rect 10229 8925 10241 8928
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 10410 8916 10416 8968
rect 10468 8956 10474 8968
rect 10870 8956 10876 8968
rect 10468 8928 10876 8956
rect 10468 8916 10474 8928
rect 10870 8916 10876 8928
rect 10928 8956 10934 8968
rect 10965 8959 11023 8965
rect 10965 8956 10977 8959
rect 10928 8928 10977 8956
rect 10928 8916 10934 8928
rect 10965 8925 10977 8928
rect 11011 8925 11023 8959
rect 13538 8956 13544 8968
rect 13499 8928 13544 8956
rect 10965 8919 11023 8925
rect 13538 8916 13544 8928
rect 13596 8916 13602 8968
rect 16393 8959 16451 8965
rect 16393 8925 16405 8959
rect 16439 8956 16451 8959
rect 16574 8956 16580 8968
rect 16439 8928 16580 8956
rect 16439 8925 16451 8928
rect 16393 8919 16451 8925
rect 16574 8916 16580 8928
rect 16632 8916 16638 8968
rect 17218 8956 17224 8968
rect 17179 8928 17224 8956
rect 17218 8916 17224 8928
rect 17276 8916 17282 8968
rect 17310 8916 17316 8968
rect 17368 8956 17374 8968
rect 17368 8928 17413 8956
rect 17368 8916 17374 8928
rect 8205 8891 8263 8897
rect 8205 8857 8217 8891
rect 8251 8888 8263 8891
rect 8386 8888 8392 8900
rect 8251 8860 8392 8888
rect 8251 8857 8263 8860
rect 8205 8851 8263 8857
rect 8386 8848 8392 8860
rect 8444 8848 8450 8900
rect 9582 8848 9588 8900
rect 9640 8888 9646 8900
rect 12986 8888 12992 8900
rect 9640 8860 9812 8888
rect 9640 8848 9646 8860
rect 2222 8780 2228 8832
rect 2280 8820 2286 8832
rect 2961 8823 3019 8829
rect 2961 8820 2973 8823
rect 2280 8792 2973 8820
rect 2280 8780 2286 8792
rect 2961 8789 2973 8792
rect 3007 8789 3019 8823
rect 2961 8783 3019 8789
rect 8294 8780 8300 8832
rect 8352 8820 8358 8832
rect 9677 8823 9735 8829
rect 9677 8820 9689 8823
rect 8352 8792 9689 8820
rect 8352 8780 8358 8792
rect 9677 8789 9689 8792
rect 9723 8789 9735 8823
rect 9784 8820 9812 8860
rect 11900 8860 12992 8888
rect 11900 8820 11928 8860
rect 12986 8848 12992 8860
rect 13044 8848 13050 8900
rect 13262 8848 13268 8900
rect 13320 8888 13326 8900
rect 17034 8888 17040 8900
rect 13320 8860 17040 8888
rect 13320 8848 13326 8860
rect 17034 8848 17040 8860
rect 17092 8848 17098 8900
rect 12342 8820 12348 8832
rect 9784 8792 11928 8820
rect 12303 8792 12348 8820
rect 9677 8783 9735 8789
rect 12342 8780 12348 8792
rect 12400 8780 12406 8832
rect 12621 8823 12679 8829
rect 12621 8789 12633 8823
rect 12667 8820 12679 8823
rect 13630 8820 13636 8832
rect 12667 8792 13636 8820
rect 12667 8789 12679 8792
rect 12621 8783 12679 8789
rect 13630 8780 13636 8792
rect 13688 8780 13694 8832
rect 14090 8780 14096 8832
rect 14148 8820 14154 8832
rect 16850 8820 16856 8832
rect 14148 8792 16856 8820
rect 14148 8780 14154 8792
rect 16850 8780 16856 8792
rect 16908 8780 16914 8832
rect 18046 8820 18052 8832
rect 18007 8792 18052 8820
rect 18046 8780 18052 8792
rect 18104 8780 18110 8832
rect 1104 8730 18860 8752
rect 1104 8678 3947 8730
rect 3999 8678 4011 8730
rect 4063 8678 4075 8730
rect 4127 8678 4139 8730
rect 4191 8678 9878 8730
rect 9930 8678 9942 8730
rect 9994 8678 10006 8730
rect 10058 8678 10070 8730
rect 10122 8678 15808 8730
rect 15860 8678 15872 8730
rect 15924 8678 15936 8730
rect 15988 8678 16000 8730
rect 16052 8678 18860 8730
rect 1104 8656 18860 8678
rect 3326 8576 3332 8628
rect 3384 8616 3390 8628
rect 3513 8619 3571 8625
rect 3513 8616 3525 8619
rect 3384 8588 3525 8616
rect 3384 8576 3390 8588
rect 3513 8585 3525 8588
rect 3559 8585 3571 8619
rect 3513 8579 3571 8585
rect 4890 8576 4896 8628
rect 4948 8616 4954 8628
rect 4985 8619 5043 8625
rect 4985 8616 4997 8619
rect 4948 8588 4997 8616
rect 4948 8576 4954 8588
rect 4985 8585 4997 8588
rect 5031 8585 5043 8619
rect 4985 8579 5043 8585
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 5445 8619 5503 8625
rect 5445 8616 5457 8619
rect 5408 8588 5457 8616
rect 5408 8576 5414 8588
rect 5445 8585 5457 8588
rect 5491 8585 5503 8619
rect 5445 8579 5503 8585
rect 5994 8576 6000 8628
rect 6052 8576 6058 8628
rect 7377 8619 7435 8625
rect 7377 8585 7389 8619
rect 7423 8616 7435 8619
rect 11698 8616 11704 8628
rect 7423 8588 11560 8616
rect 11659 8588 11704 8616
rect 7423 8585 7435 8588
rect 7377 8579 7435 8585
rect 3050 8508 3056 8560
rect 3108 8548 3114 8560
rect 3602 8548 3608 8560
rect 3108 8520 3608 8548
rect 3108 8508 3114 8520
rect 3602 8508 3608 8520
rect 3660 8508 3666 8560
rect 6012 8548 6040 8576
rect 6457 8551 6515 8557
rect 6457 8548 6469 8551
rect 6012 8520 6469 8548
rect 6457 8517 6469 8520
rect 6503 8548 6515 8551
rect 6730 8548 6736 8560
rect 6503 8520 6736 8548
rect 6503 8517 6515 8520
rect 6457 8511 6515 8517
rect 6730 8508 6736 8520
rect 6788 8508 6794 8560
rect 9769 8551 9827 8557
rect 9769 8548 9781 8551
rect 8036 8520 9781 8548
rect 3237 8483 3295 8489
rect 3237 8449 3249 8483
rect 3283 8480 3295 8483
rect 3326 8480 3332 8492
rect 3283 8452 3332 8480
rect 3283 8449 3295 8452
rect 3237 8443 3295 8449
rect 3326 8440 3332 8452
rect 3384 8440 3390 8492
rect 5994 8480 6000 8492
rect 3528 8452 3740 8480
rect 5955 8452 6000 8480
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8412 1731 8415
rect 3528 8412 3556 8452
rect 1719 8384 3556 8412
rect 3605 8415 3663 8421
rect 1719 8381 1731 8384
rect 1673 8375 1731 8381
rect 3605 8381 3617 8415
rect 3651 8381 3663 8415
rect 3712 8412 3740 8452
rect 5994 8440 6000 8452
rect 6052 8440 6058 8492
rect 5813 8415 5871 8421
rect 5813 8412 5825 8415
rect 3712 8384 5825 8412
rect 3605 8375 3663 8381
rect 5813 8381 5825 8384
rect 5859 8412 5871 8415
rect 6086 8412 6092 8424
rect 5859 8384 6092 8412
rect 5859 8381 5871 8384
rect 5813 8375 5871 8381
rect 3513 8347 3571 8353
rect 3513 8313 3525 8347
rect 3559 8344 3571 8347
rect 3620 8344 3648 8375
rect 6086 8372 6092 8384
rect 6144 8372 6150 8424
rect 6641 8415 6699 8421
rect 6641 8381 6653 8415
rect 6687 8412 6699 8415
rect 8036 8412 8064 8520
rect 9769 8517 9781 8520
rect 9815 8548 9827 8551
rect 10318 8548 10324 8560
rect 9815 8520 10324 8548
rect 9815 8517 9827 8520
rect 9769 8511 9827 8517
rect 10318 8508 10324 8520
rect 10376 8508 10382 8560
rect 8113 8483 8171 8489
rect 8113 8449 8125 8483
rect 8159 8480 8171 8483
rect 8386 8480 8392 8492
rect 8159 8452 8392 8480
rect 8159 8449 8171 8452
rect 8113 8443 8171 8449
rect 8386 8440 8392 8452
rect 8444 8480 8450 8492
rect 9490 8480 9496 8492
rect 8444 8452 9496 8480
rect 8444 8440 8450 8452
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 8478 8412 8484 8424
rect 6687 8384 8064 8412
rect 8439 8384 8484 8412
rect 6687 8381 6699 8384
rect 6641 8375 6699 8381
rect 8478 8372 8484 8384
rect 8536 8372 8542 8424
rect 9674 8372 9680 8424
rect 9732 8412 9738 8424
rect 10321 8415 10379 8421
rect 10321 8412 10333 8415
rect 9732 8384 10333 8412
rect 9732 8372 9738 8384
rect 10321 8381 10333 8384
rect 10367 8412 10379 8415
rect 10870 8412 10876 8424
rect 10367 8384 10876 8412
rect 10367 8381 10379 8384
rect 10321 8375 10379 8381
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 11532 8412 11560 8588
rect 11698 8576 11704 8588
rect 11756 8576 11762 8628
rect 12986 8576 12992 8628
rect 13044 8616 13050 8628
rect 14090 8616 14096 8628
rect 13044 8588 14096 8616
rect 13044 8576 13050 8588
rect 14090 8576 14096 8588
rect 14148 8576 14154 8628
rect 15841 8619 15899 8625
rect 14384 8588 15424 8616
rect 11716 8480 11744 8576
rect 12434 8508 12440 8560
rect 12492 8548 12498 8560
rect 14274 8548 14280 8560
rect 12492 8520 14280 8548
rect 12492 8508 12498 8520
rect 14274 8508 14280 8520
rect 14332 8508 14338 8560
rect 13446 8480 13452 8492
rect 11716 8452 13452 8480
rect 13446 8440 13452 8452
rect 13504 8440 13510 8492
rect 13265 8415 13323 8421
rect 11532 8384 13216 8412
rect 3878 8353 3884 8356
rect 3872 8344 3884 8353
rect 3559 8316 3648 8344
rect 3791 8316 3884 8344
rect 3559 8313 3571 8316
rect 3513 8307 3571 8313
rect 3872 8307 3884 8316
rect 3936 8344 3942 8356
rect 5442 8344 5448 8356
rect 3936 8316 5448 8344
rect 3878 8304 3884 8307
rect 3936 8304 3942 8316
rect 5442 8304 5448 8316
rect 5500 8304 5506 8356
rect 5905 8347 5963 8353
rect 5905 8313 5917 8347
rect 5951 8344 5963 8347
rect 6178 8344 6184 8356
rect 5951 8316 6184 8344
rect 5951 8313 5963 8316
rect 5905 8307 5963 8313
rect 6178 8304 6184 8316
rect 6236 8344 6242 8356
rect 7377 8347 7435 8353
rect 7377 8344 7389 8347
rect 6236 8316 7389 8344
rect 6236 8304 6242 8316
rect 7377 8313 7389 8316
rect 7423 8313 7435 8347
rect 7377 8307 7435 8313
rect 7742 8304 7748 8356
rect 7800 8344 7806 8356
rect 7837 8347 7895 8353
rect 7837 8344 7849 8347
rect 7800 8316 7849 8344
rect 7800 8304 7806 8316
rect 7837 8313 7849 8316
rect 7883 8313 7895 8347
rect 7837 8307 7895 8313
rect 7929 8347 7987 8353
rect 7929 8313 7941 8347
rect 7975 8344 7987 8347
rect 8202 8344 8208 8356
rect 7975 8316 8208 8344
rect 7975 8313 7987 8316
rect 7929 8307 7987 8313
rect 8202 8304 8208 8316
rect 8260 8304 8266 8356
rect 8570 8304 8576 8356
rect 8628 8344 8634 8356
rect 10410 8344 10416 8356
rect 8628 8316 10416 8344
rect 8628 8304 8634 8316
rect 10410 8304 10416 8316
rect 10468 8304 10474 8356
rect 10502 8304 10508 8356
rect 10560 8353 10566 8356
rect 10560 8347 10624 8353
rect 10560 8313 10578 8347
rect 10612 8313 10624 8347
rect 10560 8307 10624 8313
rect 10560 8304 10566 8307
rect 934 8236 940 8288
rect 992 8276 998 8288
rect 1857 8279 1915 8285
rect 1857 8276 1869 8279
rect 992 8248 1869 8276
rect 992 8236 998 8248
rect 1857 8245 1869 8248
rect 1903 8245 1915 8279
rect 1857 8239 1915 8245
rect 2498 8236 2504 8288
rect 2556 8276 2562 8288
rect 2593 8279 2651 8285
rect 2593 8276 2605 8279
rect 2556 8248 2605 8276
rect 2556 8236 2562 8248
rect 2593 8245 2605 8248
rect 2639 8245 2651 8279
rect 2958 8276 2964 8288
rect 2919 8248 2964 8276
rect 2593 8239 2651 8245
rect 2958 8236 2964 8248
rect 3016 8236 3022 8288
rect 3050 8236 3056 8288
rect 3108 8276 3114 8288
rect 6454 8276 6460 8288
rect 3108 8248 6460 8276
rect 3108 8236 3114 8248
rect 6454 8236 6460 8248
rect 6512 8236 6518 8288
rect 7466 8276 7472 8288
rect 7427 8248 7472 8276
rect 7466 8236 7472 8248
rect 7524 8236 7530 8288
rect 8938 8236 8944 8288
rect 8996 8276 9002 8288
rect 12250 8276 12256 8288
rect 8996 8248 12256 8276
rect 8996 8236 9002 8248
rect 12250 8236 12256 8248
rect 12308 8236 12314 8288
rect 12618 8236 12624 8288
rect 12676 8276 12682 8288
rect 12897 8279 12955 8285
rect 12897 8276 12909 8279
rect 12676 8248 12909 8276
rect 12676 8236 12682 8248
rect 12897 8245 12909 8248
rect 12943 8245 12955 8279
rect 13188 8276 13216 8384
rect 13265 8381 13277 8415
rect 13311 8412 13323 8415
rect 13722 8412 13728 8424
rect 13311 8384 13728 8412
rect 13311 8381 13323 8384
rect 13265 8375 13323 8381
rect 13722 8372 13728 8384
rect 13780 8412 13786 8424
rect 14384 8412 14412 8588
rect 15396 8548 15424 8588
rect 15841 8585 15853 8619
rect 15887 8616 15899 8619
rect 16114 8616 16120 8628
rect 15887 8588 16120 8616
rect 15887 8585 15899 8588
rect 15841 8579 15899 8585
rect 16114 8576 16120 8588
rect 16172 8616 16178 8628
rect 16574 8616 16580 8628
rect 16172 8588 16580 8616
rect 16172 8576 16178 8588
rect 16574 8576 16580 8588
rect 16632 8576 16638 8628
rect 16758 8616 16764 8628
rect 16719 8588 16764 8616
rect 16758 8576 16764 8588
rect 16816 8576 16822 8628
rect 17126 8548 17132 8560
rect 15396 8520 17132 8548
rect 17126 8508 17132 8520
rect 17184 8508 17190 8560
rect 16666 8480 16672 8492
rect 16040 8452 16672 8480
rect 13780 8384 14412 8412
rect 14461 8415 14519 8421
rect 13780 8372 13786 8384
rect 14461 8381 14473 8415
rect 14507 8381 14519 8415
rect 14461 8375 14519 8381
rect 14728 8415 14786 8421
rect 14728 8381 14740 8415
rect 14774 8412 14786 8415
rect 16040 8412 16068 8452
rect 16666 8440 16672 8452
rect 16724 8480 16730 8492
rect 17310 8480 17316 8492
rect 16724 8452 17316 8480
rect 16724 8440 16730 8452
rect 17310 8440 17316 8452
rect 17368 8440 17374 8492
rect 14774 8384 16068 8412
rect 14774 8381 14786 8384
rect 14728 8375 14786 8381
rect 13538 8304 13544 8356
rect 13596 8344 13602 8356
rect 14476 8344 14504 8375
rect 16114 8372 16120 8424
rect 16172 8421 16178 8424
rect 16172 8415 16210 8421
rect 16198 8381 16210 8415
rect 17126 8412 17132 8424
rect 17087 8384 17132 8412
rect 16172 8375 16210 8381
rect 16172 8372 16178 8375
rect 17126 8372 17132 8384
rect 17184 8372 17190 8424
rect 17954 8372 17960 8424
rect 18012 8412 18018 8424
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 18012 8384 18061 8412
rect 18012 8372 18018 8384
rect 18049 8381 18061 8384
rect 18095 8381 18107 8415
rect 18049 8375 18107 8381
rect 14918 8344 14924 8356
rect 13596 8316 14924 8344
rect 13596 8304 13602 8316
rect 14918 8304 14924 8316
rect 14976 8304 14982 8356
rect 15562 8304 15568 8356
rect 15620 8344 15626 8356
rect 16255 8347 16313 8353
rect 16255 8344 16267 8347
rect 15620 8316 16267 8344
rect 15620 8304 15626 8316
rect 16255 8313 16267 8316
rect 16301 8313 16313 8347
rect 16255 8307 16313 8313
rect 13357 8279 13415 8285
rect 13357 8276 13369 8279
rect 13188 8248 13369 8276
rect 12897 8239 12955 8245
rect 13357 8245 13369 8248
rect 13403 8276 13415 8279
rect 17126 8276 17132 8288
rect 13403 8248 17132 8276
rect 13403 8245 13415 8248
rect 13357 8239 13415 8245
rect 17126 8236 17132 8248
rect 17184 8276 17190 8288
rect 17221 8279 17279 8285
rect 17221 8276 17233 8279
rect 17184 8248 17233 8276
rect 17184 8236 17190 8248
rect 17221 8245 17233 8248
rect 17267 8245 17279 8279
rect 18230 8276 18236 8288
rect 18191 8248 18236 8276
rect 17221 8239 17279 8245
rect 18230 8236 18236 8248
rect 18288 8236 18294 8288
rect 1104 8186 18860 8208
rect 1104 8134 6912 8186
rect 6964 8134 6976 8186
rect 7028 8134 7040 8186
rect 7092 8134 7104 8186
rect 7156 8134 12843 8186
rect 12895 8134 12907 8186
rect 12959 8134 12971 8186
rect 13023 8134 13035 8186
rect 13087 8134 18860 8186
rect 1104 8112 18860 8134
rect 2041 8075 2099 8081
rect 2041 8041 2053 8075
rect 2087 8072 2099 8075
rect 3418 8072 3424 8084
rect 2087 8044 3424 8072
rect 2087 8041 2099 8044
rect 2041 8035 2099 8041
rect 3418 8032 3424 8044
rect 3476 8032 3482 8084
rect 4525 8075 4583 8081
rect 4525 8041 4537 8075
rect 4571 8072 4583 8075
rect 5258 8072 5264 8084
rect 4571 8044 5264 8072
rect 4571 8041 4583 8044
rect 4525 8035 4583 8041
rect 5258 8032 5264 8044
rect 5316 8032 5322 8084
rect 5442 8032 5448 8084
rect 5500 8072 5506 8084
rect 6917 8075 6975 8081
rect 6917 8072 6929 8075
rect 5500 8044 6929 8072
rect 5500 8032 5506 8044
rect 6917 8041 6929 8044
rect 6963 8041 6975 8075
rect 6917 8035 6975 8041
rect 7466 8032 7472 8084
rect 7524 8072 7530 8084
rect 8021 8075 8079 8081
rect 8021 8072 8033 8075
rect 7524 8044 8033 8072
rect 7524 8032 7530 8044
rect 8021 8041 8033 8044
rect 8067 8041 8079 8075
rect 8021 8035 8079 8041
rect 8113 8075 8171 8081
rect 8113 8041 8125 8075
rect 8159 8072 8171 8075
rect 8294 8072 8300 8084
rect 8159 8044 8300 8072
rect 8159 8041 8171 8044
rect 8113 8035 8171 8041
rect 8294 8032 8300 8044
rect 8352 8032 8358 8084
rect 12345 8075 12403 8081
rect 8680 8044 11652 8072
rect 2130 7964 2136 8016
rect 2188 8004 2194 8016
rect 3053 8007 3111 8013
rect 3053 8004 3065 8007
rect 2188 7976 3065 8004
rect 2188 7964 2194 7976
rect 3053 7973 3065 7976
rect 3099 8004 3111 8007
rect 3510 8004 3516 8016
rect 3099 7976 3516 8004
rect 3099 7973 3111 7976
rect 3053 7967 3111 7973
rect 3510 7964 3516 7976
rect 3568 7964 3574 8016
rect 5804 8007 5862 8013
rect 5804 8004 5816 8007
rect 5184 7976 5816 8004
rect 1946 7936 1952 7948
rect 1907 7908 1952 7936
rect 1946 7896 1952 7908
rect 2004 7896 2010 7948
rect 2682 7896 2688 7948
rect 2740 7936 2746 7948
rect 2961 7939 3019 7945
rect 2961 7936 2973 7939
rect 2740 7908 2973 7936
rect 2740 7896 2746 7908
rect 2961 7905 2973 7908
rect 3007 7905 3019 7939
rect 2961 7899 3019 7905
rect 4893 7939 4951 7945
rect 4893 7905 4905 7939
rect 4939 7905 4951 7939
rect 4893 7899 4951 7905
rect 2222 7868 2228 7880
rect 2183 7840 2228 7868
rect 2222 7828 2228 7840
rect 2280 7828 2286 7880
rect 3237 7871 3295 7877
rect 3237 7837 3249 7871
rect 3283 7868 3295 7871
rect 3326 7868 3332 7880
rect 3283 7840 3332 7868
rect 3283 7837 3295 7840
rect 3237 7831 3295 7837
rect 3326 7828 3332 7840
rect 3384 7868 3390 7880
rect 3878 7868 3884 7880
rect 3384 7840 3884 7868
rect 3384 7828 3390 7840
rect 3878 7828 3884 7840
rect 3936 7828 3942 7880
rect 1486 7692 1492 7744
rect 1544 7732 1550 7744
rect 1581 7735 1639 7741
rect 1581 7732 1593 7735
rect 1544 7704 1593 7732
rect 1544 7692 1550 7704
rect 1581 7701 1593 7704
rect 1627 7701 1639 7735
rect 2590 7732 2596 7744
rect 2551 7704 2596 7732
rect 1581 7695 1639 7701
rect 2590 7692 2596 7704
rect 2648 7692 2654 7744
rect 4338 7692 4344 7744
rect 4396 7732 4402 7744
rect 4908 7732 4936 7899
rect 5184 7880 5212 7976
rect 5804 7973 5816 7976
rect 5850 8004 5862 8007
rect 5994 8004 6000 8016
rect 5850 7976 6000 8004
rect 5850 7973 5862 7976
rect 5804 7967 5862 7973
rect 5994 7964 6000 7976
rect 6052 7964 6058 8016
rect 5534 7936 5540 7948
rect 5495 7908 5540 7936
rect 5534 7896 5540 7908
rect 5592 7896 5598 7948
rect 5626 7896 5632 7948
rect 5684 7936 5690 7948
rect 8680 7936 8708 8044
rect 9766 8004 9772 8016
rect 5684 7908 8708 7936
rect 8864 7976 9772 8004
rect 5684 7896 5690 7908
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7837 5043 7871
rect 5166 7868 5172 7880
rect 5079 7840 5172 7868
rect 4985 7831 5043 7837
rect 5000 7800 5028 7831
rect 5166 7828 5172 7840
rect 5224 7828 5230 7880
rect 5644 7868 5672 7896
rect 5276 7840 5672 7868
rect 8205 7871 8263 7877
rect 5276 7800 5304 7840
rect 8205 7837 8217 7871
rect 8251 7868 8263 7871
rect 8864 7868 8892 7976
rect 9766 7964 9772 7976
rect 9824 8004 9830 8016
rect 9922 8007 9980 8013
rect 9922 8004 9934 8007
rect 9824 7976 9934 8004
rect 9824 7964 9830 7976
rect 9922 7973 9934 7976
rect 9968 7973 9980 8007
rect 9922 7967 9980 7973
rect 8938 7896 8944 7948
rect 8996 7936 9002 7948
rect 8996 7908 9041 7936
rect 8996 7896 9002 7908
rect 10318 7896 10324 7948
rect 10376 7936 10382 7948
rect 11517 7939 11575 7945
rect 11517 7936 11529 7939
rect 10376 7908 11529 7936
rect 10376 7896 10382 7908
rect 11517 7905 11529 7908
rect 11563 7905 11575 7939
rect 11624 7936 11652 8044
rect 12345 8041 12357 8075
rect 12391 8072 12403 8075
rect 12618 8072 12624 8084
rect 12391 8044 12624 8072
rect 12391 8041 12403 8044
rect 12345 8035 12403 8041
rect 12618 8032 12624 8044
rect 12676 8032 12682 8084
rect 12897 8075 12955 8081
rect 12897 8041 12909 8075
rect 12943 8041 12955 8075
rect 13262 8072 13268 8084
rect 13223 8044 13268 8072
rect 12897 8035 12955 8041
rect 12253 8007 12311 8013
rect 12253 7973 12265 8007
rect 12299 8004 12311 8007
rect 12912 8004 12940 8035
rect 13262 8032 13268 8044
rect 13320 8032 13326 8084
rect 16666 8072 16672 8084
rect 16627 8044 16672 8072
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 16942 8072 16948 8084
rect 16903 8044 16948 8072
rect 16942 8032 16948 8044
rect 17000 8032 17006 8084
rect 17313 8075 17371 8081
rect 17313 8041 17325 8075
rect 17359 8072 17371 8075
rect 17770 8072 17776 8084
rect 17359 8044 17776 8072
rect 17359 8041 17371 8044
rect 17313 8035 17371 8041
rect 17770 8032 17776 8044
rect 17828 8032 17834 8084
rect 13357 8007 13415 8013
rect 13357 8004 13369 8007
rect 12299 7976 12940 8004
rect 13188 7976 13369 8004
rect 12299 7973 12311 7976
rect 12253 7967 12311 7973
rect 13188 7936 13216 7976
rect 13357 7973 13369 7976
rect 13403 8004 13415 8007
rect 16684 8004 16712 8032
rect 13403 7976 15700 8004
rect 16684 7976 17540 8004
rect 13403 7973 13415 7976
rect 13357 7967 13415 7973
rect 14274 7936 14280 7948
rect 11624 7908 13216 7936
rect 14235 7908 14280 7936
rect 11517 7899 11575 7905
rect 14274 7896 14280 7908
rect 14332 7896 14338 7948
rect 14369 7939 14427 7945
rect 14369 7905 14381 7939
rect 14415 7936 14427 7939
rect 14642 7936 14648 7948
rect 14415 7908 14648 7936
rect 14415 7905 14427 7908
rect 14369 7899 14427 7905
rect 9030 7868 9036 7880
rect 8251 7840 8892 7868
rect 8991 7840 9036 7868
rect 8251 7837 8263 7840
rect 8205 7831 8263 7837
rect 9030 7828 9036 7840
rect 9088 7828 9094 7880
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7868 9275 7871
rect 9398 7868 9404 7880
rect 9263 7840 9404 7868
rect 9263 7837 9275 7840
rect 9217 7831 9275 7837
rect 9398 7828 9404 7840
rect 9456 7828 9462 7880
rect 9674 7828 9680 7880
rect 9732 7868 9738 7880
rect 9732 7840 9777 7868
rect 10704 7840 12296 7868
rect 9732 7828 9738 7840
rect 5000 7772 5304 7800
rect 6564 7772 7788 7800
rect 5810 7732 5816 7744
rect 4396 7704 5816 7732
rect 4396 7692 4402 7704
rect 5810 7692 5816 7704
rect 5868 7732 5874 7744
rect 6564 7732 6592 7772
rect 7650 7732 7656 7744
rect 5868 7704 6592 7732
rect 7611 7704 7656 7732
rect 5868 7692 5874 7704
rect 7650 7692 7656 7704
rect 7708 7692 7714 7744
rect 7760 7732 7788 7772
rect 8294 7760 8300 7812
rect 8352 7800 8358 7812
rect 8573 7803 8631 7809
rect 8573 7800 8585 7803
rect 8352 7772 8585 7800
rect 8352 7760 8358 7772
rect 8573 7769 8585 7772
rect 8619 7769 8631 7803
rect 10704 7800 10732 7840
rect 8573 7763 8631 7769
rect 10612 7772 10732 7800
rect 11333 7803 11391 7809
rect 10612 7732 10640 7772
rect 11333 7769 11345 7803
rect 11379 7800 11391 7803
rect 11974 7800 11980 7812
rect 11379 7772 11980 7800
rect 11379 7769 11391 7772
rect 11333 7763 11391 7769
rect 11974 7760 11980 7772
rect 12032 7800 12038 7812
rect 12158 7800 12164 7812
rect 12032 7772 12164 7800
rect 12032 7760 12038 7772
rect 12158 7760 12164 7772
rect 12216 7760 12222 7812
rect 12268 7800 12296 7840
rect 12342 7828 12348 7880
rect 12400 7868 12406 7880
rect 12529 7871 12587 7877
rect 12529 7868 12541 7871
rect 12400 7840 12541 7868
rect 12400 7828 12406 7840
rect 12529 7837 12541 7840
rect 12575 7868 12587 7871
rect 13170 7868 13176 7880
rect 12575 7840 13176 7868
rect 12575 7837 12587 7840
rect 12529 7831 12587 7837
rect 13170 7828 13176 7840
rect 13228 7828 13234 7880
rect 13446 7868 13452 7880
rect 13407 7840 13452 7868
rect 13446 7828 13452 7840
rect 13504 7828 13510 7880
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 14384 7868 14412 7899
rect 14642 7896 14648 7908
rect 14700 7896 14706 7948
rect 15194 7896 15200 7948
rect 15252 7936 15258 7948
rect 15545 7939 15603 7945
rect 15545 7936 15557 7939
rect 15252 7908 15557 7936
rect 15252 7896 15258 7908
rect 15545 7905 15557 7908
rect 15591 7905 15603 7939
rect 15672 7936 15700 7976
rect 17218 7936 17224 7948
rect 15672 7908 17224 7936
rect 15545 7899 15603 7905
rect 17218 7896 17224 7908
rect 17276 7896 17282 7948
rect 17402 7936 17408 7948
rect 17363 7908 17408 7936
rect 17402 7896 17408 7908
rect 17460 7896 17466 7948
rect 13964 7840 14412 7868
rect 14461 7871 14519 7877
rect 13964 7828 13970 7840
rect 14461 7837 14473 7871
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 13262 7800 13268 7812
rect 12268 7772 13268 7800
rect 13262 7760 13268 7772
rect 13320 7760 13326 7812
rect 13464 7800 13492 7828
rect 14476 7800 14504 7831
rect 14918 7828 14924 7880
rect 14976 7868 14982 7880
rect 15289 7871 15347 7877
rect 15289 7868 15301 7871
rect 14976 7840 15301 7868
rect 14976 7828 14982 7840
rect 15289 7837 15301 7840
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 13464 7772 14504 7800
rect 17236 7800 17264 7896
rect 17512 7877 17540 7976
rect 17586 7964 17592 8016
rect 17644 8004 17650 8016
rect 17862 8004 17868 8016
rect 17644 7976 17868 8004
rect 17644 7964 17650 7976
rect 17862 7964 17868 7976
rect 17920 7964 17926 8016
rect 17957 7939 18015 7945
rect 17957 7905 17969 7939
rect 18003 7905 18015 7939
rect 17957 7899 18015 7905
rect 17497 7871 17555 7877
rect 17497 7837 17509 7871
rect 17543 7837 17555 7871
rect 17497 7831 17555 7837
rect 17972 7800 18000 7899
rect 17236 7772 18000 7800
rect 7760 7704 10640 7732
rect 10870 7692 10876 7744
rect 10928 7732 10934 7744
rect 11057 7735 11115 7741
rect 11057 7732 11069 7735
rect 10928 7704 11069 7732
rect 10928 7692 10934 7704
rect 11057 7701 11069 7704
rect 11103 7701 11115 7735
rect 11057 7695 11115 7701
rect 11790 7692 11796 7744
rect 11848 7732 11854 7744
rect 11885 7735 11943 7741
rect 11885 7732 11897 7735
rect 11848 7704 11897 7732
rect 11848 7692 11854 7704
rect 11885 7701 11897 7704
rect 11931 7701 11943 7735
rect 11885 7695 11943 7701
rect 13078 7692 13084 7744
rect 13136 7732 13142 7744
rect 13909 7735 13967 7741
rect 13909 7732 13921 7735
rect 13136 7704 13921 7732
rect 13136 7692 13142 7704
rect 13909 7701 13921 7704
rect 13955 7701 13967 7735
rect 13909 7695 13967 7701
rect 14274 7692 14280 7744
rect 14332 7732 14338 7744
rect 16482 7732 16488 7744
rect 14332 7704 16488 7732
rect 14332 7692 14338 7704
rect 16482 7692 16488 7704
rect 16540 7692 16546 7744
rect 17126 7692 17132 7744
rect 17184 7732 17190 7744
rect 17402 7732 17408 7744
rect 17184 7704 17408 7732
rect 17184 7692 17190 7704
rect 17402 7692 17408 7704
rect 17460 7692 17466 7744
rect 18141 7735 18199 7741
rect 18141 7701 18153 7735
rect 18187 7732 18199 7735
rect 18690 7732 18696 7744
rect 18187 7704 18696 7732
rect 18187 7701 18199 7704
rect 18141 7695 18199 7701
rect 18690 7692 18696 7704
rect 18748 7692 18754 7744
rect 1104 7642 18860 7664
rect 1104 7590 3947 7642
rect 3999 7590 4011 7642
rect 4063 7590 4075 7642
rect 4127 7590 4139 7642
rect 4191 7590 9878 7642
rect 9930 7590 9942 7642
rect 9994 7590 10006 7642
rect 10058 7590 10070 7642
rect 10122 7590 15808 7642
rect 15860 7590 15872 7642
rect 15924 7590 15936 7642
rect 15988 7590 16000 7642
rect 16052 7590 18860 7642
rect 1104 7568 18860 7590
rect 1762 7528 1768 7540
rect 1723 7500 1768 7528
rect 1762 7488 1768 7500
rect 1820 7488 1826 7540
rect 1946 7488 1952 7540
rect 2004 7528 2010 7540
rect 2133 7531 2191 7537
rect 2133 7528 2145 7531
rect 2004 7500 2145 7528
rect 2004 7488 2010 7500
rect 2133 7497 2145 7500
rect 2179 7497 2191 7531
rect 2133 7491 2191 7497
rect 3605 7531 3663 7537
rect 3605 7497 3617 7531
rect 3651 7528 3663 7531
rect 4246 7528 4252 7540
rect 3651 7500 4252 7528
rect 3651 7497 3663 7500
rect 3605 7491 3663 7497
rect 4246 7488 4252 7500
rect 4304 7488 4310 7540
rect 9677 7531 9735 7537
rect 9677 7528 9689 7531
rect 8312 7500 9689 7528
rect 5442 7460 5448 7472
rect 4264 7432 5448 7460
rect 1854 7352 1860 7404
rect 1912 7392 1918 7404
rect 2685 7395 2743 7401
rect 2685 7392 2697 7395
rect 1912 7364 2697 7392
rect 1912 7352 1918 7364
rect 2685 7361 2697 7364
rect 2731 7361 2743 7395
rect 2685 7355 2743 7361
rect 2958 7352 2964 7404
rect 3016 7392 3022 7404
rect 4264 7401 4292 7432
rect 5442 7420 5448 7432
rect 5500 7420 5506 7472
rect 3145 7395 3203 7401
rect 3145 7392 3157 7395
rect 3016 7364 3157 7392
rect 3016 7352 3022 7364
rect 3145 7361 3157 7364
rect 3191 7361 3203 7395
rect 3145 7355 3203 7361
rect 4249 7395 4307 7401
rect 4249 7361 4261 7395
rect 4295 7361 4307 7395
rect 5166 7392 5172 7404
rect 5127 7364 5172 7392
rect 4249 7355 4307 7361
rect 5166 7352 5172 7364
rect 5224 7352 5230 7404
rect 6178 7392 6184 7404
rect 6139 7364 6184 7392
rect 6178 7352 6184 7364
rect 6236 7352 6242 7404
rect 7742 7392 7748 7404
rect 7703 7364 7748 7392
rect 7742 7352 7748 7364
rect 7800 7352 7806 7404
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7392 7987 7395
rect 8312 7392 8340 7500
rect 9677 7497 9689 7500
rect 9723 7528 9735 7531
rect 9766 7528 9772 7540
rect 9723 7500 9772 7528
rect 9723 7497 9735 7500
rect 9677 7491 9735 7497
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 13906 7528 13912 7540
rect 9876 7500 13912 7528
rect 9876 7460 9904 7500
rect 13906 7488 13912 7500
rect 13964 7488 13970 7540
rect 14090 7488 14096 7540
rect 14148 7528 14154 7540
rect 15470 7528 15476 7540
rect 14148 7500 15476 7528
rect 14148 7488 14154 7500
rect 15470 7488 15476 7500
rect 15528 7488 15534 7540
rect 16114 7488 16120 7540
rect 16172 7528 16178 7540
rect 16298 7528 16304 7540
rect 16172 7500 16304 7528
rect 16172 7488 16178 7500
rect 16298 7488 16304 7500
rect 16356 7488 16362 7540
rect 7975 7364 8340 7392
rect 9784 7432 9904 7460
rect 7975 7361 7987 7364
rect 7929 7355 7987 7361
rect 1581 7327 1639 7333
rect 1581 7293 1593 7327
rect 1627 7324 1639 7327
rect 3050 7324 3056 7336
rect 1627 7296 3056 7324
rect 1627 7293 1639 7296
rect 1581 7287 1639 7293
rect 3050 7284 3056 7296
rect 3108 7284 3114 7336
rect 4798 7284 4804 7336
rect 4856 7324 4862 7336
rect 5077 7327 5135 7333
rect 5077 7324 5089 7327
rect 4856 7296 5089 7324
rect 4856 7284 4862 7296
rect 5077 7293 5089 7296
rect 5123 7324 5135 7327
rect 8294 7324 8300 7336
rect 5123 7296 8156 7324
rect 8255 7296 8300 7324
rect 5123 7293 5135 7296
rect 5077 7287 5135 7293
rect 2498 7256 2504 7268
rect 2459 7228 2504 7256
rect 2498 7216 2504 7228
rect 2556 7216 2562 7268
rect 2590 7216 2596 7268
rect 2648 7256 2654 7268
rect 2648 7228 2693 7256
rect 2648 7216 2654 7228
rect 3786 7216 3792 7268
rect 3844 7256 3850 7268
rect 3973 7259 4031 7265
rect 3973 7256 3985 7259
rect 3844 7228 3985 7256
rect 3844 7216 3850 7228
rect 3973 7225 3985 7228
rect 4019 7256 4031 7259
rect 7653 7259 7711 7265
rect 4019 7228 7420 7256
rect 4019 7225 4031 7228
rect 3973 7219 4031 7225
rect 4065 7191 4123 7197
rect 4065 7157 4077 7191
rect 4111 7188 4123 7191
rect 4617 7191 4675 7197
rect 4617 7188 4629 7191
rect 4111 7160 4629 7188
rect 4111 7157 4123 7160
rect 4065 7151 4123 7157
rect 4617 7157 4629 7160
rect 4663 7157 4675 7191
rect 4982 7188 4988 7200
rect 4943 7160 4988 7188
rect 4617 7151 4675 7157
rect 4982 7148 4988 7160
rect 5040 7148 5046 7200
rect 5626 7188 5632 7200
rect 5587 7160 5632 7188
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 5994 7188 6000 7200
rect 5955 7160 6000 7188
rect 5994 7148 6000 7160
rect 6052 7148 6058 7200
rect 6086 7148 6092 7200
rect 6144 7188 6150 7200
rect 7282 7188 7288 7200
rect 6144 7160 6189 7188
rect 7243 7160 7288 7188
rect 6144 7148 6150 7160
rect 7282 7148 7288 7160
rect 7340 7148 7346 7200
rect 7392 7188 7420 7228
rect 7653 7225 7665 7259
rect 7699 7256 7711 7259
rect 8018 7256 8024 7268
rect 7699 7228 8024 7256
rect 7699 7225 7711 7228
rect 7653 7219 7711 7225
rect 8018 7216 8024 7228
rect 8076 7216 8082 7268
rect 8128 7256 8156 7296
rect 8294 7284 8300 7296
rect 8352 7284 8358 7336
rect 8386 7284 8392 7336
rect 8444 7324 8450 7336
rect 8570 7333 8576 7336
rect 8553 7327 8576 7333
rect 8553 7324 8565 7327
rect 8444 7296 8565 7324
rect 8444 7284 8450 7296
rect 8553 7293 8565 7296
rect 8628 7324 8634 7336
rect 9784 7324 9812 7432
rect 10502 7420 10508 7472
rect 10560 7460 10566 7472
rect 10870 7460 10876 7472
rect 10560 7432 10876 7460
rect 10560 7420 10566 7432
rect 10870 7420 10876 7432
rect 10928 7420 10934 7472
rect 13078 7460 13084 7472
rect 12912 7432 13084 7460
rect 10965 7395 11023 7401
rect 10965 7361 10977 7395
rect 11011 7392 11023 7395
rect 11054 7392 11060 7404
rect 11011 7364 11060 7392
rect 11011 7361 11023 7364
rect 10965 7355 11023 7361
rect 11054 7352 11060 7364
rect 11112 7352 11118 7404
rect 11790 7392 11796 7404
rect 11751 7364 11796 7392
rect 11790 7352 11796 7364
rect 11848 7352 11854 7404
rect 11882 7352 11888 7404
rect 11940 7392 11946 7404
rect 12912 7401 12940 7432
rect 13078 7420 13084 7432
rect 13136 7420 13142 7472
rect 14734 7420 14740 7472
rect 14792 7460 14798 7472
rect 15010 7460 15016 7472
rect 14792 7432 15016 7460
rect 14792 7420 14798 7432
rect 15010 7420 15016 7432
rect 15068 7420 15074 7472
rect 12897 7395 12955 7401
rect 11940 7364 11985 7392
rect 11940 7352 11946 7364
rect 12897 7361 12909 7395
rect 12943 7361 12955 7395
rect 12897 7355 12955 7361
rect 12989 7395 13047 7401
rect 12989 7361 13001 7395
rect 13035 7392 13047 7395
rect 13170 7392 13176 7404
rect 13035 7364 13176 7392
rect 13035 7361 13047 7364
rect 12989 7355 13047 7361
rect 13170 7352 13176 7364
rect 13228 7352 13234 7404
rect 13538 7352 13544 7404
rect 13596 7392 13602 7404
rect 13725 7395 13783 7401
rect 13725 7392 13737 7395
rect 13596 7364 13737 7392
rect 13596 7352 13602 7364
rect 13725 7361 13737 7364
rect 13771 7361 13783 7395
rect 13725 7355 13783 7361
rect 14918 7352 14924 7404
rect 14976 7392 14982 7404
rect 16117 7395 16175 7401
rect 16117 7392 16129 7395
rect 14976 7364 16129 7392
rect 14976 7352 14982 7364
rect 16117 7361 16129 7364
rect 16163 7392 16175 7395
rect 16482 7392 16488 7404
rect 16163 7364 16488 7392
rect 16163 7361 16175 7364
rect 16117 7355 16175 7361
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7392 17187 7395
rect 17494 7392 17500 7404
rect 17175 7364 17500 7392
rect 17175 7361 17187 7364
rect 17129 7355 17187 7361
rect 17494 7352 17500 7364
rect 17552 7352 17558 7404
rect 12805 7327 12863 7333
rect 8628 7296 8701 7324
rect 9232 7296 9812 7324
rect 9876 7296 12572 7324
rect 8553 7287 8576 7293
rect 8570 7284 8576 7287
rect 8628 7284 8634 7296
rect 9232 7256 9260 7296
rect 9876 7256 9904 7296
rect 8128 7228 9260 7256
rect 9324 7228 9904 7256
rect 10689 7259 10747 7265
rect 9324 7188 9352 7228
rect 10689 7225 10701 7259
rect 10735 7256 10747 7259
rect 11238 7256 11244 7268
rect 10735 7228 11244 7256
rect 10735 7225 10747 7228
rect 10689 7219 10747 7225
rect 11238 7216 11244 7228
rect 11296 7216 11302 7268
rect 11701 7259 11759 7265
rect 11701 7225 11713 7259
rect 11747 7256 11759 7259
rect 11747 7228 12480 7256
rect 11747 7225 11759 7228
rect 11701 7219 11759 7225
rect 7392 7160 9352 7188
rect 9674 7148 9680 7200
rect 9732 7188 9738 7200
rect 12452 7197 12480 7228
rect 10321 7191 10379 7197
rect 10321 7188 10333 7191
rect 9732 7160 10333 7188
rect 9732 7148 9738 7160
rect 10321 7157 10333 7160
rect 10367 7157 10379 7191
rect 10321 7151 10379 7157
rect 10781 7191 10839 7197
rect 10781 7157 10793 7191
rect 10827 7188 10839 7191
rect 11333 7191 11391 7197
rect 11333 7188 11345 7191
rect 10827 7160 11345 7188
rect 10827 7157 10839 7160
rect 10781 7151 10839 7157
rect 11333 7157 11345 7160
rect 11379 7157 11391 7191
rect 11333 7151 11391 7157
rect 12437 7191 12495 7197
rect 12437 7157 12449 7191
rect 12483 7157 12495 7191
rect 12544 7188 12572 7296
rect 12805 7293 12817 7327
rect 12851 7324 12863 7327
rect 13262 7324 13268 7336
rect 12851 7296 13268 7324
rect 12851 7293 12863 7296
rect 12805 7287 12863 7293
rect 13262 7284 13268 7296
rect 13320 7284 13326 7336
rect 13992 7327 14050 7333
rect 13992 7293 14004 7327
rect 14038 7324 14050 7327
rect 14936 7324 14964 7352
rect 14038 7296 14964 7324
rect 14038 7293 14050 7296
rect 13992 7287 14050 7293
rect 15010 7284 15016 7336
rect 15068 7324 15074 7336
rect 16390 7324 16396 7336
rect 15068 7296 16396 7324
rect 15068 7284 15074 7296
rect 16390 7284 16396 7296
rect 16448 7284 16454 7336
rect 17218 7284 17224 7336
rect 17276 7324 17282 7336
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 17276 7296 18061 7324
rect 17276 7284 17282 7296
rect 18049 7293 18061 7296
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 12618 7216 12624 7268
rect 12676 7256 12682 7268
rect 16666 7256 16672 7268
rect 12676 7228 16672 7256
rect 12676 7216 12682 7228
rect 16666 7216 16672 7228
rect 16724 7216 16730 7268
rect 16853 7259 16911 7265
rect 16853 7225 16865 7259
rect 16899 7256 16911 7259
rect 17497 7259 17555 7265
rect 17497 7256 17509 7259
rect 16899 7228 17509 7256
rect 16899 7225 16911 7228
rect 16853 7219 16911 7225
rect 17497 7225 17509 7228
rect 17543 7225 17555 7259
rect 17497 7219 17555 7225
rect 15010 7188 15016 7200
rect 12544 7160 15016 7188
rect 12437 7151 12495 7157
rect 15010 7148 15016 7160
rect 15068 7148 15074 7200
rect 15105 7191 15163 7197
rect 15105 7157 15117 7191
rect 15151 7188 15163 7191
rect 15194 7188 15200 7200
rect 15151 7160 15200 7188
rect 15151 7157 15163 7160
rect 15105 7151 15163 7157
rect 15194 7148 15200 7160
rect 15252 7148 15258 7200
rect 15470 7188 15476 7200
rect 15431 7160 15476 7188
rect 15470 7148 15476 7160
rect 15528 7148 15534 7200
rect 15654 7148 15660 7200
rect 15712 7188 15718 7200
rect 15841 7191 15899 7197
rect 15841 7188 15853 7191
rect 15712 7160 15853 7188
rect 15712 7148 15718 7160
rect 15841 7157 15853 7160
rect 15887 7157 15899 7191
rect 15841 7151 15899 7157
rect 15933 7191 15991 7197
rect 15933 7157 15945 7191
rect 15979 7188 15991 7191
rect 16114 7188 16120 7200
rect 15979 7160 16120 7188
rect 15979 7157 15991 7160
rect 15933 7151 15991 7157
rect 16114 7148 16120 7160
rect 16172 7148 16178 7200
rect 16482 7188 16488 7200
rect 16443 7160 16488 7188
rect 16482 7148 16488 7160
rect 16540 7148 16546 7200
rect 16758 7148 16764 7200
rect 16816 7188 16822 7200
rect 16945 7191 17003 7197
rect 16945 7188 16957 7191
rect 16816 7160 16957 7188
rect 16816 7148 16822 7160
rect 16945 7157 16957 7160
rect 16991 7157 17003 7191
rect 16945 7151 17003 7157
rect 17678 7148 17684 7200
rect 17736 7188 17742 7200
rect 18233 7191 18291 7197
rect 18233 7188 18245 7191
rect 17736 7160 18245 7188
rect 17736 7148 17742 7160
rect 18233 7157 18245 7160
rect 18279 7157 18291 7191
rect 18233 7151 18291 7157
rect 1104 7098 18860 7120
rect 1104 7046 6912 7098
rect 6964 7046 6976 7098
rect 7028 7046 7040 7098
rect 7092 7046 7104 7098
rect 7156 7046 12843 7098
rect 12895 7046 12907 7098
rect 12959 7046 12971 7098
rect 13023 7046 13035 7098
rect 13087 7046 18860 7098
rect 1104 7024 18860 7046
rect 3510 6984 3516 6996
rect 3471 6956 3516 6984
rect 3510 6944 3516 6956
rect 3568 6944 3574 6996
rect 5166 6944 5172 6996
rect 5224 6984 5230 6996
rect 5445 6987 5503 6993
rect 5445 6984 5457 6987
rect 5224 6956 5457 6984
rect 5224 6944 5230 6956
rect 5445 6953 5457 6956
rect 5491 6953 5503 6987
rect 5445 6947 5503 6953
rect 5994 6944 6000 6996
rect 6052 6984 6058 6996
rect 6273 6987 6331 6993
rect 6273 6984 6285 6987
rect 6052 6956 6285 6984
rect 6052 6944 6058 6956
rect 6273 6953 6285 6956
rect 6319 6953 6331 6987
rect 6273 6947 6331 6953
rect 6564 6956 7420 6984
rect 3712 6888 4476 6916
rect 1673 6851 1731 6857
rect 1673 6817 1685 6851
rect 1719 6817 1731 6851
rect 2222 6848 2228 6860
rect 2183 6820 2228 6848
rect 1673 6811 1731 6817
rect 1688 6780 1716 6811
rect 2222 6808 2228 6820
rect 2280 6808 2286 6860
rect 2777 6851 2835 6857
rect 2777 6817 2789 6851
rect 2823 6848 2835 6851
rect 3237 6851 3295 6857
rect 3237 6848 3249 6851
rect 2823 6820 3249 6848
rect 2823 6817 2835 6820
rect 2777 6811 2835 6817
rect 3237 6817 3249 6820
rect 3283 6817 3295 6851
rect 3237 6811 3295 6817
rect 3329 6851 3387 6857
rect 3329 6817 3341 6851
rect 3375 6848 3387 6851
rect 3712 6848 3740 6888
rect 3375 6820 3740 6848
rect 3375 6817 3387 6820
rect 3329 6811 3387 6817
rect 3786 6808 3792 6860
rect 3844 6848 3850 6860
rect 4321 6851 4379 6857
rect 4321 6848 4333 6851
rect 3844 6820 4333 6848
rect 3844 6808 3850 6820
rect 4321 6817 4333 6820
rect 4367 6817 4379 6851
rect 4448 6848 4476 6888
rect 4982 6876 4988 6928
rect 5040 6916 5046 6928
rect 6564 6916 6592 6956
rect 5040 6888 6592 6916
rect 6641 6919 6699 6925
rect 5040 6876 5046 6888
rect 6641 6885 6653 6919
rect 6687 6916 6699 6919
rect 7392 6916 7420 6956
rect 7742 6944 7748 6996
rect 7800 6984 7806 6996
rect 8021 6987 8079 6993
rect 8021 6984 8033 6987
rect 7800 6956 8033 6984
rect 7800 6944 7806 6956
rect 8021 6953 8033 6956
rect 8067 6953 8079 6987
rect 8021 6947 8079 6953
rect 8389 6987 8447 6993
rect 8389 6953 8401 6987
rect 8435 6984 8447 6987
rect 8754 6984 8760 6996
rect 8435 6956 8760 6984
rect 8435 6953 8447 6956
rect 8389 6947 8447 6953
rect 8754 6944 8760 6956
rect 8812 6944 8818 6996
rect 11609 6987 11667 6993
rect 11609 6953 11621 6987
rect 11655 6984 11667 6987
rect 11882 6984 11888 6996
rect 11655 6956 11888 6984
rect 11655 6953 11667 6956
rect 11609 6947 11667 6953
rect 11882 6944 11888 6956
rect 11940 6944 11946 6996
rect 12437 6987 12495 6993
rect 12437 6953 12449 6987
rect 12483 6984 12495 6987
rect 12618 6984 12624 6996
rect 12483 6956 12624 6984
rect 12483 6953 12495 6956
rect 12437 6947 12495 6953
rect 12618 6944 12624 6956
rect 12676 6944 12682 6996
rect 13262 6944 13268 6996
rect 13320 6984 13326 6996
rect 13630 6984 13636 6996
rect 13320 6956 13636 6984
rect 13320 6944 13326 6956
rect 13630 6944 13636 6956
rect 13688 6984 13694 6996
rect 14553 6987 14611 6993
rect 13688 6956 14412 6984
rect 13688 6944 13694 6956
rect 14274 6916 14280 6928
rect 6687 6888 7328 6916
rect 7392 6888 14280 6916
rect 6687 6885 6699 6888
rect 6641 6879 6699 6885
rect 7300 6857 7328 6888
rect 14274 6876 14280 6888
rect 14332 6876 14338 6928
rect 14384 6916 14412 6956
rect 14553 6953 14565 6987
rect 14599 6984 14611 6987
rect 16482 6984 16488 6996
rect 14599 6956 16488 6984
rect 14599 6953 14611 6956
rect 14553 6947 14611 6953
rect 16482 6944 16488 6956
rect 16540 6944 16546 6996
rect 16574 6944 16580 6996
rect 16632 6984 16638 6996
rect 16669 6987 16727 6993
rect 16669 6984 16681 6987
rect 16632 6956 16681 6984
rect 16632 6944 16638 6956
rect 16669 6953 16681 6956
rect 16715 6953 16727 6987
rect 17310 6984 17316 6996
rect 17271 6956 17316 6984
rect 16669 6947 16727 6953
rect 17310 6944 17316 6956
rect 17368 6944 17374 6996
rect 17402 6916 17408 6928
rect 14384 6888 17408 6916
rect 17402 6876 17408 6888
rect 17460 6876 17466 6928
rect 6733 6851 6791 6857
rect 6733 6848 6745 6851
rect 4448 6820 6745 6848
rect 4321 6811 4379 6817
rect 6733 6817 6745 6820
rect 6779 6848 6791 6851
rect 7285 6851 7343 6857
rect 6779 6820 7236 6848
rect 6779 6817 6791 6820
rect 6733 6811 6791 6817
rect 3050 6780 3056 6792
rect 1688 6752 3056 6780
rect 3050 6740 3056 6752
rect 3108 6740 3114 6792
rect 4062 6780 4068 6792
rect 3160 6752 4068 6780
rect 2958 6712 2964 6724
rect 2919 6684 2964 6712
rect 2958 6672 2964 6684
rect 3016 6672 3022 6724
rect 1854 6644 1860 6656
rect 1815 6616 1860 6644
rect 1854 6604 1860 6616
rect 1912 6604 1918 6656
rect 2406 6644 2412 6656
rect 2367 6616 2412 6644
rect 2406 6604 2412 6616
rect 2464 6604 2470 6656
rect 2498 6604 2504 6656
rect 2556 6644 2562 6656
rect 3160 6644 3188 6752
rect 4062 6740 4068 6752
rect 4120 6740 4126 6792
rect 5994 6740 6000 6792
rect 6052 6780 6058 6792
rect 6825 6783 6883 6789
rect 6825 6780 6837 6783
rect 6052 6752 6837 6780
rect 6052 6740 6058 6752
rect 6825 6749 6837 6752
rect 6871 6749 6883 6783
rect 7208 6780 7236 6820
rect 7285 6817 7297 6851
rect 7331 6817 7343 6851
rect 10318 6848 10324 6860
rect 7285 6811 7343 6817
rect 8496 6820 10324 6848
rect 8496 6792 8524 6820
rect 10318 6808 10324 6820
rect 10376 6808 10382 6860
rect 10496 6851 10554 6857
rect 10496 6817 10508 6851
rect 10542 6848 10554 6851
rect 13170 6848 13176 6860
rect 10542 6820 13176 6848
rect 10542 6817 10554 6820
rect 10496 6811 10554 6817
rect 8110 6780 8116 6792
rect 7208 6752 8116 6780
rect 6825 6743 6883 6749
rect 8110 6740 8116 6752
rect 8168 6740 8174 6792
rect 8478 6780 8484 6792
rect 8439 6752 8484 6780
rect 8478 6740 8484 6752
rect 8536 6740 8542 6792
rect 8570 6740 8576 6792
rect 8628 6780 8634 6792
rect 8628 6752 8673 6780
rect 8628 6740 8634 6752
rect 8754 6740 8760 6792
rect 8812 6780 8818 6792
rect 9033 6783 9091 6789
rect 9033 6780 9045 6783
rect 8812 6752 9045 6780
rect 8812 6740 8818 6752
rect 9033 6749 9045 6752
rect 9079 6749 9091 6783
rect 9033 6743 9091 6749
rect 9122 6740 9128 6792
rect 9180 6780 9186 6792
rect 10226 6780 10232 6792
rect 9180 6752 10232 6780
rect 9180 6740 9186 6752
rect 10226 6740 10232 6752
rect 10284 6740 10290 6792
rect 12434 6740 12440 6792
rect 12492 6780 12498 6792
rect 12636 6789 12664 6820
rect 13170 6808 13176 6820
rect 13228 6808 13234 6860
rect 13446 6848 13452 6860
rect 13407 6820 13452 6848
rect 13446 6808 13452 6820
rect 13504 6808 13510 6860
rect 13541 6851 13599 6857
rect 13541 6817 13553 6851
rect 13587 6848 13599 6851
rect 14090 6848 14096 6860
rect 13587 6820 14096 6848
rect 13587 6817 13599 6820
rect 13541 6811 13599 6817
rect 12529 6783 12587 6789
rect 12529 6780 12541 6783
rect 12492 6752 12541 6780
rect 12492 6740 12498 6752
rect 12529 6749 12541 6752
rect 12575 6749 12587 6783
rect 12529 6743 12587 6749
rect 12621 6783 12679 6789
rect 12621 6749 12633 6783
rect 12667 6749 12679 6783
rect 13556 6780 13584 6811
rect 14090 6808 14096 6820
rect 14148 6808 14154 6860
rect 15378 6848 15384 6860
rect 14200 6820 15384 6848
rect 12621 6743 12679 6749
rect 12820 6752 13584 6780
rect 13633 6783 13691 6789
rect 8386 6672 8392 6724
rect 8444 6712 8450 6724
rect 8938 6712 8944 6724
rect 8444 6684 8944 6712
rect 8444 6672 8450 6684
rect 8938 6672 8944 6684
rect 8996 6672 9002 6724
rect 12820 6712 12848 6752
rect 13633 6749 13645 6783
rect 13679 6749 13691 6783
rect 13633 6743 13691 6749
rect 11164 6684 12848 6712
rect 2556 6616 3188 6644
rect 3237 6647 3295 6653
rect 2556 6604 2562 6616
rect 3237 6613 3249 6647
rect 3283 6644 3295 6647
rect 11164 6644 11192 6684
rect 13170 6672 13176 6724
rect 13228 6712 13234 6724
rect 13648 6712 13676 6743
rect 14200 6721 14228 6820
rect 15378 6808 15384 6820
rect 15436 6808 15442 6860
rect 15556 6851 15614 6857
rect 15556 6817 15568 6851
rect 15602 6848 15614 6851
rect 16758 6848 16764 6860
rect 15602 6820 16764 6848
rect 15602 6817 15614 6820
rect 15556 6811 15614 6817
rect 16758 6808 16764 6820
rect 16816 6808 16822 6860
rect 17954 6848 17960 6860
rect 17915 6820 17960 6848
rect 17954 6808 17960 6820
rect 18012 6808 18018 6860
rect 14645 6783 14703 6789
rect 14645 6749 14657 6783
rect 14691 6749 14703 6783
rect 14645 6743 14703 6749
rect 14829 6783 14887 6789
rect 14829 6749 14841 6783
rect 14875 6780 14887 6783
rect 14918 6780 14924 6792
rect 14875 6752 14924 6780
rect 14875 6749 14887 6752
rect 14829 6743 14887 6749
rect 13228 6684 13676 6712
rect 14185 6715 14243 6721
rect 13228 6672 13234 6684
rect 14185 6681 14197 6715
rect 14231 6681 14243 6715
rect 14185 6675 14243 6681
rect 3283 6616 11192 6644
rect 3283 6613 3295 6616
rect 3237 6607 3295 6613
rect 11790 6604 11796 6656
rect 11848 6644 11854 6656
rect 12069 6647 12127 6653
rect 12069 6644 12081 6647
rect 11848 6616 12081 6644
rect 11848 6604 11854 6616
rect 12069 6613 12081 6616
rect 12115 6613 12127 6647
rect 12069 6607 12127 6613
rect 12158 6604 12164 6656
rect 12216 6644 12222 6656
rect 13081 6647 13139 6653
rect 13081 6644 13093 6647
rect 12216 6616 13093 6644
rect 12216 6604 12222 6616
rect 13081 6613 13093 6616
rect 13127 6613 13139 6647
rect 14660 6644 14688 6743
rect 14918 6740 14924 6752
rect 14976 6740 14982 6792
rect 15010 6740 15016 6792
rect 15068 6780 15074 6792
rect 15289 6783 15347 6789
rect 15289 6780 15301 6783
rect 15068 6752 15301 6780
rect 15068 6740 15074 6752
rect 15289 6749 15301 6752
rect 15335 6749 15347 6783
rect 15289 6743 15347 6749
rect 16482 6740 16488 6792
rect 16540 6780 16546 6792
rect 17405 6783 17463 6789
rect 17405 6780 17417 6783
rect 16540 6752 17417 6780
rect 16540 6740 16546 6752
rect 17405 6749 17417 6752
rect 17451 6749 17463 6783
rect 17405 6743 17463 6749
rect 17494 6740 17500 6792
rect 17552 6780 17558 6792
rect 17552 6752 17597 6780
rect 17552 6740 17558 6752
rect 16945 6715 17003 6721
rect 16945 6712 16957 6715
rect 16224 6684 16957 6712
rect 16224 6644 16252 6684
rect 16945 6681 16957 6684
rect 16991 6681 17003 6715
rect 16945 6675 17003 6681
rect 18138 6644 18144 6656
rect 14660 6616 16252 6644
rect 18099 6616 18144 6644
rect 13081 6607 13139 6613
rect 18138 6604 18144 6616
rect 18196 6604 18202 6656
rect 1104 6554 18860 6576
rect 1104 6502 3947 6554
rect 3999 6502 4011 6554
rect 4063 6502 4075 6554
rect 4127 6502 4139 6554
rect 4191 6502 9878 6554
rect 9930 6502 9942 6554
rect 9994 6502 10006 6554
rect 10058 6502 10070 6554
rect 10122 6502 15808 6554
rect 15860 6502 15872 6554
rect 15924 6502 15936 6554
rect 15988 6502 16000 6554
rect 16052 6502 18860 6554
rect 1104 6480 18860 6502
rect 3050 6400 3056 6452
rect 3108 6440 3114 6452
rect 4614 6440 4620 6452
rect 3108 6412 4620 6440
rect 3108 6400 3114 6412
rect 4614 6400 4620 6412
rect 4672 6400 4678 6452
rect 4724 6412 5672 6440
rect 4154 6332 4160 6384
rect 4212 6372 4218 6384
rect 4338 6372 4344 6384
rect 4212 6344 4344 6372
rect 4212 6332 4218 6344
rect 4338 6332 4344 6344
rect 4396 6332 4402 6384
rect 4522 6332 4528 6384
rect 4580 6372 4586 6384
rect 4724 6372 4752 6412
rect 4580 6344 4752 6372
rect 5644 6372 5672 6412
rect 6086 6400 6092 6452
rect 6144 6440 6150 6452
rect 6825 6443 6883 6449
rect 6825 6440 6837 6443
rect 6144 6412 6837 6440
rect 6144 6400 6150 6412
rect 6825 6409 6837 6412
rect 6871 6409 6883 6443
rect 6825 6403 6883 6409
rect 7190 6400 7196 6452
rect 7248 6440 7254 6452
rect 7374 6440 7380 6452
rect 7248 6412 7380 6440
rect 7248 6400 7254 6412
rect 7374 6400 7380 6412
rect 7432 6400 7438 6452
rect 8018 6440 8024 6452
rect 7979 6412 8024 6440
rect 8018 6400 8024 6412
rect 8076 6400 8082 6452
rect 8110 6400 8116 6452
rect 8168 6440 8174 6452
rect 11146 6440 11152 6452
rect 8168 6412 11152 6440
rect 8168 6400 8174 6412
rect 11146 6400 11152 6412
rect 11204 6400 11210 6452
rect 11238 6400 11244 6452
rect 11296 6440 11302 6452
rect 11333 6443 11391 6449
rect 11333 6440 11345 6443
rect 11296 6412 11345 6440
rect 11296 6400 11302 6412
rect 11333 6409 11345 6412
rect 11379 6409 11391 6443
rect 15010 6440 15016 6452
rect 11333 6403 11391 6409
rect 14108 6412 15016 6440
rect 8386 6372 8392 6384
rect 5644 6344 8392 6372
rect 4580 6332 4586 6344
rect 8386 6332 8392 6344
rect 8444 6332 8450 6384
rect 8496 6344 9076 6372
rect 3988 6276 4844 6304
rect 1670 6236 1676 6248
rect 1631 6208 1676 6236
rect 1670 6196 1676 6208
rect 1728 6196 1734 6248
rect 2409 6239 2467 6245
rect 2409 6205 2421 6239
rect 2455 6236 2467 6239
rect 2498 6236 2504 6248
rect 2455 6208 2504 6236
rect 2455 6205 2467 6208
rect 2409 6199 2467 6205
rect 2498 6196 2504 6208
rect 2556 6196 2562 6248
rect 3988 6236 4016 6276
rect 2608 6208 4016 6236
rect 4065 6239 4123 6245
rect 2222 6128 2228 6180
rect 2280 6168 2286 6180
rect 2608 6168 2636 6208
rect 4065 6205 4077 6239
rect 4111 6236 4123 6239
rect 4154 6236 4160 6248
rect 4111 6208 4160 6236
rect 4111 6205 4123 6208
rect 4065 6199 4123 6205
rect 4154 6196 4160 6208
rect 4212 6196 4218 6248
rect 4246 6196 4252 6248
rect 4304 6236 4310 6248
rect 4709 6239 4767 6245
rect 4709 6236 4721 6239
rect 4304 6208 4721 6236
rect 4304 6196 4310 6208
rect 4709 6205 4721 6208
rect 4755 6205 4767 6239
rect 4816 6236 4844 6276
rect 5994 6264 6000 6316
rect 6052 6304 6058 6316
rect 8496 6313 8524 6344
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 6052 6276 7389 6304
rect 6052 6264 6058 6276
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 8481 6307 8539 6313
rect 8481 6304 8493 6307
rect 7377 6267 7435 6273
rect 7852 6276 8493 6304
rect 7852 6236 7880 6276
rect 8481 6273 8493 6276
rect 8527 6273 8539 6307
rect 8481 6267 8539 6273
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 8628 6276 8673 6304
rect 8628 6264 8634 6276
rect 4816 6208 7880 6236
rect 8389 6239 8447 6245
rect 4709 6199 4767 6205
rect 8389 6205 8401 6239
rect 8435 6236 8447 6239
rect 8754 6236 8760 6248
rect 8435 6208 8760 6236
rect 8435 6205 8447 6208
rect 8389 6199 8447 6205
rect 8754 6196 8760 6208
rect 8812 6196 8818 6248
rect 2280 6140 2636 6168
rect 2676 6171 2734 6177
rect 2280 6128 2286 6140
rect 2676 6137 2688 6171
rect 2722 6168 2734 6171
rect 3050 6168 3056 6180
rect 2722 6140 3056 6168
rect 2722 6137 2734 6140
rect 2676 6131 2734 6137
rect 3050 6128 3056 6140
rect 3108 6128 3114 6180
rect 3326 6128 3332 6180
rect 3384 6168 3390 6180
rect 3384 6140 4292 6168
rect 3384 6128 3390 6140
rect 1394 6060 1400 6112
rect 1452 6100 1458 6112
rect 1857 6103 1915 6109
rect 1857 6100 1869 6103
rect 1452 6072 1869 6100
rect 1452 6060 1458 6072
rect 1857 6069 1869 6072
rect 1903 6069 1915 6103
rect 1857 6063 1915 6069
rect 3142 6060 3148 6112
rect 3200 6100 3206 6112
rect 3786 6100 3792 6112
rect 3200 6072 3792 6100
rect 3200 6060 3206 6072
rect 3786 6060 3792 6072
rect 3844 6060 3850 6112
rect 4264 6109 4292 6140
rect 4614 6128 4620 6180
rect 4672 6168 4678 6180
rect 4954 6171 5012 6177
rect 4954 6168 4966 6171
rect 4672 6140 4966 6168
rect 4672 6128 4678 6140
rect 4954 6137 4966 6140
rect 5000 6168 5012 6171
rect 5994 6168 6000 6180
rect 5000 6140 6000 6168
rect 5000 6137 5012 6140
rect 4954 6131 5012 6137
rect 5994 6128 6000 6140
rect 6052 6128 6058 6180
rect 7190 6168 7196 6180
rect 7151 6140 7196 6168
rect 7190 6128 7196 6140
rect 7248 6128 7254 6180
rect 7374 6128 7380 6180
rect 7432 6168 7438 6180
rect 9048 6168 9076 6344
rect 9122 6332 9128 6384
rect 9180 6332 9186 6384
rect 13446 6372 13452 6384
rect 11624 6344 13452 6372
rect 9140 6245 9168 6332
rect 10873 6307 10931 6313
rect 10873 6273 10885 6307
rect 10919 6304 10931 6307
rect 11624 6304 11652 6344
rect 13446 6332 13452 6344
rect 13504 6332 13510 6384
rect 11790 6304 11796 6316
rect 10919 6276 11652 6304
rect 11751 6276 11796 6304
rect 10919 6273 10931 6276
rect 10873 6267 10931 6273
rect 11790 6264 11796 6276
rect 11848 6264 11854 6316
rect 11882 6264 11888 6316
rect 11940 6304 11946 6316
rect 11940 6276 11985 6304
rect 11940 6264 11946 6276
rect 12342 6264 12348 6316
rect 12400 6304 12406 6316
rect 12529 6307 12587 6313
rect 12529 6304 12541 6307
rect 12400 6276 12541 6304
rect 12400 6264 12406 6276
rect 12529 6273 12541 6276
rect 12575 6273 12587 6307
rect 13170 6304 13176 6316
rect 13131 6276 13176 6304
rect 12529 6267 12587 6273
rect 13170 6264 13176 6276
rect 13228 6264 13234 6316
rect 14108 6313 14136 6412
rect 15010 6400 15016 6412
rect 15068 6400 15074 6452
rect 16114 6440 16120 6452
rect 16075 6412 16120 6440
rect 16114 6400 16120 6412
rect 16172 6400 16178 6452
rect 17589 6443 17647 6449
rect 17589 6409 17601 6443
rect 17635 6440 17647 6443
rect 17954 6440 17960 6452
rect 17635 6412 17960 6440
rect 17635 6409 17647 6412
rect 17589 6403 17647 6409
rect 17954 6400 17960 6412
rect 18012 6400 18018 6452
rect 15473 6375 15531 6381
rect 15473 6341 15485 6375
rect 15519 6341 15531 6375
rect 15473 6335 15531 6341
rect 14093 6307 14151 6313
rect 14093 6304 14105 6307
rect 13372 6276 14105 6304
rect 9125 6239 9183 6245
rect 9125 6205 9137 6239
rect 9171 6205 9183 6239
rect 11514 6236 11520 6248
rect 9125 6199 9183 6205
rect 9324 6208 11520 6236
rect 9324 6168 9352 6208
rect 11514 6196 11520 6208
rect 11572 6196 11578 6248
rect 11701 6239 11759 6245
rect 11701 6205 11713 6239
rect 11747 6236 11759 6239
rect 12158 6236 12164 6248
rect 11747 6208 12164 6236
rect 11747 6205 11759 6208
rect 11701 6199 11759 6205
rect 12158 6196 12164 6208
rect 12216 6196 12222 6248
rect 7432 6140 8616 6168
rect 9048 6140 9352 6168
rect 9392 6171 9450 6177
rect 7432 6128 7438 6140
rect 4249 6103 4307 6109
rect 4249 6069 4261 6103
rect 4295 6069 4307 6103
rect 4249 6063 4307 6069
rect 4338 6060 4344 6112
rect 4396 6100 4402 6112
rect 6089 6103 6147 6109
rect 6089 6100 6101 6103
rect 4396 6072 6101 6100
rect 4396 6060 4402 6072
rect 6089 6069 6101 6072
rect 6135 6100 6147 6103
rect 6178 6100 6184 6112
rect 6135 6072 6184 6100
rect 6135 6069 6147 6072
rect 6089 6063 6147 6069
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 7285 6103 7343 6109
rect 7285 6069 7297 6103
rect 7331 6100 7343 6103
rect 7466 6100 7472 6112
rect 7331 6072 7472 6100
rect 7331 6069 7343 6072
rect 7285 6063 7343 6069
rect 7466 6060 7472 6072
rect 7524 6060 7530 6112
rect 8588 6100 8616 6140
rect 9392 6137 9404 6171
rect 9438 6168 9450 6171
rect 10962 6168 10968 6180
rect 9438 6140 10968 6168
rect 9438 6137 9450 6140
rect 9392 6131 9450 6137
rect 10962 6128 10968 6140
rect 11020 6128 11026 6180
rect 12342 6168 12348 6180
rect 11072 6140 12348 6168
rect 10505 6103 10563 6109
rect 10505 6100 10517 6103
rect 8588 6072 10517 6100
rect 10505 6069 10517 6072
rect 10551 6069 10563 6103
rect 10505 6063 10563 6069
rect 10594 6060 10600 6112
rect 10652 6100 10658 6112
rect 11072 6100 11100 6140
rect 12342 6128 12348 6140
rect 12400 6168 12406 6180
rect 12621 6171 12679 6177
rect 12621 6168 12633 6171
rect 12400 6140 12633 6168
rect 12400 6128 12406 6140
rect 12621 6137 12633 6140
rect 12667 6137 12679 6171
rect 12621 6131 12679 6137
rect 12710 6128 12716 6180
rect 12768 6168 12774 6180
rect 13372 6168 13400 6276
rect 14093 6273 14105 6276
rect 14139 6273 14151 6307
rect 15488 6304 15516 6335
rect 16390 6332 16396 6384
rect 16448 6372 16454 6384
rect 17862 6372 17868 6384
rect 16448 6344 17868 6372
rect 16448 6332 16454 6344
rect 17862 6332 17868 6344
rect 17920 6332 17926 6384
rect 16758 6304 16764 6316
rect 15488 6276 16764 6304
rect 14093 6267 14151 6273
rect 16758 6264 16764 6276
rect 16816 6304 16822 6316
rect 17494 6304 17500 6316
rect 16816 6276 17500 6304
rect 16816 6264 16822 6276
rect 17494 6264 17500 6276
rect 17552 6264 17558 6316
rect 15930 6196 15936 6248
rect 15988 6236 15994 6248
rect 16482 6236 16488 6248
rect 15988 6208 16488 6236
rect 15988 6196 15994 6208
rect 16482 6196 16488 6208
rect 16540 6196 16546 6248
rect 16666 6196 16672 6248
rect 16724 6236 16730 6248
rect 17405 6239 17463 6245
rect 17405 6236 17417 6239
rect 16724 6208 17417 6236
rect 16724 6196 16730 6208
rect 17405 6205 17417 6208
rect 17451 6205 17463 6239
rect 17405 6199 17463 6205
rect 18049 6239 18107 6245
rect 18049 6205 18061 6239
rect 18095 6236 18107 6239
rect 18506 6236 18512 6248
rect 18095 6208 18512 6236
rect 18095 6205 18107 6208
rect 18049 6199 18107 6205
rect 18506 6196 18512 6208
rect 18564 6196 18570 6248
rect 12768 6140 13400 6168
rect 12768 6128 12774 6140
rect 14274 6128 14280 6180
rect 14332 6177 14338 6180
rect 14332 6171 14396 6177
rect 14332 6137 14350 6171
rect 14384 6168 14396 6171
rect 17218 6168 17224 6180
rect 14384 6140 17224 6168
rect 14384 6137 14396 6140
rect 14332 6131 14396 6137
rect 14332 6128 14338 6131
rect 17218 6128 17224 6140
rect 17276 6128 17282 6180
rect 16482 6100 16488 6112
rect 10652 6072 11100 6100
rect 16443 6072 16488 6100
rect 10652 6060 10658 6072
rect 16482 6060 16488 6072
rect 16540 6060 16546 6112
rect 16574 6060 16580 6112
rect 16632 6100 16638 6112
rect 18230 6100 18236 6112
rect 16632 6072 16677 6100
rect 18191 6072 18236 6100
rect 16632 6060 16638 6072
rect 18230 6060 18236 6072
rect 18288 6060 18294 6112
rect 1104 6010 18860 6032
rect 1104 5958 6912 6010
rect 6964 5958 6976 6010
rect 7028 5958 7040 6010
rect 7092 5958 7104 6010
rect 7156 5958 12843 6010
rect 12895 5958 12907 6010
rect 12959 5958 12971 6010
rect 13023 5958 13035 6010
rect 13087 5958 18860 6010
rect 1104 5936 18860 5958
rect 2409 5899 2467 5905
rect 2409 5865 2421 5899
rect 2455 5896 2467 5899
rect 2961 5899 3019 5905
rect 2961 5896 2973 5899
rect 2455 5868 2973 5896
rect 2455 5865 2467 5868
rect 2409 5859 2467 5865
rect 2961 5865 2973 5868
rect 3007 5865 3019 5899
rect 4433 5899 4491 5905
rect 4433 5896 4445 5899
rect 2961 5859 3019 5865
rect 3160 5868 4445 5896
rect 2866 5788 2872 5840
rect 2924 5828 2930 5840
rect 3160 5828 3188 5868
rect 4433 5865 4445 5868
rect 4479 5865 4491 5899
rect 4433 5859 4491 5865
rect 4525 5899 4583 5905
rect 4525 5865 4537 5899
rect 4571 5896 4583 5899
rect 5997 5899 6055 5905
rect 5997 5896 6009 5899
rect 4571 5868 6009 5896
rect 4571 5865 4583 5868
rect 4525 5859 4583 5865
rect 5997 5865 6009 5868
rect 6043 5865 6055 5899
rect 5997 5859 6055 5865
rect 6549 5899 6607 5905
rect 6549 5865 6561 5899
rect 6595 5865 6607 5899
rect 6549 5859 6607 5865
rect 5626 5828 5632 5840
rect 2924 5800 3188 5828
rect 3252 5800 5632 5828
rect 2924 5788 2930 5800
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5760 1455 5763
rect 2130 5760 2136 5772
rect 1443 5732 2136 5760
rect 1443 5729 1455 5732
rect 1397 5723 1455 5729
rect 2130 5720 2136 5732
rect 2188 5720 2194 5772
rect 2317 5763 2375 5769
rect 2317 5729 2329 5763
rect 2363 5760 2375 5763
rect 3252 5760 3280 5800
rect 5626 5788 5632 5800
rect 5684 5788 5690 5840
rect 6564 5828 6592 5859
rect 7282 5856 7288 5908
rect 7340 5896 7346 5908
rect 7469 5899 7527 5905
rect 7469 5896 7481 5899
rect 7340 5868 7481 5896
rect 7340 5856 7346 5868
rect 7469 5865 7481 5868
rect 7515 5865 7527 5899
rect 7469 5859 7527 5865
rect 7561 5899 7619 5905
rect 7561 5865 7573 5899
rect 7607 5896 7619 5899
rect 7650 5896 7656 5908
rect 7607 5868 7656 5896
rect 7607 5865 7619 5868
rect 7561 5859 7619 5865
rect 7650 5856 7656 5868
rect 7708 5856 7714 5908
rect 10226 5856 10232 5908
rect 10284 5896 10290 5908
rect 10962 5896 10968 5908
rect 10284 5868 10968 5896
rect 10284 5856 10290 5868
rect 10962 5856 10968 5868
rect 11020 5856 11026 5908
rect 11054 5856 11060 5908
rect 11112 5896 11118 5908
rect 12529 5899 12587 5905
rect 12529 5896 12541 5899
rect 11112 5868 12541 5896
rect 11112 5856 11118 5868
rect 12529 5865 12541 5868
rect 12575 5865 12587 5899
rect 14274 5896 14280 5908
rect 14235 5868 14280 5896
rect 12529 5859 12587 5865
rect 11238 5828 11244 5840
rect 5828 5800 6592 5828
rect 6656 5800 11244 5828
rect 2363 5732 3280 5760
rect 3329 5763 3387 5769
rect 2363 5729 2375 5732
rect 2317 5723 2375 5729
rect 3329 5729 3341 5763
rect 3375 5760 3387 5763
rect 3881 5763 3939 5769
rect 3881 5760 3893 5763
rect 3375 5732 3893 5760
rect 3375 5729 3387 5732
rect 3329 5723 3387 5729
rect 3881 5729 3893 5732
rect 3927 5729 3939 5763
rect 3881 5723 3939 5729
rect 4522 5720 4528 5772
rect 4580 5760 4586 5772
rect 4893 5763 4951 5769
rect 4893 5760 4905 5763
rect 4580 5732 4905 5760
rect 4580 5720 4586 5732
rect 4893 5729 4905 5732
rect 4939 5729 4951 5763
rect 4893 5723 4951 5729
rect 5074 5720 5080 5772
rect 5132 5760 5138 5772
rect 5828 5760 5856 5800
rect 5132 5732 5856 5760
rect 5905 5763 5963 5769
rect 5132 5720 5138 5732
rect 5905 5729 5917 5763
rect 5951 5760 5963 5763
rect 6362 5760 6368 5772
rect 5951 5732 6368 5760
rect 5951 5729 5963 5732
rect 5905 5723 5963 5729
rect 6362 5720 6368 5732
rect 6420 5760 6426 5772
rect 6656 5760 6684 5800
rect 11238 5788 11244 5800
rect 11296 5788 11302 5840
rect 11416 5831 11474 5837
rect 11416 5797 11428 5831
rect 11462 5828 11474 5831
rect 11882 5828 11888 5840
rect 11462 5800 11888 5828
rect 11462 5797 11474 5800
rect 11416 5791 11474 5797
rect 11882 5788 11888 5800
rect 11940 5788 11946 5840
rect 12544 5828 12572 5859
rect 14274 5856 14280 5868
rect 14332 5856 14338 5908
rect 15654 5896 15660 5908
rect 15615 5868 15660 5896
rect 15654 5856 15660 5868
rect 15712 5856 15718 5908
rect 16482 5856 16488 5908
rect 16540 5896 16546 5908
rect 16669 5899 16727 5905
rect 16669 5896 16681 5899
rect 16540 5868 16681 5896
rect 16540 5856 16546 5868
rect 16669 5865 16681 5868
rect 16715 5865 16727 5899
rect 16669 5859 16727 5865
rect 17037 5899 17095 5905
rect 17037 5865 17049 5899
rect 17083 5896 17095 5899
rect 18598 5896 18604 5908
rect 17083 5868 18604 5896
rect 17083 5865 17095 5868
rect 17037 5859 17095 5865
rect 18598 5856 18604 5868
rect 18656 5856 18662 5908
rect 13142 5831 13200 5837
rect 13142 5828 13154 5831
rect 12544 5800 13154 5828
rect 13142 5797 13154 5800
rect 13188 5797 13200 5831
rect 16022 5828 16028 5840
rect 15983 5800 16028 5828
rect 13142 5791 13200 5797
rect 16022 5788 16028 5800
rect 16080 5828 16086 5840
rect 18046 5828 18052 5840
rect 16080 5800 18052 5828
rect 16080 5788 16086 5800
rect 18046 5788 18052 5800
rect 18104 5788 18110 5840
rect 6420 5732 6684 5760
rect 6420 5720 6426 5732
rect 6730 5720 6736 5772
rect 6788 5760 6794 5772
rect 6788 5732 6833 5760
rect 6788 5720 6794 5732
rect 9214 5720 9220 5772
rect 9272 5760 9278 5772
rect 9677 5763 9735 5769
rect 9677 5760 9689 5763
rect 9272 5732 9689 5760
rect 9272 5720 9278 5732
rect 9677 5729 9689 5732
rect 9723 5729 9735 5763
rect 9677 5723 9735 5729
rect 10045 5763 10103 5769
rect 10045 5729 10057 5763
rect 10091 5760 10103 5763
rect 10226 5760 10232 5772
rect 10091 5732 10232 5760
rect 10091 5729 10103 5732
rect 10045 5723 10103 5729
rect 10226 5720 10232 5732
rect 10284 5720 10290 5772
rect 10410 5760 10416 5772
rect 10371 5732 10416 5760
rect 10410 5720 10416 5732
rect 10468 5760 10474 5772
rect 10594 5760 10600 5772
rect 10468 5732 10600 5760
rect 10468 5720 10474 5732
rect 10594 5720 10600 5732
rect 10652 5720 10658 5772
rect 10756 5763 10814 5769
rect 10756 5729 10768 5763
rect 10802 5760 10814 5763
rect 10870 5760 10876 5772
rect 10802 5732 10876 5760
rect 10802 5729 10814 5732
rect 10756 5723 10814 5729
rect 10870 5720 10876 5732
rect 10928 5720 10934 5772
rect 10962 5720 10968 5772
rect 11020 5760 11026 5772
rect 11149 5763 11207 5769
rect 11149 5760 11161 5763
rect 11020 5732 11161 5760
rect 11020 5720 11026 5732
rect 11149 5729 11161 5732
rect 11195 5760 11207 5763
rect 12250 5760 12256 5772
rect 11195 5732 12256 5760
rect 11195 5729 11207 5732
rect 11149 5723 11207 5729
rect 12250 5720 12256 5732
rect 12308 5720 12314 5772
rect 14645 5763 14703 5769
rect 14645 5729 14657 5763
rect 14691 5760 14703 5763
rect 16117 5763 16175 5769
rect 14691 5732 16068 5760
rect 14691 5729 14703 5732
rect 14645 5723 14703 5729
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 3142 5692 3148 5704
rect 2639 5664 3148 5692
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 3142 5652 3148 5664
rect 3200 5652 3206 5704
rect 3418 5692 3424 5704
rect 3379 5664 3424 5692
rect 3418 5652 3424 5664
rect 3476 5652 3482 5704
rect 3605 5695 3663 5701
rect 3605 5661 3617 5695
rect 3651 5692 3663 5695
rect 4338 5692 4344 5704
rect 3651 5664 4344 5692
rect 3651 5661 3663 5664
rect 3605 5655 3663 5661
rect 3050 5584 3056 5636
rect 3108 5624 3114 5636
rect 3620 5624 3648 5655
rect 4338 5652 4344 5664
rect 4396 5652 4402 5704
rect 4433 5695 4491 5701
rect 4433 5661 4445 5695
rect 4479 5692 4491 5695
rect 4985 5695 5043 5701
rect 4985 5692 4997 5695
rect 4479 5664 4997 5692
rect 4479 5661 4491 5664
rect 4433 5655 4491 5661
rect 4985 5661 4997 5664
rect 5031 5661 5043 5695
rect 4985 5655 5043 5661
rect 5169 5695 5227 5701
rect 5169 5661 5181 5695
rect 5215 5692 5227 5695
rect 5442 5692 5448 5704
rect 5215 5664 5448 5692
rect 5215 5661 5227 5664
rect 5169 5655 5227 5661
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 5994 5652 6000 5704
rect 6052 5692 6058 5704
rect 6089 5695 6147 5701
rect 6089 5692 6101 5695
rect 6052 5664 6101 5692
rect 6052 5652 6058 5664
rect 6089 5661 6101 5664
rect 6135 5692 6147 5695
rect 6454 5692 6460 5704
rect 6135 5664 6460 5692
rect 6135 5661 6147 5664
rect 6089 5655 6147 5661
rect 6454 5652 6460 5664
rect 6512 5652 6518 5704
rect 7745 5695 7803 5701
rect 7745 5661 7757 5695
rect 7791 5692 7803 5695
rect 10502 5692 10508 5704
rect 7791 5664 10508 5692
rect 7791 5661 7803 5664
rect 7745 5655 7803 5661
rect 10502 5652 10508 5664
rect 10560 5652 10566 5704
rect 12710 5652 12716 5704
rect 12768 5692 12774 5704
rect 12897 5695 12955 5701
rect 12897 5692 12909 5695
rect 12768 5664 12909 5692
rect 12768 5652 12774 5664
rect 12897 5661 12909 5664
rect 12943 5661 12955 5695
rect 12897 5655 12955 5661
rect 14550 5652 14556 5704
rect 14608 5692 14614 5704
rect 15654 5692 15660 5704
rect 14608 5664 15660 5692
rect 14608 5652 14614 5664
rect 15654 5652 15660 5664
rect 15712 5652 15718 5704
rect 3108 5596 3648 5624
rect 3881 5627 3939 5633
rect 3108 5584 3114 5596
rect 3881 5593 3893 5627
rect 3927 5624 3939 5627
rect 5537 5627 5595 5633
rect 5537 5624 5549 5627
rect 3927 5596 5549 5624
rect 3927 5593 3939 5596
rect 3881 5587 3939 5593
rect 5537 5593 5549 5596
rect 5583 5593 5595 5627
rect 5537 5587 5595 5593
rect 7466 5584 7472 5636
rect 7524 5624 7530 5636
rect 15930 5624 15936 5636
rect 7524 5596 7696 5624
rect 7524 5584 7530 5596
rect 1578 5556 1584 5568
rect 1539 5528 1584 5556
rect 1578 5516 1584 5528
rect 1636 5516 1642 5568
rect 1854 5516 1860 5568
rect 1912 5556 1918 5568
rect 1949 5559 2007 5565
rect 1949 5556 1961 5559
rect 1912 5528 1961 5556
rect 1912 5516 1918 5528
rect 1949 5525 1961 5528
rect 1995 5525 2007 5559
rect 1949 5519 2007 5525
rect 2774 5516 2780 5568
rect 2832 5556 2838 5568
rect 4522 5556 4528 5568
rect 2832 5528 4528 5556
rect 2832 5516 2838 5528
rect 4522 5516 4528 5528
rect 4580 5516 4586 5568
rect 7101 5559 7159 5565
rect 7101 5525 7113 5559
rect 7147 5556 7159 5559
rect 7558 5556 7564 5568
rect 7147 5528 7564 5556
rect 7147 5525 7159 5528
rect 7101 5519 7159 5525
rect 7558 5516 7564 5528
rect 7616 5516 7622 5568
rect 7668 5556 7696 5596
rect 10704 5596 11192 5624
rect 10704 5556 10732 5596
rect 7668 5528 10732 5556
rect 10827 5559 10885 5565
rect 10827 5525 10839 5559
rect 10873 5556 10885 5559
rect 11054 5556 11060 5568
rect 10873 5528 11060 5556
rect 10873 5525 10885 5528
rect 10827 5519 10885 5525
rect 11054 5516 11060 5528
rect 11112 5516 11118 5568
rect 11164 5556 11192 5596
rect 14752 5596 15936 5624
rect 14752 5556 14780 5596
rect 15930 5584 15936 5596
rect 15988 5584 15994 5636
rect 16040 5624 16068 5732
rect 16117 5729 16129 5763
rect 16163 5760 16175 5763
rect 16666 5760 16672 5772
rect 16163 5732 16672 5760
rect 16163 5729 16175 5732
rect 16117 5723 16175 5729
rect 16666 5720 16672 5732
rect 16724 5720 16730 5772
rect 16942 5720 16948 5772
rect 17000 5760 17006 5772
rect 17129 5763 17187 5769
rect 17129 5760 17141 5763
rect 17000 5732 17141 5760
rect 17000 5720 17006 5732
rect 17129 5729 17141 5732
rect 17175 5729 17187 5763
rect 17862 5760 17868 5772
rect 17823 5732 17868 5760
rect 17129 5723 17187 5729
rect 17862 5720 17868 5732
rect 17920 5720 17926 5772
rect 16301 5695 16359 5701
rect 16301 5661 16313 5695
rect 16347 5692 16359 5695
rect 16758 5692 16764 5704
rect 16347 5664 16764 5692
rect 16347 5661 16359 5664
rect 16301 5655 16359 5661
rect 16758 5652 16764 5664
rect 16816 5652 16822 5704
rect 17218 5652 17224 5704
rect 17276 5692 17282 5704
rect 17276 5664 17321 5692
rect 17276 5652 17282 5664
rect 16482 5624 16488 5636
rect 16040 5596 16488 5624
rect 16482 5584 16488 5596
rect 16540 5584 16546 5636
rect 11164 5528 14780 5556
rect 14829 5559 14887 5565
rect 14829 5525 14841 5559
rect 14875 5556 14887 5559
rect 17770 5556 17776 5568
rect 14875 5528 17776 5556
rect 14875 5525 14887 5528
rect 14829 5519 14887 5525
rect 17770 5516 17776 5528
rect 17828 5516 17834 5568
rect 17862 5516 17868 5568
rect 17920 5556 17926 5568
rect 18049 5559 18107 5565
rect 18049 5556 18061 5559
rect 17920 5528 18061 5556
rect 17920 5516 17926 5528
rect 18049 5525 18061 5528
rect 18095 5525 18107 5559
rect 18049 5519 18107 5525
rect 1104 5466 18860 5488
rect 1104 5414 3947 5466
rect 3999 5414 4011 5466
rect 4063 5414 4075 5466
rect 4127 5414 4139 5466
rect 4191 5414 9878 5466
rect 9930 5414 9942 5466
rect 9994 5414 10006 5466
rect 10058 5414 10070 5466
rect 10122 5414 15808 5466
rect 15860 5414 15872 5466
rect 15924 5414 15936 5466
rect 15988 5414 16000 5466
rect 16052 5414 18860 5466
rect 1104 5392 18860 5414
rect 3053 5355 3111 5361
rect 3053 5321 3065 5355
rect 3099 5352 3111 5355
rect 3418 5352 3424 5364
rect 3099 5324 3424 5352
rect 3099 5321 3111 5324
rect 3053 5315 3111 5321
rect 3418 5312 3424 5324
rect 3476 5312 3482 5364
rect 6454 5352 6460 5364
rect 3528 5324 6132 5352
rect 6415 5324 6460 5352
rect 2866 5244 2872 5296
rect 2924 5284 2930 5296
rect 3528 5284 3556 5324
rect 2924 5256 3556 5284
rect 2924 5244 2930 5256
rect 4246 5244 4252 5296
rect 4304 5284 4310 5296
rect 4304 5256 5120 5284
rect 4304 5244 4310 5256
rect 5092 5228 5120 5256
rect 3697 5219 3755 5225
rect 3697 5185 3709 5219
rect 3743 5216 3755 5219
rect 4614 5216 4620 5228
rect 3743 5188 4620 5216
rect 3743 5185 3755 5188
rect 3697 5179 3755 5185
rect 4614 5176 4620 5188
rect 4672 5176 4678 5228
rect 4709 5219 4767 5225
rect 4709 5185 4721 5219
rect 4755 5185 4767 5219
rect 5074 5216 5080 5228
rect 4987 5188 5080 5216
rect 4709 5179 4767 5185
rect 1854 5148 1860 5160
rect 1815 5120 1860 5148
rect 1854 5108 1860 5120
rect 1912 5108 1918 5160
rect 4724 5148 4752 5179
rect 5074 5176 5080 5188
rect 5132 5176 5138 5228
rect 4724 5120 5387 5148
rect 198 5040 204 5092
rect 256 5080 262 5092
rect 2133 5083 2191 5089
rect 2133 5080 2145 5083
rect 256 5052 2145 5080
rect 256 5040 262 5052
rect 2133 5049 2145 5052
rect 2179 5049 2191 5083
rect 2133 5043 2191 5049
rect 3421 5083 3479 5089
rect 3421 5049 3433 5083
rect 3467 5080 3479 5083
rect 4525 5083 4583 5089
rect 3467 5052 4108 5080
rect 3467 5049 3479 5052
rect 3421 5043 3479 5049
rect 3510 5012 3516 5024
rect 3471 4984 3516 5012
rect 3510 4972 3516 4984
rect 3568 4972 3574 5024
rect 4080 5021 4108 5052
rect 4525 5049 4537 5083
rect 4571 5080 4583 5083
rect 4706 5080 4712 5092
rect 4571 5052 4712 5080
rect 4571 5049 4583 5052
rect 4525 5043 4583 5049
rect 4706 5040 4712 5052
rect 4764 5040 4770 5092
rect 5359 5089 5387 5120
rect 5344 5083 5402 5089
rect 5344 5049 5356 5083
rect 5390 5080 5402 5083
rect 5442 5080 5448 5092
rect 5390 5052 5448 5080
rect 5390 5049 5402 5052
rect 5344 5043 5402 5049
rect 5442 5040 5448 5052
rect 5500 5040 5506 5092
rect 4065 5015 4123 5021
rect 4065 4981 4077 5015
rect 4111 4981 4123 5015
rect 4065 4975 4123 4981
rect 4246 4972 4252 5024
rect 4304 5012 4310 5024
rect 4433 5015 4491 5021
rect 4433 5012 4445 5015
rect 4304 4984 4445 5012
rect 4304 4972 4310 4984
rect 4433 4981 4445 4984
rect 4479 5012 4491 5015
rect 5258 5012 5264 5024
rect 4479 4984 5264 5012
rect 4479 4981 4491 4984
rect 4433 4975 4491 4981
rect 5258 4972 5264 4984
rect 5316 4972 5322 5024
rect 6104 5012 6132 5324
rect 6454 5312 6460 5324
rect 6512 5312 6518 5364
rect 9214 5352 9220 5364
rect 6932 5324 9220 5352
rect 6932 5293 6960 5324
rect 9214 5312 9220 5324
rect 9272 5312 9278 5364
rect 9306 5312 9312 5364
rect 9364 5352 9370 5364
rect 10870 5352 10876 5364
rect 9364 5324 10876 5352
rect 9364 5312 9370 5324
rect 10870 5312 10876 5324
rect 10928 5352 10934 5364
rect 12618 5352 12624 5364
rect 10928 5324 12624 5352
rect 10928 5312 10934 5324
rect 12618 5312 12624 5324
rect 12676 5312 12682 5364
rect 14660 5324 15884 5352
rect 6917 5287 6975 5293
rect 6917 5253 6929 5287
rect 6963 5253 6975 5287
rect 14660 5284 14688 5324
rect 6917 5247 6975 5253
rect 11808 5256 14688 5284
rect 7285 5151 7343 5157
rect 7285 5117 7297 5151
rect 7331 5148 7343 5151
rect 7374 5148 7380 5160
rect 7331 5120 7380 5148
rect 7331 5117 7343 5120
rect 7285 5111 7343 5117
rect 7374 5108 7380 5120
rect 7432 5108 7438 5160
rect 8297 5151 8355 5157
rect 8297 5117 8309 5151
rect 8343 5148 8355 5151
rect 8386 5148 8392 5160
rect 8343 5120 8392 5148
rect 8343 5117 8355 5120
rect 8297 5111 8355 5117
rect 8386 5108 8392 5120
rect 8444 5108 8450 5160
rect 9950 5148 9956 5160
rect 9911 5120 9956 5148
rect 9950 5108 9956 5120
rect 10008 5108 10014 5160
rect 11330 5108 11336 5160
rect 11388 5108 11394 5160
rect 11808 5157 11836 5256
rect 15194 5244 15200 5296
rect 15252 5284 15258 5296
rect 15856 5284 15884 5324
rect 16574 5312 16580 5364
rect 16632 5352 16638 5364
rect 16669 5355 16727 5361
rect 16669 5352 16681 5355
rect 16632 5324 16681 5352
rect 16632 5312 16638 5324
rect 16669 5321 16681 5324
rect 16715 5321 16727 5355
rect 16669 5315 16727 5321
rect 16758 5284 16764 5296
rect 15252 5256 15792 5284
rect 15856 5256 16764 5284
rect 15252 5244 15258 5256
rect 12342 5176 12348 5228
rect 12400 5216 12406 5228
rect 12400 5188 14780 5216
rect 12400 5176 12406 5188
rect 11793 5151 11851 5157
rect 11793 5117 11805 5151
rect 11839 5117 11851 5151
rect 14752 5148 14780 5188
rect 14826 5176 14832 5228
rect 14884 5216 14890 5228
rect 14884 5188 14929 5216
rect 14884 5176 14890 5188
rect 15470 5176 15476 5228
rect 15528 5216 15534 5228
rect 15764 5225 15792 5256
rect 16758 5244 16764 5256
rect 16816 5244 16822 5296
rect 15657 5219 15715 5225
rect 15657 5216 15669 5219
rect 15528 5188 15669 5216
rect 15528 5176 15534 5188
rect 15657 5185 15669 5188
rect 15703 5185 15715 5219
rect 15657 5179 15715 5185
rect 15749 5219 15807 5225
rect 15749 5185 15761 5219
rect 15795 5185 15807 5219
rect 17218 5216 17224 5228
rect 17179 5188 17224 5216
rect 15749 5179 15807 5185
rect 17218 5176 17224 5188
rect 17276 5176 17282 5228
rect 16244 5151 16302 5157
rect 16244 5148 16256 5151
rect 14752 5120 16256 5148
rect 11793 5111 11851 5117
rect 16244 5117 16256 5120
rect 16290 5117 16302 5151
rect 17034 5148 17040 5160
rect 16995 5120 17040 5148
rect 16244 5111 16302 5117
rect 17034 5108 17040 5120
rect 17092 5108 17098 5160
rect 18046 5148 18052 5160
rect 18007 5120 18052 5148
rect 18046 5108 18052 5120
rect 18104 5108 18110 5160
rect 7653 5083 7711 5089
rect 7653 5049 7665 5083
rect 7699 5080 7711 5083
rect 7834 5080 7840 5092
rect 7699 5052 7840 5080
rect 7699 5049 7711 5052
rect 7653 5043 7711 5049
rect 7834 5040 7840 5052
rect 7892 5040 7898 5092
rect 8564 5083 8622 5089
rect 8564 5049 8576 5083
rect 8610 5080 8622 5083
rect 8938 5080 8944 5092
rect 8610 5052 8944 5080
rect 8610 5049 8622 5052
rect 8564 5043 8622 5049
rect 8938 5040 8944 5052
rect 8996 5040 9002 5092
rect 10226 5089 10232 5092
rect 10198 5083 10232 5089
rect 10198 5080 10210 5083
rect 9692 5052 10210 5080
rect 9398 5012 9404 5024
rect 6104 4984 9404 5012
rect 9398 4972 9404 4984
rect 9456 4972 9462 5024
rect 9692 5021 9720 5052
rect 10198 5049 10210 5052
rect 10284 5080 10290 5092
rect 11348 5080 11376 5108
rect 12529 5083 12587 5089
rect 12529 5080 12541 5083
rect 10284 5052 10346 5080
rect 11348 5052 12541 5080
rect 10198 5043 10232 5049
rect 10226 5040 10232 5043
rect 10284 5040 10290 5052
rect 12529 5049 12541 5052
rect 12575 5049 12587 5083
rect 12529 5043 12587 5049
rect 12618 5040 12624 5092
rect 12676 5080 12682 5092
rect 13541 5083 13599 5089
rect 12676 5052 12721 5080
rect 12676 5040 12682 5052
rect 13541 5049 13553 5083
rect 13587 5080 13599 5083
rect 13630 5080 13636 5092
rect 13587 5052 13636 5080
rect 13587 5049 13599 5052
rect 13541 5043 13599 5049
rect 13630 5040 13636 5052
rect 13688 5040 13694 5092
rect 13909 5083 13967 5089
rect 13909 5080 13921 5083
rect 13832 5052 13921 5080
rect 13832 5024 13860 5052
rect 13909 5049 13921 5052
rect 13955 5049 13967 5083
rect 13909 5043 13967 5049
rect 14001 5083 14059 5089
rect 14001 5049 14013 5083
rect 14047 5080 14059 5083
rect 16347 5083 16405 5089
rect 16347 5080 16359 5083
rect 14047 5052 16359 5080
rect 14047 5049 14059 5052
rect 14001 5043 14059 5049
rect 16347 5049 16359 5052
rect 16393 5049 16405 5083
rect 16347 5043 16405 5049
rect 9677 5015 9735 5021
rect 9677 4981 9689 5015
rect 9723 4981 9735 5015
rect 9677 4975 9735 4981
rect 10318 4972 10324 5024
rect 10376 5012 10382 5024
rect 11333 5015 11391 5021
rect 11333 5012 11345 5015
rect 10376 4984 11345 5012
rect 10376 4972 10382 4984
rect 11333 4981 11345 4984
rect 11379 4981 11391 5015
rect 11333 4975 11391 4981
rect 11977 5015 12035 5021
rect 11977 4981 11989 5015
rect 12023 5012 12035 5015
rect 13722 5012 13728 5024
rect 12023 4984 13728 5012
rect 12023 4981 12035 4984
rect 11977 4975 12035 4981
rect 13722 4972 13728 4984
rect 13780 4972 13786 5024
rect 13814 4972 13820 5024
rect 13872 4972 13878 5024
rect 15194 5012 15200 5024
rect 15155 4984 15200 5012
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 15378 4972 15384 5024
rect 15436 5012 15442 5024
rect 15565 5015 15623 5021
rect 15565 5012 15577 5015
rect 15436 4984 15577 5012
rect 15436 4972 15442 4984
rect 15565 4981 15577 4984
rect 15611 4981 15623 5015
rect 15565 4975 15623 4981
rect 16850 4972 16856 5024
rect 16908 5012 16914 5024
rect 17129 5015 17187 5021
rect 17129 5012 17141 5015
rect 16908 4984 17141 5012
rect 16908 4972 16914 4984
rect 17129 4981 17141 4984
rect 17175 5012 17187 5015
rect 17494 5012 17500 5024
rect 17175 4984 17500 5012
rect 17175 4981 17187 4984
rect 17129 4975 17187 4981
rect 17494 4972 17500 4984
rect 17552 4972 17558 5024
rect 18230 5012 18236 5024
rect 18191 4984 18236 5012
rect 18230 4972 18236 4984
rect 18288 4972 18294 5024
rect 1104 4922 18860 4944
rect 1104 4870 6912 4922
rect 6964 4870 6976 4922
rect 7028 4870 7040 4922
rect 7092 4870 7104 4922
rect 7156 4870 12843 4922
rect 12895 4870 12907 4922
rect 12959 4870 12971 4922
rect 13023 4870 13035 4922
rect 13087 4870 18860 4922
rect 1104 4848 18860 4870
rect 2406 4808 2412 4820
rect 2367 4780 2412 4808
rect 2406 4768 2412 4780
rect 2464 4768 2470 4820
rect 3510 4768 3516 4820
rect 3568 4808 3574 4820
rect 4525 4811 4583 4817
rect 4525 4808 4537 4811
rect 3568 4780 4537 4808
rect 3568 4768 3574 4780
rect 4525 4777 4537 4780
rect 4571 4777 4583 4811
rect 4525 4771 4583 4777
rect 4985 4811 5043 4817
rect 4985 4777 4997 4811
rect 5031 4808 5043 4811
rect 5166 4808 5172 4820
rect 5031 4780 5172 4808
rect 5031 4777 5043 4780
rect 4985 4771 5043 4777
rect 5166 4768 5172 4780
rect 5224 4768 5230 4820
rect 6181 4811 6239 4817
rect 6181 4777 6193 4811
rect 6227 4808 6239 4811
rect 7466 4808 7472 4820
rect 6227 4780 7472 4808
rect 6227 4777 6239 4780
rect 6181 4771 6239 4777
rect 7466 4768 7472 4780
rect 7524 4768 7530 4820
rect 15194 4808 15200 4820
rect 7760 4780 15200 4808
rect 7760 4740 7788 4780
rect 15194 4768 15200 4780
rect 15252 4768 15258 4820
rect 16666 4808 16672 4820
rect 16627 4780 16672 4808
rect 16666 4768 16672 4780
rect 16724 4768 16730 4820
rect 17037 4811 17095 4817
rect 17037 4777 17049 4811
rect 17083 4808 17095 4811
rect 17954 4808 17960 4820
rect 17083 4780 17960 4808
rect 17083 4777 17095 4780
rect 17037 4771 17095 4777
rect 17954 4768 17960 4780
rect 18012 4768 18018 4820
rect 9306 4740 9312 4752
rect 3068 4712 7788 4740
rect 9267 4712 9312 4740
rect 3068 4681 3096 4712
rect 9306 4700 9312 4712
rect 9364 4700 9370 4752
rect 10318 4749 10324 4752
rect 10312 4740 10324 4749
rect 10279 4712 10324 4740
rect 10312 4703 10324 4712
rect 10318 4700 10324 4703
rect 10376 4700 10382 4752
rect 11054 4700 11060 4752
rect 11112 4740 11118 4752
rect 13081 4743 13139 4749
rect 13081 4740 13093 4743
rect 11112 4712 13093 4740
rect 11112 4700 11118 4712
rect 13081 4709 13093 4712
rect 13127 4709 13139 4743
rect 13998 4740 14004 4752
rect 13959 4712 14004 4740
rect 13081 4703 13139 4709
rect 13998 4700 14004 4712
rect 14056 4700 14062 4752
rect 15473 4743 15531 4749
rect 15473 4709 15485 4743
rect 15519 4740 15531 4743
rect 15562 4740 15568 4752
rect 15519 4712 15568 4740
rect 15519 4709 15531 4712
rect 15473 4703 15531 4709
rect 15562 4700 15568 4712
rect 15620 4700 15626 4752
rect 1673 4675 1731 4681
rect 1673 4641 1685 4675
rect 1719 4641 1731 4675
rect 1673 4635 1731 4641
rect 2133 4675 2191 4681
rect 2133 4641 2145 4675
rect 2179 4672 2191 4675
rect 2225 4675 2283 4681
rect 2225 4672 2237 4675
rect 2179 4644 2237 4672
rect 2179 4641 2191 4644
rect 2133 4635 2191 4641
rect 2225 4641 2237 4644
rect 2271 4641 2283 4675
rect 2225 4635 2283 4641
rect 3053 4675 3111 4681
rect 3053 4641 3065 4675
rect 3099 4641 3111 4675
rect 3053 4635 3111 4641
rect 1688 4536 1716 4635
rect 3786 4632 3792 4684
rect 3844 4672 3850 4684
rect 4893 4675 4951 4681
rect 4893 4672 4905 4675
rect 3844 4644 4905 4672
rect 3844 4632 3850 4644
rect 4893 4641 4905 4644
rect 4939 4641 4951 4675
rect 4893 4635 4951 4641
rect 5074 4632 5080 4684
rect 5132 4672 5138 4684
rect 6273 4675 6331 4681
rect 6273 4672 6285 4675
rect 5132 4644 6285 4672
rect 5132 4632 5138 4644
rect 6273 4641 6285 4644
rect 6319 4641 6331 4675
rect 6273 4635 6331 4641
rect 6540 4675 6598 4681
rect 6540 4641 6552 4675
rect 6586 4672 6598 4675
rect 7374 4672 7380 4684
rect 6586 4644 7380 4672
rect 6586 4641 6598 4644
rect 6540 4635 6598 4641
rect 7374 4632 7380 4644
rect 7432 4632 7438 4684
rect 8938 4672 8944 4684
rect 8899 4644 8944 4672
rect 8938 4632 8944 4644
rect 8996 4632 9002 4684
rect 11701 4675 11759 4681
rect 9048 4644 11100 4672
rect 3142 4564 3148 4616
rect 3200 4604 3206 4616
rect 3237 4607 3295 4613
rect 3237 4604 3249 4607
rect 3200 4576 3249 4604
rect 3200 4564 3206 4576
rect 3237 4573 3249 4576
rect 3283 4573 3295 4607
rect 3237 4567 3295 4573
rect 5169 4607 5227 4613
rect 5169 4573 5181 4607
rect 5215 4604 5227 4607
rect 5442 4604 5448 4616
rect 5215 4576 5448 4604
rect 5215 4573 5227 4576
rect 5169 4567 5227 4573
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 9048 4604 9076 4644
rect 7576 4576 9076 4604
rect 7576 4536 7604 4576
rect 9950 4564 9956 4616
rect 10008 4604 10014 4616
rect 10045 4607 10103 4613
rect 10045 4604 10057 4607
rect 10008 4576 10057 4604
rect 10008 4564 10014 4576
rect 10045 4573 10057 4576
rect 10091 4573 10103 4607
rect 11072 4604 11100 4644
rect 11701 4641 11713 4675
rect 11747 4672 11759 4675
rect 11790 4672 11796 4684
rect 11747 4644 11796 4672
rect 11747 4641 11759 4644
rect 11701 4635 11759 4641
rect 11790 4632 11796 4644
rect 11848 4632 11854 4684
rect 12345 4675 12403 4681
rect 12345 4641 12357 4675
rect 12391 4641 12403 4675
rect 12345 4635 12403 4641
rect 14645 4675 14703 4681
rect 14645 4641 14657 4675
rect 14691 4672 14703 4675
rect 15194 4672 15200 4684
rect 14691 4644 15200 4672
rect 14691 4641 14703 4644
rect 14645 4635 14703 4641
rect 11072 4576 12020 4604
rect 10045 4567 10103 4573
rect 8570 4536 8576 4548
rect 1688 4508 6316 4536
rect 1854 4468 1860 4480
rect 1815 4440 1860 4468
rect 1854 4428 1860 4440
rect 1912 4428 1918 4480
rect 2133 4471 2191 4477
rect 2133 4437 2145 4471
rect 2179 4468 2191 4471
rect 6181 4471 6239 4477
rect 6181 4468 6193 4471
rect 2179 4440 6193 4468
rect 2179 4437 2191 4440
rect 2133 4431 2191 4437
rect 6181 4437 6193 4440
rect 6227 4437 6239 4471
rect 6288 4468 6316 4508
rect 7208 4508 7604 4536
rect 8483 4508 8576 4536
rect 7208 4468 7236 4508
rect 8570 4496 8576 4508
rect 8628 4536 8634 4548
rect 9214 4536 9220 4548
rect 8628 4508 9220 4536
rect 8628 4496 8634 4508
rect 9214 4496 9220 4508
rect 9272 4496 9278 4548
rect 7650 4468 7656 4480
rect 6288 4440 7236 4468
rect 7611 4440 7656 4468
rect 6181 4431 6239 4437
rect 7650 4428 7656 4440
rect 7708 4428 7714 4480
rect 10060 4468 10088 4567
rect 10962 4468 10968 4480
rect 10060 4440 10968 4468
rect 10962 4428 10968 4440
rect 11020 4428 11026 4480
rect 11422 4468 11428 4480
rect 11383 4440 11428 4468
rect 11422 4428 11428 4440
rect 11480 4428 11486 4480
rect 11882 4468 11888 4480
rect 11843 4440 11888 4468
rect 11882 4428 11888 4440
rect 11940 4428 11946 4480
rect 11992 4468 12020 4576
rect 12360 4536 12388 4635
rect 15194 4632 15200 4644
rect 15252 4632 15258 4684
rect 17402 4632 17408 4684
rect 17460 4672 17466 4684
rect 17865 4675 17923 4681
rect 17865 4672 17877 4675
rect 17460 4644 17877 4672
rect 17460 4632 17466 4644
rect 17865 4641 17877 4644
rect 17911 4641 17923 4675
rect 17865 4635 17923 4641
rect 12989 4607 13047 4613
rect 12989 4573 13001 4607
rect 13035 4604 13047 4607
rect 13262 4604 13268 4616
rect 13035 4576 13268 4604
rect 13035 4573 13047 4576
rect 12989 4567 13047 4573
rect 13262 4564 13268 4576
rect 13320 4564 13326 4616
rect 14550 4564 14556 4616
rect 14608 4604 14614 4616
rect 15381 4607 15439 4613
rect 15381 4604 15393 4607
rect 14608 4576 15393 4604
rect 14608 4564 14614 4576
rect 15381 4573 15393 4576
rect 15427 4573 15439 4607
rect 16206 4604 16212 4616
rect 16167 4576 16212 4604
rect 15381 4567 15439 4573
rect 16206 4564 16212 4576
rect 16264 4564 16270 4616
rect 17126 4604 17132 4616
rect 17087 4576 17132 4604
rect 17126 4564 17132 4576
rect 17184 4564 17190 4616
rect 17218 4564 17224 4616
rect 17276 4604 17282 4616
rect 17276 4576 17321 4604
rect 17276 4564 17282 4576
rect 16850 4536 16856 4548
rect 12360 4508 16856 4536
rect 16850 4496 16856 4508
rect 16908 4496 16914 4548
rect 12434 4468 12440 4480
rect 11992 4440 12440 4468
rect 12434 4428 12440 4440
rect 12492 4428 12498 4480
rect 12529 4471 12587 4477
rect 12529 4437 12541 4471
rect 12575 4468 12587 4471
rect 12710 4468 12716 4480
rect 12575 4440 12716 4468
rect 12575 4437 12587 4440
rect 12529 4431 12587 4437
rect 12710 4428 12716 4440
rect 12768 4428 12774 4480
rect 14829 4471 14887 4477
rect 14829 4437 14841 4471
rect 14875 4468 14887 4471
rect 16206 4468 16212 4480
rect 14875 4440 16212 4468
rect 14875 4437 14887 4440
rect 14829 4431 14887 4437
rect 16206 4428 16212 4440
rect 16264 4428 16270 4480
rect 17862 4428 17868 4480
rect 17920 4468 17926 4480
rect 18049 4471 18107 4477
rect 18049 4468 18061 4471
rect 17920 4440 18061 4468
rect 17920 4428 17926 4440
rect 18049 4437 18061 4440
rect 18095 4437 18107 4471
rect 18049 4431 18107 4437
rect 1104 4378 18860 4400
rect 1104 4326 3947 4378
rect 3999 4326 4011 4378
rect 4063 4326 4075 4378
rect 4127 4326 4139 4378
rect 4191 4326 9878 4378
rect 9930 4326 9942 4378
rect 9994 4326 10006 4378
rect 10058 4326 10070 4378
rect 10122 4326 15808 4378
rect 15860 4326 15872 4378
rect 15924 4326 15936 4378
rect 15988 4326 16000 4378
rect 16052 4326 18860 4378
rect 1104 4304 18860 4326
rect 4338 4264 4344 4276
rect 4080 4236 4344 4264
rect 4080 4137 4108 4236
rect 4338 4224 4344 4236
rect 4396 4224 4402 4276
rect 5442 4264 5448 4276
rect 5403 4236 5448 4264
rect 5442 4224 5448 4236
rect 5500 4224 5506 4276
rect 8386 4264 8392 4276
rect 7760 4236 8392 4264
rect 5074 4156 5080 4208
rect 5132 4196 5138 4208
rect 7760 4196 7788 4236
rect 8386 4224 8392 4236
rect 8444 4224 8450 4276
rect 8938 4224 8944 4276
rect 8996 4264 9002 4276
rect 9125 4267 9183 4273
rect 9125 4264 9137 4267
rect 8996 4236 9137 4264
rect 8996 4224 9002 4236
rect 9125 4233 9137 4236
rect 9171 4233 9183 4267
rect 9125 4227 9183 4233
rect 9398 4224 9404 4276
rect 9456 4264 9462 4276
rect 17126 4264 17132 4276
rect 9456 4236 17132 4264
rect 9456 4224 9462 4236
rect 17126 4224 17132 4236
rect 17184 4224 17190 4276
rect 5132 4168 7788 4196
rect 5132 4156 5138 4168
rect 4065 4131 4123 4137
rect 4065 4097 4077 4131
rect 4111 4097 4123 4131
rect 4065 4091 4123 4097
rect 5626 4088 5632 4140
rect 5684 4128 5690 4140
rect 6546 4128 6552 4140
rect 5684 4100 6552 4128
rect 5684 4088 5690 4100
rect 6546 4088 6552 4100
rect 6604 4088 6610 4140
rect 7760 4137 7788 4168
rect 9766 4156 9772 4208
rect 9824 4196 9830 4208
rect 12621 4199 12679 4205
rect 12621 4196 12633 4199
rect 9824 4168 12633 4196
rect 9824 4156 9830 4168
rect 12621 4165 12633 4168
rect 12667 4165 12679 4199
rect 15746 4196 15752 4208
rect 12621 4159 12679 4165
rect 14971 4168 15752 4196
rect 7745 4131 7803 4137
rect 7745 4097 7757 4131
rect 7791 4097 7803 4131
rect 7745 4091 7803 4097
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 9582 4128 9588 4140
rect 9272 4100 9588 4128
rect 9272 4088 9278 4100
rect 9582 4088 9588 4100
rect 9640 4128 9646 4140
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 9640 4100 10057 4128
rect 9640 4088 9646 4100
rect 10045 4097 10057 4100
rect 10091 4128 10103 4131
rect 10781 4131 10839 4137
rect 10091 4100 10548 4128
rect 10091 4097 10103 4100
rect 10045 4091 10103 4097
rect 1581 4063 1639 4069
rect 1581 4029 1593 4063
rect 1627 4060 1639 4063
rect 2317 4063 2375 4069
rect 1627 4032 2268 4060
rect 1627 4029 1639 4032
rect 1581 4023 1639 4029
rect 1857 3995 1915 4001
rect 1857 3961 1869 3995
rect 1903 3992 1915 3995
rect 2130 3992 2136 4004
rect 1903 3964 2136 3992
rect 1903 3961 1915 3964
rect 1857 3955 1915 3961
rect 2130 3952 2136 3964
rect 2188 3952 2194 4004
rect 2240 3992 2268 4032
rect 2317 4029 2329 4063
rect 2363 4060 2375 4063
rect 8478 4060 8484 4072
rect 2363 4032 8484 4060
rect 2363 4029 2375 4032
rect 2317 4023 2375 4029
rect 8478 4020 8484 4032
rect 8536 4020 8542 4072
rect 9306 4020 9312 4072
rect 9364 4060 9370 4072
rect 9401 4063 9459 4069
rect 9401 4060 9413 4063
rect 9364 4032 9413 4060
rect 9364 4020 9370 4032
rect 9401 4029 9413 4032
rect 9447 4029 9459 4063
rect 9401 4023 9459 4029
rect 10318 4020 10324 4072
rect 10376 4060 10382 4072
rect 10413 4063 10471 4069
rect 10413 4060 10425 4063
rect 10376 4032 10425 4060
rect 10376 4020 10382 4032
rect 10413 4029 10425 4032
rect 10459 4029 10471 4063
rect 10520 4060 10548 4100
rect 10781 4097 10793 4131
rect 10827 4128 10839 4131
rect 14971 4128 14999 4168
rect 15746 4156 15752 4168
rect 15804 4156 15810 4208
rect 16482 4156 16488 4208
rect 16540 4196 16546 4208
rect 16540 4168 16620 4196
rect 16540 4156 16546 4168
rect 15102 4128 15108 4140
rect 10827 4100 12388 4128
rect 10827 4097 10839 4100
rect 10781 4091 10839 4097
rect 11057 4063 11115 4069
rect 11057 4060 11069 4063
rect 10520 4032 11069 4060
rect 10413 4023 10471 4029
rect 11057 4029 11069 4032
rect 11103 4029 11115 4063
rect 11422 4060 11428 4072
rect 11383 4032 11428 4060
rect 11057 4023 11115 4029
rect 11422 4020 11428 4032
rect 11480 4020 11486 4072
rect 11790 4060 11796 4072
rect 11751 4032 11796 4060
rect 11790 4020 11796 4032
rect 11848 4020 11854 4072
rect 12253 4063 12311 4069
rect 12253 4029 12265 4063
rect 12299 4029 12311 4063
rect 12253 4023 12311 4029
rect 4332 3995 4390 4001
rect 2240 3964 4292 3992
rect 2498 3924 2504 3936
rect 2459 3896 2504 3924
rect 2498 3884 2504 3896
rect 2556 3884 2562 3936
rect 4264 3924 4292 3964
rect 4332 3961 4344 3995
rect 4378 3992 4390 3995
rect 4614 3992 4620 4004
rect 4378 3964 4620 3992
rect 4378 3961 4390 3964
rect 4332 3955 4390 3961
rect 4614 3952 4620 3964
rect 4672 3952 4678 4004
rect 8012 3995 8070 4001
rect 8012 3961 8024 3995
rect 8058 3992 8070 3995
rect 8294 3992 8300 4004
rect 8058 3964 8300 3992
rect 8058 3961 8070 3964
rect 8012 3955 8070 3961
rect 8294 3952 8300 3964
rect 8352 3952 8358 4004
rect 11974 3952 11980 4004
rect 12032 3992 12038 4004
rect 12268 3992 12296 4023
rect 12032 3964 12296 3992
rect 12360 3992 12388 4100
rect 12452 4100 14999 4128
rect 15063 4100 15108 4128
rect 12452 4069 12480 4100
rect 15102 4088 15108 4100
rect 15160 4088 15166 4140
rect 15286 4088 15292 4140
rect 15344 4128 15350 4140
rect 16592 4137 16620 4168
rect 15657 4131 15715 4137
rect 15657 4128 15669 4131
rect 15344 4100 15669 4128
rect 15344 4088 15350 4100
rect 15657 4097 15669 4100
rect 15703 4097 15715 4131
rect 15657 4091 15715 4097
rect 16577 4131 16635 4137
rect 16577 4097 16589 4131
rect 16623 4097 16635 4131
rect 17586 4128 17592 4140
rect 16577 4091 16635 4097
rect 17420 4100 17592 4128
rect 12437 4063 12495 4069
rect 12437 4029 12449 4063
rect 12483 4029 12495 4063
rect 12437 4023 12495 4029
rect 13081 4063 13139 4069
rect 13081 4029 13093 4063
rect 13127 4060 13139 4063
rect 13170 4060 13176 4072
rect 13127 4032 13176 4060
rect 13127 4029 13139 4032
rect 13081 4023 13139 4029
rect 12452 3992 12480 4023
rect 13170 4020 13176 4032
rect 13228 4020 13234 4072
rect 13630 4060 13636 4072
rect 13591 4032 13636 4060
rect 13630 4020 13636 4032
rect 13688 4020 13694 4072
rect 17420 4069 17448 4100
rect 17586 4088 17592 4100
rect 17644 4088 17650 4140
rect 17770 4088 17776 4140
rect 17828 4128 17834 4140
rect 18506 4128 18512 4140
rect 17828 4100 18512 4128
rect 17828 4088 17834 4100
rect 18506 4088 18512 4100
rect 18564 4088 18570 4140
rect 16980 4063 17038 4069
rect 16980 4060 16992 4063
rect 16500 4032 16992 4060
rect 14274 3992 14280 4004
rect 12360 3964 12480 3992
rect 14235 3964 14280 3992
rect 12032 3952 12038 3964
rect 14274 3952 14280 3964
rect 14332 3952 14338 4004
rect 14369 3995 14427 4001
rect 14369 3961 14381 3995
rect 14415 3992 14427 3995
rect 14415 3964 15424 3992
rect 14415 3961 14427 3964
rect 14369 3955 14427 3961
rect 7926 3924 7932 3936
rect 4264 3896 7932 3924
rect 7926 3884 7932 3896
rect 7984 3884 7990 3936
rect 8754 3884 8760 3936
rect 8812 3924 8818 3936
rect 9585 3927 9643 3933
rect 9585 3924 9597 3927
rect 8812 3896 9597 3924
rect 8812 3884 8818 3896
rect 9585 3893 9597 3896
rect 9631 3893 9643 3927
rect 9585 3887 9643 3893
rect 10962 3884 10968 3936
rect 11020 3924 11026 3936
rect 12069 3927 12127 3933
rect 12069 3924 12081 3927
rect 11020 3896 12081 3924
rect 11020 3884 11026 3896
rect 12069 3893 12081 3896
rect 12115 3893 12127 3927
rect 12069 3887 12127 3893
rect 13265 3927 13323 3933
rect 13265 3893 13277 3927
rect 13311 3924 13323 3927
rect 13446 3924 13452 3936
rect 13311 3896 13452 3924
rect 13311 3893 13323 3896
rect 13265 3887 13323 3893
rect 13446 3884 13452 3896
rect 13504 3884 13510 3936
rect 13817 3927 13875 3933
rect 13817 3893 13829 3927
rect 13863 3924 13875 3927
rect 13998 3924 14004 3936
rect 13863 3896 14004 3924
rect 13863 3893 13875 3896
rect 13817 3887 13875 3893
rect 13998 3884 14004 3896
rect 14056 3884 14062 3936
rect 15396 3924 15424 3964
rect 15746 3952 15752 4004
rect 15804 3992 15810 4004
rect 16500 3992 16528 4032
rect 16980 4029 16992 4032
rect 17026 4029 17038 4063
rect 16980 4023 17038 4029
rect 17405 4063 17463 4069
rect 17405 4029 17417 4063
rect 17451 4029 17463 4063
rect 17405 4023 17463 4029
rect 17494 4020 17500 4072
rect 17552 4060 17558 4072
rect 18049 4063 18107 4069
rect 18049 4060 18061 4063
rect 17552 4032 18061 4060
rect 17552 4020 17558 4032
rect 18049 4029 18061 4032
rect 18095 4029 18107 4063
rect 18049 4023 18107 4029
rect 15804 3964 16528 3992
rect 15804 3952 15810 3964
rect 16574 3952 16580 4004
rect 16632 3992 16638 4004
rect 19610 3992 19616 4004
rect 16632 3964 19616 3992
rect 16632 3952 16638 3964
rect 19610 3952 19616 3964
rect 19668 3952 19674 4004
rect 17083 3927 17141 3933
rect 17083 3924 17095 3927
rect 15396 3896 17095 3924
rect 17083 3893 17095 3896
rect 17129 3893 17141 3927
rect 17586 3924 17592 3936
rect 17547 3896 17592 3924
rect 17083 3887 17141 3893
rect 17586 3884 17592 3896
rect 17644 3884 17650 3936
rect 18230 3924 18236 3936
rect 18191 3896 18236 3924
rect 18230 3884 18236 3896
rect 18288 3884 18294 3936
rect 1104 3834 18860 3856
rect 1104 3782 6912 3834
rect 6964 3782 6976 3834
rect 7028 3782 7040 3834
rect 7092 3782 7104 3834
rect 7156 3782 12843 3834
rect 12895 3782 12907 3834
rect 12959 3782 12971 3834
rect 13023 3782 13035 3834
rect 13087 3782 18860 3834
rect 1104 3760 18860 3782
rect 6641 3723 6699 3729
rect 1688 3692 3924 3720
rect 1688 3593 1716 3692
rect 3786 3652 3792 3664
rect 2240 3624 3792 3652
rect 2240 3593 2268 3624
rect 3786 3612 3792 3624
rect 3844 3612 3850 3664
rect 3896 3652 3924 3692
rect 6641 3689 6653 3723
rect 6687 3720 6699 3723
rect 6825 3723 6883 3729
rect 6825 3720 6837 3723
rect 6687 3692 6837 3720
rect 6687 3689 6699 3692
rect 6641 3683 6699 3689
rect 6825 3689 6837 3692
rect 6871 3689 6883 3723
rect 8294 3720 8300 3732
rect 8255 3692 8300 3720
rect 6825 3683 6883 3689
rect 8294 3680 8300 3692
rect 8352 3680 8358 3732
rect 15010 3720 15016 3732
rect 10152 3692 11560 3720
rect 5350 3652 5356 3664
rect 3896 3624 5356 3652
rect 5350 3612 5356 3624
rect 5408 3612 5414 3664
rect 5528 3655 5586 3661
rect 5528 3621 5540 3655
rect 5574 3652 5586 3655
rect 7650 3652 7656 3664
rect 5574 3624 7656 3652
rect 5574 3621 5586 3624
rect 5528 3615 5586 3621
rect 7650 3612 7656 3624
rect 7708 3612 7714 3664
rect 1673 3587 1731 3593
rect 1673 3553 1685 3587
rect 1719 3553 1731 3587
rect 1673 3547 1731 3553
rect 2225 3587 2283 3593
rect 2225 3553 2237 3587
rect 2271 3553 2283 3587
rect 2225 3547 2283 3553
rect 2774 3544 2780 3596
rect 2832 3584 2838 3596
rect 2832 3556 2877 3584
rect 2832 3544 2838 3556
rect 4338 3544 4344 3596
rect 4396 3584 4402 3596
rect 5261 3587 5319 3593
rect 5261 3584 5273 3587
rect 4396 3556 5273 3584
rect 4396 3544 4402 3556
rect 5261 3553 5273 3556
rect 5307 3584 5319 3587
rect 6825 3587 6883 3593
rect 5307 3556 6500 3584
rect 5307 3553 5319 3556
rect 5261 3547 5319 3553
rect 2130 3476 2136 3528
rect 2188 3516 2194 3528
rect 3050 3516 3056 3528
rect 2188 3488 3056 3516
rect 2188 3476 2194 3488
rect 3050 3476 3056 3488
rect 3108 3476 3114 3528
rect 6472 3516 6500 3556
rect 6825 3553 6837 3587
rect 6871 3584 6883 3587
rect 7173 3587 7231 3593
rect 7173 3584 7185 3587
rect 6871 3556 7185 3584
rect 6871 3553 6883 3556
rect 6825 3547 6883 3553
rect 7173 3553 7185 3556
rect 7219 3584 7231 3587
rect 7466 3584 7472 3596
rect 7219 3556 7472 3584
rect 7219 3553 7231 3556
rect 7173 3547 7231 3553
rect 7466 3544 7472 3556
rect 7524 3544 7530 3596
rect 8312 3584 8340 3680
rect 8386 3612 8392 3664
rect 8444 3652 8450 3664
rect 9674 3652 9680 3664
rect 8444 3624 9680 3652
rect 8444 3612 8450 3624
rect 9674 3612 9680 3624
rect 9732 3612 9738 3664
rect 8941 3587 8999 3593
rect 8941 3584 8953 3587
rect 8312 3556 8953 3584
rect 8941 3553 8953 3556
rect 8987 3553 8999 3587
rect 8941 3547 8999 3553
rect 9582 3544 9588 3596
rect 9640 3584 9646 3596
rect 10152 3593 10180 3692
rect 11048 3655 11106 3661
rect 11048 3621 11060 3655
rect 11094 3652 11106 3655
rect 11422 3652 11428 3664
rect 11094 3624 11428 3652
rect 11094 3621 11106 3624
rect 11048 3615 11106 3621
rect 11422 3612 11428 3624
rect 11480 3612 11486 3664
rect 11532 3652 11560 3692
rect 12636 3692 15016 3720
rect 12636 3661 12664 3692
rect 15010 3680 15016 3692
rect 15068 3680 15074 3732
rect 12253 3655 12311 3661
rect 12253 3652 12265 3655
rect 11532 3624 12265 3652
rect 12253 3621 12265 3624
rect 12299 3621 12311 3655
rect 12253 3615 12311 3621
rect 12621 3655 12679 3661
rect 12621 3621 12633 3655
rect 12667 3621 12679 3655
rect 13538 3652 13544 3664
rect 13499 3624 13544 3652
rect 12621 3615 12679 3621
rect 13538 3612 13544 3624
rect 13596 3612 13602 3664
rect 13906 3612 13912 3664
rect 13964 3652 13970 3664
rect 15427 3655 15485 3661
rect 15427 3652 15439 3655
rect 13964 3624 15439 3652
rect 13964 3612 13970 3624
rect 15427 3621 15439 3624
rect 15473 3621 15485 3655
rect 15427 3615 15485 3621
rect 15654 3612 15660 3664
rect 15712 3652 15718 3664
rect 15841 3655 15899 3661
rect 15841 3652 15853 3655
rect 15712 3624 15853 3652
rect 15712 3612 15718 3624
rect 15841 3621 15853 3624
rect 15887 3621 15899 3655
rect 15841 3615 15899 3621
rect 15933 3655 15991 3661
rect 15933 3621 15945 3655
rect 15979 3652 15991 3655
rect 16298 3652 16304 3664
rect 15979 3624 16304 3652
rect 15979 3621 15991 3624
rect 15933 3615 15991 3621
rect 16298 3612 16304 3624
rect 16356 3612 16362 3664
rect 16850 3652 16856 3664
rect 16811 3624 16856 3652
rect 16850 3612 16856 3624
rect 16908 3612 16914 3664
rect 17034 3612 17040 3664
rect 17092 3652 17098 3664
rect 17092 3624 17908 3652
rect 17092 3612 17098 3624
rect 9769 3587 9827 3593
rect 9769 3584 9781 3587
rect 9640 3556 9781 3584
rect 9640 3544 9646 3556
rect 9769 3553 9781 3556
rect 9815 3553 9827 3587
rect 9769 3547 9827 3553
rect 10137 3587 10195 3593
rect 10137 3553 10149 3587
rect 10183 3553 10195 3587
rect 10137 3547 10195 3553
rect 6917 3519 6975 3525
rect 6917 3516 6929 3519
rect 6472 3488 6929 3516
rect 6917 3485 6929 3488
rect 6963 3485 6975 3519
rect 8570 3516 8576 3528
rect 8531 3488 8576 3516
rect 6917 3479 6975 3485
rect 8570 3476 8576 3488
rect 8628 3476 8634 3528
rect 10152 3516 10180 3547
rect 10226 3544 10232 3596
rect 10284 3584 10290 3596
rect 11882 3584 11888 3596
rect 10284 3556 11888 3584
rect 10284 3544 10290 3556
rect 11882 3544 11888 3556
rect 11940 3544 11946 3596
rect 14090 3584 14096 3596
rect 14051 3556 14096 3584
rect 14090 3544 14096 3556
rect 14148 3544 14154 3596
rect 14461 3587 14519 3593
rect 14461 3553 14473 3587
rect 14507 3584 14519 3587
rect 14645 3587 14703 3593
rect 14645 3584 14657 3587
rect 14507 3556 14657 3584
rect 14507 3553 14519 3556
rect 14461 3547 14519 3553
rect 14645 3553 14657 3556
rect 14691 3553 14703 3587
rect 14645 3547 14703 3553
rect 15102 3544 15108 3596
rect 15160 3584 15166 3596
rect 17880 3593 17908 3624
rect 15324 3587 15382 3593
rect 15324 3584 15336 3587
rect 15160 3556 15336 3584
rect 15160 3544 15166 3556
rect 15324 3553 15336 3556
rect 15370 3553 15382 3587
rect 15324 3547 15382 3553
rect 17129 3587 17187 3593
rect 17129 3553 17141 3587
rect 17175 3553 17187 3587
rect 17129 3547 17187 3553
rect 17865 3587 17923 3593
rect 17865 3553 17877 3587
rect 17911 3553 17923 3587
rect 17865 3547 17923 3553
rect 10778 3516 10784 3528
rect 8864 3488 10180 3516
rect 10739 3488 10784 3516
rect 1854 3448 1860 3460
rect 1815 3420 1860 3448
rect 1854 3408 1860 3420
rect 1912 3408 1918 3460
rect 1210 3340 1216 3392
rect 1268 3380 1274 3392
rect 2409 3383 2467 3389
rect 2409 3380 2421 3383
rect 1268 3352 2421 3380
rect 1268 3340 1274 3352
rect 2409 3349 2421 3352
rect 2455 3349 2467 3383
rect 2958 3380 2964 3392
rect 2919 3352 2964 3380
rect 2409 3343 2467 3349
rect 2958 3340 2964 3352
rect 3016 3340 3022 3392
rect 5166 3340 5172 3392
rect 5224 3380 5230 3392
rect 8864 3380 8892 3488
rect 10778 3476 10784 3488
rect 10836 3476 10842 3528
rect 12158 3476 12164 3528
rect 12216 3516 12222 3528
rect 12529 3519 12587 3525
rect 12529 3516 12541 3519
rect 12216 3488 12541 3516
rect 12216 3476 12222 3488
rect 12529 3485 12541 3488
rect 12575 3485 12587 3519
rect 12529 3479 12587 3485
rect 14001 3519 14059 3525
rect 14001 3485 14013 3519
rect 14047 3516 14059 3519
rect 17144 3516 17172 3547
rect 14047 3488 17172 3516
rect 14047 3485 14059 3488
rect 14001 3479 14059 3485
rect 10318 3448 10324 3460
rect 10279 3420 10324 3448
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 14461 3451 14519 3457
rect 14461 3448 14473 3451
rect 11716 3420 14473 3448
rect 9030 3380 9036 3392
rect 5224 3352 8892 3380
rect 8991 3352 9036 3380
rect 5224 3340 5230 3352
rect 9030 3340 9036 3352
rect 9088 3340 9094 3392
rect 9674 3340 9680 3392
rect 9732 3380 9738 3392
rect 11716 3380 11744 3420
rect 14461 3417 14473 3420
rect 14507 3417 14519 3451
rect 14461 3411 14519 3417
rect 14829 3451 14887 3457
rect 14829 3417 14841 3451
rect 14875 3448 14887 3451
rect 15654 3448 15660 3460
rect 14875 3420 15660 3448
rect 14875 3417 14887 3420
rect 14829 3411 14887 3417
rect 15654 3408 15660 3420
rect 15712 3408 15718 3460
rect 16666 3448 16672 3460
rect 16040 3420 16672 3448
rect 9732 3352 11744 3380
rect 12161 3383 12219 3389
rect 9732 3340 9738 3352
rect 12161 3349 12173 3383
rect 12207 3380 12219 3383
rect 12253 3383 12311 3389
rect 12253 3380 12265 3383
rect 12207 3352 12265 3380
rect 12207 3349 12219 3352
rect 12161 3343 12219 3349
rect 12253 3349 12265 3352
rect 12299 3349 12311 3383
rect 12253 3343 12311 3349
rect 12342 3340 12348 3392
rect 12400 3380 12406 3392
rect 14001 3383 14059 3389
rect 14001 3380 14013 3383
rect 12400 3352 14013 3380
rect 12400 3340 12406 3352
rect 14001 3349 14013 3352
rect 14047 3349 14059 3383
rect 14001 3343 14059 3349
rect 14277 3383 14335 3389
rect 14277 3349 14289 3383
rect 14323 3380 14335 3383
rect 16040 3380 16068 3420
rect 16666 3408 16672 3420
rect 16724 3408 16730 3460
rect 14323 3352 16068 3380
rect 14323 3349 14335 3352
rect 14277 3343 14335 3349
rect 16114 3340 16120 3392
rect 16172 3380 16178 3392
rect 17313 3383 17371 3389
rect 17313 3380 17325 3383
rect 16172 3352 17325 3380
rect 16172 3340 16178 3352
rect 17313 3349 17325 3352
rect 17359 3349 17371 3383
rect 18046 3380 18052 3392
rect 18007 3352 18052 3380
rect 17313 3343 17371 3349
rect 18046 3340 18052 3352
rect 18104 3340 18110 3392
rect 1104 3290 18860 3312
rect 1104 3238 3947 3290
rect 3999 3238 4011 3290
rect 4063 3238 4075 3290
rect 4127 3238 4139 3290
rect 4191 3238 9878 3290
rect 9930 3238 9942 3290
rect 9994 3238 10006 3290
rect 10058 3238 10070 3290
rect 10122 3238 15808 3290
rect 15860 3238 15872 3290
rect 15924 3238 15936 3290
rect 15988 3238 16000 3290
rect 16052 3238 18860 3290
rect 1104 3216 18860 3238
rect 2130 3136 2136 3188
rect 2188 3176 2194 3188
rect 5718 3176 5724 3188
rect 2188 3148 5724 3176
rect 2188 3136 2194 3148
rect 5718 3136 5724 3148
rect 5776 3136 5782 3188
rect 8386 3176 8392 3188
rect 7208 3148 8392 3176
rect 2406 3108 2412 3120
rect 2367 3080 2412 3108
rect 2406 3068 2412 3080
rect 2464 3068 2470 3120
rect 4982 3108 4988 3120
rect 2884 3080 4988 3108
rect 2884 3040 2912 3080
rect 4982 3068 4988 3080
rect 5040 3068 5046 3120
rect 7208 3040 7236 3148
rect 8386 3136 8392 3148
rect 8444 3136 8450 3188
rect 9030 3136 9036 3188
rect 9088 3176 9094 3188
rect 11790 3176 11796 3188
rect 9088 3148 11796 3176
rect 9088 3136 9094 3148
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 7282 3068 7288 3120
rect 7340 3108 7346 3120
rect 8113 3111 8171 3117
rect 8113 3108 8125 3111
rect 7340 3080 8125 3108
rect 7340 3068 7346 3080
rect 8113 3077 8125 3080
rect 8159 3077 8171 3111
rect 10778 3108 10784 3120
rect 8113 3071 8171 3077
rect 8496 3080 10784 3108
rect 1688 3012 2912 3040
rect 2976 3012 7236 3040
rect 7561 3043 7619 3049
rect 1688 2981 1716 3012
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2941 1731 2975
rect 1673 2935 1731 2941
rect 2225 2975 2283 2981
rect 2225 2941 2237 2975
rect 2271 2972 2283 2975
rect 2774 2972 2780 2984
rect 2271 2944 2780 2972
rect 2271 2941 2283 2944
rect 2225 2935 2283 2941
rect 2774 2932 2780 2944
rect 2832 2932 2838 2984
rect 2976 2981 3004 3012
rect 7561 3009 7573 3043
rect 7607 3040 7619 3043
rect 7607 3012 7972 3040
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 2961 2975 3019 2981
rect 2961 2941 2973 2975
rect 3007 2941 3019 2975
rect 2961 2935 3019 2941
rect 3697 2975 3755 2981
rect 3697 2941 3709 2975
rect 3743 2972 3755 2975
rect 4246 2972 4252 2984
rect 3743 2944 4252 2972
rect 3743 2941 3755 2944
rect 3697 2935 3755 2941
rect 4246 2932 4252 2944
rect 4304 2932 4310 2984
rect 6308 2975 6366 2981
rect 6308 2972 6320 2975
rect 6288 2941 6320 2972
rect 6354 2941 6366 2975
rect 6288 2935 6366 2941
rect 2682 2864 2688 2916
rect 2740 2904 2746 2916
rect 3237 2907 3295 2913
rect 3237 2904 3249 2907
rect 2740 2876 3249 2904
rect 2740 2864 2746 2876
rect 3237 2873 3249 2876
rect 3283 2873 3295 2907
rect 3237 2867 3295 2873
rect 1854 2836 1860 2848
rect 1815 2808 1860 2836
rect 1854 2796 1860 2808
rect 1912 2796 1918 2848
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 3881 2839 3939 2845
rect 3881 2836 3893 2839
rect 2832 2808 3893 2836
rect 2832 2796 2838 2808
rect 3881 2805 3893 2808
rect 3927 2805 3939 2839
rect 6288 2836 6316 2935
rect 6730 2932 6736 2984
rect 6788 2972 6794 2984
rect 6917 2975 6975 2981
rect 6917 2972 6929 2975
rect 6788 2944 6929 2972
rect 6788 2932 6794 2944
rect 6917 2941 6929 2944
rect 6963 2941 6975 2975
rect 6917 2935 6975 2941
rect 7285 2975 7343 2981
rect 7285 2941 7297 2975
rect 7331 2972 7343 2975
rect 7650 2972 7656 2984
rect 7331 2944 7656 2972
rect 7331 2941 7343 2944
rect 7285 2935 7343 2941
rect 7650 2932 7656 2944
rect 7708 2932 7714 2984
rect 7944 2981 7972 3012
rect 7929 2975 7987 2981
rect 7929 2941 7941 2975
rect 7975 2972 7987 2975
rect 8496 2972 8524 3080
rect 10778 3068 10784 3080
rect 10836 3068 10842 3120
rect 12250 3108 12256 3120
rect 10888 3080 12256 3108
rect 8662 3040 8668 3052
rect 8623 3012 8668 3040
rect 8662 3000 8668 3012
rect 8720 3000 8726 3052
rect 9122 3000 9128 3052
rect 9180 3040 9186 3052
rect 9674 3040 9680 3052
rect 9180 3012 9536 3040
rect 9635 3012 9680 3040
rect 9180 3000 9186 3012
rect 7975 2944 8524 2972
rect 9508 2972 9536 3012
rect 9674 3000 9680 3012
rect 9732 3000 9738 3052
rect 10888 3040 10916 3080
rect 12250 3068 12256 3080
rect 12308 3068 12314 3120
rect 12526 3068 12532 3120
rect 12584 3108 12590 3120
rect 12584 3080 18092 3108
rect 12584 3068 12590 3080
rect 9784 3012 10916 3040
rect 11701 3043 11759 3049
rect 9784 2972 9812 3012
rect 11701 3009 11713 3043
rect 11747 3040 11759 3043
rect 12342 3040 12348 3052
rect 11747 3012 12348 3040
rect 11747 3009 11759 3012
rect 11701 3003 11759 3009
rect 12342 3000 12348 3012
rect 12400 3000 12406 3052
rect 12618 3000 12624 3052
rect 12676 3040 12682 3052
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12676 3012 13001 3040
rect 12676 3000 12682 3012
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 14001 3043 14059 3049
rect 14001 3009 14013 3043
rect 14047 3040 14059 3043
rect 14090 3040 14096 3052
rect 14047 3012 14096 3040
rect 14047 3009 14059 3012
rect 14001 3003 14059 3009
rect 14090 3000 14096 3012
rect 14148 3000 14154 3052
rect 14366 3040 14372 3052
rect 14327 3012 14372 3040
rect 14366 3000 14372 3012
rect 14424 3000 14430 3052
rect 14734 3000 14740 3052
rect 14792 3040 14798 3052
rect 15841 3043 15899 3049
rect 15841 3040 15853 3043
rect 14792 3012 15853 3040
rect 14792 3000 14798 3012
rect 15841 3009 15853 3012
rect 15887 3009 15899 3043
rect 15841 3003 15899 3009
rect 16206 3000 16212 3052
rect 16264 3040 16270 3052
rect 17126 3040 17132 3052
rect 16264 3012 17132 3040
rect 16264 3000 16270 3012
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 9508 2944 9812 2972
rect 9953 2975 10011 2981
rect 7975 2941 7987 2944
rect 7929 2935 7987 2941
rect 9953 2941 9965 2975
rect 9999 2972 10011 2975
rect 10410 2972 10416 2984
rect 9999 2944 10416 2972
rect 9999 2941 10011 2944
rect 9953 2935 10011 2941
rect 10410 2932 10416 2944
rect 10468 2932 10474 2984
rect 12472 2975 12530 2981
rect 12472 2972 12484 2975
rect 11716 2944 12484 2972
rect 6411 2907 6469 2913
rect 6411 2873 6423 2907
rect 6457 2904 6469 2907
rect 8202 2904 8208 2916
rect 6457 2876 8208 2904
rect 6457 2873 6469 2876
rect 6411 2867 6469 2873
rect 8202 2864 8208 2876
rect 8260 2864 8266 2916
rect 8757 2907 8815 2913
rect 8757 2873 8769 2907
rect 8803 2873 8815 2907
rect 8757 2867 8815 2873
rect 7834 2836 7840 2848
rect 6288 2808 7840 2836
rect 3881 2799 3939 2805
rect 7834 2796 7840 2808
rect 7892 2836 7898 2848
rect 8772 2836 8800 2867
rect 9490 2864 9496 2916
rect 9548 2904 9554 2916
rect 10689 2907 10747 2913
rect 10689 2904 10701 2907
rect 9548 2876 10701 2904
rect 9548 2864 9554 2876
rect 10689 2873 10701 2876
rect 10735 2873 10747 2907
rect 10689 2867 10747 2873
rect 10778 2864 10784 2916
rect 10836 2904 10842 2916
rect 10836 2876 10929 2904
rect 10836 2864 10842 2876
rect 7892 2808 8800 2836
rect 7892 2796 7898 2808
rect 9122 2796 9128 2848
rect 9180 2836 9186 2848
rect 10137 2839 10195 2845
rect 10137 2836 10149 2839
rect 9180 2808 10149 2836
rect 9180 2796 9186 2808
rect 10137 2805 10149 2808
rect 10183 2805 10195 2839
rect 10796 2836 10824 2864
rect 11716 2836 11744 2944
rect 12472 2941 12484 2944
rect 12518 2941 12530 2975
rect 12472 2935 12530 2941
rect 17218 2932 17224 2984
rect 17276 2972 17282 2984
rect 18064 2981 18092 3080
rect 17405 2975 17463 2981
rect 17405 2972 17417 2975
rect 17276 2944 17417 2972
rect 17276 2932 17282 2944
rect 17405 2941 17417 2944
rect 17451 2941 17463 2975
rect 17405 2935 17463 2941
rect 18049 2975 18107 2981
rect 18049 2941 18061 2975
rect 18095 2941 18107 2975
rect 18049 2935 18107 2941
rect 11790 2864 11796 2916
rect 11848 2904 11854 2916
rect 13081 2907 13139 2913
rect 11848 2876 13032 2904
rect 11848 2864 11854 2876
rect 10796 2808 11744 2836
rect 10137 2799 10195 2805
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 12575 2839 12633 2845
rect 12575 2836 12587 2839
rect 12492 2808 12587 2836
rect 12492 2796 12498 2808
rect 12575 2805 12587 2808
rect 12621 2805 12633 2839
rect 13004 2836 13032 2876
rect 13081 2873 13093 2907
rect 13127 2904 13139 2907
rect 13170 2904 13176 2916
rect 13127 2876 13176 2904
rect 13127 2873 13139 2876
rect 13081 2867 13139 2873
rect 13170 2864 13176 2876
rect 13228 2864 13234 2916
rect 14461 2907 14519 2913
rect 14461 2873 14473 2907
rect 14507 2873 14519 2907
rect 14461 2867 14519 2873
rect 15381 2907 15439 2913
rect 15381 2873 15393 2907
rect 15427 2873 15439 2907
rect 15381 2867 15439 2873
rect 14476 2836 14504 2867
rect 15102 2836 15108 2848
rect 13004 2808 15108 2836
rect 12575 2799 12633 2805
rect 15102 2796 15108 2808
rect 15160 2796 15166 2848
rect 15194 2796 15200 2848
rect 15252 2836 15258 2848
rect 15396 2836 15424 2867
rect 15930 2864 15936 2916
rect 15988 2904 15994 2916
rect 15988 2876 16033 2904
rect 15988 2864 15994 2876
rect 16758 2864 16764 2916
rect 16816 2904 16822 2916
rect 16853 2907 16911 2913
rect 16853 2904 16865 2907
rect 16816 2876 16865 2904
rect 16816 2864 16822 2876
rect 16853 2873 16865 2876
rect 16899 2873 16911 2907
rect 16853 2867 16911 2873
rect 17586 2836 17592 2848
rect 15252 2808 15424 2836
rect 17547 2808 17592 2836
rect 15252 2796 15258 2808
rect 17586 2796 17592 2808
rect 17644 2796 17650 2848
rect 17862 2796 17868 2848
rect 17920 2836 17926 2848
rect 18233 2839 18291 2845
rect 18233 2836 18245 2839
rect 17920 2808 18245 2836
rect 17920 2796 17926 2808
rect 18233 2805 18245 2808
rect 18279 2805 18291 2839
rect 18233 2799 18291 2805
rect 1104 2746 18860 2768
rect 1104 2694 6912 2746
rect 6964 2694 6976 2746
rect 7028 2694 7040 2746
rect 7092 2694 7104 2746
rect 7156 2694 12843 2746
rect 12895 2694 12907 2746
rect 12959 2694 12971 2746
rect 13023 2694 13035 2746
rect 13087 2694 18860 2746
rect 1104 2672 18860 2694
rect 6638 2592 6644 2644
rect 6696 2632 6702 2644
rect 8113 2635 8171 2641
rect 8113 2632 8125 2635
rect 6696 2604 8125 2632
rect 6696 2592 6702 2604
rect 8113 2601 8125 2604
rect 8159 2601 8171 2635
rect 8113 2595 8171 2601
rect 8849 2635 8907 2641
rect 8849 2601 8861 2635
rect 8895 2632 8907 2635
rect 8895 2604 13124 2632
rect 8895 2601 8907 2604
rect 8849 2595 8907 2601
rect 13096 2576 13124 2604
rect 15010 2592 15016 2644
rect 15068 2641 15074 2644
rect 15068 2635 15117 2641
rect 15068 2601 15071 2635
rect 15105 2601 15117 2635
rect 15068 2595 15117 2601
rect 15212 2604 17172 2632
rect 15068 2592 15074 2595
rect 1670 2524 1676 2576
rect 1728 2564 1734 2576
rect 3329 2567 3387 2573
rect 3329 2564 3341 2567
rect 1728 2536 3341 2564
rect 1728 2524 1734 2536
rect 3329 2533 3341 2536
rect 3375 2533 3387 2567
rect 3329 2527 3387 2533
rect 5718 2524 5724 2576
rect 5776 2564 5782 2576
rect 6273 2567 6331 2573
rect 6273 2564 6285 2567
rect 5776 2536 6285 2564
rect 5776 2524 5782 2536
rect 6273 2533 6285 2536
rect 6319 2533 6331 2567
rect 7558 2564 7564 2576
rect 6273 2527 6331 2533
rect 7208 2536 7564 2564
rect 1486 2456 1492 2508
rect 1544 2496 1550 2508
rect 1581 2499 1639 2505
rect 1581 2496 1593 2499
rect 1544 2468 1593 2496
rect 1544 2456 1550 2468
rect 1581 2465 1593 2468
rect 1627 2465 1639 2499
rect 1581 2459 1639 2465
rect 2317 2499 2375 2505
rect 2317 2465 2329 2499
rect 2363 2496 2375 2499
rect 3053 2499 3111 2505
rect 2363 2468 3004 2496
rect 2363 2465 2375 2468
rect 2317 2459 2375 2465
rect 658 2388 664 2440
rect 716 2428 722 2440
rect 1765 2431 1823 2437
rect 1765 2428 1777 2431
rect 716 2400 1777 2428
rect 716 2388 722 2400
rect 1765 2397 1777 2400
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2397 2559 2431
rect 2976 2428 3004 2468
rect 3053 2465 3065 2499
rect 3099 2496 3111 2499
rect 3418 2496 3424 2508
rect 3099 2468 3424 2496
rect 3099 2465 3111 2468
rect 3053 2459 3111 2465
rect 3418 2456 3424 2468
rect 3476 2456 3482 2508
rect 4065 2499 4123 2505
rect 4065 2465 4077 2499
rect 4111 2496 4123 2499
rect 5442 2496 5448 2508
rect 4111 2468 5448 2496
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 5442 2456 5448 2468
rect 5500 2456 5506 2508
rect 5604 2499 5662 2505
rect 5604 2465 5616 2499
rect 5650 2496 5662 2499
rect 5810 2496 5816 2508
rect 5650 2468 5816 2496
rect 5650 2465 5662 2468
rect 5604 2459 5662 2465
rect 5810 2456 5816 2468
rect 5868 2456 5874 2508
rect 5997 2499 6055 2505
rect 5997 2465 6009 2499
rect 6043 2496 6055 2499
rect 7208 2496 7236 2536
rect 7558 2524 7564 2536
rect 7616 2524 7622 2576
rect 7653 2567 7711 2573
rect 7653 2533 7665 2567
rect 7699 2564 7711 2567
rect 7699 2536 8156 2564
rect 7699 2533 7711 2536
rect 7653 2527 7711 2533
rect 6043 2468 7236 2496
rect 7285 2499 7343 2505
rect 6043 2465 6055 2468
rect 5997 2459 6055 2465
rect 7285 2465 7297 2499
rect 7331 2496 7343 2499
rect 7466 2496 7472 2508
rect 7331 2468 7472 2496
rect 7331 2465 7343 2468
rect 7285 2459 7343 2465
rect 7466 2456 7472 2468
rect 7524 2456 7530 2508
rect 7834 2456 7840 2508
rect 7892 2496 7898 2508
rect 7929 2499 7987 2505
rect 7929 2496 7941 2499
rect 7892 2468 7941 2496
rect 7892 2456 7898 2468
rect 7929 2465 7941 2468
rect 7975 2465 7987 2499
rect 8128 2496 8156 2536
rect 8202 2524 8208 2576
rect 8260 2564 8266 2576
rect 9953 2567 10011 2573
rect 9953 2564 9965 2567
rect 8260 2536 9965 2564
rect 8260 2524 8266 2536
rect 9953 2533 9965 2536
rect 9999 2533 10011 2567
rect 9953 2527 10011 2533
rect 10686 2524 10692 2576
rect 10744 2564 10750 2576
rect 10873 2567 10931 2573
rect 10873 2564 10885 2567
rect 10744 2536 10885 2564
rect 10744 2524 10750 2536
rect 10873 2533 10885 2536
rect 10919 2533 10931 2567
rect 10873 2527 10931 2533
rect 11333 2567 11391 2573
rect 11333 2533 11345 2567
rect 11379 2564 11391 2567
rect 12434 2564 12440 2576
rect 11379 2536 12440 2564
rect 11379 2533 11391 2536
rect 11333 2527 11391 2533
rect 12434 2524 12440 2536
rect 12492 2524 12498 2576
rect 13078 2524 13084 2576
rect 13136 2524 13142 2576
rect 13173 2567 13231 2573
rect 13173 2533 13185 2567
rect 13219 2564 13231 2567
rect 13906 2564 13912 2576
rect 13219 2536 13912 2564
rect 13219 2533 13231 2536
rect 13173 2527 13231 2533
rect 13906 2524 13912 2536
rect 13964 2524 13970 2576
rect 14093 2567 14151 2573
rect 14093 2533 14105 2567
rect 14139 2564 14151 2567
rect 14182 2564 14188 2576
rect 14139 2536 14188 2564
rect 14139 2533 14151 2536
rect 14093 2527 14151 2533
rect 14182 2524 14188 2536
rect 14240 2524 14246 2576
rect 14737 2567 14795 2573
rect 14737 2564 14749 2567
rect 14384 2536 14749 2564
rect 8481 2499 8539 2505
rect 8481 2496 8493 2499
rect 8128 2468 8493 2496
rect 7929 2459 7987 2465
rect 8481 2465 8493 2468
rect 8527 2496 8539 2499
rect 8849 2499 8907 2505
rect 8849 2496 8861 2499
rect 8527 2468 8861 2496
rect 8527 2465 8539 2468
rect 8481 2459 8539 2465
rect 8849 2465 8861 2468
rect 8895 2465 8907 2499
rect 9030 2496 9036 2508
rect 8991 2468 9036 2496
rect 8849 2459 8907 2465
rect 9030 2456 9036 2468
rect 9088 2456 9094 2508
rect 14384 2505 14412 2536
rect 14737 2533 14749 2536
rect 14783 2533 14795 2567
rect 14737 2527 14795 2533
rect 14826 2524 14832 2576
rect 14884 2564 14890 2576
rect 15212 2564 15240 2604
rect 14884 2536 15240 2564
rect 14884 2524 14890 2536
rect 15286 2524 15292 2576
rect 15344 2564 15350 2576
rect 15657 2567 15715 2573
rect 15657 2564 15669 2567
rect 15344 2536 15669 2564
rect 15344 2524 15350 2536
rect 15657 2533 15669 2536
rect 15703 2533 15715 2567
rect 15657 2527 15715 2533
rect 17144 2505 17172 2604
rect 14369 2499 14427 2505
rect 14369 2465 14381 2499
rect 14415 2465 14427 2499
rect 14956 2499 15014 2505
rect 14956 2496 14968 2499
rect 14369 2459 14427 2465
rect 14476 2468 14968 2496
rect 3234 2428 3240 2440
rect 2976 2400 3240 2428
rect 2501 2391 2559 2397
rect 1118 2320 1124 2372
rect 1176 2360 1182 2372
rect 2516 2360 2544 2391
rect 3234 2388 3240 2400
rect 3292 2388 3298 2440
rect 3602 2388 3608 2440
rect 3660 2428 3666 2440
rect 4249 2431 4307 2437
rect 4249 2428 4261 2431
rect 3660 2400 4261 2428
rect 3660 2388 3666 2400
rect 4249 2397 4261 2400
rect 4295 2397 4307 2431
rect 4249 2391 4307 2397
rect 6730 2388 6736 2440
rect 6788 2428 6794 2440
rect 6917 2431 6975 2437
rect 6917 2428 6929 2431
rect 6788 2400 6929 2428
rect 6788 2388 6794 2400
rect 6917 2397 6929 2400
rect 6963 2428 6975 2431
rect 8570 2428 8576 2440
rect 6963 2400 8576 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 8570 2388 8576 2400
rect 8628 2388 8634 2440
rect 9861 2431 9919 2437
rect 9861 2397 9873 2431
rect 9907 2428 9919 2431
rect 11054 2428 11060 2440
rect 9907 2400 11060 2428
rect 9907 2397 9919 2400
rect 9861 2391 9919 2397
rect 11054 2388 11060 2400
rect 11112 2388 11118 2440
rect 11241 2431 11299 2437
rect 11241 2397 11253 2431
rect 11287 2428 11299 2431
rect 11606 2428 11612 2440
rect 11287 2400 11612 2428
rect 11287 2397 11299 2400
rect 11241 2391 11299 2397
rect 11606 2388 11612 2400
rect 11664 2388 11670 2440
rect 12066 2428 12072 2440
rect 12027 2400 12072 2428
rect 12066 2388 12072 2400
rect 12124 2388 12130 2440
rect 12618 2388 12624 2440
rect 12676 2428 12682 2440
rect 13081 2431 13139 2437
rect 13081 2428 13093 2431
rect 12676 2400 13093 2428
rect 12676 2388 12682 2400
rect 13081 2397 13093 2400
rect 13127 2397 13139 2431
rect 13081 2391 13139 2397
rect 13170 2388 13176 2440
rect 13228 2428 13234 2440
rect 14476 2428 14504 2468
rect 14956 2465 14968 2468
rect 15002 2465 15014 2499
rect 14956 2459 15014 2465
rect 17129 2499 17187 2505
rect 17129 2465 17141 2499
rect 17175 2465 17187 2499
rect 17681 2499 17739 2505
rect 17681 2496 17693 2499
rect 17129 2459 17187 2465
rect 17420 2468 17693 2496
rect 13228 2400 14504 2428
rect 13228 2388 13234 2400
rect 15102 2388 15108 2440
rect 15160 2428 15166 2440
rect 15565 2431 15623 2437
rect 15565 2428 15577 2431
rect 15160 2400 15577 2428
rect 15160 2388 15166 2400
rect 15565 2397 15577 2400
rect 15611 2397 15623 2431
rect 15838 2428 15844 2440
rect 15799 2400 15844 2428
rect 15565 2391 15623 2397
rect 15838 2388 15844 2400
rect 15896 2388 15902 2440
rect 16942 2388 16948 2440
rect 17000 2428 17006 2440
rect 17420 2428 17448 2468
rect 17681 2465 17693 2468
rect 17727 2465 17739 2499
rect 17681 2459 17739 2465
rect 17000 2400 17448 2428
rect 17000 2388 17006 2400
rect 17586 2388 17592 2440
rect 17644 2428 17650 2440
rect 17862 2428 17868 2440
rect 17644 2400 17868 2428
rect 17644 2388 17650 2400
rect 17862 2388 17868 2400
rect 17920 2388 17926 2440
rect 1176 2332 2544 2360
rect 1176 2320 1182 2332
rect 7650 2320 7656 2372
rect 7708 2360 7714 2372
rect 8665 2363 8723 2369
rect 8665 2360 8677 2363
rect 7708 2332 8677 2360
rect 7708 2320 7714 2332
rect 8665 2329 8677 2332
rect 8711 2329 8723 2363
rect 8665 2323 8723 2329
rect 10318 2320 10324 2372
rect 10376 2360 10382 2372
rect 10376 2332 14780 2360
rect 10376 2320 10382 2332
rect 5675 2295 5733 2301
rect 5675 2261 5687 2295
rect 5721 2292 5733 2295
rect 8110 2292 8116 2304
rect 5721 2264 8116 2292
rect 5721 2261 5733 2264
rect 5675 2255 5733 2261
rect 8110 2252 8116 2264
rect 8168 2252 8174 2304
rect 8202 2252 8208 2304
rect 8260 2292 8266 2304
rect 9217 2295 9275 2301
rect 9217 2292 9229 2295
rect 8260 2264 9229 2292
rect 8260 2252 8266 2264
rect 9217 2261 9229 2264
rect 9263 2261 9275 2295
rect 9217 2255 9275 2261
rect 10594 2252 10600 2304
rect 10652 2292 10658 2304
rect 14752 2301 14780 2332
rect 15930 2320 15936 2372
rect 15988 2320 15994 2372
rect 14553 2295 14611 2301
rect 14553 2292 14565 2295
rect 10652 2264 14565 2292
rect 10652 2252 10658 2264
rect 14553 2261 14565 2264
rect 14599 2261 14611 2295
rect 14553 2255 14611 2261
rect 14737 2295 14795 2301
rect 14737 2261 14749 2295
rect 14783 2292 14795 2295
rect 15948 2292 15976 2320
rect 17310 2292 17316 2304
rect 14783 2264 15976 2292
rect 17271 2264 17316 2292
rect 14783 2261 14795 2264
rect 14737 2255 14795 2261
rect 17310 2252 17316 2264
rect 17368 2252 17374 2304
rect 17862 2292 17868 2304
rect 17823 2264 17868 2292
rect 17862 2252 17868 2264
rect 17920 2252 17926 2304
rect 1104 2202 18860 2224
rect 1104 2150 3947 2202
rect 3999 2150 4011 2202
rect 4063 2150 4075 2202
rect 4127 2150 4139 2202
rect 4191 2150 9878 2202
rect 9930 2150 9942 2202
rect 9994 2150 10006 2202
rect 10058 2150 10070 2202
rect 10122 2150 15808 2202
rect 15860 2150 15872 2202
rect 15924 2150 15936 2202
rect 15988 2150 16000 2202
rect 16052 2150 18860 2202
rect 1104 2128 18860 2150
rect 5442 2048 5448 2100
rect 5500 2088 5506 2100
rect 14458 2088 14464 2100
rect 5500 2060 14464 2088
rect 5500 2048 5506 2060
rect 14458 2048 14464 2060
rect 14516 2048 14522 2100
rect 8110 1980 8116 2032
rect 8168 2020 8174 2032
rect 15286 2020 15292 2032
rect 8168 1992 15292 2020
rect 8168 1980 8174 1992
rect 15286 1980 15292 1992
rect 15344 1980 15350 2032
rect 5810 1912 5816 1964
rect 5868 1952 5874 1964
rect 10318 1952 10324 1964
rect 5868 1924 10324 1952
rect 5868 1912 5874 1924
rect 10318 1912 10324 1924
rect 10376 1912 10382 1964
rect 13446 1912 13452 1964
rect 13504 1952 13510 1964
rect 18138 1952 18144 1964
rect 13504 1924 18144 1952
rect 13504 1912 13510 1924
rect 18138 1912 18144 1924
rect 18196 1912 18202 1964
rect 13998 1708 14004 1760
rect 14056 1748 14062 1760
rect 17586 1748 17592 1760
rect 14056 1720 17592 1748
rect 14056 1708 14062 1720
rect 17586 1708 17592 1720
rect 17644 1708 17650 1760
rect 12710 1640 12716 1692
rect 12768 1680 12774 1692
rect 19150 1680 19156 1692
rect 12768 1652 19156 1680
rect 12768 1640 12774 1652
rect 19150 1640 19156 1652
rect 19208 1640 19214 1692
<< via1 >>
rect 3608 15240 3660 15292
rect 4344 15240 4396 15292
rect 4068 15172 4120 15224
rect 7288 15172 7340 15224
rect 6912 14662 6964 14714
rect 6976 14662 7028 14714
rect 7040 14662 7092 14714
rect 7104 14662 7156 14714
rect 12843 14662 12895 14714
rect 12907 14662 12959 14714
rect 12971 14662 13023 14714
rect 13035 14662 13087 14714
rect 1584 14560 1636 14612
rect 13912 14492 13964 14544
rect 18328 14492 18380 14544
rect 2596 14356 2648 14408
rect 11060 14424 11112 14476
rect 9956 14356 10008 14408
rect 12440 14356 12492 14408
rect 3332 14288 3384 14340
rect 14004 14288 14056 14340
rect 2780 14220 2832 14272
rect 14188 14220 14240 14272
rect 3947 14118 3999 14170
rect 4011 14118 4063 14170
rect 4075 14118 4127 14170
rect 4139 14118 4191 14170
rect 9878 14118 9930 14170
rect 9942 14118 9994 14170
rect 10006 14118 10058 14170
rect 10070 14118 10122 14170
rect 15808 14118 15860 14170
rect 15872 14118 15924 14170
rect 15936 14118 15988 14170
rect 16000 14118 16052 14170
rect 296 14016 348 14068
rect 940 13948 992 14000
rect 2872 14016 2924 14068
rect 6920 14016 6972 14068
rect 2228 13948 2280 14000
rect 6276 13948 6328 14000
rect 13544 13948 13596 14000
rect 15660 13948 15712 14000
rect 10692 13880 10744 13932
rect 2596 13812 2648 13864
rect 2780 13855 2832 13864
rect 2780 13821 2789 13855
rect 2789 13821 2823 13855
rect 2823 13821 2832 13855
rect 3332 13855 3384 13864
rect 2780 13812 2832 13821
rect 3332 13821 3341 13855
rect 3341 13821 3375 13855
rect 3375 13821 3384 13855
rect 3332 13812 3384 13821
rect 6092 13812 6144 13864
rect 6552 13812 6604 13864
rect 14372 13812 14424 13864
rect 15016 13812 15068 13864
rect 16212 13880 16264 13932
rect 15384 13812 15436 13864
rect 16396 13812 16448 13864
rect 7380 13744 7432 13796
rect 9220 13744 9272 13796
rect 14832 13744 14884 13796
rect 3516 13676 3568 13728
rect 15292 13719 15344 13728
rect 15292 13685 15301 13719
rect 15301 13685 15335 13719
rect 15335 13685 15344 13719
rect 15292 13676 15344 13685
rect 15844 13719 15896 13728
rect 15844 13685 15853 13719
rect 15853 13685 15887 13719
rect 15887 13685 15896 13719
rect 15844 13676 15896 13685
rect 6912 13574 6964 13626
rect 6976 13574 7028 13626
rect 7040 13574 7092 13626
rect 7104 13574 7156 13626
rect 12843 13574 12895 13626
rect 12907 13574 12959 13626
rect 12971 13574 13023 13626
rect 13035 13574 13087 13626
rect 4804 13472 4856 13524
rect 15292 13472 15344 13524
rect 4252 13404 4304 13456
rect 13544 13404 13596 13456
rect 14188 13404 14240 13456
rect 18972 13404 19024 13456
rect 2228 13379 2280 13388
rect 2228 13345 2237 13379
rect 2237 13345 2271 13379
rect 2271 13345 2280 13379
rect 2228 13336 2280 13345
rect 5448 13336 5500 13388
rect 15844 13336 15896 13388
rect 2320 13311 2372 13320
rect 2320 13277 2329 13311
rect 2329 13277 2363 13311
rect 2363 13277 2372 13311
rect 2320 13268 2372 13277
rect 2504 13311 2556 13320
rect 2504 13277 2513 13311
rect 2513 13277 2547 13311
rect 2547 13277 2556 13311
rect 2504 13268 2556 13277
rect 10692 13268 10744 13320
rect 17040 13268 17092 13320
rect 3424 13200 3476 13252
rect 10876 13200 10928 13252
rect 11060 13200 11112 13252
rect 12072 13200 12124 13252
rect 3608 13132 3660 13184
rect 13820 13200 13872 13252
rect 15016 13200 15068 13252
rect 17684 13132 17736 13184
rect 3947 13030 3999 13082
rect 4011 13030 4063 13082
rect 4075 13030 4127 13082
rect 4139 13030 4191 13082
rect 9878 13030 9930 13082
rect 9942 13030 9994 13082
rect 10006 13030 10058 13082
rect 10070 13030 10122 13082
rect 15808 13030 15860 13082
rect 15872 13030 15924 13082
rect 15936 13030 15988 13082
rect 16000 13030 16052 13082
rect 2320 12928 2372 12980
rect 5264 12928 5316 12980
rect 14004 12928 14056 12980
rect 19616 12928 19668 12980
rect 3516 12860 3568 12912
rect 6368 12860 6420 12912
rect 2596 12792 2648 12844
rect 4620 12792 4672 12844
rect 4712 12792 4764 12844
rect 7656 12792 7708 12844
rect 3608 12767 3660 12776
rect 3608 12733 3617 12767
rect 3617 12733 3651 12767
rect 3651 12733 3660 12767
rect 3608 12724 3660 12733
rect 4896 12767 4948 12776
rect 4896 12733 4905 12767
rect 4905 12733 4939 12767
rect 4939 12733 4948 12767
rect 4896 12724 4948 12733
rect 3424 12656 3476 12708
rect 13728 12792 13780 12844
rect 15200 12724 15252 12776
rect 15568 12724 15620 12776
rect 2780 12588 2832 12640
rect 3148 12588 3200 12640
rect 3700 12631 3752 12640
rect 3700 12597 3709 12631
rect 3709 12597 3743 12631
rect 3743 12597 3752 12631
rect 3700 12588 3752 12597
rect 4068 12588 4120 12640
rect 10600 12656 10652 12708
rect 14372 12656 14424 12708
rect 6912 12486 6964 12538
rect 6976 12486 7028 12538
rect 7040 12486 7092 12538
rect 7104 12486 7156 12538
rect 12843 12486 12895 12538
rect 12907 12486 12959 12538
rect 12971 12486 13023 12538
rect 13035 12486 13087 12538
rect 2320 12384 2372 12436
rect 2504 12384 2556 12436
rect 2596 12359 2648 12368
rect 2596 12325 2630 12359
rect 2630 12325 2648 12359
rect 2596 12316 2648 12325
rect 2688 12316 2740 12368
rect 3608 12248 3660 12300
rect 3792 12248 3844 12300
rect 4620 12316 4672 12368
rect 15568 12384 15620 12436
rect 6184 12316 6236 12368
rect 15384 12316 15436 12368
rect 1860 12223 1912 12232
rect 1860 12189 1869 12223
rect 1869 12189 1903 12223
rect 1903 12189 1912 12223
rect 1860 12180 1912 12189
rect 5448 12180 5500 12232
rect 2688 12044 2740 12096
rect 3792 12044 3844 12096
rect 7748 12112 7800 12164
rect 13176 12248 13228 12300
rect 14556 12248 14608 12300
rect 12164 12180 12216 12232
rect 16396 12180 16448 12232
rect 16580 12112 16632 12164
rect 7380 12044 7432 12096
rect 10600 12044 10652 12096
rect 16488 12044 16540 12096
rect 3947 11942 3999 11994
rect 4011 11942 4063 11994
rect 4075 11942 4127 11994
rect 4139 11942 4191 11994
rect 9878 11942 9930 11994
rect 9942 11942 9994 11994
rect 10006 11942 10058 11994
rect 10070 11942 10122 11994
rect 15808 11942 15860 11994
rect 15872 11942 15924 11994
rect 15936 11942 15988 11994
rect 16000 11942 16052 11994
rect 2228 11883 2280 11892
rect 2228 11849 2237 11883
rect 2237 11849 2271 11883
rect 2271 11849 2280 11883
rect 2228 11840 2280 11849
rect 3792 11840 3844 11892
rect 2596 11772 2648 11824
rect 2688 11772 2740 11824
rect 4620 11840 4672 11892
rect 4988 11840 5040 11892
rect 5816 11840 5868 11892
rect 17776 11840 17828 11892
rect 6092 11772 6144 11824
rect 17316 11772 17368 11824
rect 5264 11704 5316 11756
rect 8116 11704 8168 11756
rect 1860 11636 1912 11688
rect 3056 11636 3108 11688
rect 5356 11636 5408 11688
rect 2320 11568 2372 11620
rect 1768 11500 1820 11552
rect 5540 11568 5592 11620
rect 7840 11679 7892 11688
rect 7840 11645 7849 11679
rect 7849 11645 7883 11679
rect 7883 11645 7892 11679
rect 7840 11636 7892 11645
rect 10324 11704 10376 11756
rect 10968 11704 11020 11756
rect 9680 11636 9732 11688
rect 11152 11636 11204 11688
rect 9036 11568 9088 11620
rect 9404 11568 9456 11620
rect 10784 11568 10836 11620
rect 15476 11568 15528 11620
rect 7840 11500 7892 11552
rect 8300 11500 8352 11552
rect 12532 11500 12584 11552
rect 13176 11500 13228 11552
rect 6912 11398 6964 11450
rect 6976 11398 7028 11450
rect 7040 11398 7092 11450
rect 7104 11398 7156 11450
rect 12843 11398 12895 11450
rect 12907 11398 12959 11450
rect 12971 11398 13023 11450
rect 13035 11398 13087 11450
rect 3700 11296 3752 11348
rect 5080 11296 5132 11348
rect 6092 11339 6144 11348
rect 6092 11305 6101 11339
rect 6101 11305 6135 11339
rect 6135 11305 6144 11339
rect 6092 11296 6144 11305
rect 2412 11228 2464 11280
rect 2688 11228 2740 11280
rect 2780 11228 2832 11280
rect 10784 11296 10836 11348
rect 6736 11228 6788 11280
rect 2044 11203 2096 11212
rect 2044 11169 2053 11203
rect 2053 11169 2087 11203
rect 2087 11169 2096 11203
rect 2044 11160 2096 11169
rect 3056 11203 3108 11212
rect 3056 11169 3065 11203
rect 3065 11169 3099 11203
rect 3099 11169 3108 11203
rect 3056 11160 3108 11169
rect 4988 11203 5040 11212
rect 4988 11169 4997 11203
rect 4997 11169 5031 11203
rect 5031 11169 5040 11203
rect 4988 11160 5040 11169
rect 5908 11160 5960 11212
rect 2136 11135 2188 11144
rect 2136 11101 2145 11135
rect 2145 11101 2179 11135
rect 2179 11101 2188 11135
rect 2136 11092 2188 11101
rect 2320 11135 2372 11144
rect 2320 11101 2329 11135
rect 2329 11101 2363 11135
rect 2363 11101 2372 11135
rect 2320 11092 2372 11101
rect 2504 11092 2556 11144
rect 1676 11024 1728 11076
rect 2780 11024 2832 11076
rect 2964 11092 3016 11144
rect 3424 11092 3476 11144
rect 5264 11135 5316 11144
rect 5264 11101 5273 11135
rect 5273 11101 5307 11135
rect 5307 11101 5316 11135
rect 5264 11092 5316 11101
rect 5816 11092 5868 11144
rect 7380 11160 7432 11212
rect 9772 11160 9824 11212
rect 10324 11160 10376 11212
rect 12624 11160 12676 11212
rect 13268 11160 13320 11212
rect 18052 11160 18104 11212
rect 6184 11135 6236 11144
rect 6184 11101 6193 11135
rect 6193 11101 6227 11135
rect 6227 11101 6236 11135
rect 6184 11092 6236 11101
rect 6644 11092 6696 11144
rect 12348 11135 12400 11144
rect 12348 11101 12357 11135
rect 12357 11101 12391 11135
rect 12391 11101 12400 11135
rect 12348 11092 12400 11101
rect 12440 11092 12492 11144
rect 15200 11092 15252 11144
rect 15476 11092 15528 11144
rect 5448 11024 5500 11076
rect 10968 11024 11020 11076
rect 1860 10956 1912 11008
rect 5632 10999 5684 11008
rect 5632 10965 5641 10999
rect 5641 10965 5675 10999
rect 5675 10965 5684 10999
rect 5632 10956 5684 10965
rect 8116 10999 8168 11008
rect 8116 10965 8125 10999
rect 8125 10965 8159 10999
rect 8159 10965 8168 10999
rect 8116 10956 8168 10965
rect 8208 10956 8260 11008
rect 11520 10999 11572 11008
rect 11520 10965 11529 10999
rect 11529 10965 11563 10999
rect 11563 10965 11572 10999
rect 11520 10956 11572 10965
rect 12164 10956 12216 11008
rect 13636 10956 13688 11008
rect 14280 10956 14332 11008
rect 15568 10956 15620 11008
rect 17868 10956 17920 11008
rect 3947 10854 3999 10906
rect 4011 10854 4063 10906
rect 4075 10854 4127 10906
rect 4139 10854 4191 10906
rect 9878 10854 9930 10906
rect 9942 10854 9994 10906
rect 10006 10854 10058 10906
rect 10070 10854 10122 10906
rect 15808 10854 15860 10906
rect 15872 10854 15924 10906
rect 15936 10854 15988 10906
rect 16000 10854 16052 10906
rect 2044 10752 2096 10804
rect 4988 10752 5040 10804
rect 7656 10752 7708 10804
rect 9404 10795 9456 10804
rect 9404 10761 9413 10795
rect 9413 10761 9447 10795
rect 9447 10761 9456 10795
rect 9404 10752 9456 10761
rect 5540 10684 5592 10736
rect 1860 10659 1912 10668
rect 1860 10625 1869 10659
rect 1869 10625 1903 10659
rect 1903 10625 1912 10659
rect 1860 10616 1912 10625
rect 2044 10659 2096 10668
rect 2044 10625 2053 10659
rect 2053 10625 2087 10659
rect 2087 10625 2096 10659
rect 2044 10616 2096 10625
rect 2412 10591 2464 10600
rect 2412 10557 2421 10591
rect 2421 10557 2455 10591
rect 2455 10557 2464 10591
rect 2412 10548 2464 10557
rect 1584 10480 1636 10532
rect 2688 10523 2740 10532
rect 2688 10489 2722 10523
rect 2722 10489 2740 10523
rect 2688 10480 2740 10489
rect 3424 10480 3476 10532
rect 3608 10548 3660 10600
rect 4804 10548 4856 10600
rect 5632 10616 5684 10668
rect 7380 10616 7432 10668
rect 10324 10616 10376 10668
rect 12624 10795 12676 10804
rect 12624 10761 12633 10795
rect 12633 10761 12667 10795
rect 12667 10761 12676 10795
rect 12624 10752 12676 10761
rect 11428 10684 11480 10736
rect 13636 10684 13688 10736
rect 13268 10659 13320 10668
rect 13268 10625 13277 10659
rect 13277 10625 13311 10659
rect 13311 10625 13320 10659
rect 13268 10616 13320 10625
rect 13544 10616 13596 10668
rect 15660 10684 15712 10736
rect 16488 10659 16540 10668
rect 16488 10625 16497 10659
rect 16497 10625 16531 10659
rect 16531 10625 16540 10659
rect 16488 10616 16540 10625
rect 17592 10659 17644 10668
rect 17592 10625 17601 10659
rect 17601 10625 17635 10659
rect 17635 10625 17644 10659
rect 17592 10616 17644 10625
rect 6644 10548 6696 10600
rect 8116 10548 8168 10600
rect 9772 10548 9824 10600
rect 10416 10591 10468 10600
rect 10416 10557 10425 10591
rect 10425 10557 10459 10591
rect 10459 10557 10468 10591
rect 10416 10548 10468 10557
rect 12440 10548 12492 10600
rect 13452 10548 13504 10600
rect 13636 10548 13688 10600
rect 2044 10412 2096 10464
rect 2596 10412 2648 10464
rect 4344 10412 4396 10464
rect 4712 10455 4764 10464
rect 4712 10421 4721 10455
rect 4721 10421 4755 10455
rect 4755 10421 4764 10455
rect 4712 10412 4764 10421
rect 4896 10412 4948 10464
rect 5448 10480 5500 10532
rect 6736 10412 6788 10464
rect 7748 10412 7800 10464
rect 9588 10412 9640 10464
rect 9772 10455 9824 10464
rect 9772 10421 9781 10455
rect 9781 10421 9815 10455
rect 9815 10421 9824 10455
rect 9772 10412 9824 10421
rect 10508 10412 10560 10464
rect 11336 10480 11388 10532
rect 18512 10548 18564 10600
rect 14924 10480 14976 10532
rect 15476 10412 15528 10464
rect 16396 10455 16448 10464
rect 16396 10421 16405 10455
rect 16405 10421 16439 10455
rect 16439 10421 16448 10455
rect 16396 10412 16448 10421
rect 6912 10310 6964 10362
rect 6976 10310 7028 10362
rect 7040 10310 7092 10362
rect 7104 10310 7156 10362
rect 12843 10310 12895 10362
rect 12907 10310 12959 10362
rect 12971 10310 13023 10362
rect 13035 10310 13087 10362
rect 2136 10208 2188 10260
rect 3608 10208 3660 10260
rect 4620 10208 4672 10260
rect 4896 10208 4948 10260
rect 9680 10251 9732 10260
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 3056 10072 3108 10124
rect 3516 10072 3568 10124
rect 2596 10047 2648 10056
rect 2596 10013 2605 10047
rect 2605 10013 2639 10047
rect 2639 10013 2648 10047
rect 2596 10004 2648 10013
rect 3424 10004 3476 10056
rect 4068 10072 4120 10124
rect 4436 10115 4488 10124
rect 4436 10081 4445 10115
rect 4445 10081 4479 10115
rect 4479 10081 4488 10115
rect 4436 10072 4488 10081
rect 4528 10047 4580 10056
rect 4528 10013 4537 10047
rect 4537 10013 4571 10047
rect 4571 10013 4580 10047
rect 4528 10004 4580 10013
rect 5816 10140 5868 10192
rect 6184 10140 6236 10192
rect 7656 10140 7708 10192
rect 6000 10072 6052 10124
rect 5632 10004 5684 10056
rect 6644 10072 6696 10124
rect 9680 10217 9689 10251
rect 9689 10217 9723 10251
rect 9723 10217 9732 10251
rect 9680 10208 9732 10217
rect 10048 10251 10100 10260
rect 10048 10217 10057 10251
rect 10057 10217 10091 10251
rect 10091 10217 10100 10251
rect 10048 10208 10100 10217
rect 12440 10208 12492 10260
rect 14924 10251 14976 10260
rect 12624 10140 12676 10192
rect 13452 10140 13504 10192
rect 14924 10217 14933 10251
rect 14933 10217 14967 10251
rect 14967 10217 14976 10251
rect 14924 10208 14976 10217
rect 16396 10208 16448 10260
rect 17500 10251 17552 10260
rect 17500 10217 17509 10251
rect 17509 10217 17543 10251
rect 17543 10217 17552 10251
rect 17500 10208 17552 10217
rect 10600 10072 10652 10124
rect 11060 10115 11112 10124
rect 11060 10081 11069 10115
rect 11069 10081 11103 10115
rect 11103 10081 11112 10115
rect 11060 10072 11112 10081
rect 12716 10115 12768 10124
rect 12716 10081 12725 10115
rect 12725 10081 12759 10115
rect 12759 10081 12768 10115
rect 12716 10072 12768 10081
rect 13636 10072 13688 10124
rect 15200 10072 15252 10124
rect 16120 10072 16172 10124
rect 17592 10140 17644 10192
rect 17224 10072 17276 10124
rect 7472 10004 7524 10056
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 11152 10047 11204 10056
rect 11152 10013 11161 10047
rect 11161 10013 11195 10047
rect 11195 10013 11204 10047
rect 11152 10004 11204 10013
rect 11336 10047 11388 10056
rect 11336 10013 11345 10047
rect 11345 10013 11379 10047
rect 11379 10013 11388 10047
rect 12808 10047 12860 10056
rect 11336 10004 11388 10013
rect 12808 10013 12817 10047
rect 12817 10013 12851 10047
rect 12851 10013 12860 10047
rect 12808 10004 12860 10013
rect 18052 10115 18104 10124
rect 18052 10081 18061 10115
rect 18061 10081 18095 10115
rect 18095 10081 18104 10115
rect 18052 10072 18104 10081
rect 4712 9936 4764 9988
rect 1400 9868 1452 9920
rect 4252 9868 4304 9920
rect 5540 9868 5592 9920
rect 7196 9868 7248 9920
rect 8852 9868 8904 9920
rect 9772 9936 9824 9988
rect 11888 9936 11940 9988
rect 12256 9936 12308 9988
rect 12348 9936 12400 9988
rect 10600 9868 10652 9920
rect 15200 9868 15252 9920
rect 16488 9868 16540 9920
rect 18420 9868 18472 9920
rect 3947 9766 3999 9818
rect 4011 9766 4063 9818
rect 4075 9766 4127 9818
rect 4139 9766 4191 9818
rect 9878 9766 9930 9818
rect 9942 9766 9994 9818
rect 10006 9766 10058 9818
rect 10070 9766 10122 9818
rect 15808 9766 15860 9818
rect 15872 9766 15924 9818
rect 15936 9766 15988 9818
rect 16000 9766 16052 9818
rect 2688 9664 2740 9716
rect 3424 9664 3476 9716
rect 5908 9596 5960 9648
rect 7840 9639 7892 9648
rect 3792 9528 3844 9580
rect 4068 9528 4120 9580
rect 6184 9528 6236 9580
rect 1768 9460 1820 9512
rect 1952 9503 2004 9512
rect 1952 9469 1961 9503
rect 1961 9469 1995 9503
rect 1995 9469 2004 9503
rect 1952 9460 2004 9469
rect 7840 9605 7849 9639
rect 7849 9605 7883 9639
rect 7883 9605 7892 9639
rect 7840 9596 7892 9605
rect 8484 9664 8536 9716
rect 9036 9664 9088 9716
rect 10508 9664 10560 9716
rect 8300 9596 8352 9648
rect 8576 9596 8628 9648
rect 9496 9596 9548 9648
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 9404 9571 9456 9580
rect 7196 9503 7248 9512
rect 7196 9469 7205 9503
rect 7205 9469 7239 9503
rect 7239 9469 7248 9503
rect 7196 9460 7248 9469
rect 7472 9460 7524 9512
rect 9404 9537 9413 9571
rect 9413 9537 9447 9571
rect 9447 9537 9456 9571
rect 9404 9528 9456 9537
rect 10784 9528 10836 9580
rect 10600 9460 10652 9512
rect 10876 9460 10928 9512
rect 11336 9664 11388 9716
rect 12348 9664 12400 9716
rect 12440 9664 12492 9716
rect 12808 9664 12860 9716
rect 15384 9664 15436 9716
rect 17500 9664 17552 9716
rect 11612 9571 11664 9580
rect 11612 9537 11621 9571
rect 11621 9537 11655 9571
rect 11655 9537 11664 9571
rect 11612 9528 11664 9537
rect 13544 9571 13596 9580
rect 13544 9537 13553 9571
rect 13553 9537 13587 9571
rect 13587 9537 13596 9571
rect 14924 9571 14976 9580
rect 13544 9528 13596 9537
rect 14924 9537 14933 9571
rect 14933 9537 14967 9571
rect 14967 9537 14976 9571
rect 14924 9528 14976 9537
rect 15200 9528 15252 9580
rect 16120 9528 16172 9580
rect 17224 9528 17276 9580
rect 17960 9528 18012 9580
rect 15476 9460 15528 9512
rect 16580 9460 16632 9512
rect 2228 9435 2280 9444
rect 2228 9401 2262 9435
rect 2262 9401 2280 9435
rect 2228 9392 2280 9401
rect 2412 9392 2464 9444
rect 3332 9392 3384 9444
rect 4160 9392 4212 9444
rect 4436 9392 4488 9444
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 3424 9324 3476 9376
rect 4252 9367 4304 9376
rect 4252 9333 4261 9367
rect 4261 9333 4295 9367
rect 4295 9333 4304 9367
rect 4252 9324 4304 9333
rect 4344 9367 4396 9376
rect 4344 9333 4353 9367
rect 4353 9333 4387 9367
rect 4387 9333 4396 9367
rect 4344 9324 4396 9333
rect 4528 9324 4580 9376
rect 5080 9324 5132 9376
rect 6092 9367 6144 9376
rect 6092 9333 6101 9367
rect 6101 9333 6135 9367
rect 6135 9333 6144 9367
rect 6092 9324 6144 9333
rect 6184 9367 6236 9376
rect 6184 9333 6193 9367
rect 6193 9333 6227 9367
rect 6227 9333 6236 9367
rect 6184 9324 6236 9333
rect 6460 9324 6512 9376
rect 12164 9392 12216 9444
rect 12808 9392 12860 9444
rect 7564 9324 7616 9376
rect 8208 9324 8260 9376
rect 8392 9324 8444 9376
rect 8668 9324 8720 9376
rect 9036 9324 9088 9376
rect 9128 9324 9180 9376
rect 11980 9324 12032 9376
rect 12348 9324 12400 9376
rect 14096 9324 14148 9376
rect 14464 9324 14516 9376
rect 15660 9367 15712 9376
rect 15660 9333 15669 9367
rect 15669 9333 15703 9367
rect 15703 9333 15712 9367
rect 15660 9324 15712 9333
rect 16672 9367 16724 9376
rect 16672 9333 16681 9367
rect 16681 9333 16715 9367
rect 16715 9333 16724 9367
rect 16672 9324 16724 9333
rect 16764 9367 16816 9376
rect 16764 9333 16773 9367
rect 16773 9333 16807 9367
rect 16807 9333 16816 9367
rect 17592 9367 17644 9376
rect 16764 9324 16816 9333
rect 17592 9333 17601 9367
rect 17601 9333 17635 9367
rect 17635 9333 17644 9367
rect 17592 9324 17644 9333
rect 18328 9324 18380 9376
rect 6912 9222 6964 9274
rect 6976 9222 7028 9274
rect 7040 9222 7092 9274
rect 7104 9222 7156 9274
rect 12843 9222 12895 9274
rect 12907 9222 12959 9274
rect 12971 9222 13023 9274
rect 13035 9222 13087 9274
rect 4344 9120 4396 9172
rect 11888 9120 11940 9172
rect 12256 9120 12308 9172
rect 12716 9120 12768 9172
rect 13176 9120 13228 9172
rect 15292 9120 15344 9172
rect 15660 9120 15712 9172
rect 16396 9120 16448 9172
rect 16672 9120 16724 9172
rect 17132 9163 17184 9172
rect 17132 9129 17141 9163
rect 17141 9129 17175 9163
rect 17175 9129 17184 9163
rect 17132 9120 17184 9129
rect 1952 9052 2004 9104
rect 1860 9027 1912 9036
rect 1860 8993 1894 9027
rect 1894 8993 1912 9027
rect 1860 8984 1912 8993
rect 4068 8984 4120 9036
rect 4896 8984 4948 9036
rect 3056 8916 3108 8968
rect 9036 9052 9088 9104
rect 9128 9052 9180 9104
rect 13084 9052 13136 9104
rect 18604 9052 18656 9104
rect 5264 9027 5316 9036
rect 5264 8993 5273 9027
rect 5273 8993 5307 9027
rect 5307 8993 5316 9027
rect 5264 8984 5316 8993
rect 5540 8984 5592 9036
rect 6644 8984 6696 9036
rect 5356 8959 5408 8968
rect 5356 8925 5365 8959
rect 5365 8925 5399 8959
rect 5399 8925 5408 8959
rect 5356 8916 5408 8925
rect 5448 8959 5500 8968
rect 5448 8925 5457 8959
rect 5457 8925 5491 8959
rect 5491 8925 5500 8959
rect 5448 8916 5500 8925
rect 8944 8916 8996 8968
rect 9036 8959 9088 8968
rect 9036 8925 9045 8959
rect 9045 8925 9079 8959
rect 9079 8925 9088 8959
rect 9404 8984 9456 9036
rect 9588 8984 9640 9036
rect 11060 8984 11112 9036
rect 11704 8984 11756 9036
rect 12164 8984 12216 9036
rect 12992 8984 13044 9036
rect 14740 8984 14792 9036
rect 16948 8984 17000 9036
rect 17960 8984 18012 9036
rect 9036 8916 9088 8925
rect 9496 8916 9548 8968
rect 10416 8916 10468 8968
rect 10876 8916 10928 8968
rect 13544 8959 13596 8968
rect 13544 8925 13553 8959
rect 13553 8925 13587 8959
rect 13587 8925 13596 8959
rect 13544 8916 13596 8925
rect 16580 8916 16632 8968
rect 17224 8959 17276 8968
rect 17224 8925 17233 8959
rect 17233 8925 17267 8959
rect 17267 8925 17276 8959
rect 17224 8916 17276 8925
rect 17316 8959 17368 8968
rect 17316 8925 17325 8959
rect 17325 8925 17359 8959
rect 17359 8925 17368 8959
rect 17316 8916 17368 8925
rect 8392 8848 8444 8900
rect 9588 8848 9640 8900
rect 2228 8780 2280 8832
rect 8300 8780 8352 8832
rect 12992 8848 13044 8900
rect 13268 8848 13320 8900
rect 17040 8848 17092 8900
rect 12348 8823 12400 8832
rect 12348 8789 12357 8823
rect 12357 8789 12391 8823
rect 12391 8789 12400 8823
rect 12348 8780 12400 8789
rect 13636 8780 13688 8832
rect 14096 8780 14148 8832
rect 16856 8780 16908 8832
rect 18052 8823 18104 8832
rect 18052 8789 18061 8823
rect 18061 8789 18095 8823
rect 18095 8789 18104 8823
rect 18052 8780 18104 8789
rect 3947 8678 3999 8730
rect 4011 8678 4063 8730
rect 4075 8678 4127 8730
rect 4139 8678 4191 8730
rect 9878 8678 9930 8730
rect 9942 8678 9994 8730
rect 10006 8678 10058 8730
rect 10070 8678 10122 8730
rect 15808 8678 15860 8730
rect 15872 8678 15924 8730
rect 15936 8678 15988 8730
rect 16000 8678 16052 8730
rect 3332 8576 3384 8628
rect 4896 8576 4948 8628
rect 5356 8576 5408 8628
rect 6000 8576 6052 8628
rect 11704 8619 11756 8628
rect 3056 8508 3108 8560
rect 3608 8508 3660 8560
rect 6736 8508 6788 8560
rect 3332 8440 3384 8492
rect 6000 8483 6052 8492
rect 6000 8449 6009 8483
rect 6009 8449 6043 8483
rect 6043 8449 6052 8483
rect 6000 8440 6052 8449
rect 6092 8372 6144 8424
rect 10324 8508 10376 8560
rect 8392 8440 8444 8492
rect 9496 8440 9548 8492
rect 8484 8415 8536 8424
rect 8484 8381 8493 8415
rect 8493 8381 8527 8415
rect 8527 8381 8536 8415
rect 8484 8372 8536 8381
rect 9680 8372 9732 8424
rect 10876 8372 10928 8424
rect 11704 8585 11713 8619
rect 11713 8585 11747 8619
rect 11747 8585 11756 8619
rect 11704 8576 11756 8585
rect 12992 8576 13044 8628
rect 14096 8576 14148 8628
rect 12440 8508 12492 8560
rect 14280 8508 14332 8560
rect 13452 8483 13504 8492
rect 13452 8449 13461 8483
rect 13461 8449 13495 8483
rect 13495 8449 13504 8483
rect 13452 8440 13504 8449
rect 3884 8347 3936 8356
rect 3884 8313 3918 8347
rect 3918 8313 3936 8347
rect 3884 8304 3936 8313
rect 5448 8304 5500 8356
rect 6184 8304 6236 8356
rect 7748 8304 7800 8356
rect 8208 8304 8260 8356
rect 8576 8304 8628 8356
rect 10416 8304 10468 8356
rect 10508 8304 10560 8356
rect 940 8236 992 8288
rect 2504 8236 2556 8288
rect 2964 8279 3016 8288
rect 2964 8245 2973 8279
rect 2973 8245 3007 8279
rect 3007 8245 3016 8279
rect 2964 8236 3016 8245
rect 3056 8279 3108 8288
rect 3056 8245 3065 8279
rect 3065 8245 3099 8279
rect 3099 8245 3108 8279
rect 3056 8236 3108 8245
rect 6460 8236 6512 8288
rect 7472 8279 7524 8288
rect 7472 8245 7481 8279
rect 7481 8245 7515 8279
rect 7515 8245 7524 8279
rect 7472 8236 7524 8245
rect 8944 8236 8996 8288
rect 12256 8236 12308 8288
rect 12624 8236 12676 8288
rect 13728 8372 13780 8424
rect 16120 8576 16172 8628
rect 16580 8576 16632 8628
rect 16764 8619 16816 8628
rect 16764 8585 16773 8619
rect 16773 8585 16807 8619
rect 16807 8585 16816 8619
rect 16764 8576 16816 8585
rect 17132 8508 17184 8560
rect 16672 8440 16724 8492
rect 17316 8483 17368 8492
rect 17316 8449 17325 8483
rect 17325 8449 17359 8483
rect 17359 8449 17368 8483
rect 17316 8440 17368 8449
rect 13544 8304 13596 8356
rect 16120 8415 16172 8424
rect 16120 8381 16164 8415
rect 16164 8381 16172 8415
rect 17132 8415 17184 8424
rect 16120 8372 16172 8381
rect 17132 8381 17141 8415
rect 17141 8381 17175 8415
rect 17175 8381 17184 8415
rect 17132 8372 17184 8381
rect 17960 8372 18012 8424
rect 14924 8304 14976 8356
rect 15568 8304 15620 8356
rect 17132 8236 17184 8288
rect 18236 8279 18288 8288
rect 18236 8245 18245 8279
rect 18245 8245 18279 8279
rect 18279 8245 18288 8279
rect 18236 8236 18288 8245
rect 6912 8134 6964 8186
rect 6976 8134 7028 8186
rect 7040 8134 7092 8186
rect 7104 8134 7156 8186
rect 12843 8134 12895 8186
rect 12907 8134 12959 8186
rect 12971 8134 13023 8186
rect 13035 8134 13087 8186
rect 3424 8032 3476 8084
rect 5264 8032 5316 8084
rect 5448 8032 5500 8084
rect 7472 8032 7524 8084
rect 8300 8032 8352 8084
rect 2136 7964 2188 8016
rect 3516 7964 3568 8016
rect 1952 7939 2004 7948
rect 1952 7905 1961 7939
rect 1961 7905 1995 7939
rect 1995 7905 2004 7939
rect 1952 7896 2004 7905
rect 2688 7896 2740 7948
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 3332 7828 3384 7880
rect 3884 7828 3936 7880
rect 1492 7692 1544 7744
rect 2596 7735 2648 7744
rect 2596 7701 2605 7735
rect 2605 7701 2639 7735
rect 2639 7701 2648 7735
rect 2596 7692 2648 7701
rect 4344 7692 4396 7744
rect 6000 7964 6052 8016
rect 5540 7939 5592 7948
rect 5540 7905 5549 7939
rect 5549 7905 5583 7939
rect 5583 7905 5592 7939
rect 5540 7896 5592 7905
rect 5632 7896 5684 7948
rect 5172 7871 5224 7880
rect 5172 7837 5181 7871
rect 5181 7837 5215 7871
rect 5215 7837 5224 7871
rect 5172 7828 5224 7837
rect 9772 7964 9824 8016
rect 8944 7939 8996 7948
rect 8944 7905 8953 7939
rect 8953 7905 8987 7939
rect 8987 7905 8996 7939
rect 8944 7896 8996 7905
rect 10324 7896 10376 7948
rect 12624 8032 12676 8084
rect 13268 8075 13320 8084
rect 13268 8041 13277 8075
rect 13277 8041 13311 8075
rect 13311 8041 13320 8075
rect 13268 8032 13320 8041
rect 16672 8075 16724 8084
rect 16672 8041 16681 8075
rect 16681 8041 16715 8075
rect 16715 8041 16724 8075
rect 16672 8032 16724 8041
rect 16948 8075 17000 8084
rect 16948 8041 16957 8075
rect 16957 8041 16991 8075
rect 16991 8041 17000 8075
rect 16948 8032 17000 8041
rect 17776 8032 17828 8084
rect 14280 7939 14332 7948
rect 14280 7905 14289 7939
rect 14289 7905 14323 7939
rect 14323 7905 14332 7939
rect 14280 7896 14332 7905
rect 9036 7871 9088 7880
rect 9036 7837 9045 7871
rect 9045 7837 9079 7871
rect 9079 7837 9088 7871
rect 9036 7828 9088 7837
rect 9404 7828 9456 7880
rect 9680 7871 9732 7880
rect 9680 7837 9689 7871
rect 9689 7837 9723 7871
rect 9723 7837 9732 7871
rect 9680 7828 9732 7837
rect 5816 7692 5868 7744
rect 7656 7735 7708 7744
rect 7656 7701 7665 7735
rect 7665 7701 7699 7735
rect 7699 7701 7708 7735
rect 7656 7692 7708 7701
rect 8300 7760 8352 7812
rect 11980 7760 12032 7812
rect 12164 7760 12216 7812
rect 12348 7828 12400 7880
rect 13176 7828 13228 7880
rect 13452 7871 13504 7880
rect 13452 7837 13461 7871
rect 13461 7837 13495 7871
rect 13495 7837 13504 7871
rect 13452 7828 13504 7837
rect 13912 7828 13964 7880
rect 14648 7896 14700 7948
rect 15200 7896 15252 7948
rect 17224 7896 17276 7948
rect 17408 7939 17460 7948
rect 17408 7905 17417 7939
rect 17417 7905 17451 7939
rect 17451 7905 17460 7939
rect 17408 7896 17460 7905
rect 13268 7760 13320 7812
rect 14924 7828 14976 7880
rect 17592 7964 17644 8016
rect 17868 7964 17920 8016
rect 10876 7692 10928 7744
rect 11796 7692 11848 7744
rect 13084 7692 13136 7744
rect 14280 7692 14332 7744
rect 16488 7692 16540 7744
rect 17132 7692 17184 7744
rect 17408 7692 17460 7744
rect 18696 7692 18748 7744
rect 3947 7590 3999 7642
rect 4011 7590 4063 7642
rect 4075 7590 4127 7642
rect 4139 7590 4191 7642
rect 9878 7590 9930 7642
rect 9942 7590 9994 7642
rect 10006 7590 10058 7642
rect 10070 7590 10122 7642
rect 15808 7590 15860 7642
rect 15872 7590 15924 7642
rect 15936 7590 15988 7642
rect 16000 7590 16052 7642
rect 1768 7531 1820 7540
rect 1768 7497 1777 7531
rect 1777 7497 1811 7531
rect 1811 7497 1820 7531
rect 1768 7488 1820 7497
rect 1952 7488 2004 7540
rect 4252 7488 4304 7540
rect 1860 7352 1912 7404
rect 2964 7352 3016 7404
rect 5448 7420 5500 7472
rect 5172 7395 5224 7404
rect 5172 7361 5181 7395
rect 5181 7361 5215 7395
rect 5215 7361 5224 7395
rect 5172 7352 5224 7361
rect 6184 7395 6236 7404
rect 6184 7361 6193 7395
rect 6193 7361 6227 7395
rect 6227 7361 6236 7395
rect 6184 7352 6236 7361
rect 7748 7395 7800 7404
rect 7748 7361 7757 7395
rect 7757 7361 7791 7395
rect 7791 7361 7800 7395
rect 7748 7352 7800 7361
rect 9772 7488 9824 7540
rect 13912 7488 13964 7540
rect 14096 7488 14148 7540
rect 15476 7488 15528 7540
rect 16120 7488 16172 7540
rect 16304 7488 16356 7540
rect 3056 7284 3108 7336
rect 4804 7284 4856 7336
rect 8300 7327 8352 7336
rect 2504 7259 2556 7268
rect 2504 7225 2513 7259
rect 2513 7225 2547 7259
rect 2547 7225 2556 7259
rect 2504 7216 2556 7225
rect 2596 7259 2648 7268
rect 2596 7225 2605 7259
rect 2605 7225 2639 7259
rect 2639 7225 2648 7259
rect 2596 7216 2648 7225
rect 3792 7216 3844 7268
rect 4988 7191 5040 7200
rect 4988 7157 4997 7191
rect 4997 7157 5031 7191
rect 5031 7157 5040 7191
rect 4988 7148 5040 7157
rect 5632 7191 5684 7200
rect 5632 7157 5641 7191
rect 5641 7157 5675 7191
rect 5675 7157 5684 7191
rect 5632 7148 5684 7157
rect 6000 7191 6052 7200
rect 6000 7157 6009 7191
rect 6009 7157 6043 7191
rect 6043 7157 6052 7191
rect 6000 7148 6052 7157
rect 6092 7191 6144 7200
rect 6092 7157 6101 7191
rect 6101 7157 6135 7191
rect 6135 7157 6144 7191
rect 7288 7191 7340 7200
rect 6092 7148 6144 7157
rect 7288 7157 7297 7191
rect 7297 7157 7331 7191
rect 7331 7157 7340 7191
rect 7288 7148 7340 7157
rect 8024 7216 8076 7268
rect 8300 7293 8309 7327
rect 8309 7293 8343 7327
rect 8343 7293 8352 7327
rect 8300 7284 8352 7293
rect 8392 7284 8444 7336
rect 8576 7327 8628 7336
rect 8576 7293 8599 7327
rect 8599 7293 8628 7327
rect 10508 7420 10560 7472
rect 10876 7420 10928 7472
rect 11060 7352 11112 7404
rect 11796 7395 11848 7404
rect 11796 7361 11805 7395
rect 11805 7361 11839 7395
rect 11839 7361 11848 7395
rect 11796 7352 11848 7361
rect 11888 7395 11940 7404
rect 11888 7361 11897 7395
rect 11897 7361 11931 7395
rect 11931 7361 11940 7395
rect 13084 7420 13136 7472
rect 14740 7420 14792 7472
rect 15016 7420 15068 7472
rect 11888 7352 11940 7361
rect 13176 7352 13228 7404
rect 13544 7352 13596 7404
rect 14924 7352 14976 7404
rect 16488 7352 16540 7404
rect 17500 7352 17552 7404
rect 8576 7284 8628 7293
rect 11244 7216 11296 7268
rect 9680 7148 9732 7200
rect 13268 7284 13320 7336
rect 15016 7284 15068 7336
rect 16396 7284 16448 7336
rect 17224 7284 17276 7336
rect 12624 7216 12676 7268
rect 16672 7216 16724 7268
rect 15016 7148 15068 7200
rect 15200 7148 15252 7200
rect 15476 7191 15528 7200
rect 15476 7157 15485 7191
rect 15485 7157 15519 7191
rect 15519 7157 15528 7191
rect 15476 7148 15528 7157
rect 15660 7148 15712 7200
rect 16120 7148 16172 7200
rect 16488 7191 16540 7200
rect 16488 7157 16497 7191
rect 16497 7157 16531 7191
rect 16531 7157 16540 7191
rect 16488 7148 16540 7157
rect 16764 7148 16816 7200
rect 17684 7148 17736 7200
rect 6912 7046 6964 7098
rect 6976 7046 7028 7098
rect 7040 7046 7092 7098
rect 7104 7046 7156 7098
rect 12843 7046 12895 7098
rect 12907 7046 12959 7098
rect 12971 7046 13023 7098
rect 13035 7046 13087 7098
rect 3516 6987 3568 6996
rect 3516 6953 3525 6987
rect 3525 6953 3559 6987
rect 3559 6953 3568 6987
rect 3516 6944 3568 6953
rect 5172 6944 5224 6996
rect 6000 6944 6052 6996
rect 2228 6851 2280 6860
rect 2228 6817 2237 6851
rect 2237 6817 2271 6851
rect 2271 6817 2280 6851
rect 2228 6808 2280 6817
rect 3792 6808 3844 6860
rect 4988 6876 5040 6928
rect 7748 6944 7800 6996
rect 8760 6944 8812 6996
rect 11888 6944 11940 6996
rect 12624 6944 12676 6996
rect 13268 6944 13320 6996
rect 13636 6944 13688 6996
rect 14280 6876 14332 6928
rect 16488 6944 16540 6996
rect 16580 6944 16632 6996
rect 17316 6987 17368 6996
rect 17316 6953 17325 6987
rect 17325 6953 17359 6987
rect 17359 6953 17368 6987
rect 17316 6944 17368 6953
rect 17408 6876 17460 6928
rect 3056 6740 3108 6792
rect 4068 6783 4120 6792
rect 2964 6715 3016 6724
rect 2964 6681 2973 6715
rect 2973 6681 3007 6715
rect 3007 6681 3016 6715
rect 2964 6672 3016 6681
rect 1860 6647 1912 6656
rect 1860 6613 1869 6647
rect 1869 6613 1903 6647
rect 1903 6613 1912 6647
rect 1860 6604 1912 6613
rect 2412 6647 2464 6656
rect 2412 6613 2421 6647
rect 2421 6613 2455 6647
rect 2455 6613 2464 6647
rect 2412 6604 2464 6613
rect 2504 6604 2556 6656
rect 4068 6749 4077 6783
rect 4077 6749 4111 6783
rect 4111 6749 4120 6783
rect 4068 6740 4120 6749
rect 6000 6740 6052 6792
rect 10324 6808 10376 6860
rect 8116 6740 8168 6792
rect 8484 6783 8536 6792
rect 8484 6749 8493 6783
rect 8493 6749 8527 6783
rect 8527 6749 8536 6783
rect 8484 6740 8536 6749
rect 8576 6783 8628 6792
rect 8576 6749 8585 6783
rect 8585 6749 8619 6783
rect 8619 6749 8628 6783
rect 8576 6740 8628 6749
rect 8760 6740 8812 6792
rect 9128 6740 9180 6792
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 10232 6740 10284 6749
rect 12440 6740 12492 6792
rect 13176 6808 13228 6860
rect 13452 6851 13504 6860
rect 13452 6817 13461 6851
rect 13461 6817 13495 6851
rect 13495 6817 13504 6851
rect 13452 6808 13504 6817
rect 14096 6808 14148 6860
rect 8392 6672 8444 6724
rect 8944 6672 8996 6724
rect 13176 6672 13228 6724
rect 15384 6808 15436 6860
rect 16764 6808 16816 6860
rect 17960 6851 18012 6860
rect 17960 6817 17969 6851
rect 17969 6817 18003 6851
rect 18003 6817 18012 6851
rect 17960 6808 18012 6817
rect 11796 6604 11848 6656
rect 12164 6604 12216 6656
rect 14924 6740 14976 6792
rect 15016 6740 15068 6792
rect 16488 6740 16540 6792
rect 17500 6783 17552 6792
rect 17500 6749 17509 6783
rect 17509 6749 17543 6783
rect 17543 6749 17552 6783
rect 17500 6740 17552 6749
rect 18144 6647 18196 6656
rect 18144 6613 18153 6647
rect 18153 6613 18187 6647
rect 18187 6613 18196 6647
rect 18144 6604 18196 6613
rect 3947 6502 3999 6554
rect 4011 6502 4063 6554
rect 4075 6502 4127 6554
rect 4139 6502 4191 6554
rect 9878 6502 9930 6554
rect 9942 6502 9994 6554
rect 10006 6502 10058 6554
rect 10070 6502 10122 6554
rect 15808 6502 15860 6554
rect 15872 6502 15924 6554
rect 15936 6502 15988 6554
rect 16000 6502 16052 6554
rect 3056 6400 3108 6452
rect 4620 6400 4672 6452
rect 4160 6332 4212 6384
rect 4344 6332 4396 6384
rect 4528 6332 4580 6384
rect 6092 6400 6144 6452
rect 7196 6400 7248 6452
rect 7380 6400 7432 6452
rect 8024 6443 8076 6452
rect 8024 6409 8033 6443
rect 8033 6409 8067 6443
rect 8067 6409 8076 6443
rect 8024 6400 8076 6409
rect 8116 6400 8168 6452
rect 11152 6400 11204 6452
rect 11244 6400 11296 6452
rect 8392 6332 8444 6384
rect 1676 6239 1728 6248
rect 1676 6205 1685 6239
rect 1685 6205 1719 6239
rect 1719 6205 1728 6239
rect 1676 6196 1728 6205
rect 2504 6196 2556 6248
rect 2228 6128 2280 6180
rect 4160 6196 4212 6248
rect 4252 6196 4304 6248
rect 6000 6264 6052 6316
rect 8576 6307 8628 6316
rect 8576 6273 8585 6307
rect 8585 6273 8619 6307
rect 8619 6273 8628 6307
rect 8576 6264 8628 6273
rect 8760 6196 8812 6248
rect 3056 6128 3108 6180
rect 3332 6128 3384 6180
rect 1400 6060 1452 6112
rect 3148 6060 3200 6112
rect 3792 6103 3844 6112
rect 3792 6069 3801 6103
rect 3801 6069 3835 6103
rect 3835 6069 3844 6103
rect 3792 6060 3844 6069
rect 4620 6128 4672 6180
rect 6000 6128 6052 6180
rect 7196 6171 7248 6180
rect 7196 6137 7205 6171
rect 7205 6137 7239 6171
rect 7239 6137 7248 6171
rect 7196 6128 7248 6137
rect 7380 6128 7432 6180
rect 9128 6332 9180 6384
rect 13452 6332 13504 6384
rect 11796 6307 11848 6316
rect 11796 6273 11805 6307
rect 11805 6273 11839 6307
rect 11839 6273 11848 6307
rect 11796 6264 11848 6273
rect 11888 6307 11940 6316
rect 11888 6273 11897 6307
rect 11897 6273 11931 6307
rect 11931 6273 11940 6307
rect 11888 6264 11940 6273
rect 12348 6264 12400 6316
rect 13176 6307 13228 6316
rect 13176 6273 13185 6307
rect 13185 6273 13219 6307
rect 13219 6273 13228 6307
rect 13176 6264 13228 6273
rect 15016 6400 15068 6452
rect 16120 6443 16172 6452
rect 16120 6409 16129 6443
rect 16129 6409 16163 6443
rect 16163 6409 16172 6443
rect 16120 6400 16172 6409
rect 17960 6400 18012 6452
rect 11520 6196 11572 6248
rect 12164 6196 12216 6248
rect 4344 6060 4396 6112
rect 6184 6060 6236 6112
rect 7472 6060 7524 6112
rect 10968 6128 11020 6180
rect 10600 6060 10652 6112
rect 12348 6128 12400 6180
rect 12716 6128 12768 6180
rect 16396 6332 16448 6384
rect 17868 6332 17920 6384
rect 16764 6307 16816 6316
rect 16764 6273 16773 6307
rect 16773 6273 16807 6307
rect 16807 6273 16816 6307
rect 16764 6264 16816 6273
rect 17500 6264 17552 6316
rect 15936 6196 15988 6248
rect 16488 6196 16540 6248
rect 16672 6196 16724 6248
rect 18512 6196 18564 6248
rect 14280 6128 14332 6180
rect 17224 6128 17276 6180
rect 16488 6103 16540 6112
rect 16488 6069 16497 6103
rect 16497 6069 16531 6103
rect 16531 6069 16540 6103
rect 16488 6060 16540 6069
rect 16580 6103 16632 6112
rect 16580 6069 16589 6103
rect 16589 6069 16623 6103
rect 16623 6069 16632 6103
rect 18236 6103 18288 6112
rect 16580 6060 16632 6069
rect 18236 6069 18245 6103
rect 18245 6069 18279 6103
rect 18279 6069 18288 6103
rect 18236 6060 18288 6069
rect 6912 5958 6964 6010
rect 6976 5958 7028 6010
rect 7040 5958 7092 6010
rect 7104 5958 7156 6010
rect 12843 5958 12895 6010
rect 12907 5958 12959 6010
rect 12971 5958 13023 6010
rect 13035 5958 13087 6010
rect 2872 5788 2924 5840
rect 2136 5720 2188 5772
rect 5632 5788 5684 5840
rect 7288 5856 7340 5908
rect 7656 5856 7708 5908
rect 10232 5856 10284 5908
rect 10968 5856 11020 5908
rect 11060 5856 11112 5908
rect 14280 5899 14332 5908
rect 4528 5720 4580 5772
rect 5080 5720 5132 5772
rect 6368 5720 6420 5772
rect 11244 5788 11296 5840
rect 11888 5788 11940 5840
rect 14280 5865 14289 5899
rect 14289 5865 14323 5899
rect 14323 5865 14332 5899
rect 14280 5856 14332 5865
rect 15660 5899 15712 5908
rect 15660 5865 15669 5899
rect 15669 5865 15703 5899
rect 15703 5865 15712 5899
rect 15660 5856 15712 5865
rect 16488 5856 16540 5908
rect 18604 5856 18656 5908
rect 16028 5831 16080 5840
rect 16028 5797 16037 5831
rect 16037 5797 16071 5831
rect 16071 5797 16080 5831
rect 16028 5788 16080 5797
rect 18052 5788 18104 5840
rect 6736 5763 6788 5772
rect 6736 5729 6745 5763
rect 6745 5729 6779 5763
rect 6779 5729 6788 5763
rect 6736 5720 6788 5729
rect 9220 5720 9272 5772
rect 10232 5720 10284 5772
rect 10416 5763 10468 5772
rect 10416 5729 10425 5763
rect 10425 5729 10459 5763
rect 10459 5729 10468 5763
rect 10416 5720 10468 5729
rect 10600 5720 10652 5772
rect 10876 5720 10928 5772
rect 10968 5720 11020 5772
rect 12256 5720 12308 5772
rect 3148 5652 3200 5704
rect 3424 5695 3476 5704
rect 3424 5661 3433 5695
rect 3433 5661 3467 5695
rect 3467 5661 3476 5695
rect 3424 5652 3476 5661
rect 3056 5584 3108 5636
rect 4344 5652 4396 5704
rect 5448 5652 5500 5704
rect 6000 5652 6052 5704
rect 6460 5652 6512 5704
rect 10508 5652 10560 5704
rect 12716 5652 12768 5704
rect 14556 5652 14608 5704
rect 15660 5652 15712 5704
rect 7472 5584 7524 5636
rect 1584 5559 1636 5568
rect 1584 5525 1593 5559
rect 1593 5525 1627 5559
rect 1627 5525 1636 5559
rect 1584 5516 1636 5525
rect 1860 5516 1912 5568
rect 2780 5516 2832 5568
rect 4528 5516 4580 5568
rect 7564 5516 7616 5568
rect 11060 5516 11112 5568
rect 15936 5584 15988 5636
rect 16672 5720 16724 5772
rect 16948 5720 17000 5772
rect 17868 5763 17920 5772
rect 17868 5729 17877 5763
rect 17877 5729 17911 5763
rect 17911 5729 17920 5763
rect 17868 5720 17920 5729
rect 16764 5652 16816 5704
rect 17224 5695 17276 5704
rect 17224 5661 17233 5695
rect 17233 5661 17267 5695
rect 17267 5661 17276 5695
rect 17224 5652 17276 5661
rect 16488 5584 16540 5636
rect 17776 5516 17828 5568
rect 17868 5516 17920 5568
rect 3947 5414 3999 5466
rect 4011 5414 4063 5466
rect 4075 5414 4127 5466
rect 4139 5414 4191 5466
rect 9878 5414 9930 5466
rect 9942 5414 9994 5466
rect 10006 5414 10058 5466
rect 10070 5414 10122 5466
rect 15808 5414 15860 5466
rect 15872 5414 15924 5466
rect 15936 5414 15988 5466
rect 16000 5414 16052 5466
rect 3424 5312 3476 5364
rect 6460 5355 6512 5364
rect 2872 5244 2924 5296
rect 4252 5244 4304 5296
rect 4620 5176 4672 5228
rect 5080 5219 5132 5228
rect 1860 5151 1912 5160
rect 1860 5117 1869 5151
rect 1869 5117 1903 5151
rect 1903 5117 1912 5151
rect 1860 5108 1912 5117
rect 5080 5185 5089 5219
rect 5089 5185 5123 5219
rect 5123 5185 5132 5219
rect 5080 5176 5132 5185
rect 204 5040 256 5092
rect 3516 5015 3568 5024
rect 3516 4981 3525 5015
rect 3525 4981 3559 5015
rect 3559 4981 3568 5015
rect 3516 4972 3568 4981
rect 4712 5040 4764 5092
rect 5448 5040 5500 5092
rect 4252 4972 4304 5024
rect 5264 4972 5316 5024
rect 6460 5321 6469 5355
rect 6469 5321 6503 5355
rect 6503 5321 6512 5355
rect 6460 5312 6512 5321
rect 9220 5312 9272 5364
rect 9312 5312 9364 5364
rect 10876 5312 10928 5364
rect 12624 5312 12676 5364
rect 7380 5108 7432 5160
rect 8392 5108 8444 5160
rect 9956 5151 10008 5160
rect 9956 5117 9965 5151
rect 9965 5117 9999 5151
rect 9999 5117 10008 5151
rect 9956 5108 10008 5117
rect 11336 5108 11388 5160
rect 15200 5244 15252 5296
rect 16580 5312 16632 5364
rect 12348 5176 12400 5228
rect 14832 5219 14884 5228
rect 14832 5185 14841 5219
rect 14841 5185 14875 5219
rect 14875 5185 14884 5219
rect 14832 5176 14884 5185
rect 15476 5176 15528 5228
rect 16764 5244 16816 5296
rect 17224 5219 17276 5228
rect 17224 5185 17233 5219
rect 17233 5185 17267 5219
rect 17267 5185 17276 5219
rect 17224 5176 17276 5185
rect 17040 5151 17092 5160
rect 17040 5117 17049 5151
rect 17049 5117 17083 5151
rect 17083 5117 17092 5151
rect 17040 5108 17092 5117
rect 18052 5151 18104 5160
rect 18052 5117 18061 5151
rect 18061 5117 18095 5151
rect 18095 5117 18104 5151
rect 18052 5108 18104 5117
rect 7840 5040 7892 5092
rect 8944 5040 8996 5092
rect 10232 5083 10284 5092
rect 9404 4972 9456 5024
rect 10232 5049 10244 5083
rect 10244 5049 10284 5083
rect 10232 5040 10284 5049
rect 12624 5083 12676 5092
rect 12624 5049 12633 5083
rect 12633 5049 12667 5083
rect 12667 5049 12676 5083
rect 12624 5040 12676 5049
rect 13636 5040 13688 5092
rect 10324 4972 10376 5024
rect 13728 4972 13780 5024
rect 13820 4972 13872 5024
rect 15200 5015 15252 5024
rect 15200 4981 15209 5015
rect 15209 4981 15243 5015
rect 15243 4981 15252 5015
rect 15200 4972 15252 4981
rect 15384 4972 15436 5024
rect 16856 4972 16908 5024
rect 17500 4972 17552 5024
rect 18236 5015 18288 5024
rect 18236 4981 18245 5015
rect 18245 4981 18279 5015
rect 18279 4981 18288 5015
rect 18236 4972 18288 4981
rect 6912 4870 6964 4922
rect 6976 4870 7028 4922
rect 7040 4870 7092 4922
rect 7104 4870 7156 4922
rect 12843 4870 12895 4922
rect 12907 4870 12959 4922
rect 12971 4870 13023 4922
rect 13035 4870 13087 4922
rect 2412 4811 2464 4820
rect 2412 4777 2421 4811
rect 2421 4777 2455 4811
rect 2455 4777 2464 4811
rect 2412 4768 2464 4777
rect 3516 4768 3568 4820
rect 5172 4768 5224 4820
rect 7472 4768 7524 4820
rect 15200 4768 15252 4820
rect 16672 4811 16724 4820
rect 16672 4777 16681 4811
rect 16681 4777 16715 4811
rect 16715 4777 16724 4811
rect 16672 4768 16724 4777
rect 17960 4768 18012 4820
rect 9312 4743 9364 4752
rect 9312 4709 9321 4743
rect 9321 4709 9355 4743
rect 9355 4709 9364 4743
rect 9312 4700 9364 4709
rect 10324 4743 10376 4752
rect 10324 4709 10358 4743
rect 10358 4709 10376 4743
rect 10324 4700 10376 4709
rect 11060 4700 11112 4752
rect 14004 4743 14056 4752
rect 14004 4709 14013 4743
rect 14013 4709 14047 4743
rect 14047 4709 14056 4743
rect 14004 4700 14056 4709
rect 15568 4700 15620 4752
rect 3792 4632 3844 4684
rect 5080 4632 5132 4684
rect 7380 4632 7432 4684
rect 8944 4675 8996 4684
rect 8944 4641 8953 4675
rect 8953 4641 8987 4675
rect 8987 4641 8996 4675
rect 8944 4632 8996 4641
rect 3148 4564 3200 4616
rect 5448 4564 5500 4616
rect 9956 4564 10008 4616
rect 11796 4632 11848 4684
rect 8576 4539 8628 4548
rect 1860 4471 1912 4480
rect 1860 4437 1869 4471
rect 1869 4437 1903 4471
rect 1903 4437 1912 4471
rect 1860 4428 1912 4437
rect 8576 4505 8585 4539
rect 8585 4505 8619 4539
rect 8619 4505 8628 4539
rect 8576 4496 8628 4505
rect 9220 4496 9272 4548
rect 7656 4471 7708 4480
rect 7656 4437 7665 4471
rect 7665 4437 7699 4471
rect 7699 4437 7708 4471
rect 7656 4428 7708 4437
rect 10968 4428 11020 4480
rect 11428 4471 11480 4480
rect 11428 4437 11437 4471
rect 11437 4437 11471 4471
rect 11471 4437 11480 4471
rect 11428 4428 11480 4437
rect 11888 4471 11940 4480
rect 11888 4437 11897 4471
rect 11897 4437 11931 4471
rect 11931 4437 11940 4471
rect 11888 4428 11940 4437
rect 15200 4632 15252 4684
rect 17408 4632 17460 4684
rect 13268 4564 13320 4616
rect 14556 4564 14608 4616
rect 16212 4607 16264 4616
rect 16212 4573 16221 4607
rect 16221 4573 16255 4607
rect 16255 4573 16264 4607
rect 16212 4564 16264 4573
rect 17132 4607 17184 4616
rect 17132 4573 17141 4607
rect 17141 4573 17175 4607
rect 17175 4573 17184 4607
rect 17132 4564 17184 4573
rect 17224 4607 17276 4616
rect 17224 4573 17233 4607
rect 17233 4573 17267 4607
rect 17267 4573 17276 4607
rect 17224 4564 17276 4573
rect 16856 4496 16908 4548
rect 12440 4428 12492 4480
rect 12716 4428 12768 4480
rect 16212 4428 16264 4480
rect 17868 4428 17920 4480
rect 3947 4326 3999 4378
rect 4011 4326 4063 4378
rect 4075 4326 4127 4378
rect 4139 4326 4191 4378
rect 9878 4326 9930 4378
rect 9942 4326 9994 4378
rect 10006 4326 10058 4378
rect 10070 4326 10122 4378
rect 15808 4326 15860 4378
rect 15872 4326 15924 4378
rect 15936 4326 15988 4378
rect 16000 4326 16052 4378
rect 4344 4224 4396 4276
rect 5448 4267 5500 4276
rect 5448 4233 5457 4267
rect 5457 4233 5491 4267
rect 5491 4233 5500 4267
rect 5448 4224 5500 4233
rect 5080 4156 5132 4208
rect 8392 4224 8444 4276
rect 8944 4224 8996 4276
rect 9404 4224 9456 4276
rect 17132 4224 17184 4276
rect 5632 4088 5684 4140
rect 6552 4088 6604 4140
rect 9772 4156 9824 4208
rect 9220 4088 9272 4140
rect 9588 4088 9640 4140
rect 2136 3952 2188 4004
rect 8484 4020 8536 4072
rect 9312 4020 9364 4072
rect 10324 4020 10376 4072
rect 15752 4156 15804 4208
rect 16488 4156 16540 4208
rect 15108 4131 15160 4140
rect 11428 4063 11480 4072
rect 11428 4029 11437 4063
rect 11437 4029 11471 4063
rect 11471 4029 11480 4063
rect 11428 4020 11480 4029
rect 11796 4063 11848 4072
rect 11796 4029 11805 4063
rect 11805 4029 11839 4063
rect 11839 4029 11848 4063
rect 11796 4020 11848 4029
rect 2504 3927 2556 3936
rect 2504 3893 2513 3927
rect 2513 3893 2547 3927
rect 2547 3893 2556 3927
rect 2504 3884 2556 3893
rect 4620 3952 4672 4004
rect 8300 3952 8352 4004
rect 11980 3952 12032 4004
rect 15108 4097 15117 4131
rect 15117 4097 15151 4131
rect 15151 4097 15160 4131
rect 15108 4088 15160 4097
rect 15292 4088 15344 4140
rect 13176 4020 13228 4072
rect 13636 4063 13688 4072
rect 13636 4029 13645 4063
rect 13645 4029 13679 4063
rect 13679 4029 13688 4063
rect 13636 4020 13688 4029
rect 17592 4088 17644 4140
rect 17776 4088 17828 4140
rect 18512 4088 18564 4140
rect 14280 3995 14332 4004
rect 14280 3961 14289 3995
rect 14289 3961 14323 3995
rect 14323 3961 14332 3995
rect 14280 3952 14332 3961
rect 7932 3884 7984 3936
rect 8760 3884 8812 3936
rect 10968 3884 11020 3936
rect 13452 3884 13504 3936
rect 14004 3884 14056 3936
rect 15752 3995 15804 4004
rect 15752 3961 15761 3995
rect 15761 3961 15795 3995
rect 15795 3961 15804 3995
rect 17500 4020 17552 4072
rect 15752 3952 15804 3961
rect 16580 3952 16632 4004
rect 19616 3952 19668 4004
rect 17592 3927 17644 3936
rect 17592 3893 17601 3927
rect 17601 3893 17635 3927
rect 17635 3893 17644 3927
rect 17592 3884 17644 3893
rect 18236 3927 18288 3936
rect 18236 3893 18245 3927
rect 18245 3893 18279 3927
rect 18279 3893 18288 3927
rect 18236 3884 18288 3893
rect 6912 3782 6964 3834
rect 6976 3782 7028 3834
rect 7040 3782 7092 3834
rect 7104 3782 7156 3834
rect 12843 3782 12895 3834
rect 12907 3782 12959 3834
rect 12971 3782 13023 3834
rect 13035 3782 13087 3834
rect 3792 3612 3844 3664
rect 8300 3723 8352 3732
rect 8300 3689 8309 3723
rect 8309 3689 8343 3723
rect 8343 3689 8352 3723
rect 8300 3680 8352 3689
rect 5356 3612 5408 3664
rect 7656 3612 7708 3664
rect 2780 3587 2832 3596
rect 2780 3553 2789 3587
rect 2789 3553 2823 3587
rect 2823 3553 2832 3587
rect 2780 3544 2832 3553
rect 4344 3544 4396 3596
rect 2136 3476 2188 3528
rect 3056 3476 3108 3528
rect 7472 3544 7524 3596
rect 8392 3612 8444 3664
rect 9680 3612 9732 3664
rect 9588 3544 9640 3596
rect 11428 3612 11480 3664
rect 15016 3680 15068 3732
rect 13544 3655 13596 3664
rect 13544 3621 13553 3655
rect 13553 3621 13587 3655
rect 13587 3621 13596 3655
rect 13544 3612 13596 3621
rect 13912 3612 13964 3664
rect 15660 3612 15712 3664
rect 16304 3612 16356 3664
rect 16856 3655 16908 3664
rect 16856 3621 16865 3655
rect 16865 3621 16899 3655
rect 16899 3621 16908 3655
rect 16856 3612 16908 3621
rect 17040 3612 17092 3664
rect 8576 3519 8628 3528
rect 8576 3485 8585 3519
rect 8585 3485 8619 3519
rect 8619 3485 8628 3519
rect 8576 3476 8628 3485
rect 10232 3544 10284 3596
rect 11888 3544 11940 3596
rect 14096 3587 14148 3596
rect 14096 3553 14105 3587
rect 14105 3553 14139 3587
rect 14139 3553 14148 3587
rect 14096 3544 14148 3553
rect 15108 3544 15160 3596
rect 10784 3519 10836 3528
rect 1860 3451 1912 3460
rect 1860 3417 1869 3451
rect 1869 3417 1903 3451
rect 1903 3417 1912 3451
rect 1860 3408 1912 3417
rect 1216 3340 1268 3392
rect 2964 3383 3016 3392
rect 2964 3349 2973 3383
rect 2973 3349 3007 3383
rect 3007 3349 3016 3383
rect 2964 3340 3016 3349
rect 5172 3340 5224 3392
rect 10784 3485 10793 3519
rect 10793 3485 10827 3519
rect 10827 3485 10836 3519
rect 10784 3476 10836 3485
rect 12164 3476 12216 3528
rect 10324 3451 10376 3460
rect 10324 3417 10333 3451
rect 10333 3417 10367 3451
rect 10367 3417 10376 3451
rect 10324 3408 10376 3417
rect 9036 3383 9088 3392
rect 9036 3349 9045 3383
rect 9045 3349 9079 3383
rect 9079 3349 9088 3383
rect 9036 3340 9088 3349
rect 9680 3340 9732 3392
rect 15660 3408 15712 3460
rect 12348 3340 12400 3392
rect 16672 3408 16724 3460
rect 16120 3340 16172 3392
rect 18052 3383 18104 3392
rect 18052 3349 18061 3383
rect 18061 3349 18095 3383
rect 18095 3349 18104 3383
rect 18052 3340 18104 3349
rect 3947 3238 3999 3290
rect 4011 3238 4063 3290
rect 4075 3238 4127 3290
rect 4139 3238 4191 3290
rect 9878 3238 9930 3290
rect 9942 3238 9994 3290
rect 10006 3238 10058 3290
rect 10070 3238 10122 3290
rect 15808 3238 15860 3290
rect 15872 3238 15924 3290
rect 15936 3238 15988 3290
rect 16000 3238 16052 3290
rect 2136 3136 2188 3188
rect 5724 3136 5776 3188
rect 2412 3111 2464 3120
rect 2412 3077 2421 3111
rect 2421 3077 2455 3111
rect 2455 3077 2464 3111
rect 2412 3068 2464 3077
rect 4988 3068 5040 3120
rect 8392 3136 8444 3188
rect 9036 3136 9088 3188
rect 11796 3136 11848 3188
rect 7288 3068 7340 3120
rect 2780 2932 2832 2984
rect 4252 2932 4304 2984
rect 2688 2864 2740 2916
rect 1860 2839 1912 2848
rect 1860 2805 1869 2839
rect 1869 2805 1903 2839
rect 1903 2805 1912 2839
rect 1860 2796 1912 2805
rect 2780 2796 2832 2848
rect 6736 2932 6788 2984
rect 7656 2932 7708 2984
rect 10784 3068 10836 3120
rect 8668 3043 8720 3052
rect 8668 3009 8677 3043
rect 8677 3009 8711 3043
rect 8711 3009 8720 3043
rect 8668 3000 8720 3009
rect 9128 3000 9180 3052
rect 9680 3043 9732 3052
rect 9680 3009 9689 3043
rect 9689 3009 9723 3043
rect 9723 3009 9732 3043
rect 9680 3000 9732 3009
rect 12256 3068 12308 3120
rect 12532 3068 12584 3120
rect 12348 3000 12400 3052
rect 12624 3000 12676 3052
rect 14096 3000 14148 3052
rect 14372 3043 14424 3052
rect 14372 3009 14381 3043
rect 14381 3009 14415 3043
rect 14415 3009 14424 3043
rect 14372 3000 14424 3009
rect 14740 3000 14792 3052
rect 16212 3000 16264 3052
rect 17132 3000 17184 3052
rect 10416 2932 10468 2984
rect 8208 2864 8260 2916
rect 7840 2796 7892 2848
rect 9496 2864 9548 2916
rect 10784 2907 10836 2916
rect 10784 2873 10793 2907
rect 10793 2873 10827 2907
rect 10827 2873 10836 2907
rect 10784 2864 10836 2873
rect 9128 2796 9180 2848
rect 17224 2932 17276 2984
rect 11796 2864 11848 2916
rect 12440 2796 12492 2848
rect 13176 2864 13228 2916
rect 15108 2796 15160 2848
rect 15200 2796 15252 2848
rect 15936 2907 15988 2916
rect 15936 2873 15945 2907
rect 15945 2873 15979 2907
rect 15979 2873 15988 2907
rect 15936 2864 15988 2873
rect 16764 2864 16816 2916
rect 17592 2839 17644 2848
rect 17592 2805 17601 2839
rect 17601 2805 17635 2839
rect 17635 2805 17644 2839
rect 17592 2796 17644 2805
rect 17868 2796 17920 2848
rect 6912 2694 6964 2746
rect 6976 2694 7028 2746
rect 7040 2694 7092 2746
rect 7104 2694 7156 2746
rect 12843 2694 12895 2746
rect 12907 2694 12959 2746
rect 12971 2694 13023 2746
rect 13035 2694 13087 2746
rect 6644 2592 6696 2644
rect 15016 2592 15068 2644
rect 1676 2524 1728 2576
rect 5724 2524 5776 2576
rect 1492 2456 1544 2508
rect 664 2388 716 2440
rect 3424 2456 3476 2508
rect 5448 2456 5500 2508
rect 5816 2456 5868 2508
rect 7564 2524 7616 2576
rect 7472 2456 7524 2508
rect 7840 2456 7892 2508
rect 8208 2524 8260 2576
rect 10692 2524 10744 2576
rect 12440 2524 12492 2576
rect 13084 2524 13136 2576
rect 13912 2524 13964 2576
rect 14188 2524 14240 2576
rect 9036 2499 9088 2508
rect 9036 2465 9045 2499
rect 9045 2465 9079 2499
rect 9079 2465 9088 2499
rect 9036 2456 9088 2465
rect 14832 2524 14884 2576
rect 15292 2524 15344 2576
rect 1124 2320 1176 2372
rect 3240 2388 3292 2440
rect 3608 2388 3660 2440
rect 6736 2388 6788 2440
rect 8576 2388 8628 2440
rect 11060 2388 11112 2440
rect 11612 2388 11664 2440
rect 12072 2431 12124 2440
rect 12072 2397 12081 2431
rect 12081 2397 12115 2431
rect 12115 2397 12124 2431
rect 12072 2388 12124 2397
rect 12624 2388 12676 2440
rect 13176 2388 13228 2440
rect 15108 2388 15160 2440
rect 15844 2431 15896 2440
rect 15844 2397 15853 2431
rect 15853 2397 15887 2431
rect 15887 2397 15896 2431
rect 15844 2388 15896 2397
rect 16948 2388 17000 2440
rect 17592 2388 17644 2440
rect 17868 2388 17920 2440
rect 7656 2320 7708 2372
rect 10324 2320 10376 2372
rect 8116 2252 8168 2304
rect 8208 2252 8260 2304
rect 10600 2252 10652 2304
rect 15936 2320 15988 2372
rect 17316 2295 17368 2304
rect 17316 2261 17325 2295
rect 17325 2261 17359 2295
rect 17359 2261 17368 2295
rect 17316 2252 17368 2261
rect 17868 2295 17920 2304
rect 17868 2261 17877 2295
rect 17877 2261 17911 2295
rect 17911 2261 17920 2295
rect 17868 2252 17920 2261
rect 3947 2150 3999 2202
rect 4011 2150 4063 2202
rect 4075 2150 4127 2202
rect 4139 2150 4191 2202
rect 9878 2150 9930 2202
rect 9942 2150 9994 2202
rect 10006 2150 10058 2202
rect 10070 2150 10122 2202
rect 15808 2150 15860 2202
rect 15872 2150 15924 2202
rect 15936 2150 15988 2202
rect 16000 2150 16052 2202
rect 5448 2048 5500 2100
rect 14464 2048 14516 2100
rect 8116 1980 8168 2032
rect 15292 1980 15344 2032
rect 5816 1912 5868 1964
rect 10324 1912 10376 1964
rect 13452 1912 13504 1964
rect 18144 1912 18196 1964
rect 14004 1708 14056 1760
rect 17592 1708 17644 1760
rect 12716 1640 12768 1692
rect 19156 1640 19208 1692
<< metal2 >>
rect 294 16200 350 17000
rect 938 16200 994 17000
rect 1582 16200 1638 17000
rect 2226 16200 2282 17000
rect 2870 16200 2926 17000
rect 3422 16280 3478 16289
rect 3422 16215 3478 16224
rect 308 14074 336 16200
rect 296 14068 348 14074
rect 296 14010 348 14016
rect 952 14006 980 16200
rect 1596 14618 1624 16200
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 2240 14006 2268 16200
rect 2596 14408 2648 14414
rect 2596 14350 2648 14356
rect 2410 14240 2466 14249
rect 2410 14175 2466 14184
rect 940 14000 992 14006
rect 940 13942 992 13948
rect 2228 14000 2280 14006
rect 2228 13942 2280 13948
rect 1582 13832 1638 13841
rect 1582 13767 1638 13776
rect 1596 10538 1624 13767
rect 2228 13388 2280 13394
rect 2228 13330 2280 13336
rect 1860 12232 1912 12238
rect 1860 12174 1912 12180
rect 1872 11694 1900 12174
rect 2240 11898 2268 13330
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2332 12986 2360 13262
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2228 11892 2280 11898
rect 2228 11834 2280 11840
rect 1860 11688 1912 11694
rect 1860 11630 1912 11636
rect 2332 11626 2360 12378
rect 2320 11620 2372 11626
rect 2320 11562 2372 11568
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 1676 11076 1728 11082
rect 1676 11018 1728 11024
rect 1584 10532 1636 10538
rect 1584 10474 1636 10480
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1412 10033 1440 10066
rect 1398 10024 1454 10033
rect 1398 9959 1454 9968
rect 1400 9920 1452 9926
rect 1400 9862 1452 9868
rect 1412 8401 1440 9862
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1398 8392 1454 8401
rect 1398 8327 1454 8336
rect 940 8288 992 8294
rect 940 8230 992 8236
rect 204 5092 256 5098
rect 204 5034 256 5040
rect 216 800 244 5034
rect 664 2440 716 2446
rect 664 2382 716 2388
rect 676 800 704 2382
rect 952 1057 980 8230
rect 1596 7993 1624 9318
rect 1582 7984 1638 7993
rect 1582 7919 1638 7928
rect 1492 7744 1544 7750
rect 1492 7686 1544 7692
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 1412 5545 1440 6054
rect 1398 5536 1454 5545
rect 1398 5471 1454 5480
rect 1216 3392 1268 3398
rect 1216 3334 1268 3340
rect 1124 2372 1176 2378
rect 1124 2314 1176 2320
rect 938 1048 994 1057
rect 938 983 994 992
rect 1136 800 1164 2314
rect 202 0 258 800
rect 662 0 718 800
rect 1122 0 1178 800
rect 1228 649 1256 3334
rect 1504 2514 1532 7686
rect 1688 6254 1716 11018
rect 1780 9518 1808 11494
rect 2044 11212 2096 11218
rect 2044 11154 2096 11160
rect 1860 11008 1912 11014
rect 1860 10950 1912 10956
rect 1872 10674 1900 10950
rect 2056 10810 2084 11154
rect 2332 11150 2360 11562
rect 2424 11370 2452 14175
rect 2608 13870 2636 14350
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 2792 13870 2820 14214
rect 2884 14074 2912 16200
rect 3238 15872 3294 15881
rect 3238 15807 3294 15816
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2516 12442 2544 13262
rect 2596 12844 2648 12850
rect 2596 12786 2648 12792
rect 2504 12436 2556 12442
rect 2504 12378 2556 12384
rect 2608 12374 2636 12786
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 2596 12368 2648 12374
rect 2596 12310 2648 12316
rect 2688 12368 2740 12374
rect 2688 12310 2740 12316
rect 2608 11830 2636 12310
rect 2700 12102 2728 12310
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 2700 11830 2728 12038
rect 2596 11824 2648 11830
rect 2596 11766 2648 11772
rect 2688 11824 2740 11830
rect 2688 11766 2740 11772
rect 2424 11342 2544 11370
rect 2412 11280 2464 11286
rect 2412 11222 2464 11228
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2044 10804 2096 10810
rect 2044 10746 2096 10752
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 2056 10470 2084 10610
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 2148 10266 2176 11086
rect 2424 10606 2452 11222
rect 2516 11150 2544 11342
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 1768 9512 1820 9518
rect 1768 9454 1820 9460
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 1964 9110 1992 9454
rect 2424 9450 2452 10542
rect 2608 10470 2636 11766
rect 2700 11286 2728 11766
rect 2792 11286 2820 12582
rect 3056 11688 3108 11694
rect 3056 11630 3108 11636
rect 2962 11384 3018 11393
rect 2962 11319 3018 11328
rect 2688 11280 2740 11286
rect 2688 11222 2740 11228
rect 2780 11280 2832 11286
rect 2780 11222 2832 11228
rect 2792 11082 2820 11222
rect 2976 11150 3004 11319
rect 3068 11218 3096 11630
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 2976 10690 3004 11086
rect 2792 10662 3004 10690
rect 2688 10532 2740 10538
rect 2688 10474 2740 10480
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2608 10062 2636 10406
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2700 9722 2728 10474
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2686 9616 2742 9625
rect 2686 9551 2742 9560
rect 2228 9444 2280 9450
rect 2228 9386 2280 9392
rect 2412 9444 2464 9450
rect 2412 9386 2464 9392
rect 1952 9104 2004 9110
rect 1952 9046 2004 9052
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 1766 7576 1822 7585
rect 1766 7511 1768 7520
rect 1820 7511 1822 7520
rect 1768 7482 1820 7488
rect 1872 7410 1900 8978
rect 2240 8838 2268 9386
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 2136 8016 2188 8022
rect 2136 7958 2188 7964
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 1964 7546 1992 7890
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1872 5953 1900 6598
rect 1858 5944 1914 5953
rect 1858 5879 1914 5888
rect 2148 5778 2176 7958
rect 2240 7886 2268 8774
rect 2504 8288 2556 8294
rect 2504 8230 2556 8236
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2516 7274 2544 8230
rect 2700 7954 2728 9551
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2596 7744 2648 7750
rect 2596 7686 2648 7692
rect 2608 7274 2636 7686
rect 2504 7268 2556 7274
rect 2504 7210 2556 7216
rect 2596 7268 2648 7274
rect 2596 7210 2648 7216
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 2240 6186 2268 6802
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2424 6361 2452 6598
rect 2410 6352 2466 6361
rect 2410 6287 2466 6296
rect 2516 6254 2544 6598
rect 2504 6248 2556 6254
rect 2504 6190 2556 6196
rect 2228 6180 2280 6186
rect 2228 6122 2280 6128
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 2792 5692 2820 10662
rect 2870 10568 2926 10577
rect 2870 10503 2926 10512
rect 2884 7449 2912 10503
rect 3068 10248 3096 11154
rect 2976 10220 3096 10248
rect 2976 8378 3004 10220
rect 3056 10124 3108 10130
rect 3056 10066 3108 10072
rect 3068 8974 3096 10066
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 3068 8566 3096 8910
rect 3056 8560 3108 8566
rect 3056 8502 3108 8508
rect 3160 8514 3188 12582
rect 3252 9625 3280 15807
rect 3332 14340 3384 14346
rect 3332 14282 3384 14288
rect 3344 13870 3372 14282
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 3330 13424 3386 13433
rect 3330 13359 3386 13368
rect 3344 9704 3372 13359
rect 3436 13258 3464 16215
rect 3514 16200 3570 17000
rect 3606 16688 3662 16697
rect 3606 16623 3662 16632
rect 3528 13734 3556 16200
rect 3620 15298 3648 16623
rect 4158 16200 4214 17000
rect 4802 16200 4858 17000
rect 5446 16200 5502 17000
rect 6090 16200 6146 17000
rect 6734 16200 6790 17000
rect 7378 16200 7434 17000
rect 8022 16200 8078 17000
rect 8666 16200 8722 17000
rect 9310 16200 9366 17000
rect 9954 16200 10010 17000
rect 10322 16280 10378 16289
rect 10322 16215 10378 16224
rect 4066 15464 4122 15473
rect 4066 15399 4122 15408
rect 3608 15292 3660 15298
rect 3608 15234 3660 15240
rect 4080 15230 4108 15399
rect 4068 15224 4120 15230
rect 4068 15166 4120 15172
rect 3790 15056 3846 15065
rect 3790 14991 3846 15000
rect 3516 13728 3568 13734
rect 3516 13670 3568 13676
rect 3424 13252 3476 13258
rect 3424 13194 3476 13200
rect 3436 12714 3464 13194
rect 3608 13184 3660 13190
rect 3608 13126 3660 13132
rect 3514 13016 3570 13025
rect 3514 12951 3570 12960
rect 3528 12918 3556 12951
rect 3516 12912 3568 12918
rect 3516 12854 3568 12860
rect 3620 12782 3648 13126
rect 3608 12776 3660 12782
rect 3608 12718 3660 12724
rect 3424 12708 3476 12714
rect 3424 12650 3476 12656
rect 3700 12640 3752 12646
rect 3700 12582 3752 12588
rect 3608 12300 3660 12306
rect 3608 12242 3660 12248
rect 3620 11234 3648 12242
rect 3712 11354 3740 12582
rect 3804 12306 3832 14991
rect 4172 14362 4200 16200
rect 4344 15292 4396 15298
rect 4344 15234 4396 15240
rect 4172 14334 4292 14362
rect 3921 14172 4217 14192
rect 3977 14170 4001 14172
rect 4057 14170 4081 14172
rect 4137 14170 4161 14172
rect 3999 14118 4001 14170
rect 4063 14118 4075 14170
rect 4137 14118 4139 14170
rect 3977 14116 4001 14118
rect 4057 14116 4081 14118
rect 4137 14116 4161 14118
rect 3921 14096 4217 14116
rect 4264 13462 4292 14334
rect 4252 13456 4304 13462
rect 4252 13398 4304 13404
rect 3921 13084 4217 13104
rect 3977 13082 4001 13084
rect 4057 13082 4081 13084
rect 4137 13082 4161 13084
rect 3999 13030 4001 13082
rect 4063 13030 4075 13082
rect 4137 13030 4139 13082
rect 3977 13028 4001 13030
rect 4057 13028 4081 13030
rect 4137 13028 4161 13030
rect 3921 13008 4217 13028
rect 4068 12640 4120 12646
rect 4066 12608 4068 12617
rect 4120 12608 4122 12617
rect 4066 12543 4122 12552
rect 3792 12300 3844 12306
rect 3792 12242 3844 12248
rect 3790 12200 3846 12209
rect 3790 12135 3846 12144
rect 3804 12102 3832 12135
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3921 11996 4217 12016
rect 3977 11994 4001 11996
rect 4057 11994 4081 11996
rect 4137 11994 4161 11996
rect 3999 11942 4001 11994
rect 4063 11942 4075 11994
rect 4137 11942 4139 11994
rect 3977 11940 4001 11942
rect 4057 11940 4081 11942
rect 4137 11940 4161 11942
rect 3921 11920 4217 11940
rect 3792 11892 3844 11898
rect 3792 11834 3844 11840
rect 3804 11801 3832 11834
rect 3790 11792 3846 11801
rect 3790 11727 3846 11736
rect 3700 11348 3752 11354
rect 3700 11290 3752 11296
rect 3620 11206 3740 11234
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3436 10538 3464 11086
rect 3606 10976 3662 10985
rect 3606 10911 3662 10920
rect 3620 10606 3648 10911
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 3424 10532 3476 10538
rect 3424 10474 3476 10480
rect 3436 10062 3464 10474
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3528 9761 3556 10066
rect 3514 9752 3570 9761
rect 3424 9716 3476 9722
rect 3344 9676 3424 9704
rect 3514 9687 3570 9696
rect 3424 9658 3476 9664
rect 3238 9616 3294 9625
rect 3238 9551 3294 9560
rect 3332 9444 3384 9450
rect 3332 9386 3384 9392
rect 3344 8634 3372 9386
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3160 8486 3280 8514
rect 2976 8350 3188 8378
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 2870 7440 2926 7449
rect 2976 7410 3004 8230
rect 2870 7375 2926 7384
rect 2964 7404 3016 7410
rect 2884 5846 2912 7375
rect 2964 7346 3016 7352
rect 3068 7342 3096 8230
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 3056 6792 3108 6798
rect 2962 6760 3018 6769
rect 3056 6734 3108 6740
rect 2962 6695 2964 6704
rect 3016 6695 3018 6704
rect 2964 6666 3016 6672
rect 3068 6458 3096 6734
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 3160 6338 3188 8350
rect 2976 6310 3188 6338
rect 2872 5840 2924 5846
rect 2872 5782 2924 5788
rect 2792 5664 2912 5692
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 1860 5568 1912 5574
rect 1860 5510 1912 5516
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 1596 5137 1624 5510
rect 1872 5166 1900 5510
rect 1860 5160 1912 5166
rect 1582 5128 1638 5137
rect 1860 5102 1912 5108
rect 1582 5063 1638 5072
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2424 4729 2452 4762
rect 2410 4720 2466 4729
rect 2410 4655 2466 4664
rect 1860 4480 1912 4486
rect 1860 4422 1912 4428
rect 1872 4321 1900 4422
rect 1858 4312 1914 4321
rect 1858 4247 1914 4256
rect 2136 4004 2188 4010
rect 2136 3946 2188 3952
rect 2148 3534 2176 3946
rect 2504 3936 2556 3942
rect 2502 3904 2504 3913
rect 2556 3904 2558 3913
rect 2502 3839 2558 3848
rect 2792 3602 2820 5510
rect 2884 5302 2912 5664
rect 2872 5296 2924 5302
rect 2872 5238 2924 5244
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 2136 3528 2188 3534
rect 1858 3496 1914 3505
rect 2976 3482 3004 6310
rect 3056 6180 3108 6186
rect 3056 6122 3108 6128
rect 3068 5642 3096 6122
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3160 5710 3188 6054
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 3056 5636 3108 5642
rect 3056 5578 3108 5584
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 2136 3470 2188 3476
rect 1858 3431 1860 3440
rect 1912 3431 1914 3440
rect 2792 3454 3004 3482
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 1860 3402 1912 3408
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 1860 2848 1912 2854
rect 1860 2790 1912 2796
rect 1872 2689 1900 2790
rect 1858 2680 1914 2689
rect 1858 2615 1914 2624
rect 1676 2576 1728 2582
rect 1676 2518 1728 2524
rect 1492 2508 1544 2514
rect 1492 2450 1544 2456
rect 1688 800 1716 2518
rect 2148 800 2176 3130
rect 2412 3120 2464 3126
rect 2410 3088 2412 3097
rect 2464 3088 2466 3097
rect 2410 3023 2466 3032
rect 2792 2990 2820 3454
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2780 2984 2832 2990
rect 2780 2926 2832 2932
rect 2688 2916 2740 2922
rect 2688 2858 2740 2864
rect 2700 800 2728 2858
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2792 1465 2820 2790
rect 2976 2281 3004 3334
rect 2962 2272 3018 2281
rect 2962 2207 3018 2216
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 1214 640 1270 649
rect 1214 575 1270 584
rect 1674 0 1730 800
rect 2134 0 2190 800
rect 2686 0 2742 800
rect 3068 241 3096 3470
rect 3160 800 3188 4558
rect 3252 2446 3280 8486
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3344 7886 3372 8434
rect 3436 8090 3464 9318
rect 3514 9072 3570 9081
rect 3514 9007 3570 9016
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3528 8022 3556 9007
rect 3620 8945 3648 10202
rect 3606 8936 3662 8945
rect 3606 8871 3662 8880
rect 3608 8560 3660 8566
rect 3608 8502 3660 8508
rect 3516 8016 3568 8022
rect 3516 7958 3568 7964
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3514 7168 3570 7177
rect 3514 7103 3570 7112
rect 3528 7002 3556 7103
rect 3516 6996 3568 7002
rect 3516 6938 3568 6944
rect 3514 6760 3570 6769
rect 3514 6695 3570 6704
rect 3332 6180 3384 6186
rect 3332 6122 3384 6128
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3344 1873 3372 6122
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 3436 5370 3464 5646
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3528 5250 3556 6695
rect 3436 5222 3556 5250
rect 3436 2514 3464 5222
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3528 4826 3556 4966
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3620 4672 3648 8502
rect 3712 7857 3740 11206
rect 3921 10908 4217 10928
rect 3977 10906 4001 10908
rect 4057 10906 4081 10908
rect 4137 10906 4161 10908
rect 3999 10854 4001 10906
rect 4063 10854 4075 10906
rect 4137 10854 4139 10906
rect 3977 10852 4001 10854
rect 4057 10852 4081 10854
rect 4137 10852 4161 10854
rect 3921 10832 4217 10852
rect 4356 10470 4384 15234
rect 4816 13530 4844 16200
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 5460 13394 5488 16200
rect 6104 13870 6132 16200
rect 6748 14396 6776 16200
rect 7288 15224 7340 15230
rect 7288 15166 7340 15172
rect 6886 14716 7182 14736
rect 6942 14714 6966 14716
rect 7022 14714 7046 14716
rect 7102 14714 7126 14716
rect 6964 14662 6966 14714
rect 7028 14662 7040 14714
rect 7102 14662 7104 14714
rect 6942 14660 6966 14662
rect 7022 14660 7046 14662
rect 7102 14660 7126 14662
rect 6886 14640 7182 14660
rect 6748 14368 6960 14396
rect 6932 14074 6960 14368
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 6276 14000 6328 14006
rect 6276 13942 6328 13948
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 4724 12850 5028 12866
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4712 12844 5028 12850
rect 4764 12838 5028 12844
rect 4712 12786 4764 12792
rect 4632 12374 4660 12786
rect 4896 12776 4948 12782
rect 4896 12718 4948 12724
rect 4620 12368 4672 12374
rect 4620 12310 4672 12316
rect 4632 11898 4660 12310
rect 4908 11914 4936 12718
rect 5000 12050 5028 12838
rect 5000 12022 5120 12050
rect 4908 11898 5028 11914
rect 4620 11892 4672 11898
rect 4908 11892 5040 11898
rect 4908 11886 4988 11892
rect 4620 11834 4672 11840
rect 4988 11834 5040 11840
rect 5092 11354 5120 12022
rect 5276 11880 5304 12922
rect 6184 12368 6236 12374
rect 6184 12310 6236 12316
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5184 11852 5304 11880
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 5000 10810 5028 11154
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4066 10160 4122 10169
rect 4066 10095 4068 10104
rect 4120 10095 4122 10104
rect 4436 10124 4488 10130
rect 4068 10066 4120 10072
rect 4436 10066 4488 10072
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 3921 9820 4217 9840
rect 3977 9818 4001 9820
rect 4057 9818 4081 9820
rect 4137 9818 4161 9820
rect 3999 9766 4001 9818
rect 4063 9766 4075 9818
rect 4137 9766 4139 9818
rect 3977 9764 4001 9766
rect 4057 9764 4081 9766
rect 4137 9764 4161 9766
rect 3921 9744 4217 9764
rect 4264 9704 4292 9862
rect 4448 9761 4476 10066
rect 4528 10056 4580 10062
rect 4528 9998 4580 10004
rect 4172 9676 4292 9704
rect 4434 9752 4490 9761
rect 4434 9687 4490 9696
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 3698 7848 3754 7857
rect 3698 7783 3754 7792
rect 3804 7274 3832 9522
rect 4080 9042 4108 9522
rect 4172 9450 4200 9676
rect 4540 9489 4568 9998
rect 4526 9480 4582 9489
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 4436 9444 4488 9450
rect 4526 9415 4582 9424
rect 4436 9386 4488 9392
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 3921 8732 4217 8752
rect 3977 8730 4001 8732
rect 4057 8730 4081 8732
rect 4137 8730 4161 8732
rect 3999 8678 4001 8730
rect 4063 8678 4075 8730
rect 4137 8678 4139 8730
rect 3977 8676 4001 8678
rect 4057 8676 4081 8678
rect 4137 8676 4161 8678
rect 3921 8656 4217 8676
rect 3884 8356 3936 8362
rect 3884 8298 3936 8304
rect 3896 7886 3924 8298
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 3921 7644 4217 7664
rect 3977 7642 4001 7644
rect 4057 7642 4081 7644
rect 4137 7642 4161 7644
rect 3999 7590 4001 7642
rect 4063 7590 4075 7642
rect 4137 7590 4139 7642
rect 3977 7588 4001 7590
rect 4057 7588 4081 7590
rect 4137 7588 4161 7590
rect 3921 7568 4217 7588
rect 4264 7546 4292 9318
rect 4356 9178 4384 9318
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 3792 7268 3844 7274
rect 3792 7210 3844 7216
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 3804 6118 3832 6802
rect 4068 6792 4120 6798
rect 4120 6752 4292 6780
rect 4068 6734 4120 6740
rect 3921 6556 4217 6576
rect 3977 6554 4001 6556
rect 4057 6554 4081 6556
rect 4137 6554 4161 6556
rect 3999 6502 4001 6554
rect 4063 6502 4075 6554
rect 4137 6502 4139 6554
rect 3977 6500 4001 6502
rect 4057 6500 4081 6502
rect 4137 6500 4161 6502
rect 3921 6480 4217 6500
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 4172 6254 4200 6326
rect 4264 6254 4292 6752
rect 4356 6390 4384 7686
rect 4344 6384 4396 6390
rect 4344 6326 4396 6332
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3921 5468 4217 5488
rect 3977 5466 4001 5468
rect 4057 5466 4081 5468
rect 4137 5466 4161 5468
rect 3999 5414 4001 5466
rect 4063 5414 4075 5466
rect 4137 5414 4139 5466
rect 3977 5412 4001 5414
rect 4057 5412 4081 5414
rect 4137 5412 4161 5414
rect 3921 5392 4217 5412
rect 4264 5302 4292 6190
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4356 5710 4384 6054
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 4252 5296 4304 5302
rect 4304 5244 4384 5250
rect 4252 5238 4384 5244
rect 4264 5222 4384 5238
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 3792 4684 3844 4690
rect 3620 4644 3792 4672
rect 3792 4626 3844 4632
rect 3804 3670 3832 4626
rect 3921 4380 4217 4400
rect 3977 4378 4001 4380
rect 4057 4378 4081 4380
rect 4137 4378 4161 4380
rect 3999 4326 4001 4378
rect 4063 4326 4075 4378
rect 4137 4326 4139 4378
rect 3977 4324 4001 4326
rect 4057 4324 4081 4326
rect 4137 4324 4161 4326
rect 3921 4304 4217 4324
rect 3792 3664 3844 3670
rect 3792 3606 3844 3612
rect 3921 3292 4217 3312
rect 3977 3290 4001 3292
rect 4057 3290 4081 3292
rect 4137 3290 4161 3292
rect 3999 3238 4001 3290
rect 4063 3238 4075 3290
rect 4137 3238 4139 3290
rect 3977 3236 4001 3238
rect 4057 3236 4081 3238
rect 4137 3236 4161 3238
rect 3921 3216 4217 3236
rect 4264 2990 4292 4966
rect 4356 4282 4384 5222
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4356 3602 4384 4218
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4252 2984 4304 2990
rect 4252 2926 4304 2932
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 3330 1864 3386 1873
rect 3330 1799 3386 1808
rect 3620 800 3648 2382
rect 3921 2204 4217 2224
rect 3977 2202 4001 2204
rect 4057 2202 4081 2204
rect 4137 2202 4161 2204
rect 3999 2150 4001 2202
rect 4063 2150 4075 2202
rect 4137 2150 4139 2202
rect 3977 2148 4001 2150
rect 4057 2148 4081 2150
rect 4137 2148 4161 2150
rect 3921 2128 4217 2148
rect 4448 1306 4476 9386
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4540 6769 4568 9318
rect 4526 6760 4582 6769
rect 4526 6695 4582 6704
rect 4632 6458 4660 10202
rect 4724 9994 4752 10406
rect 4712 9988 4764 9994
rect 4712 9930 4764 9936
rect 4710 9480 4766 9489
rect 4710 9415 4766 9424
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4528 6384 4580 6390
rect 4528 6326 4580 6332
rect 4540 5778 4568 6326
rect 4620 6180 4672 6186
rect 4620 6122 4672 6128
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4540 5574 4568 5714
rect 4528 5568 4580 5574
rect 4528 5510 4580 5516
rect 4632 5234 4660 6122
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4724 5098 4752 9415
rect 4816 7342 4844 10542
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4908 10266 4936 10406
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 5080 9376 5132 9382
rect 5184 9364 5212 11852
rect 5460 11778 5488 12174
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5368 11750 5488 11778
rect 5276 11150 5304 11698
rect 5368 11694 5396 11750
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 5540 11620 5592 11626
rect 5540 11562 5592 11568
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5460 10538 5488 11018
rect 5552 10742 5580 11562
rect 5828 11150 5856 11834
rect 6092 11824 6144 11830
rect 6092 11766 6144 11772
rect 6104 11354 6132 11766
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 5644 10674 5672 10950
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 5828 10418 5856 11086
rect 5736 10390 5856 10418
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5262 9752 5318 9761
rect 5262 9687 5318 9696
rect 5132 9336 5212 9364
rect 5080 9318 5132 9324
rect 5276 9160 5304 9687
rect 5184 9132 5304 9160
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 4908 8634 4936 8978
rect 5078 8936 5134 8945
rect 5078 8871 5134 8880
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 5000 6934 5028 7142
rect 4988 6928 5040 6934
rect 4988 6870 5040 6876
rect 4712 5092 4764 5098
rect 4712 5034 4764 5040
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4172 1278 4476 1306
rect 4172 800 4200 1278
rect 4632 800 4660 3946
rect 5000 3126 5028 6870
rect 5092 5896 5120 8871
rect 5184 7970 5212 9132
rect 5552 9042 5580 9862
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5276 8090 5304 8978
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5368 8634 5396 8910
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5460 8362 5488 8910
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5460 8090 5488 8298
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5184 7942 5304 7970
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5184 7410 5212 7822
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5184 7002 5212 7346
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 5092 5868 5212 5896
rect 5080 5772 5132 5778
rect 5080 5714 5132 5720
rect 5092 5234 5120 5714
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 5092 4690 5120 5170
rect 5184 4826 5212 5868
rect 5276 5030 5304 7942
rect 5460 7478 5488 8026
rect 5552 7954 5580 8978
rect 5644 7954 5672 9998
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5736 7834 5764 10390
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 5552 7806 5764 7834
rect 5448 7472 5500 7478
rect 5448 7414 5500 7420
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5460 5098 5488 5646
rect 5448 5092 5500 5098
rect 5448 5034 5500 5040
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 5092 4214 5120 4626
rect 5460 4622 5488 5034
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5460 4282 5488 4558
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5080 4208 5132 4214
rect 5080 4150 5132 4156
rect 5552 3754 5580 7806
rect 5828 7750 5856 10134
rect 5920 9654 5948 11154
rect 6196 11150 6224 12310
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6196 10198 6224 11086
rect 6184 10192 6236 10198
rect 6184 10134 6236 10140
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 6012 8634 6040 10066
rect 6196 9586 6224 10134
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6092 9376 6144 9382
rect 6184 9376 6236 9382
rect 6092 9318 6144 9324
rect 6182 9344 6184 9353
rect 6236 9344 6238 9353
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 6012 8022 6040 8434
rect 6104 8430 6132 9318
rect 6182 9279 6238 9288
rect 6092 8424 6144 8430
rect 6090 8392 6092 8401
rect 6144 8392 6146 8401
rect 6196 8362 6224 9279
rect 6090 8327 6146 8336
rect 6184 8356 6236 8362
rect 6184 8298 6236 8304
rect 6000 8016 6052 8022
rect 6000 7958 6052 7964
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 5644 5846 5672 7142
rect 6012 7002 6040 7142
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 6012 6322 6040 6734
rect 6104 6458 6132 7142
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 6012 6186 6040 6258
rect 6000 6180 6052 6186
rect 6000 6122 6052 6128
rect 5632 5840 5684 5846
rect 5632 5782 5684 5788
rect 6012 5710 6040 6122
rect 6196 6118 6224 7346
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 6288 4842 6316 13942
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 6368 12912 6420 12918
rect 6368 12854 6420 12860
rect 6380 5778 6408 12854
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6472 8294 6500 9318
rect 6460 8288 6512 8294
rect 6460 8230 6512 8236
rect 6368 5772 6420 5778
rect 6368 5714 6420 5720
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6472 5370 6500 5646
rect 6460 5364 6512 5370
rect 6460 5306 6512 5312
rect 6196 4814 6316 4842
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5368 3726 5580 3754
rect 5368 3670 5396 3726
rect 5356 3664 5408 3670
rect 5356 3606 5408 3612
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 4988 3120 5040 3126
rect 4988 3062 5040 3068
rect 5184 800 5212 3334
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5460 2106 5488 2450
rect 5448 2100 5500 2106
rect 5448 2042 5500 2048
rect 5644 800 5672 4082
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5736 2582 5764 3130
rect 5724 2576 5776 2582
rect 5724 2518 5776 2524
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 5828 1970 5856 2450
rect 5816 1964 5868 1970
rect 5816 1906 5868 1912
rect 6196 800 6224 4814
rect 6564 4146 6592 13806
rect 6886 13628 7182 13648
rect 6942 13626 6966 13628
rect 7022 13626 7046 13628
rect 7102 13626 7126 13628
rect 6964 13574 6966 13626
rect 7028 13574 7040 13626
rect 7102 13574 7104 13626
rect 6942 13572 6966 13574
rect 7022 13572 7046 13574
rect 7102 13572 7126 13574
rect 6886 13552 7182 13572
rect 6886 12540 7182 12560
rect 6942 12538 6966 12540
rect 7022 12538 7046 12540
rect 7102 12538 7126 12540
rect 6964 12486 6966 12538
rect 7028 12486 7040 12538
rect 7102 12486 7104 12538
rect 6942 12484 6966 12486
rect 7022 12484 7046 12486
rect 7102 12484 7126 12486
rect 6886 12464 7182 12484
rect 6886 11452 7182 11472
rect 6942 11450 6966 11452
rect 7022 11450 7046 11452
rect 7102 11450 7126 11452
rect 6964 11398 6966 11450
rect 7028 11398 7040 11450
rect 7102 11398 7104 11450
rect 6942 11396 6966 11398
rect 7022 11396 7046 11398
rect 7102 11396 7126 11398
rect 6886 11376 7182 11396
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6656 10606 6684 11086
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6656 10130 6684 10542
rect 6748 10470 6776 11222
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6886 10364 7182 10384
rect 6942 10362 6966 10364
rect 7022 10362 7046 10364
rect 7102 10362 7126 10364
rect 6964 10310 6966 10362
rect 7028 10310 7040 10362
rect 7102 10310 7104 10362
rect 6942 10308 6966 10310
rect 7022 10308 7046 10310
rect 7102 10308 7126 10310
rect 6886 10288 7182 10308
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6656 9042 6684 10066
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7208 9518 7236 9862
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 6886 9276 7182 9296
rect 6942 9274 6966 9276
rect 7022 9274 7046 9276
rect 7102 9274 7126 9276
rect 6964 9222 6966 9274
rect 7028 9222 7040 9274
rect 7102 9222 7104 9274
rect 6942 9220 6966 9222
rect 7022 9220 7046 9222
rect 7102 9220 7126 9222
rect 6886 9200 7182 9220
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6736 8560 6788 8566
rect 6736 8502 6788 8508
rect 6748 5778 6776 8502
rect 6886 8188 7182 8208
rect 6942 8186 6966 8188
rect 7022 8186 7046 8188
rect 7102 8186 7126 8188
rect 6964 8134 6966 8186
rect 7028 8134 7040 8186
rect 7102 8134 7104 8186
rect 6942 8132 6966 8134
rect 7022 8132 7046 8134
rect 7102 8132 7126 8134
rect 6886 8112 7182 8132
rect 7300 7993 7328 15166
rect 7392 13802 7420 16200
rect 7380 13796 7432 13802
rect 7380 13738 7432 13744
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7392 11218 7420 12038
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 7392 10674 7420 11154
rect 7668 10810 7696 12786
rect 8036 12594 8064 16200
rect 7852 12566 8064 12594
rect 7748 12164 7800 12170
rect 7748 12106 7800 12112
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7392 9586 7420 10610
rect 7668 10198 7696 10746
rect 7760 10470 7788 12106
rect 7852 11694 7880 12566
rect 8116 11756 8168 11762
rect 8116 11698 8168 11704
rect 7840 11688 7892 11694
rect 7892 11648 7972 11676
rect 7840 11630 7892 11636
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7562 10024 7618 10033
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7484 9518 7512 9998
rect 7562 9959 7618 9968
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7576 9382 7604 9959
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7760 8362 7788 10406
rect 7852 9654 7880 11494
rect 7840 9648 7892 9654
rect 7840 9590 7892 9596
rect 7748 8356 7800 8362
rect 7748 8298 7800 8304
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7484 8090 7512 8230
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7286 7984 7342 7993
rect 7286 7919 7342 7928
rect 7300 7290 7328 7919
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7300 7262 7420 7290
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 6886 7100 7182 7120
rect 6942 7098 6966 7100
rect 7022 7098 7046 7100
rect 7102 7098 7126 7100
rect 6964 7046 6966 7098
rect 7028 7046 7040 7098
rect 7102 7046 7104 7098
rect 6942 7044 6966 7046
rect 7022 7044 7046 7046
rect 7102 7044 7126 7046
rect 6886 7024 7182 7044
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7208 6186 7236 6394
rect 7196 6180 7248 6186
rect 7196 6122 7248 6128
rect 6886 6012 7182 6032
rect 6942 6010 6966 6012
rect 7022 6010 7046 6012
rect 7102 6010 7126 6012
rect 6964 5958 6966 6010
rect 7028 5958 7040 6010
rect 7102 5958 7104 6010
rect 6942 5956 6966 5958
rect 7022 5956 7046 5958
rect 7102 5956 7126 5958
rect 6886 5936 7182 5956
rect 7300 5914 7328 7142
rect 7392 6458 7420 7262
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7380 6180 7432 6186
rect 7380 6122 7432 6128
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 7392 5166 7420 6122
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7484 5642 7512 6054
rect 7668 5914 7696 7686
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7760 7002 7788 7346
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7472 5636 7524 5642
rect 7472 5578 7524 5584
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 6886 4924 7182 4944
rect 6942 4922 6966 4924
rect 7022 4922 7046 4924
rect 7102 4922 7126 4924
rect 6964 4870 6966 4922
rect 7028 4870 7040 4922
rect 7102 4870 7104 4922
rect 6942 4868 6966 4870
rect 7022 4868 7046 4870
rect 7102 4868 7126 4870
rect 6886 4848 7182 4868
rect 7392 4690 7420 5102
rect 7484 4826 7512 5578
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6886 3836 7182 3856
rect 6942 3834 6966 3836
rect 7022 3834 7046 3836
rect 7102 3834 7126 3836
rect 6964 3782 6966 3834
rect 7028 3782 7040 3834
rect 7102 3782 7104 3834
rect 6942 3780 6966 3782
rect 7022 3780 7046 3782
rect 7102 3780 7126 3782
rect 6886 3760 7182 3780
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 6656 800 6684 2586
rect 6748 2446 6776 2926
rect 6886 2748 7182 2768
rect 6942 2746 6966 2748
rect 7022 2746 7046 2748
rect 7102 2746 7126 2748
rect 6964 2694 6966 2746
rect 7028 2694 7040 2746
rect 7102 2694 7104 2746
rect 6942 2692 6966 2694
rect 7022 2692 7046 2694
rect 7102 2692 7126 2694
rect 6886 2672 7182 2692
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 7300 1442 7328 3062
rect 7484 2514 7512 3538
rect 7576 2582 7604 5510
rect 7840 5092 7892 5098
rect 7840 5034 7892 5040
rect 7656 4480 7708 4486
rect 7656 4422 7708 4428
rect 7668 3670 7696 4422
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7668 2990 7696 3606
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7852 2854 7880 5034
rect 7944 3942 7972 11648
rect 8128 11014 8156 11698
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8128 10606 8156 10950
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 8220 9382 8248 10950
rect 8312 9654 8340 11494
rect 8680 10010 8708 16200
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 9036 11620 9088 11626
rect 9036 11562 9088 11568
rect 8404 9982 8708 10010
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 8404 9382 8432 9982
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8574 9752 8630 9761
rect 8484 9716 8536 9722
rect 8574 9687 8630 9696
rect 8484 9658 8536 9664
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8392 8900 8444 8906
rect 8392 8842 8444 8848
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8220 7970 8248 8298
rect 8312 8090 8340 8774
rect 8404 8498 8432 8842
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8220 7942 8340 7970
rect 8312 7818 8340 7942
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 8404 7342 8432 8434
rect 8496 8430 8524 9658
rect 8588 9654 8616 9687
rect 8576 9648 8628 9654
rect 8864 9636 8892 9862
rect 9048 9722 9076 11562
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 8864 9608 8984 9636
rect 8576 9590 8628 9596
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8850 9344 8906 9353
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 8574 8392 8630 8401
rect 8574 8327 8576 8336
rect 8628 8327 8630 8336
rect 8576 8298 8628 8304
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8024 7268 8076 7274
rect 8024 7210 8076 7216
rect 8036 6458 8064 7210
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8128 6458 8156 6734
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8312 5692 8340 7278
rect 8588 6798 8616 7278
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8392 6724 8444 6730
rect 8392 6666 8444 6672
rect 8404 6390 8432 6666
rect 8392 6384 8444 6390
rect 8392 6326 8444 6332
rect 8312 5664 8432 5692
rect 8404 5166 8432 5664
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8404 4282 8432 5102
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8496 4078 8524 6734
rect 8588 6322 8616 6734
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8576 4548 8628 4554
rect 8576 4490 8628 4496
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 8300 4004 8352 4010
rect 8300 3946 8352 3952
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 8312 3738 8340 3946
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 8404 3194 8432 3606
rect 8588 3534 8616 4490
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8208 2916 8260 2922
rect 8208 2858 8260 2864
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 7564 2576 7616 2582
rect 7564 2518 7616 2524
rect 7852 2514 7880 2790
rect 8220 2582 8248 2858
rect 8208 2576 8260 2582
rect 8208 2518 8260 2524
rect 7472 2508 7524 2514
rect 7472 2450 7524 2456
rect 7840 2508 7892 2514
rect 7840 2450 7892 2456
rect 8588 2446 8616 3470
rect 8680 3058 8708 9318
rect 8850 9279 8906 9288
rect 8758 7304 8814 7313
rect 8864 7290 8892 9279
rect 8956 8974 8984 9608
rect 9126 9480 9182 9489
rect 9126 9415 9182 9424
rect 9140 9382 9168 9415
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 9048 9194 9076 9318
rect 9048 9166 9168 9194
rect 9140 9110 9168 9166
rect 9036 9104 9088 9110
rect 9034 9072 9036 9081
rect 9128 9104 9180 9110
rect 9088 9072 9090 9081
rect 9128 9046 9180 9052
rect 9034 9007 9090 9016
rect 8944 8968 8996 8974
rect 9036 8968 9088 8974
rect 8944 8910 8996 8916
rect 9034 8936 9036 8945
rect 9088 8936 9090 8945
rect 9034 8871 9090 8880
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 8956 7954 8984 8230
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 8814 7262 8892 7290
rect 8758 7239 8814 7248
rect 8772 7002 8800 7239
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8772 6254 8800 6734
rect 8956 6730 8984 7890
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 9048 7449 9076 7822
rect 9034 7440 9090 7449
rect 9034 7375 9090 7384
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 8944 5092 8996 5098
rect 8944 5034 8996 5040
rect 8956 4690 8984 5034
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 8956 4282 8984 4626
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 7656 2372 7708 2378
rect 7656 2314 7708 2320
rect 7116 1414 7328 1442
rect 7116 800 7144 1414
rect 7668 800 7696 2314
rect 8116 2304 8168 2310
rect 8116 2246 8168 2252
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 8128 2038 8156 2246
rect 8116 2032 8168 2038
rect 8116 1974 8168 1980
rect 8220 1170 8248 2246
rect 8772 1442 8800 3878
rect 9048 3482 9076 7375
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9140 6390 9168 6734
rect 9128 6384 9180 6390
rect 9128 6326 9180 6332
rect 9232 5778 9260 13738
rect 9324 6610 9352 16200
rect 9968 14414 9996 16200
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9852 14172 10148 14192
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 9930 14118 9932 14170
rect 9994 14118 10006 14170
rect 10068 14118 10070 14170
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 9852 14096 10148 14116
rect 9852 13084 10148 13104
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 9930 13030 9932 13082
rect 9994 13030 10006 13082
rect 10068 13030 10070 13082
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 9852 13008 10148 13028
rect 9852 11996 10148 12016
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 9930 11942 9932 11994
rect 9994 11942 10006 11994
rect 10068 11942 10070 11994
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 9852 11920 10148 11940
rect 10336 11762 10364 16215
rect 10598 16200 10654 17000
rect 11242 16200 11298 17000
rect 11886 16200 11942 17000
rect 12530 16200 12586 17000
rect 13174 16200 13230 17000
rect 13818 16200 13874 17000
rect 14462 16200 14518 17000
rect 15106 16200 15162 17000
rect 15750 16200 15806 17000
rect 16302 16688 16358 16697
rect 16302 16623 16358 16632
rect 10612 12714 10640 16200
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10704 13326 10732 13874
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10600 12708 10652 12714
rect 10600 12650 10652 12656
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9404 11620 9456 11626
rect 9404 11562 9456 11568
rect 9416 10810 9444 11562
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9586 10704 9642 10713
rect 9586 10639 9642 10648
rect 9600 10470 9628 10639
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9692 10266 9720 11630
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 10324 11212 10376 11218
rect 10324 11154 10376 11160
rect 9784 10606 9812 11154
rect 9852 10908 10148 10928
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 9930 10854 9932 10906
rect 9994 10854 10006 10906
rect 10068 10854 10070 10906
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 9852 10832 10148 10852
rect 10336 10674 10364 11154
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9784 9994 9812 10406
rect 10046 10296 10102 10305
rect 10046 10231 10048 10240
rect 10100 10231 10102 10240
rect 10048 10202 10100 10208
rect 10336 10062 10364 10610
rect 10416 10600 10468 10606
rect 10416 10542 10468 10548
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9852 9820 10148 9840
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 9930 9766 9932 9818
rect 9994 9766 10006 9818
rect 10068 9766 10070 9818
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 9852 9744 10148 9764
rect 9496 9648 9548 9654
rect 9496 9590 9548 9596
rect 9586 9616 9642 9625
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 9416 9042 9444 9522
rect 9508 9217 9536 9590
rect 9586 9551 9642 9560
rect 9494 9208 9550 9217
rect 9494 9143 9550 9152
rect 9600 9042 9628 9551
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9416 7886 9444 8978
rect 10428 8974 10456 10542
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10520 9722 10548 10406
rect 10612 10130 10640 12038
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10598 10024 10654 10033
rect 10598 9959 10654 9968
rect 10612 9926 10640 9959
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 9496 8968 9548 8974
rect 10416 8968 10468 8974
rect 9496 8910 9548 8916
rect 9586 8936 9642 8945
rect 9508 8498 9536 8910
rect 10416 8910 10468 8916
rect 9586 8871 9588 8880
rect 9640 8871 9642 8880
rect 9588 8842 9640 8848
rect 10612 8809 10640 9454
rect 10598 8800 10654 8809
rect 9852 8732 10148 8752
rect 10598 8735 10654 8744
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 9930 8678 9932 8730
rect 9994 8678 10006 8730
rect 10068 8678 10070 8730
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 9852 8656 10148 8676
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9692 7886 9720 8366
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9784 7546 9812 7958
rect 10336 7954 10364 8502
rect 10414 8392 10470 8401
rect 10414 8327 10416 8336
rect 10468 8327 10470 8336
rect 10508 8356 10560 8362
rect 10416 8298 10468 8304
rect 10508 8298 10560 8304
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 9852 7644 10148 7664
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 9930 7590 9932 7642
rect 9994 7590 10006 7642
rect 10068 7590 10070 7642
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 9852 7568 10148 7588
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 10520 7478 10548 8298
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9324 6582 9536 6610
rect 9220 5772 9272 5778
rect 9220 5714 9272 5720
rect 9232 5370 9260 5714
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 9232 4554 9260 5306
rect 9324 4758 9352 5306
rect 9404 5024 9456 5030
rect 9404 4966 9456 4972
rect 9312 4752 9364 4758
rect 9312 4694 9364 4700
rect 9220 4548 9272 4554
rect 9220 4490 9272 4496
rect 9232 4146 9260 4490
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9324 4078 9352 4694
rect 9416 4282 9444 4966
rect 9404 4276 9456 4282
rect 9404 4218 9456 4224
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9048 3454 9168 3482
rect 9036 3392 9088 3398
rect 9036 3334 9088 3340
rect 9048 3194 9076 3334
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 9048 2514 9076 3130
rect 9140 3058 9168 3454
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 9508 2922 9536 6582
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9600 3602 9628 4082
rect 9692 3670 9720 7142
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10232 6792 10284 6798
rect 10336 6769 10364 6802
rect 10232 6734 10284 6740
rect 10322 6760 10378 6769
rect 9852 6556 10148 6576
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 9930 6502 9932 6554
rect 9994 6502 10006 6554
rect 10068 6502 10070 6554
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 9852 6480 10148 6500
rect 10244 5914 10272 6734
rect 10322 6695 10378 6704
rect 10232 5908 10284 5914
rect 10232 5850 10284 5856
rect 10232 5772 10284 5778
rect 10232 5714 10284 5720
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 9852 5468 10148 5488
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 9930 5414 9932 5466
rect 9994 5414 10006 5466
rect 10068 5414 10070 5466
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 9852 5392 10148 5412
rect 9956 5160 10008 5166
rect 9956 5102 10008 5108
rect 9968 4622 9996 5102
rect 10244 5098 10272 5714
rect 10232 5092 10284 5098
rect 10232 5034 10284 5040
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 10336 4758 10364 4966
rect 10324 4752 10376 4758
rect 10324 4694 10376 4700
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 9852 4380 10148 4400
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 9930 4326 9932 4378
rect 9994 4326 10006 4378
rect 10068 4326 10070 4378
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 9852 4304 10148 4324
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9692 3058 9720 3334
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9496 2916 9548 2922
rect 9496 2858 9548 2864
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 9036 2508 9088 2514
rect 9036 2450 9088 2456
rect 8128 1142 8248 1170
rect 8680 1414 8800 1442
rect 8128 800 8156 1142
rect 8680 800 8708 1414
rect 9140 800 9168 2790
rect 9784 1986 9812 4150
rect 10336 4078 10364 4694
rect 10324 4072 10376 4078
rect 10324 4014 10376 4020
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 9852 3292 10148 3312
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 9930 3238 9932 3290
rect 9994 3238 10006 3290
rect 10068 3238 10070 3290
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 9852 3216 10148 3236
rect 9852 2204 10148 2224
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 9930 2150 9932 2202
rect 9994 2150 10006 2202
rect 10068 2150 10070 2202
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 9852 2128 10148 2148
rect 9692 1958 9812 1986
rect 9692 800 9720 1958
rect 10244 1306 10272 3538
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 10336 2378 10364 3402
rect 10428 2990 10456 5714
rect 10520 5710 10548 7414
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10612 5778 10640 6054
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10416 2984 10468 2990
rect 10416 2926 10468 2932
rect 10704 2582 10732 13262
rect 11072 13258 11100 14418
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 11060 13252 11112 13258
rect 11060 13194 11112 13200
rect 10784 11620 10836 11626
rect 10784 11562 10836 11568
rect 10796 11354 10824 11562
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 10796 9586 10824 11290
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10888 9518 10916 13194
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 10980 11082 11008 11698
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10876 9512 10928 9518
rect 10874 9480 10876 9489
rect 10928 9480 10930 9489
rect 10874 9415 10930 9424
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10888 8430 10916 8910
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10888 7478 10916 7686
rect 10876 7472 10928 7478
rect 10876 7414 10928 7420
rect 10980 6186 11008 11018
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 11072 9897 11100 10066
rect 11164 10062 11192 11630
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11058 9888 11114 9897
rect 11058 9823 11114 9832
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 11072 8537 11100 8978
rect 11256 8786 11284 16200
rect 11520 11008 11572 11014
rect 11520 10950 11572 10956
rect 11428 10736 11480 10742
rect 11426 10704 11428 10713
rect 11480 10704 11482 10713
rect 11426 10639 11482 10648
rect 11336 10532 11388 10538
rect 11336 10474 11388 10480
rect 11348 10062 11376 10474
rect 11532 10305 11560 10950
rect 11518 10296 11574 10305
rect 11518 10231 11574 10240
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11348 9722 11376 9998
rect 11900 9994 11928 16200
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12072 13252 12124 13258
rect 12072 13194 12124 13200
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 11610 9888 11666 9897
rect 11610 9823 11666 9832
rect 11336 9716 11388 9722
rect 11336 9658 11388 9664
rect 11518 9616 11574 9625
rect 11624 9586 11652 9823
rect 11518 9551 11574 9560
rect 11612 9580 11664 9586
rect 11256 8758 11376 8786
rect 11058 8528 11114 8537
rect 11058 8463 11114 8472
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 10968 6180 11020 6186
rect 10968 6122 11020 6128
rect 11072 5914 11100 7346
rect 11244 7268 11296 7274
rect 11244 7210 11296 7216
rect 11150 6896 11206 6905
rect 11150 6831 11206 6840
rect 11164 6458 11192 6831
rect 11256 6458 11284 7210
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 10980 5778 11008 5850
rect 11244 5840 11296 5846
rect 11244 5782 11296 5788
rect 10876 5772 10928 5778
rect 10876 5714 10928 5720
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10888 5370 10916 5714
rect 10876 5364 10928 5370
rect 10876 5306 10928 5312
rect 10980 4486 11008 5714
rect 11256 5681 11284 5782
rect 11242 5672 11298 5681
rect 11242 5607 11298 5616
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 11072 4758 11100 5510
rect 11348 5166 11376 8758
rect 11532 6254 11560 9551
rect 11612 9522 11664 9528
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 11992 9217 12020 9318
rect 11978 9208 12034 9217
rect 11888 9172 11940 9178
rect 11978 9143 12034 9152
rect 11888 9114 11940 9120
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11716 8634 11744 8978
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11808 7410 11836 7686
rect 11900 7585 11928 9114
rect 11980 7812 12032 7818
rect 11980 7754 12032 7760
rect 11886 7576 11942 7585
rect 11886 7511 11942 7520
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 11900 7002 11928 7346
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11808 6322 11836 6598
rect 11900 6322 11928 6938
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11900 5846 11928 6258
rect 11888 5840 11940 5846
rect 11888 5782 11940 5788
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11060 4752 11112 4758
rect 11060 4694 11112 4700
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 11428 4480 11480 4486
rect 11428 4422 11480 4428
rect 10980 3942 11008 4422
rect 11440 4078 11468 4422
rect 11808 4078 11836 4626
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11428 4072 11480 4078
rect 11796 4072 11848 4078
rect 11428 4014 11480 4020
rect 11794 4040 11796 4049
rect 11848 4040 11850 4049
rect 10968 3936 11020 3942
rect 10796 3896 10968 3924
rect 10796 3534 10824 3896
rect 10968 3878 11020 3884
rect 11440 3670 11468 4014
rect 11794 3975 11850 3984
rect 11428 3664 11480 3670
rect 11428 3606 11480 3612
rect 11900 3602 11928 4422
rect 11992 4010 12020 7754
rect 11980 4004 12032 4010
rect 11980 3946 12032 3952
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 10784 3120 10836 3126
rect 10784 3062 10836 3068
rect 10796 2922 10824 3062
rect 11808 2922 11836 3130
rect 10784 2916 10836 2922
rect 10784 2858 10836 2864
rect 11796 2916 11848 2922
rect 11796 2858 11848 2864
rect 10692 2576 10744 2582
rect 10692 2518 10744 2524
rect 12084 2446 12112 13194
rect 12164 12232 12216 12238
rect 12164 12174 12216 12180
rect 12176 11014 12204 12174
rect 12452 11370 12480 14350
rect 12544 11558 12572 16200
rect 12817 14716 13113 14736
rect 12873 14714 12897 14716
rect 12953 14714 12977 14716
rect 13033 14714 13057 14716
rect 12895 14662 12897 14714
rect 12959 14662 12971 14714
rect 13033 14662 13035 14714
rect 12873 14660 12897 14662
rect 12953 14660 12977 14662
rect 13033 14660 13057 14662
rect 12817 14640 13113 14660
rect 12817 13628 13113 13648
rect 12873 13626 12897 13628
rect 12953 13626 12977 13628
rect 13033 13626 13057 13628
rect 12895 13574 12897 13626
rect 12959 13574 12971 13626
rect 13033 13574 13035 13626
rect 12873 13572 12897 13574
rect 12953 13572 12977 13574
rect 13033 13572 13057 13574
rect 12817 13552 13113 13572
rect 12817 12540 13113 12560
rect 12873 12538 12897 12540
rect 12953 12538 12977 12540
rect 13033 12538 13057 12540
rect 12895 12486 12897 12538
rect 12959 12486 12971 12538
rect 13033 12486 13035 12538
rect 12873 12484 12897 12486
rect 12953 12484 12977 12486
rect 13033 12484 13057 12486
rect 12817 12464 13113 12484
rect 13188 12306 13216 16200
rect 13544 14000 13596 14006
rect 13544 13942 13596 13948
rect 13556 13462 13584 13942
rect 13544 13456 13596 13462
rect 13544 13398 13596 13404
rect 13832 13258 13860 16200
rect 13912 14544 13964 14550
rect 13912 14486 13964 14492
rect 13820 13252 13872 13258
rect 13820 13194 13872 13200
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 13450 11792 13506 11801
rect 13450 11727 13506 11736
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 12817 11452 13113 11472
rect 12873 11450 12897 11452
rect 12953 11450 12977 11452
rect 13033 11450 13057 11452
rect 12895 11398 12897 11450
rect 12959 11398 12971 11450
rect 13033 11398 13035 11450
rect 12873 11396 12897 11398
rect 12953 11396 12977 11398
rect 13033 11396 13057 11398
rect 12817 11376 13113 11396
rect 12452 11342 12572 11370
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 12162 10568 12218 10577
rect 12162 10503 12218 10512
rect 12176 9450 12204 10503
rect 12360 9994 12388 11086
rect 12452 10606 12480 11086
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12452 10266 12480 10542
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12256 9988 12308 9994
rect 12256 9930 12308 9936
rect 12348 9988 12400 9994
rect 12348 9930 12400 9936
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 12268 9178 12296 9930
rect 12360 9722 12388 9930
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12256 9172 12308 9178
rect 12256 9114 12308 9120
rect 12360 9081 12388 9318
rect 12346 9072 12402 9081
rect 12164 9036 12216 9042
rect 12346 9007 12402 9016
rect 12164 8978 12216 8984
rect 12176 7818 12204 8978
rect 12452 8922 12480 9658
rect 12268 8894 12480 8922
rect 12268 8294 12296 8894
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12256 8288 12308 8294
rect 12256 8230 12308 8236
rect 12360 7886 12388 8774
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12164 7812 12216 7818
rect 12164 7754 12216 7760
rect 12346 7576 12402 7585
rect 12346 7511 12402 7520
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12176 6254 12204 6598
rect 12360 6322 12388 7511
rect 12452 6798 12480 8502
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 12348 6180 12400 6186
rect 12348 6122 12400 6128
rect 12254 5808 12310 5817
rect 12254 5743 12256 5752
rect 12308 5743 12310 5752
rect 12256 5714 12308 5720
rect 12360 5234 12388 6122
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 12452 4486 12480 6734
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 11060 2440 11112 2446
rect 11612 2440 11664 2446
rect 11112 2400 11192 2428
rect 11060 2382 11112 2388
rect 10324 2372 10376 2378
rect 10324 2314 10376 2320
rect 10336 1970 10364 2314
rect 10600 2304 10652 2310
rect 10600 2246 10652 2252
rect 10324 1964 10376 1970
rect 10324 1906 10376 1912
rect 10152 1278 10272 1306
rect 10152 800 10180 1278
rect 10612 800 10640 2246
rect 11164 800 11192 2400
rect 11612 2382 11664 2388
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 11624 800 11652 2382
rect 12176 800 12204 3470
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12256 3120 12308 3126
rect 12254 3088 12256 3097
rect 12308 3088 12310 3097
rect 12360 3058 12388 3334
rect 12544 3210 12572 11342
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12636 10810 12664 11154
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12817 10364 13113 10384
rect 12873 10362 12897 10364
rect 12953 10362 12977 10364
rect 13033 10362 13057 10364
rect 12895 10310 12897 10362
rect 12959 10310 12971 10362
rect 13033 10310 13035 10362
rect 12873 10308 12897 10310
rect 12953 10308 12977 10310
rect 13033 10308 13057 10310
rect 12817 10288 13113 10308
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12636 8378 12664 10134
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 12728 9178 12756 10066
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12820 9722 12848 9998
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 13188 9636 13216 11494
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13280 10674 13308 11154
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13464 10606 13492 11727
rect 13636 11008 13688 11014
rect 13636 10950 13688 10956
rect 13648 10742 13676 10950
rect 13636 10736 13688 10742
rect 13636 10678 13688 10684
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13464 10198 13492 10542
rect 13452 10192 13504 10198
rect 13452 10134 13504 10140
rect 13157 9608 13216 9636
rect 12806 9480 12862 9489
rect 13157 9466 13185 9608
rect 13556 9586 13584 10610
rect 13636 10600 13688 10606
rect 13636 10542 13688 10548
rect 13648 10130 13676 10542
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13157 9438 13216 9466
rect 12806 9415 12808 9424
rect 12860 9415 12862 9424
rect 12808 9386 12860 9392
rect 12817 9276 13113 9296
rect 12873 9274 12897 9276
rect 12953 9274 12977 9276
rect 13033 9274 13057 9276
rect 12895 9222 12897 9274
rect 12959 9222 12971 9274
rect 13033 9222 13035 9274
rect 12873 9220 12897 9222
rect 12953 9220 12977 9222
rect 13033 9220 13057 9222
rect 12817 9200 13113 9220
rect 13188 9178 13216 9438
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13084 9104 13136 9110
rect 12990 9072 13046 9081
rect 13084 9046 13136 9052
rect 12990 9007 12992 9016
rect 13044 9007 13046 9016
rect 12992 8978 13044 8984
rect 12992 8900 13044 8906
rect 12992 8842 13044 8848
rect 13004 8634 13032 8842
rect 13096 8809 13124 9046
rect 13556 8974 13584 9522
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 13082 8800 13138 8809
rect 13082 8735 13138 8744
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 12636 8350 12756 8378
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12636 8090 12664 8230
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12622 7848 12678 7857
rect 12622 7783 12678 7792
rect 12636 7274 12664 7783
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 12636 7002 12664 7210
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12728 6769 12756 8350
rect 12817 8188 13113 8208
rect 12873 8186 12897 8188
rect 12953 8186 12977 8188
rect 13033 8186 13057 8188
rect 12895 8134 12897 8186
rect 12959 8134 12971 8186
rect 13033 8134 13035 8186
rect 12873 8132 12897 8134
rect 12953 8132 12977 8134
rect 13033 8132 13057 8134
rect 12817 8112 13113 8132
rect 13280 8090 13308 8842
rect 13648 8838 13676 10066
rect 13740 9602 13768 12786
rect 13740 9574 13860 9602
rect 13832 9364 13860 9574
rect 13740 9336 13860 9364
rect 13636 8832 13688 8838
rect 13556 8792 13636 8820
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 13096 7478 13124 7686
rect 13084 7472 13136 7478
rect 13084 7414 13136 7420
rect 13188 7410 13216 7822
rect 13280 7818 13308 8026
rect 13464 7886 13492 8434
rect 13556 8362 13584 8792
rect 13636 8774 13688 8780
rect 13740 8514 13768 9336
rect 13924 9194 13952 14486
rect 14004 14340 14056 14346
rect 14004 14282 14056 14288
rect 14016 12986 14044 14282
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 14200 13462 14228 14214
rect 14476 13954 14504 16200
rect 15120 13954 15148 16200
rect 15566 15872 15622 15881
rect 15566 15807 15622 15816
rect 15198 15464 15254 15473
rect 15198 15399 15254 15408
rect 14384 13926 14504 13954
rect 15028 13926 15148 13954
rect 14384 13870 14412 13926
rect 15028 13870 15056 13926
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 14832 13796 14884 13802
rect 14832 13738 14884 13744
rect 14188 13456 14240 13462
rect 14188 13398 14240 13404
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 13648 8486 13768 8514
rect 13832 9166 13952 9194
rect 13544 8356 13596 8362
rect 13544 8298 13596 8304
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13268 7812 13320 7818
rect 13268 7754 13320 7760
rect 13556 7410 13584 8298
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 12817 7100 13113 7120
rect 12873 7098 12897 7100
rect 12953 7098 12977 7100
rect 13033 7098 13057 7100
rect 12895 7046 12897 7098
rect 12959 7046 12971 7098
rect 13033 7046 13035 7098
rect 12873 7044 12897 7046
rect 12953 7044 12977 7046
rect 13033 7044 13057 7046
rect 12817 7024 13113 7044
rect 13188 6866 13216 7346
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 13280 7002 13308 7278
rect 13648 7002 13676 8486
rect 13728 8424 13780 8430
rect 13726 8392 13728 8401
rect 13780 8392 13782 8401
rect 13726 8327 13782 8336
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13176 6860 13228 6866
rect 13176 6802 13228 6808
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 12714 6760 12770 6769
rect 13188 6730 13216 6802
rect 12714 6695 12770 6704
rect 13176 6724 13228 6730
rect 13176 6666 13228 6672
rect 13464 6390 13492 6802
rect 13832 6780 13860 9166
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13924 7546 13952 7822
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 13556 6752 13860 6780
rect 13452 6384 13504 6390
rect 13452 6326 13504 6332
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 12716 6180 12768 6186
rect 12716 6122 12768 6128
rect 12728 5817 12756 6122
rect 12817 6012 13113 6032
rect 12873 6010 12897 6012
rect 12953 6010 12977 6012
rect 13033 6010 13057 6012
rect 12895 5958 12897 6010
rect 12959 5958 12971 6010
rect 13033 5958 13035 6010
rect 12873 5956 12897 5958
rect 12953 5956 12977 5958
rect 13033 5956 13057 5958
rect 12817 5936 13113 5956
rect 12714 5808 12770 5817
rect 12714 5743 12770 5752
rect 12728 5710 12756 5743
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12636 5098 12664 5306
rect 12624 5092 12676 5098
rect 12624 5034 12676 5040
rect 12817 4924 13113 4944
rect 12873 4922 12897 4924
rect 12953 4922 12977 4924
rect 13033 4922 13057 4924
rect 12895 4870 12897 4922
rect 12959 4870 12971 4922
rect 13033 4870 13035 4922
rect 12873 4868 12897 4870
rect 12953 4868 12977 4870
rect 13033 4868 13057 4870
rect 12817 4848 13113 4868
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 12544 3182 12664 3210
rect 12532 3120 12584 3126
rect 12530 3088 12532 3097
rect 12584 3088 12586 3097
rect 12254 3023 12310 3032
rect 12348 3052 12400 3058
rect 12636 3058 12664 3182
rect 12530 3023 12586 3032
rect 12624 3052 12676 3058
rect 12348 2994 12400 3000
rect 12624 2994 12676 3000
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12452 2582 12480 2790
rect 12440 2576 12492 2582
rect 12440 2518 12492 2524
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 12636 800 12664 2382
rect 12728 1698 12756 4422
rect 13188 4078 13216 6258
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 12817 3836 13113 3856
rect 12873 3834 12897 3836
rect 12953 3834 12977 3836
rect 13033 3834 13057 3836
rect 12895 3782 12897 3834
rect 12959 3782 12971 3834
rect 13033 3782 13035 3834
rect 12873 3780 12897 3782
rect 12953 3780 12977 3782
rect 13033 3780 13057 3782
rect 12817 3760 13113 3780
rect 13176 2916 13228 2922
rect 13176 2858 13228 2864
rect 12817 2748 13113 2768
rect 12873 2746 12897 2748
rect 12953 2746 12977 2748
rect 13033 2746 13057 2748
rect 12895 2694 12897 2746
rect 12959 2694 12971 2746
rect 13033 2694 13035 2746
rect 12873 2692 12897 2694
rect 12953 2692 12977 2694
rect 13033 2692 13057 2694
rect 12817 2672 13113 2692
rect 13084 2576 13136 2582
rect 13188 2530 13216 2858
rect 13136 2524 13216 2530
rect 13084 2518 13216 2524
rect 13096 2502 13216 2518
rect 13188 2446 13216 2502
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 12716 1692 12768 1698
rect 12716 1634 12768 1640
rect 13280 898 13308 4558
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13464 1970 13492 3878
rect 13556 3670 13584 6752
rect 13636 5092 13688 5098
rect 13636 5034 13688 5040
rect 13648 4078 13676 5034
rect 13728 5024 13780 5030
rect 13726 4992 13728 5001
rect 13820 5024 13872 5030
rect 13780 4992 13782 5001
rect 13820 4966 13872 4972
rect 13726 4927 13782 4936
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 13832 2564 13860 4966
rect 14016 4758 14044 12922
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14108 8838 14136 9318
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 14108 8634 14136 8774
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 14108 6866 14136 7482
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 14004 4752 14056 4758
rect 14004 4694 14056 4700
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 13912 3664 13964 3670
rect 13912 3606 13964 3612
rect 13924 2582 13952 3606
rect 13648 2536 13860 2564
rect 13912 2576 13964 2582
rect 13452 1964 13504 1970
rect 13452 1906 13504 1912
rect 13188 870 13308 898
rect 13188 800 13216 870
rect 13648 800 13676 2536
rect 13912 2518 13964 2524
rect 14016 1766 14044 3878
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 14108 3058 14136 3538
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 14200 2582 14228 13398
rect 14372 12708 14424 12714
rect 14372 12650 14424 12656
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14292 8566 14320 10950
rect 14280 8560 14332 8566
rect 14280 8502 14332 8508
rect 14280 7948 14332 7954
rect 14280 7890 14332 7896
rect 14292 7750 14320 7890
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 14292 6934 14320 7686
rect 14280 6928 14332 6934
rect 14280 6870 14332 6876
rect 14280 6180 14332 6186
rect 14280 6122 14332 6128
rect 14292 5914 14320 6122
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 14280 4004 14332 4010
rect 14280 3946 14332 3952
rect 14188 2576 14240 2582
rect 14188 2518 14240 2524
rect 14004 1760 14056 1766
rect 14004 1702 14056 1708
rect 14292 1442 14320 3946
rect 14384 3058 14412 12650
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 14476 2106 14504 9318
rect 14568 5710 14596 12242
rect 14740 9036 14792 9042
rect 14740 8978 14792 8984
rect 14648 7948 14700 7954
rect 14648 7890 14700 7896
rect 14556 5704 14608 5710
rect 14556 5646 14608 5652
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14568 2360 14596 4558
rect 14660 2938 14688 7890
rect 14752 7857 14780 8978
rect 14738 7848 14794 7857
rect 14738 7783 14794 7792
rect 14740 7472 14792 7478
rect 14740 7414 14792 7420
rect 14752 3058 14780 7414
rect 14844 5234 14872 13738
rect 15016 13252 15068 13258
rect 15016 13194 15068 13200
rect 14924 10532 14976 10538
rect 14924 10474 14976 10480
rect 14936 10266 14964 10474
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 14936 9586 14964 10202
rect 14924 9580 14976 9586
rect 14924 9522 14976 9528
rect 14924 8356 14976 8362
rect 14924 8298 14976 8304
rect 14936 7886 14964 8298
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 15028 7478 15056 13194
rect 15016 7472 15068 7478
rect 15016 7414 15068 7420
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 14936 6798 14964 7346
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 15028 7206 15056 7278
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 15028 6458 15056 6734
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 15120 4146 15148 13926
rect 15212 12782 15240 15399
rect 15290 15056 15346 15065
rect 15290 14991 15346 15000
rect 15304 13841 15332 14991
rect 15384 13864 15436 13870
rect 15290 13832 15346 13841
rect 15384 13806 15436 13812
rect 15474 13832 15530 13841
rect 15290 13767 15346 13776
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15304 13530 15332 13670
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15290 13424 15346 13433
rect 15290 13359 15346 13368
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15304 12594 15332 13359
rect 15212 12566 15332 12594
rect 15212 11150 15240 12566
rect 15396 12458 15424 13806
rect 15474 13767 15530 13776
rect 15304 12430 15424 12458
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 15212 9926 15240 10066
rect 15200 9920 15252 9926
rect 15200 9862 15252 9868
rect 15212 9586 15240 9862
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15304 9489 15332 12430
rect 15384 12368 15436 12374
rect 15384 12310 15436 12316
rect 15396 10713 15424 12310
rect 15488 11626 15516 13767
rect 15580 12866 15608 15807
rect 15764 14362 15792 16200
rect 16118 14648 16174 14657
rect 16118 14583 16174 14592
rect 15672 14334 15792 14362
rect 15672 14006 15700 14334
rect 15782 14172 16078 14192
rect 15838 14170 15862 14172
rect 15918 14170 15942 14172
rect 15998 14170 16022 14172
rect 15860 14118 15862 14170
rect 15924 14118 15936 14170
rect 15998 14118 16000 14170
rect 15838 14116 15862 14118
rect 15918 14116 15942 14118
rect 15998 14116 16022 14118
rect 15782 14096 16078 14116
rect 15660 14000 15712 14006
rect 15660 13942 15712 13948
rect 15844 13728 15896 13734
rect 15844 13670 15896 13676
rect 15856 13394 15884 13670
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15782 13084 16078 13104
rect 15838 13082 15862 13084
rect 15918 13082 15942 13084
rect 15998 13082 16022 13084
rect 15860 13030 15862 13082
rect 15924 13030 15936 13082
rect 15998 13030 16000 13082
rect 15838 13028 15862 13030
rect 15918 13028 15942 13030
rect 15998 13028 16022 13030
rect 15782 13008 16078 13028
rect 15580 12838 15792 12866
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 15580 12442 15608 12718
rect 15658 12472 15714 12481
rect 15568 12436 15620 12442
rect 15658 12407 15714 12416
rect 15568 12378 15620 12384
rect 15672 12322 15700 12407
rect 15580 12294 15700 12322
rect 15476 11620 15528 11626
rect 15476 11562 15528 11568
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15382 10704 15438 10713
rect 15382 10639 15438 10648
rect 15488 10554 15516 11086
rect 15580 11014 15608 12294
rect 15764 12186 15792 12838
rect 15672 12158 15792 12186
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15672 10742 15700 12158
rect 15782 11996 16078 12016
rect 15838 11994 15862 11996
rect 15918 11994 15942 11996
rect 15998 11994 16022 11996
rect 15860 11942 15862 11994
rect 15924 11942 15936 11994
rect 15998 11942 16000 11994
rect 15838 11940 15862 11942
rect 15918 11940 15942 11942
rect 15998 11940 16022 11942
rect 15782 11920 16078 11940
rect 15782 10908 16078 10928
rect 15838 10906 15862 10908
rect 15918 10906 15942 10908
rect 15998 10906 16022 10908
rect 15860 10854 15862 10906
rect 15924 10854 15936 10906
rect 15998 10854 16000 10906
rect 15838 10852 15862 10854
rect 15918 10852 15942 10854
rect 15998 10852 16022 10854
rect 15782 10832 16078 10852
rect 15660 10736 15712 10742
rect 15660 10678 15712 10684
rect 15672 10577 15700 10678
rect 15658 10568 15714 10577
rect 15488 10526 15608 10554
rect 15476 10464 15528 10470
rect 15382 10432 15438 10441
rect 15476 10406 15528 10412
rect 15382 10367 15438 10376
rect 15396 9722 15424 10367
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15488 9518 15516 10406
rect 15476 9512 15528 9518
rect 15290 9480 15346 9489
rect 15476 9454 15528 9460
rect 15290 9415 15346 9424
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15200 7948 15252 7954
rect 15200 7890 15252 7896
rect 15212 7206 15240 7890
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15212 5302 15240 7142
rect 15200 5296 15252 5302
rect 15200 5238 15252 5244
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15212 4826 15240 4966
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 15016 3732 15068 3738
rect 15016 3674 15068 3680
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14660 2910 14872 2938
rect 14844 2582 14872 2910
rect 15028 2650 15056 3674
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 15120 2854 15148 3538
rect 15212 2854 15240 4626
rect 15304 4146 15332 9114
rect 15580 8514 15608 10526
rect 15658 10503 15714 10512
rect 16132 10282 16160 14583
rect 16212 13932 16264 13938
rect 16212 13874 16264 13880
rect 15672 10254 16160 10282
rect 15672 9625 15700 10254
rect 16120 10124 16172 10130
rect 16120 10066 16172 10072
rect 15782 9820 16078 9840
rect 15838 9818 15862 9820
rect 15918 9818 15942 9820
rect 15998 9818 16022 9820
rect 15860 9766 15862 9818
rect 15924 9766 15936 9818
rect 15998 9766 16000 9818
rect 15838 9764 15862 9766
rect 15918 9764 15942 9766
rect 15998 9764 16022 9766
rect 15782 9744 16078 9764
rect 15658 9616 15714 9625
rect 16132 9586 16160 10066
rect 15658 9551 15714 9560
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 15672 9178 15700 9318
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 15782 8732 16078 8752
rect 15838 8730 15862 8732
rect 15918 8730 15942 8732
rect 15998 8730 16022 8732
rect 15860 8678 15862 8730
rect 15924 8678 15936 8730
rect 15998 8678 16000 8730
rect 15838 8676 15862 8678
rect 15918 8676 15942 8678
rect 15998 8676 16022 8678
rect 15782 8656 16078 8676
rect 16132 8634 16160 9522
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 15488 8486 15608 8514
rect 15488 7546 15516 8486
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 15568 8356 15620 8362
rect 15568 8298 15620 8304
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15396 5030 15424 6802
rect 15488 5234 15516 7142
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15580 4758 15608 8298
rect 15782 7644 16078 7664
rect 15838 7642 15862 7644
rect 15918 7642 15942 7644
rect 15998 7642 16022 7644
rect 15860 7590 15862 7642
rect 15924 7590 15936 7642
rect 15998 7590 16000 7642
rect 15838 7588 15862 7590
rect 15918 7588 15942 7590
rect 15998 7588 16022 7590
rect 15782 7568 16078 7588
rect 16132 7546 16160 8366
rect 16120 7540 16172 7546
rect 16120 7482 16172 7488
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 15672 5914 15700 7142
rect 15782 6556 16078 6576
rect 15838 6554 15862 6556
rect 15918 6554 15942 6556
rect 15998 6554 16022 6556
rect 15860 6502 15862 6554
rect 15924 6502 15936 6554
rect 15998 6502 16000 6554
rect 15838 6500 15862 6502
rect 15918 6500 15942 6502
rect 15998 6500 16022 6502
rect 15782 6480 16078 6500
rect 16132 6458 16160 7142
rect 16120 6452 16172 6458
rect 16120 6394 16172 6400
rect 15936 6248 15988 6254
rect 15936 6190 15988 6196
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15568 4752 15620 4758
rect 15568 4694 15620 4700
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15672 3670 15700 5646
rect 15948 5642 15976 6190
rect 16028 5840 16080 5846
rect 16028 5782 16080 5788
rect 16040 5681 16068 5782
rect 16026 5672 16082 5681
rect 15936 5636 15988 5642
rect 16026 5607 16082 5616
rect 15936 5578 15988 5584
rect 15782 5468 16078 5488
rect 15838 5466 15862 5468
rect 15918 5466 15942 5468
rect 15998 5466 16022 5468
rect 15860 5414 15862 5466
rect 15924 5414 15936 5466
rect 15998 5414 16000 5466
rect 15838 5412 15862 5414
rect 15918 5412 15942 5414
rect 15998 5412 16022 5414
rect 15782 5392 16078 5412
rect 16224 4622 16252 13874
rect 16316 13682 16344 16623
rect 16394 16200 16450 17000
rect 17038 16200 17094 17000
rect 17682 16200 17738 17000
rect 18326 16200 18382 17000
rect 18970 16200 19026 17000
rect 19614 16200 19670 17000
rect 16408 13870 16436 16200
rect 16486 14240 16542 14249
rect 16486 14175 16542 14184
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 16316 13654 16436 13682
rect 16302 12880 16358 12889
rect 16302 12815 16358 12824
rect 16316 12050 16344 12815
rect 16408 12238 16436 13654
rect 16396 12232 16448 12238
rect 16396 12174 16448 12180
rect 16500 12102 16528 14175
rect 17052 13326 17080 16200
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 17498 13288 17554 13297
rect 17498 13223 17554 13232
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16488 12096 16540 12102
rect 16316 12022 16436 12050
rect 16488 12038 16540 12044
rect 16408 10985 16436 12022
rect 16592 11257 16620 12106
rect 17316 11824 17368 11830
rect 17316 11766 17368 11772
rect 16578 11248 16634 11257
rect 16578 11183 16634 11192
rect 16394 10976 16450 10985
rect 16394 10911 16450 10920
rect 16670 10840 16726 10849
rect 16670 10775 16726 10784
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16408 10266 16436 10406
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16394 10160 16450 10169
rect 16394 10095 16450 10104
rect 16408 9330 16436 10095
rect 16500 9926 16528 10610
rect 16684 10169 16712 10775
rect 16670 10160 16726 10169
rect 16670 10095 16726 10104
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 16578 10024 16634 10033
rect 16578 9959 16634 9968
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16592 9518 16620 9959
rect 17130 9888 17186 9897
rect 17130 9823 17186 9832
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 16672 9376 16724 9382
rect 16408 9302 16528 9330
rect 16672 9318 16724 9324
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 15782 4380 16078 4400
rect 15838 4378 15862 4380
rect 15918 4378 15942 4380
rect 15998 4378 16022 4380
rect 15860 4326 15862 4378
rect 15924 4326 15936 4378
rect 15998 4326 16000 4378
rect 15838 4324 15862 4326
rect 15918 4324 15942 4326
rect 15998 4324 16022 4326
rect 15782 4304 16078 4324
rect 15752 4208 15804 4214
rect 15752 4150 15804 4156
rect 15764 4010 15792 4150
rect 15752 4004 15804 4010
rect 15752 3946 15804 3952
rect 15660 3664 15712 3670
rect 15660 3606 15712 3612
rect 15660 3460 15712 3466
rect 15660 3402 15712 3408
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 15016 2644 15068 2650
rect 15016 2586 15068 2592
rect 14832 2576 14884 2582
rect 14832 2518 14884 2524
rect 15292 2576 15344 2582
rect 15292 2518 15344 2524
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 14568 2332 14688 2360
rect 14464 2100 14516 2106
rect 14464 2042 14516 2048
rect 14108 1414 14320 1442
rect 14108 800 14136 1414
rect 14660 800 14688 2332
rect 15120 800 15148 2382
rect 15304 2038 15332 2518
rect 15292 2032 15344 2038
rect 15292 1974 15344 1980
rect 15672 800 15700 3402
rect 16120 3392 16172 3398
rect 16120 3334 16172 3340
rect 15782 3292 16078 3312
rect 15838 3290 15862 3292
rect 15918 3290 15942 3292
rect 15998 3290 16022 3292
rect 15860 3238 15862 3290
rect 15924 3238 15936 3290
rect 15998 3238 16000 3290
rect 15838 3236 15862 3238
rect 15918 3236 15942 3238
rect 15998 3236 16022 3238
rect 15782 3216 16078 3236
rect 15936 2916 15988 2922
rect 15936 2858 15988 2864
rect 15842 2544 15898 2553
rect 15842 2479 15898 2488
rect 15856 2446 15884 2479
rect 15844 2440 15896 2446
rect 15844 2382 15896 2388
rect 15948 2378 15976 2858
rect 15936 2372 15988 2378
rect 15936 2314 15988 2320
rect 15782 2204 16078 2224
rect 15838 2202 15862 2204
rect 15918 2202 15942 2204
rect 15998 2202 16022 2204
rect 15860 2150 15862 2202
rect 15924 2150 15936 2202
rect 15998 2150 16000 2202
rect 15838 2148 15862 2150
rect 15918 2148 15942 2150
rect 15998 2148 16022 2150
rect 15782 2128 16078 2148
rect 16132 800 16160 3334
rect 16224 3058 16252 4422
rect 16316 4049 16344 7482
rect 16408 7342 16436 9114
rect 16500 7750 16528 9302
rect 16684 9178 16712 9318
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16592 8634 16620 8910
rect 16776 8634 16804 9318
rect 17144 9178 17172 9823
rect 17236 9586 17264 10066
rect 17224 9580 17276 9586
rect 17224 9522 17276 9528
rect 17132 9172 17184 9178
rect 17052 9132 17132 9160
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16684 8090 16712 8434
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16396 7336 16448 7342
rect 16396 7278 16448 7284
rect 16500 7290 16528 7346
rect 16408 6390 16436 7278
rect 16500 7262 16620 7290
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16500 7002 16528 7142
rect 16592 7002 16620 7262
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 16580 6996 16632 7002
rect 16580 6938 16632 6944
rect 16486 6896 16542 6905
rect 16486 6831 16542 6840
rect 16500 6798 16528 6831
rect 16488 6792 16540 6798
rect 16488 6734 16540 6740
rect 16396 6384 16448 6390
rect 16396 6326 16448 6332
rect 16500 6254 16528 6734
rect 16684 6254 16712 7210
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16776 7041 16804 7142
rect 16762 7032 16818 7041
rect 16762 6967 16818 6976
rect 16764 6860 16816 6866
rect 16764 6802 16816 6808
rect 16776 6322 16804 6802
rect 16764 6316 16816 6322
rect 16764 6258 16816 6264
rect 16488 6248 16540 6254
rect 16488 6190 16540 6196
rect 16672 6248 16724 6254
rect 16672 6190 16724 6196
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 16500 5914 16528 6054
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16488 5636 16540 5642
rect 16488 5578 16540 5584
rect 16500 4214 16528 5578
rect 16592 5370 16620 6054
rect 16672 5772 16724 5778
rect 16672 5714 16724 5720
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 16578 4992 16634 5001
rect 16578 4927 16634 4936
rect 16488 4208 16540 4214
rect 16488 4150 16540 4156
rect 16302 4040 16358 4049
rect 16592 4010 16620 4927
rect 16684 4826 16712 5714
rect 16776 5710 16804 6258
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 16764 5296 16816 5302
rect 16764 5238 16816 5244
rect 16672 4820 16724 4826
rect 16672 4762 16724 4768
rect 16302 3975 16358 3984
rect 16580 4004 16632 4010
rect 16316 3670 16344 3975
rect 16580 3946 16632 3952
rect 16304 3664 16356 3670
rect 16304 3606 16356 3612
rect 16672 3460 16724 3466
rect 16672 3402 16724 3408
rect 16212 3052 16264 3058
rect 16212 2994 16264 3000
rect 16684 800 16712 3402
rect 16776 2922 16804 5238
rect 16868 5030 16896 8774
rect 16960 8090 16988 8978
rect 17052 8906 17080 9132
rect 17132 9114 17184 9120
rect 17130 9072 17186 9081
rect 17328 9058 17356 11766
rect 17406 11248 17462 11257
rect 17406 11183 17462 11192
rect 17420 9602 17448 11183
rect 17512 10266 17540 13223
rect 17696 13190 17724 16200
rect 18340 14550 18368 16200
rect 18328 14544 18380 14550
rect 18328 14486 18380 14492
rect 18984 13462 19012 16200
rect 18972 13456 19024 13462
rect 18972 13398 19024 13404
rect 17684 13184 17736 13190
rect 17684 13126 17736 13132
rect 19628 12986 19656 16200
rect 19616 12980 19668 12986
rect 19616 12922 19668 12928
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17788 11665 17816 11834
rect 17774 11656 17830 11665
rect 17774 11591 17830 11600
rect 17592 10668 17644 10674
rect 17592 10610 17644 10616
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17512 9722 17540 10202
rect 17604 10198 17632 10610
rect 17592 10192 17644 10198
rect 17592 10134 17644 10140
rect 17500 9716 17552 9722
rect 17500 9658 17552 9664
rect 17420 9574 17724 9602
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17328 9030 17448 9058
rect 17130 9007 17186 9016
rect 17040 8900 17092 8906
rect 17040 8842 17092 8848
rect 17038 8664 17094 8673
rect 17038 8599 17094 8608
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 16946 7848 17002 7857
rect 16946 7783 17002 7792
rect 16960 5778 16988 7783
rect 16948 5772 17000 5778
rect 16948 5714 17000 5720
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16856 4548 16908 4554
rect 16856 4490 16908 4496
rect 16868 3670 16896 4490
rect 16856 3664 16908 3670
rect 16856 3606 16908 3612
rect 16764 2916 16816 2922
rect 16764 2858 16816 2864
rect 16960 2446 16988 5714
rect 17052 5166 17080 8599
rect 17144 8566 17172 9007
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17144 8430 17172 8502
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 17132 8288 17184 8294
rect 17132 8230 17184 8236
rect 17144 7834 17172 8230
rect 17236 7954 17264 8910
rect 17328 8498 17356 8910
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 17314 7984 17370 7993
rect 17224 7948 17276 7954
rect 17420 7954 17448 9030
rect 17604 8265 17632 9318
rect 17590 8256 17646 8265
rect 17590 8191 17646 8200
rect 17592 8016 17644 8022
rect 17592 7958 17644 7964
rect 17314 7919 17370 7928
rect 17408 7948 17460 7954
rect 17224 7890 17276 7896
rect 17144 7806 17264 7834
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 17040 5160 17092 5166
rect 17040 5102 17092 5108
rect 17144 4706 17172 7686
rect 17236 7342 17264 7806
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 17328 7002 17356 7919
rect 17408 7890 17460 7896
rect 17420 7750 17448 7890
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 17500 7404 17552 7410
rect 17500 7346 17552 7352
rect 17316 6996 17368 7002
rect 17316 6938 17368 6944
rect 17408 6928 17460 6934
rect 17408 6870 17460 6876
rect 17224 6180 17276 6186
rect 17224 6122 17276 6128
rect 17236 5710 17264 6122
rect 17224 5704 17276 5710
rect 17224 5646 17276 5652
rect 17236 5234 17264 5646
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 17052 4678 17172 4706
rect 17052 3670 17080 4678
rect 17236 4622 17264 5170
rect 17420 4690 17448 6870
rect 17512 6798 17540 7346
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17512 6322 17540 6734
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 17408 4684 17460 4690
rect 17408 4626 17460 4632
rect 17132 4616 17184 4622
rect 17132 4558 17184 4564
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 17144 4282 17172 4558
rect 17132 4276 17184 4282
rect 17132 4218 17184 4224
rect 17144 3720 17172 4218
rect 17512 4078 17540 4966
rect 17604 4146 17632 7958
rect 17696 7290 17724 9574
rect 17788 8090 17816 11591
rect 18052 11212 18104 11218
rect 18052 11154 18104 11160
rect 17868 11008 17920 11014
rect 17868 10950 17920 10956
rect 17776 8084 17828 8090
rect 17776 8026 17828 8032
rect 17880 8022 17908 10950
rect 18064 10130 18092 11154
rect 18512 10600 18564 10606
rect 18512 10542 18564 10548
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 17972 9042 18000 9522
rect 18328 9376 18380 9382
rect 18328 9318 18380 9324
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 17972 8537 18000 8978
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 17958 8528 18014 8537
rect 17958 8463 18014 8472
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 17868 8016 17920 8022
rect 17972 7993 18000 8366
rect 17868 7958 17920 7964
rect 17958 7984 18014 7993
rect 17958 7919 18014 7928
rect 18064 7449 18092 8774
rect 18236 8288 18288 8294
rect 18236 8230 18288 8236
rect 18050 7440 18106 7449
rect 18050 7375 18106 7384
rect 17958 7304 18014 7313
rect 17696 7262 17816 7290
rect 17684 7200 17736 7206
rect 17684 7142 17736 7148
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17500 4072 17552 4078
rect 17500 4014 17552 4020
rect 17592 3936 17644 3942
rect 17592 3878 17644 3884
rect 17144 3692 17264 3720
rect 17040 3664 17092 3670
rect 17040 3606 17092 3612
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 17144 800 17172 2994
rect 17236 2990 17264 3692
rect 17604 3641 17632 3878
rect 17590 3632 17646 3641
rect 17590 3567 17646 3576
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 17592 2848 17644 2854
rect 17592 2790 17644 2796
rect 17604 2689 17632 2790
rect 17590 2680 17646 2689
rect 17590 2615 17646 2624
rect 17592 2440 17644 2446
rect 17592 2382 17644 2388
rect 17316 2304 17368 2310
rect 17314 2272 17316 2281
rect 17368 2272 17370 2281
rect 17314 2207 17370 2216
rect 17604 1873 17632 2382
rect 17590 1864 17646 1873
rect 17590 1799 17646 1808
rect 17592 1760 17644 1766
rect 17592 1702 17644 1708
rect 17604 800 17632 1702
rect 3054 232 3110 241
rect 3054 167 3110 176
rect 3146 0 3202 800
rect 3606 0 3662 800
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 5170 0 5226 800
rect 5630 0 5686 800
rect 6182 0 6238 800
rect 6642 0 6698 800
rect 7102 0 7158 800
rect 7654 0 7710 800
rect 8114 0 8170 800
rect 8666 0 8722 800
rect 9126 0 9182 800
rect 9678 0 9734 800
rect 10138 0 10194 800
rect 10598 0 10654 800
rect 11150 0 11206 800
rect 11610 0 11666 800
rect 12162 0 12218 800
rect 12622 0 12678 800
rect 13174 0 13230 800
rect 13634 0 13690 800
rect 14094 0 14150 800
rect 14646 0 14702 800
rect 15106 0 15162 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16670 0 16726 800
rect 17130 0 17186 800
rect 17590 0 17646 800
rect 17696 649 17724 7142
rect 17788 5658 17816 7262
rect 17958 7239 18014 7248
rect 17972 6866 18000 7239
rect 18248 7041 18276 8230
rect 18340 7857 18368 9318
rect 18326 7848 18382 7857
rect 18326 7783 18382 7792
rect 18234 7032 18290 7041
rect 18234 6967 18290 6976
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 17958 6488 18014 6497
rect 17958 6423 17960 6432
rect 18012 6423 18014 6432
rect 17960 6394 18012 6400
rect 17868 6384 17920 6390
rect 17868 6326 17920 6332
rect 17880 5778 17908 6326
rect 18156 6089 18184 6598
rect 18236 6112 18288 6118
rect 18142 6080 18198 6089
rect 18236 6054 18288 6060
rect 18142 6015 18198 6024
rect 18052 5840 18104 5846
rect 18052 5782 18104 5788
rect 17868 5772 17920 5778
rect 17868 5714 17920 5720
rect 17788 5630 18000 5658
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 17788 4146 17816 5510
rect 17880 4865 17908 5510
rect 17866 4856 17922 4865
rect 17972 4826 18000 5630
rect 18064 5166 18092 5782
rect 18248 5681 18276 6054
rect 18234 5672 18290 5681
rect 18234 5607 18290 5616
rect 18432 5273 18460 9862
rect 18524 6254 18552 10542
rect 18602 9480 18658 9489
rect 18602 9415 18658 9424
rect 18616 9110 18644 9415
rect 18604 9104 18656 9110
rect 18604 9046 18656 9052
rect 18512 6248 18564 6254
rect 18512 6190 18564 6196
rect 18616 5914 18644 9046
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18418 5264 18474 5273
rect 18418 5199 18474 5208
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 17866 4791 17922 4800
rect 17960 4820 18012 4826
rect 17960 4762 18012 4768
rect 17868 4480 17920 4486
rect 18248 4457 18276 4966
rect 17868 4422 17920 4428
rect 18234 4448 18290 4457
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 17880 4049 17908 4422
rect 18234 4383 18290 4392
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 17866 4040 17922 4049
rect 17866 3975 17922 3984
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 18064 3097 18092 3334
rect 18050 3088 18106 3097
rect 18050 3023 18106 3032
rect 17868 2848 17920 2854
rect 17868 2790 17920 2796
rect 17880 2446 17908 2790
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 17868 2304 17920 2310
rect 17868 2246 17920 2252
rect 17880 1057 17908 2246
rect 18144 1964 18196 1970
rect 18144 1906 18196 1912
rect 17866 1048 17922 1057
rect 17866 983 17922 992
rect 18156 800 18184 1906
rect 17682 640 17738 649
rect 17682 575 17738 584
rect 18142 0 18198 800
rect 18248 241 18276 3878
rect 18524 1306 18552 4082
rect 18708 1465 18736 7686
rect 19616 4004 19668 4010
rect 19616 3946 19668 3952
rect 19156 1692 19208 1698
rect 19156 1634 19208 1640
rect 18694 1456 18750 1465
rect 18694 1391 18750 1400
rect 18524 1278 18644 1306
rect 18616 800 18644 1278
rect 19168 800 19196 1634
rect 19628 800 19656 3946
rect 18234 232 18290 241
rect 18234 167 18290 176
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19614 0 19670 800
<< via2 >>
rect 3422 16224 3478 16280
rect 2410 14184 2466 14240
rect 1582 13776 1638 13832
rect 1398 9968 1454 10024
rect 1398 8336 1454 8392
rect 1582 7928 1638 7984
rect 1398 5480 1454 5536
rect 938 992 994 1048
rect 3238 15816 3294 15872
rect 2962 11328 3018 11384
rect 2686 9560 2742 9616
rect 1766 7540 1822 7576
rect 1766 7520 1768 7540
rect 1768 7520 1820 7540
rect 1820 7520 1822 7540
rect 1858 5888 1914 5944
rect 2410 6296 2466 6352
rect 2870 10512 2926 10568
rect 3330 13368 3386 13424
rect 3606 16632 3662 16688
rect 10322 16224 10378 16280
rect 4066 15408 4122 15464
rect 3790 15000 3846 15056
rect 3514 12960 3570 13016
rect 3921 14170 3977 14172
rect 4001 14170 4057 14172
rect 4081 14170 4137 14172
rect 4161 14170 4217 14172
rect 3921 14118 3947 14170
rect 3947 14118 3977 14170
rect 4001 14118 4011 14170
rect 4011 14118 4057 14170
rect 4081 14118 4127 14170
rect 4127 14118 4137 14170
rect 4161 14118 4191 14170
rect 4191 14118 4217 14170
rect 3921 14116 3977 14118
rect 4001 14116 4057 14118
rect 4081 14116 4137 14118
rect 4161 14116 4217 14118
rect 3921 13082 3977 13084
rect 4001 13082 4057 13084
rect 4081 13082 4137 13084
rect 4161 13082 4217 13084
rect 3921 13030 3947 13082
rect 3947 13030 3977 13082
rect 4001 13030 4011 13082
rect 4011 13030 4057 13082
rect 4081 13030 4127 13082
rect 4127 13030 4137 13082
rect 4161 13030 4191 13082
rect 4191 13030 4217 13082
rect 3921 13028 3977 13030
rect 4001 13028 4057 13030
rect 4081 13028 4137 13030
rect 4161 13028 4217 13030
rect 4066 12588 4068 12608
rect 4068 12588 4120 12608
rect 4120 12588 4122 12608
rect 4066 12552 4122 12588
rect 3790 12144 3846 12200
rect 3921 11994 3977 11996
rect 4001 11994 4057 11996
rect 4081 11994 4137 11996
rect 4161 11994 4217 11996
rect 3921 11942 3947 11994
rect 3947 11942 3977 11994
rect 4001 11942 4011 11994
rect 4011 11942 4057 11994
rect 4081 11942 4127 11994
rect 4127 11942 4137 11994
rect 4161 11942 4191 11994
rect 4191 11942 4217 11994
rect 3921 11940 3977 11942
rect 4001 11940 4057 11942
rect 4081 11940 4137 11942
rect 4161 11940 4217 11942
rect 3790 11736 3846 11792
rect 3606 10920 3662 10976
rect 3514 9696 3570 9752
rect 3238 9560 3294 9616
rect 2870 7384 2926 7440
rect 2962 6724 3018 6760
rect 2962 6704 2964 6724
rect 2964 6704 3016 6724
rect 3016 6704 3018 6724
rect 1582 5072 1638 5128
rect 2410 4664 2466 4720
rect 1858 4256 1914 4312
rect 2502 3884 2504 3904
rect 2504 3884 2556 3904
rect 2556 3884 2558 3904
rect 2502 3848 2558 3884
rect 1858 3460 1914 3496
rect 1858 3440 1860 3460
rect 1860 3440 1912 3460
rect 1912 3440 1914 3460
rect 1858 2624 1914 2680
rect 2410 3068 2412 3088
rect 2412 3068 2464 3088
rect 2464 3068 2466 3088
rect 2410 3032 2466 3068
rect 2962 2216 3018 2272
rect 2778 1400 2834 1456
rect 1214 584 1270 640
rect 3514 9016 3570 9072
rect 3606 8880 3662 8936
rect 3514 7112 3570 7168
rect 3514 6704 3570 6760
rect 3921 10906 3977 10908
rect 4001 10906 4057 10908
rect 4081 10906 4137 10908
rect 4161 10906 4217 10908
rect 3921 10854 3947 10906
rect 3947 10854 3977 10906
rect 4001 10854 4011 10906
rect 4011 10854 4057 10906
rect 4081 10854 4127 10906
rect 4127 10854 4137 10906
rect 4161 10854 4191 10906
rect 4191 10854 4217 10906
rect 3921 10852 3977 10854
rect 4001 10852 4057 10854
rect 4081 10852 4137 10854
rect 4161 10852 4217 10854
rect 6886 14714 6942 14716
rect 6966 14714 7022 14716
rect 7046 14714 7102 14716
rect 7126 14714 7182 14716
rect 6886 14662 6912 14714
rect 6912 14662 6942 14714
rect 6966 14662 6976 14714
rect 6976 14662 7022 14714
rect 7046 14662 7092 14714
rect 7092 14662 7102 14714
rect 7126 14662 7156 14714
rect 7156 14662 7182 14714
rect 6886 14660 6942 14662
rect 6966 14660 7022 14662
rect 7046 14660 7102 14662
rect 7126 14660 7182 14662
rect 4066 10124 4122 10160
rect 4066 10104 4068 10124
rect 4068 10104 4120 10124
rect 4120 10104 4122 10124
rect 3921 9818 3977 9820
rect 4001 9818 4057 9820
rect 4081 9818 4137 9820
rect 4161 9818 4217 9820
rect 3921 9766 3947 9818
rect 3947 9766 3977 9818
rect 4001 9766 4011 9818
rect 4011 9766 4057 9818
rect 4081 9766 4127 9818
rect 4127 9766 4137 9818
rect 4161 9766 4191 9818
rect 4191 9766 4217 9818
rect 3921 9764 3977 9766
rect 4001 9764 4057 9766
rect 4081 9764 4137 9766
rect 4161 9764 4217 9766
rect 4434 9696 4490 9752
rect 3698 7792 3754 7848
rect 4526 9424 4582 9480
rect 3921 8730 3977 8732
rect 4001 8730 4057 8732
rect 4081 8730 4137 8732
rect 4161 8730 4217 8732
rect 3921 8678 3947 8730
rect 3947 8678 3977 8730
rect 4001 8678 4011 8730
rect 4011 8678 4057 8730
rect 4081 8678 4127 8730
rect 4127 8678 4137 8730
rect 4161 8678 4191 8730
rect 4191 8678 4217 8730
rect 3921 8676 3977 8678
rect 4001 8676 4057 8678
rect 4081 8676 4137 8678
rect 4161 8676 4217 8678
rect 3921 7642 3977 7644
rect 4001 7642 4057 7644
rect 4081 7642 4137 7644
rect 4161 7642 4217 7644
rect 3921 7590 3947 7642
rect 3947 7590 3977 7642
rect 4001 7590 4011 7642
rect 4011 7590 4057 7642
rect 4081 7590 4127 7642
rect 4127 7590 4137 7642
rect 4161 7590 4191 7642
rect 4191 7590 4217 7642
rect 3921 7588 3977 7590
rect 4001 7588 4057 7590
rect 4081 7588 4137 7590
rect 4161 7588 4217 7590
rect 3921 6554 3977 6556
rect 4001 6554 4057 6556
rect 4081 6554 4137 6556
rect 4161 6554 4217 6556
rect 3921 6502 3947 6554
rect 3947 6502 3977 6554
rect 4001 6502 4011 6554
rect 4011 6502 4057 6554
rect 4081 6502 4127 6554
rect 4127 6502 4137 6554
rect 4161 6502 4191 6554
rect 4191 6502 4217 6554
rect 3921 6500 3977 6502
rect 4001 6500 4057 6502
rect 4081 6500 4137 6502
rect 4161 6500 4217 6502
rect 3921 5466 3977 5468
rect 4001 5466 4057 5468
rect 4081 5466 4137 5468
rect 4161 5466 4217 5468
rect 3921 5414 3947 5466
rect 3947 5414 3977 5466
rect 4001 5414 4011 5466
rect 4011 5414 4057 5466
rect 4081 5414 4127 5466
rect 4127 5414 4137 5466
rect 4161 5414 4191 5466
rect 4191 5414 4217 5466
rect 3921 5412 3977 5414
rect 4001 5412 4057 5414
rect 4081 5412 4137 5414
rect 4161 5412 4217 5414
rect 3921 4378 3977 4380
rect 4001 4378 4057 4380
rect 4081 4378 4137 4380
rect 4161 4378 4217 4380
rect 3921 4326 3947 4378
rect 3947 4326 3977 4378
rect 4001 4326 4011 4378
rect 4011 4326 4057 4378
rect 4081 4326 4127 4378
rect 4127 4326 4137 4378
rect 4161 4326 4191 4378
rect 4191 4326 4217 4378
rect 3921 4324 3977 4326
rect 4001 4324 4057 4326
rect 4081 4324 4137 4326
rect 4161 4324 4217 4326
rect 3921 3290 3977 3292
rect 4001 3290 4057 3292
rect 4081 3290 4137 3292
rect 4161 3290 4217 3292
rect 3921 3238 3947 3290
rect 3947 3238 3977 3290
rect 4001 3238 4011 3290
rect 4011 3238 4057 3290
rect 4081 3238 4127 3290
rect 4127 3238 4137 3290
rect 4161 3238 4191 3290
rect 4191 3238 4217 3290
rect 3921 3236 3977 3238
rect 4001 3236 4057 3238
rect 4081 3236 4137 3238
rect 4161 3236 4217 3238
rect 3330 1808 3386 1864
rect 3921 2202 3977 2204
rect 4001 2202 4057 2204
rect 4081 2202 4137 2204
rect 4161 2202 4217 2204
rect 3921 2150 3947 2202
rect 3947 2150 3977 2202
rect 4001 2150 4011 2202
rect 4011 2150 4057 2202
rect 4081 2150 4127 2202
rect 4127 2150 4137 2202
rect 4161 2150 4191 2202
rect 4191 2150 4217 2202
rect 3921 2148 3977 2150
rect 4001 2148 4057 2150
rect 4081 2148 4137 2150
rect 4161 2148 4217 2150
rect 4526 6704 4582 6760
rect 4710 9424 4766 9480
rect 5262 9696 5318 9752
rect 5078 8880 5134 8936
rect 6182 9324 6184 9344
rect 6184 9324 6236 9344
rect 6236 9324 6238 9344
rect 6182 9288 6238 9324
rect 6090 8372 6092 8392
rect 6092 8372 6144 8392
rect 6144 8372 6146 8392
rect 6090 8336 6146 8372
rect 6886 13626 6942 13628
rect 6966 13626 7022 13628
rect 7046 13626 7102 13628
rect 7126 13626 7182 13628
rect 6886 13574 6912 13626
rect 6912 13574 6942 13626
rect 6966 13574 6976 13626
rect 6976 13574 7022 13626
rect 7046 13574 7092 13626
rect 7092 13574 7102 13626
rect 7126 13574 7156 13626
rect 7156 13574 7182 13626
rect 6886 13572 6942 13574
rect 6966 13572 7022 13574
rect 7046 13572 7102 13574
rect 7126 13572 7182 13574
rect 6886 12538 6942 12540
rect 6966 12538 7022 12540
rect 7046 12538 7102 12540
rect 7126 12538 7182 12540
rect 6886 12486 6912 12538
rect 6912 12486 6942 12538
rect 6966 12486 6976 12538
rect 6976 12486 7022 12538
rect 7046 12486 7092 12538
rect 7092 12486 7102 12538
rect 7126 12486 7156 12538
rect 7156 12486 7182 12538
rect 6886 12484 6942 12486
rect 6966 12484 7022 12486
rect 7046 12484 7102 12486
rect 7126 12484 7182 12486
rect 6886 11450 6942 11452
rect 6966 11450 7022 11452
rect 7046 11450 7102 11452
rect 7126 11450 7182 11452
rect 6886 11398 6912 11450
rect 6912 11398 6942 11450
rect 6966 11398 6976 11450
rect 6976 11398 7022 11450
rect 7046 11398 7092 11450
rect 7092 11398 7102 11450
rect 7126 11398 7156 11450
rect 7156 11398 7182 11450
rect 6886 11396 6942 11398
rect 6966 11396 7022 11398
rect 7046 11396 7102 11398
rect 7126 11396 7182 11398
rect 6886 10362 6942 10364
rect 6966 10362 7022 10364
rect 7046 10362 7102 10364
rect 7126 10362 7182 10364
rect 6886 10310 6912 10362
rect 6912 10310 6942 10362
rect 6966 10310 6976 10362
rect 6976 10310 7022 10362
rect 7046 10310 7092 10362
rect 7092 10310 7102 10362
rect 7126 10310 7156 10362
rect 7156 10310 7182 10362
rect 6886 10308 6942 10310
rect 6966 10308 7022 10310
rect 7046 10308 7102 10310
rect 7126 10308 7182 10310
rect 6886 9274 6942 9276
rect 6966 9274 7022 9276
rect 7046 9274 7102 9276
rect 7126 9274 7182 9276
rect 6886 9222 6912 9274
rect 6912 9222 6942 9274
rect 6966 9222 6976 9274
rect 6976 9222 7022 9274
rect 7046 9222 7092 9274
rect 7092 9222 7102 9274
rect 7126 9222 7156 9274
rect 7156 9222 7182 9274
rect 6886 9220 6942 9222
rect 6966 9220 7022 9222
rect 7046 9220 7102 9222
rect 7126 9220 7182 9222
rect 6886 8186 6942 8188
rect 6966 8186 7022 8188
rect 7046 8186 7102 8188
rect 7126 8186 7182 8188
rect 6886 8134 6912 8186
rect 6912 8134 6942 8186
rect 6966 8134 6976 8186
rect 6976 8134 7022 8186
rect 7046 8134 7092 8186
rect 7092 8134 7102 8186
rect 7126 8134 7156 8186
rect 7156 8134 7182 8186
rect 6886 8132 6942 8134
rect 6966 8132 7022 8134
rect 7046 8132 7102 8134
rect 7126 8132 7182 8134
rect 7562 9968 7618 10024
rect 7286 7928 7342 7984
rect 6886 7098 6942 7100
rect 6966 7098 7022 7100
rect 7046 7098 7102 7100
rect 7126 7098 7182 7100
rect 6886 7046 6912 7098
rect 6912 7046 6942 7098
rect 6966 7046 6976 7098
rect 6976 7046 7022 7098
rect 7046 7046 7092 7098
rect 7092 7046 7102 7098
rect 7126 7046 7156 7098
rect 7156 7046 7182 7098
rect 6886 7044 6942 7046
rect 6966 7044 7022 7046
rect 7046 7044 7102 7046
rect 7126 7044 7182 7046
rect 6886 6010 6942 6012
rect 6966 6010 7022 6012
rect 7046 6010 7102 6012
rect 7126 6010 7182 6012
rect 6886 5958 6912 6010
rect 6912 5958 6942 6010
rect 6966 5958 6976 6010
rect 6976 5958 7022 6010
rect 7046 5958 7092 6010
rect 7092 5958 7102 6010
rect 7126 5958 7156 6010
rect 7156 5958 7182 6010
rect 6886 5956 6942 5958
rect 6966 5956 7022 5958
rect 7046 5956 7102 5958
rect 7126 5956 7182 5958
rect 6886 4922 6942 4924
rect 6966 4922 7022 4924
rect 7046 4922 7102 4924
rect 7126 4922 7182 4924
rect 6886 4870 6912 4922
rect 6912 4870 6942 4922
rect 6966 4870 6976 4922
rect 6976 4870 7022 4922
rect 7046 4870 7092 4922
rect 7092 4870 7102 4922
rect 7126 4870 7156 4922
rect 7156 4870 7182 4922
rect 6886 4868 6942 4870
rect 6966 4868 7022 4870
rect 7046 4868 7102 4870
rect 7126 4868 7182 4870
rect 6886 3834 6942 3836
rect 6966 3834 7022 3836
rect 7046 3834 7102 3836
rect 7126 3834 7182 3836
rect 6886 3782 6912 3834
rect 6912 3782 6942 3834
rect 6966 3782 6976 3834
rect 6976 3782 7022 3834
rect 7046 3782 7092 3834
rect 7092 3782 7102 3834
rect 7126 3782 7156 3834
rect 7156 3782 7182 3834
rect 6886 3780 6942 3782
rect 6966 3780 7022 3782
rect 7046 3780 7102 3782
rect 7126 3780 7182 3782
rect 6886 2746 6942 2748
rect 6966 2746 7022 2748
rect 7046 2746 7102 2748
rect 7126 2746 7182 2748
rect 6886 2694 6912 2746
rect 6912 2694 6942 2746
rect 6966 2694 6976 2746
rect 6976 2694 7022 2746
rect 7046 2694 7092 2746
rect 7092 2694 7102 2746
rect 7126 2694 7156 2746
rect 7156 2694 7182 2746
rect 6886 2692 6942 2694
rect 6966 2692 7022 2694
rect 7046 2692 7102 2694
rect 7126 2692 7182 2694
rect 8574 9696 8630 9752
rect 8574 8356 8630 8392
rect 8574 8336 8576 8356
rect 8576 8336 8628 8356
rect 8628 8336 8630 8356
rect 8850 9288 8906 9344
rect 8758 7248 8814 7304
rect 9126 9424 9182 9480
rect 9034 9052 9036 9072
rect 9036 9052 9088 9072
rect 9088 9052 9090 9072
rect 9034 9016 9090 9052
rect 9034 8916 9036 8936
rect 9036 8916 9088 8936
rect 9088 8916 9090 8936
rect 9034 8880 9090 8916
rect 9034 7384 9090 7440
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9878 14170
rect 9878 14118 9908 14170
rect 9932 14118 9942 14170
rect 9942 14118 9988 14170
rect 10012 14118 10058 14170
rect 10058 14118 10068 14170
rect 10092 14118 10122 14170
rect 10122 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9878 13082
rect 9878 13030 9908 13082
rect 9932 13030 9942 13082
rect 9942 13030 9988 13082
rect 10012 13030 10058 13082
rect 10058 13030 10068 13082
rect 10092 13030 10122 13082
rect 10122 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9878 11994
rect 9878 11942 9908 11994
rect 9932 11942 9942 11994
rect 9942 11942 9988 11994
rect 10012 11942 10058 11994
rect 10058 11942 10068 11994
rect 10092 11942 10122 11994
rect 10122 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 16302 16632 16358 16688
rect 9586 10648 9642 10704
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9878 10906
rect 9878 10854 9908 10906
rect 9932 10854 9942 10906
rect 9942 10854 9988 10906
rect 10012 10854 10058 10906
rect 10058 10854 10068 10906
rect 10092 10854 10122 10906
rect 10122 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 10046 10260 10102 10296
rect 10046 10240 10048 10260
rect 10048 10240 10100 10260
rect 10100 10240 10102 10260
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9878 9818
rect 9878 9766 9908 9818
rect 9932 9766 9942 9818
rect 9942 9766 9988 9818
rect 10012 9766 10058 9818
rect 10058 9766 10068 9818
rect 10092 9766 10122 9818
rect 10122 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 9586 9560 9642 9616
rect 9494 9152 9550 9208
rect 10598 9968 10654 10024
rect 9586 8900 9642 8936
rect 9586 8880 9588 8900
rect 9588 8880 9640 8900
rect 9640 8880 9642 8900
rect 10598 8744 10654 8800
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9878 8730
rect 9878 8678 9908 8730
rect 9932 8678 9942 8730
rect 9942 8678 9988 8730
rect 10012 8678 10058 8730
rect 10058 8678 10068 8730
rect 10092 8678 10122 8730
rect 10122 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 10414 8356 10470 8392
rect 10414 8336 10416 8356
rect 10416 8336 10468 8356
rect 10468 8336 10470 8356
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9878 7642
rect 9878 7590 9908 7642
rect 9932 7590 9942 7642
rect 9942 7590 9988 7642
rect 10012 7590 10058 7642
rect 10058 7590 10068 7642
rect 10092 7590 10122 7642
rect 10122 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9878 6554
rect 9878 6502 9908 6554
rect 9932 6502 9942 6554
rect 9942 6502 9988 6554
rect 10012 6502 10058 6554
rect 10058 6502 10068 6554
rect 10092 6502 10122 6554
rect 10122 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 10322 6704 10378 6760
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9878 5466
rect 9878 5414 9908 5466
rect 9932 5414 9942 5466
rect 9942 5414 9988 5466
rect 10012 5414 10058 5466
rect 10058 5414 10068 5466
rect 10092 5414 10122 5466
rect 10122 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9878 4378
rect 9878 4326 9908 4378
rect 9932 4326 9942 4378
rect 9942 4326 9988 4378
rect 10012 4326 10058 4378
rect 10058 4326 10068 4378
rect 10092 4326 10122 4378
rect 10122 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9878 3290
rect 9878 3238 9908 3290
rect 9932 3238 9942 3290
rect 9942 3238 9988 3290
rect 10012 3238 10058 3290
rect 10058 3238 10068 3290
rect 10092 3238 10122 3290
rect 10122 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9878 2202
rect 9878 2150 9908 2202
rect 9932 2150 9942 2202
rect 9942 2150 9988 2202
rect 10012 2150 10058 2202
rect 10058 2150 10068 2202
rect 10092 2150 10122 2202
rect 10122 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 10874 9460 10876 9480
rect 10876 9460 10928 9480
rect 10928 9460 10930 9480
rect 10874 9424 10930 9460
rect 11058 9832 11114 9888
rect 11426 10684 11428 10704
rect 11428 10684 11480 10704
rect 11480 10684 11482 10704
rect 11426 10648 11482 10684
rect 11518 10240 11574 10296
rect 11610 9832 11666 9888
rect 11518 9560 11574 9616
rect 11058 8472 11114 8528
rect 11150 6840 11206 6896
rect 11242 5616 11298 5672
rect 11978 9152 12034 9208
rect 11886 7520 11942 7576
rect 11794 4020 11796 4040
rect 11796 4020 11848 4040
rect 11848 4020 11850 4040
rect 11794 3984 11850 4020
rect 12817 14714 12873 14716
rect 12897 14714 12953 14716
rect 12977 14714 13033 14716
rect 13057 14714 13113 14716
rect 12817 14662 12843 14714
rect 12843 14662 12873 14714
rect 12897 14662 12907 14714
rect 12907 14662 12953 14714
rect 12977 14662 13023 14714
rect 13023 14662 13033 14714
rect 13057 14662 13087 14714
rect 13087 14662 13113 14714
rect 12817 14660 12873 14662
rect 12897 14660 12953 14662
rect 12977 14660 13033 14662
rect 13057 14660 13113 14662
rect 12817 13626 12873 13628
rect 12897 13626 12953 13628
rect 12977 13626 13033 13628
rect 13057 13626 13113 13628
rect 12817 13574 12843 13626
rect 12843 13574 12873 13626
rect 12897 13574 12907 13626
rect 12907 13574 12953 13626
rect 12977 13574 13023 13626
rect 13023 13574 13033 13626
rect 13057 13574 13087 13626
rect 13087 13574 13113 13626
rect 12817 13572 12873 13574
rect 12897 13572 12953 13574
rect 12977 13572 13033 13574
rect 13057 13572 13113 13574
rect 12817 12538 12873 12540
rect 12897 12538 12953 12540
rect 12977 12538 13033 12540
rect 13057 12538 13113 12540
rect 12817 12486 12843 12538
rect 12843 12486 12873 12538
rect 12897 12486 12907 12538
rect 12907 12486 12953 12538
rect 12977 12486 13023 12538
rect 13023 12486 13033 12538
rect 13057 12486 13087 12538
rect 13087 12486 13113 12538
rect 12817 12484 12873 12486
rect 12897 12484 12953 12486
rect 12977 12484 13033 12486
rect 13057 12484 13113 12486
rect 13450 11736 13506 11792
rect 12817 11450 12873 11452
rect 12897 11450 12953 11452
rect 12977 11450 13033 11452
rect 13057 11450 13113 11452
rect 12817 11398 12843 11450
rect 12843 11398 12873 11450
rect 12897 11398 12907 11450
rect 12907 11398 12953 11450
rect 12977 11398 13023 11450
rect 13023 11398 13033 11450
rect 13057 11398 13087 11450
rect 13087 11398 13113 11450
rect 12817 11396 12873 11398
rect 12897 11396 12953 11398
rect 12977 11396 13033 11398
rect 13057 11396 13113 11398
rect 12162 10512 12218 10568
rect 12346 9016 12402 9072
rect 12346 7520 12402 7576
rect 12254 5772 12310 5808
rect 12254 5752 12256 5772
rect 12256 5752 12308 5772
rect 12308 5752 12310 5772
rect 12254 3068 12256 3088
rect 12256 3068 12308 3088
rect 12308 3068 12310 3088
rect 12254 3032 12310 3068
rect 12817 10362 12873 10364
rect 12897 10362 12953 10364
rect 12977 10362 13033 10364
rect 13057 10362 13113 10364
rect 12817 10310 12843 10362
rect 12843 10310 12873 10362
rect 12897 10310 12907 10362
rect 12907 10310 12953 10362
rect 12977 10310 13023 10362
rect 13023 10310 13033 10362
rect 13057 10310 13087 10362
rect 13087 10310 13113 10362
rect 12817 10308 12873 10310
rect 12897 10308 12953 10310
rect 12977 10308 13033 10310
rect 13057 10308 13113 10310
rect 12806 9444 12862 9480
rect 12806 9424 12808 9444
rect 12808 9424 12860 9444
rect 12860 9424 12862 9444
rect 12817 9274 12873 9276
rect 12897 9274 12953 9276
rect 12977 9274 13033 9276
rect 13057 9274 13113 9276
rect 12817 9222 12843 9274
rect 12843 9222 12873 9274
rect 12897 9222 12907 9274
rect 12907 9222 12953 9274
rect 12977 9222 13023 9274
rect 13023 9222 13033 9274
rect 13057 9222 13087 9274
rect 13087 9222 13113 9274
rect 12817 9220 12873 9222
rect 12897 9220 12953 9222
rect 12977 9220 13033 9222
rect 13057 9220 13113 9222
rect 12990 9036 13046 9072
rect 12990 9016 12992 9036
rect 12992 9016 13044 9036
rect 13044 9016 13046 9036
rect 13082 8744 13138 8800
rect 12622 7792 12678 7848
rect 12817 8186 12873 8188
rect 12897 8186 12953 8188
rect 12977 8186 13033 8188
rect 13057 8186 13113 8188
rect 12817 8134 12843 8186
rect 12843 8134 12873 8186
rect 12897 8134 12907 8186
rect 12907 8134 12953 8186
rect 12977 8134 13023 8186
rect 13023 8134 13033 8186
rect 13057 8134 13087 8186
rect 13087 8134 13113 8186
rect 12817 8132 12873 8134
rect 12897 8132 12953 8134
rect 12977 8132 13033 8134
rect 13057 8132 13113 8134
rect 15566 15816 15622 15872
rect 15198 15408 15254 15464
rect 12817 7098 12873 7100
rect 12897 7098 12953 7100
rect 12977 7098 13033 7100
rect 13057 7098 13113 7100
rect 12817 7046 12843 7098
rect 12843 7046 12873 7098
rect 12897 7046 12907 7098
rect 12907 7046 12953 7098
rect 12977 7046 13023 7098
rect 13023 7046 13033 7098
rect 13057 7046 13087 7098
rect 13087 7046 13113 7098
rect 12817 7044 12873 7046
rect 12897 7044 12953 7046
rect 12977 7044 13033 7046
rect 13057 7044 13113 7046
rect 13726 8372 13728 8392
rect 13728 8372 13780 8392
rect 13780 8372 13782 8392
rect 13726 8336 13782 8372
rect 12714 6704 12770 6760
rect 12817 6010 12873 6012
rect 12897 6010 12953 6012
rect 12977 6010 13033 6012
rect 13057 6010 13113 6012
rect 12817 5958 12843 6010
rect 12843 5958 12873 6010
rect 12897 5958 12907 6010
rect 12907 5958 12953 6010
rect 12977 5958 13023 6010
rect 13023 5958 13033 6010
rect 13057 5958 13087 6010
rect 13087 5958 13113 6010
rect 12817 5956 12873 5958
rect 12897 5956 12953 5958
rect 12977 5956 13033 5958
rect 13057 5956 13113 5958
rect 12714 5752 12770 5808
rect 12817 4922 12873 4924
rect 12897 4922 12953 4924
rect 12977 4922 13033 4924
rect 13057 4922 13113 4924
rect 12817 4870 12843 4922
rect 12843 4870 12873 4922
rect 12897 4870 12907 4922
rect 12907 4870 12953 4922
rect 12977 4870 13023 4922
rect 13023 4870 13033 4922
rect 13057 4870 13087 4922
rect 13087 4870 13113 4922
rect 12817 4868 12873 4870
rect 12897 4868 12953 4870
rect 12977 4868 13033 4870
rect 13057 4868 13113 4870
rect 12530 3068 12532 3088
rect 12532 3068 12584 3088
rect 12584 3068 12586 3088
rect 12530 3032 12586 3068
rect 12817 3834 12873 3836
rect 12897 3834 12953 3836
rect 12977 3834 13033 3836
rect 13057 3834 13113 3836
rect 12817 3782 12843 3834
rect 12843 3782 12873 3834
rect 12897 3782 12907 3834
rect 12907 3782 12953 3834
rect 12977 3782 13023 3834
rect 13023 3782 13033 3834
rect 13057 3782 13087 3834
rect 13087 3782 13113 3834
rect 12817 3780 12873 3782
rect 12897 3780 12953 3782
rect 12977 3780 13033 3782
rect 13057 3780 13113 3782
rect 12817 2746 12873 2748
rect 12897 2746 12953 2748
rect 12977 2746 13033 2748
rect 13057 2746 13113 2748
rect 12817 2694 12843 2746
rect 12843 2694 12873 2746
rect 12897 2694 12907 2746
rect 12907 2694 12953 2746
rect 12977 2694 13023 2746
rect 13023 2694 13033 2746
rect 13057 2694 13087 2746
rect 13087 2694 13113 2746
rect 12817 2692 12873 2694
rect 12897 2692 12953 2694
rect 12977 2692 13033 2694
rect 13057 2692 13113 2694
rect 13726 4972 13728 4992
rect 13728 4972 13780 4992
rect 13780 4972 13782 4992
rect 13726 4936 13782 4972
rect 14738 7792 14794 7848
rect 15290 15000 15346 15056
rect 15290 13776 15346 13832
rect 15290 13368 15346 13424
rect 15474 13776 15530 13832
rect 16118 14592 16174 14648
rect 15782 14170 15838 14172
rect 15862 14170 15918 14172
rect 15942 14170 15998 14172
rect 16022 14170 16078 14172
rect 15782 14118 15808 14170
rect 15808 14118 15838 14170
rect 15862 14118 15872 14170
rect 15872 14118 15918 14170
rect 15942 14118 15988 14170
rect 15988 14118 15998 14170
rect 16022 14118 16052 14170
rect 16052 14118 16078 14170
rect 15782 14116 15838 14118
rect 15862 14116 15918 14118
rect 15942 14116 15998 14118
rect 16022 14116 16078 14118
rect 15782 13082 15838 13084
rect 15862 13082 15918 13084
rect 15942 13082 15998 13084
rect 16022 13082 16078 13084
rect 15782 13030 15808 13082
rect 15808 13030 15838 13082
rect 15862 13030 15872 13082
rect 15872 13030 15918 13082
rect 15942 13030 15988 13082
rect 15988 13030 15998 13082
rect 16022 13030 16052 13082
rect 16052 13030 16078 13082
rect 15782 13028 15838 13030
rect 15862 13028 15918 13030
rect 15942 13028 15998 13030
rect 16022 13028 16078 13030
rect 15658 12416 15714 12472
rect 15382 10648 15438 10704
rect 15782 11994 15838 11996
rect 15862 11994 15918 11996
rect 15942 11994 15998 11996
rect 16022 11994 16078 11996
rect 15782 11942 15808 11994
rect 15808 11942 15838 11994
rect 15862 11942 15872 11994
rect 15872 11942 15918 11994
rect 15942 11942 15988 11994
rect 15988 11942 15998 11994
rect 16022 11942 16052 11994
rect 16052 11942 16078 11994
rect 15782 11940 15838 11942
rect 15862 11940 15918 11942
rect 15942 11940 15998 11942
rect 16022 11940 16078 11942
rect 15782 10906 15838 10908
rect 15862 10906 15918 10908
rect 15942 10906 15998 10908
rect 16022 10906 16078 10908
rect 15782 10854 15808 10906
rect 15808 10854 15838 10906
rect 15862 10854 15872 10906
rect 15872 10854 15918 10906
rect 15942 10854 15988 10906
rect 15988 10854 15998 10906
rect 16022 10854 16052 10906
rect 16052 10854 16078 10906
rect 15782 10852 15838 10854
rect 15862 10852 15918 10854
rect 15942 10852 15998 10854
rect 16022 10852 16078 10854
rect 15382 10376 15438 10432
rect 15290 9424 15346 9480
rect 15658 10512 15714 10568
rect 15782 9818 15838 9820
rect 15862 9818 15918 9820
rect 15942 9818 15998 9820
rect 16022 9818 16078 9820
rect 15782 9766 15808 9818
rect 15808 9766 15838 9818
rect 15862 9766 15872 9818
rect 15872 9766 15918 9818
rect 15942 9766 15988 9818
rect 15988 9766 15998 9818
rect 16022 9766 16052 9818
rect 16052 9766 16078 9818
rect 15782 9764 15838 9766
rect 15862 9764 15918 9766
rect 15942 9764 15998 9766
rect 16022 9764 16078 9766
rect 15658 9560 15714 9616
rect 15782 8730 15838 8732
rect 15862 8730 15918 8732
rect 15942 8730 15998 8732
rect 16022 8730 16078 8732
rect 15782 8678 15808 8730
rect 15808 8678 15838 8730
rect 15862 8678 15872 8730
rect 15872 8678 15918 8730
rect 15942 8678 15988 8730
rect 15988 8678 15998 8730
rect 16022 8678 16052 8730
rect 16052 8678 16078 8730
rect 15782 8676 15838 8678
rect 15862 8676 15918 8678
rect 15942 8676 15998 8678
rect 16022 8676 16078 8678
rect 15782 7642 15838 7644
rect 15862 7642 15918 7644
rect 15942 7642 15998 7644
rect 16022 7642 16078 7644
rect 15782 7590 15808 7642
rect 15808 7590 15838 7642
rect 15862 7590 15872 7642
rect 15872 7590 15918 7642
rect 15942 7590 15988 7642
rect 15988 7590 15998 7642
rect 16022 7590 16052 7642
rect 16052 7590 16078 7642
rect 15782 7588 15838 7590
rect 15862 7588 15918 7590
rect 15942 7588 15998 7590
rect 16022 7588 16078 7590
rect 15782 6554 15838 6556
rect 15862 6554 15918 6556
rect 15942 6554 15998 6556
rect 16022 6554 16078 6556
rect 15782 6502 15808 6554
rect 15808 6502 15838 6554
rect 15862 6502 15872 6554
rect 15872 6502 15918 6554
rect 15942 6502 15988 6554
rect 15988 6502 15998 6554
rect 16022 6502 16052 6554
rect 16052 6502 16078 6554
rect 15782 6500 15838 6502
rect 15862 6500 15918 6502
rect 15942 6500 15998 6502
rect 16022 6500 16078 6502
rect 16026 5616 16082 5672
rect 15782 5466 15838 5468
rect 15862 5466 15918 5468
rect 15942 5466 15998 5468
rect 16022 5466 16078 5468
rect 15782 5414 15808 5466
rect 15808 5414 15838 5466
rect 15862 5414 15872 5466
rect 15872 5414 15918 5466
rect 15942 5414 15988 5466
rect 15988 5414 15998 5466
rect 16022 5414 16052 5466
rect 16052 5414 16078 5466
rect 15782 5412 15838 5414
rect 15862 5412 15918 5414
rect 15942 5412 15998 5414
rect 16022 5412 16078 5414
rect 16486 14184 16542 14240
rect 16302 12824 16358 12880
rect 17498 13232 17554 13288
rect 16578 11192 16634 11248
rect 16394 10920 16450 10976
rect 16670 10784 16726 10840
rect 16394 10104 16450 10160
rect 16670 10104 16726 10160
rect 16578 9968 16634 10024
rect 17130 9832 17186 9888
rect 15782 4378 15838 4380
rect 15862 4378 15918 4380
rect 15942 4378 15998 4380
rect 16022 4378 16078 4380
rect 15782 4326 15808 4378
rect 15808 4326 15838 4378
rect 15862 4326 15872 4378
rect 15872 4326 15918 4378
rect 15942 4326 15988 4378
rect 15988 4326 15998 4378
rect 16022 4326 16052 4378
rect 16052 4326 16078 4378
rect 15782 4324 15838 4326
rect 15862 4324 15918 4326
rect 15942 4324 15998 4326
rect 16022 4324 16078 4326
rect 15782 3290 15838 3292
rect 15862 3290 15918 3292
rect 15942 3290 15998 3292
rect 16022 3290 16078 3292
rect 15782 3238 15808 3290
rect 15808 3238 15838 3290
rect 15862 3238 15872 3290
rect 15872 3238 15918 3290
rect 15942 3238 15988 3290
rect 15988 3238 15998 3290
rect 16022 3238 16052 3290
rect 16052 3238 16078 3290
rect 15782 3236 15838 3238
rect 15862 3236 15918 3238
rect 15942 3236 15998 3238
rect 16022 3236 16078 3238
rect 15842 2488 15898 2544
rect 15782 2202 15838 2204
rect 15862 2202 15918 2204
rect 15942 2202 15998 2204
rect 16022 2202 16078 2204
rect 15782 2150 15808 2202
rect 15808 2150 15838 2202
rect 15862 2150 15872 2202
rect 15872 2150 15918 2202
rect 15942 2150 15988 2202
rect 15988 2150 15998 2202
rect 16022 2150 16052 2202
rect 16052 2150 16078 2202
rect 15782 2148 15838 2150
rect 15862 2148 15918 2150
rect 15942 2148 15998 2150
rect 16022 2148 16078 2150
rect 16486 6840 16542 6896
rect 16762 6976 16818 7032
rect 16578 4936 16634 4992
rect 16302 3984 16358 4040
rect 17130 9016 17186 9072
rect 17406 11192 17462 11248
rect 17774 11600 17830 11656
rect 17038 8608 17094 8664
rect 16946 7792 17002 7848
rect 17314 7928 17370 7984
rect 17590 8200 17646 8256
rect 17958 8472 18014 8528
rect 17958 7928 18014 7984
rect 18050 7384 18106 7440
rect 17590 3576 17646 3632
rect 17590 2624 17646 2680
rect 17314 2252 17316 2272
rect 17316 2252 17368 2272
rect 17368 2252 17370 2272
rect 17314 2216 17370 2252
rect 17590 1808 17646 1864
rect 3054 176 3110 232
rect 17958 7248 18014 7304
rect 18326 7792 18382 7848
rect 18234 6976 18290 7032
rect 17958 6452 18014 6488
rect 17958 6432 17960 6452
rect 17960 6432 18012 6452
rect 18012 6432 18014 6452
rect 18142 6024 18198 6080
rect 17866 4800 17922 4856
rect 18234 5616 18290 5672
rect 18602 9424 18658 9480
rect 18418 5208 18474 5264
rect 18234 4392 18290 4448
rect 17866 3984 17922 4040
rect 18050 3032 18106 3088
rect 17866 992 17922 1048
rect 17682 584 17738 640
rect 18694 1400 18750 1456
rect 18234 176 18290 232
<< metal3 >>
rect 0 16690 800 16720
rect 3601 16690 3667 16693
rect 0 16688 3667 16690
rect 0 16632 3606 16688
rect 3662 16632 3667 16688
rect 0 16630 3667 16632
rect 0 16600 800 16630
rect 3601 16627 3667 16630
rect 16297 16690 16363 16693
rect 19200 16690 20000 16720
rect 16297 16688 20000 16690
rect 16297 16632 16302 16688
rect 16358 16632 20000 16688
rect 16297 16630 20000 16632
rect 16297 16627 16363 16630
rect 19200 16600 20000 16630
rect 0 16282 800 16312
rect 3417 16282 3483 16285
rect 0 16280 3483 16282
rect 0 16224 3422 16280
rect 3478 16224 3483 16280
rect 0 16222 3483 16224
rect 0 16192 800 16222
rect 3417 16219 3483 16222
rect 10317 16282 10383 16285
rect 19200 16282 20000 16312
rect 10317 16280 20000 16282
rect 10317 16224 10322 16280
rect 10378 16224 20000 16280
rect 10317 16222 20000 16224
rect 10317 16219 10383 16222
rect 19200 16192 20000 16222
rect 0 15874 800 15904
rect 3233 15874 3299 15877
rect 0 15872 3299 15874
rect 0 15816 3238 15872
rect 3294 15816 3299 15872
rect 0 15814 3299 15816
rect 0 15784 800 15814
rect 3233 15811 3299 15814
rect 15561 15874 15627 15877
rect 19200 15874 20000 15904
rect 15561 15872 20000 15874
rect 15561 15816 15566 15872
rect 15622 15816 20000 15872
rect 15561 15814 20000 15816
rect 15561 15811 15627 15814
rect 19200 15784 20000 15814
rect 0 15466 800 15496
rect 4061 15466 4127 15469
rect 0 15464 4127 15466
rect 0 15408 4066 15464
rect 4122 15408 4127 15464
rect 0 15406 4127 15408
rect 0 15376 800 15406
rect 4061 15403 4127 15406
rect 15193 15466 15259 15469
rect 19200 15466 20000 15496
rect 15193 15464 20000 15466
rect 15193 15408 15198 15464
rect 15254 15408 20000 15464
rect 15193 15406 20000 15408
rect 15193 15403 15259 15406
rect 19200 15376 20000 15406
rect 0 15058 800 15088
rect 3785 15058 3851 15061
rect 0 15056 3851 15058
rect 0 15000 3790 15056
rect 3846 15000 3851 15056
rect 0 14998 3851 15000
rect 0 14968 800 14998
rect 3785 14995 3851 14998
rect 15285 15058 15351 15061
rect 19200 15058 20000 15088
rect 15285 15056 20000 15058
rect 15285 15000 15290 15056
rect 15346 15000 20000 15056
rect 15285 14998 20000 15000
rect 15285 14995 15351 14998
rect 19200 14968 20000 14998
rect 6874 14720 7194 14721
rect 0 14650 800 14680
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7194 14720
rect 6874 14655 7194 14656
rect 12805 14720 13125 14721
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 14655 13125 14656
rect 16113 14650 16179 14653
rect 19200 14650 20000 14680
rect 0 14590 6746 14650
rect 0 14560 800 14590
rect 6686 14514 6746 14590
rect 16113 14648 20000 14650
rect 16113 14592 16118 14648
rect 16174 14592 20000 14648
rect 16113 14590 20000 14592
rect 16113 14587 16179 14590
rect 19200 14560 20000 14590
rect 8518 14514 8524 14516
rect 6686 14454 8524 14514
rect 8518 14452 8524 14454
rect 8588 14452 8594 14516
rect 0 14242 800 14272
rect 2405 14242 2471 14245
rect 0 14240 2471 14242
rect 0 14184 2410 14240
rect 2466 14184 2471 14240
rect 0 14182 2471 14184
rect 0 14152 800 14182
rect 2405 14179 2471 14182
rect 16481 14242 16547 14245
rect 19200 14242 20000 14272
rect 16481 14240 20000 14242
rect 16481 14184 16486 14240
rect 16542 14184 20000 14240
rect 16481 14182 20000 14184
rect 16481 14179 16547 14182
rect 3909 14176 4229 14177
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 14111 4229 14112
rect 9840 14176 10160 14177
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 14111 10160 14112
rect 15770 14176 16090 14177
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 19200 14152 20000 14182
rect 15770 14111 16090 14112
rect 0 13834 800 13864
rect 1577 13834 1643 13837
rect 0 13832 1643 13834
rect 0 13776 1582 13832
rect 1638 13776 1643 13832
rect 0 13774 1643 13776
rect 0 13744 800 13774
rect 1577 13771 1643 13774
rect 15285 13834 15351 13837
rect 15469 13834 15535 13837
rect 19200 13834 20000 13864
rect 15285 13832 15394 13834
rect 15285 13776 15290 13832
rect 15346 13776 15394 13832
rect 15285 13771 15394 13776
rect 15469 13832 20000 13834
rect 15469 13776 15474 13832
rect 15530 13776 20000 13832
rect 15469 13774 20000 13776
rect 15469 13771 15535 13774
rect 6874 13632 7194 13633
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7194 13632
rect 6874 13567 7194 13568
rect 12805 13632 13125 13633
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 13567 13125 13568
rect 0 13426 800 13456
rect 15334 13429 15394 13771
rect 19200 13744 20000 13774
rect 3325 13426 3391 13429
rect 0 13424 3391 13426
rect 0 13368 3330 13424
rect 3386 13368 3391 13424
rect 0 13366 3391 13368
rect 0 13336 800 13366
rect 3325 13363 3391 13366
rect 15285 13424 15394 13429
rect 15285 13368 15290 13424
rect 15346 13368 15394 13424
rect 15285 13366 15394 13368
rect 15285 13363 15351 13366
rect 17493 13290 17559 13293
rect 19200 13290 20000 13320
rect 17493 13288 20000 13290
rect 17493 13232 17498 13288
rect 17554 13232 20000 13288
rect 17493 13230 20000 13232
rect 17493 13227 17559 13230
rect 19200 13200 20000 13230
rect 3909 13088 4229 13089
rect 0 13018 800 13048
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 13023 4229 13024
rect 9840 13088 10160 13089
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 13023 10160 13024
rect 15770 13088 16090 13089
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 15770 13023 16090 13024
rect 3509 13018 3575 13021
rect 0 13016 3575 13018
rect 0 12960 3514 13016
rect 3570 12960 3575 13016
rect 0 12958 3575 12960
rect 0 12928 800 12958
rect 3509 12955 3575 12958
rect 16297 12882 16363 12885
rect 19200 12882 20000 12912
rect 16297 12880 20000 12882
rect 16297 12824 16302 12880
rect 16358 12824 20000 12880
rect 16297 12822 20000 12824
rect 16297 12819 16363 12822
rect 19200 12792 20000 12822
rect 0 12610 800 12640
rect 4061 12610 4127 12613
rect 0 12608 4127 12610
rect 0 12552 4066 12608
rect 4122 12552 4127 12608
rect 0 12550 4127 12552
rect 0 12520 800 12550
rect 4061 12547 4127 12550
rect 6874 12544 7194 12545
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7194 12544
rect 6874 12479 7194 12480
rect 12805 12544 13125 12545
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 12479 13125 12480
rect 15653 12474 15719 12477
rect 19200 12474 20000 12504
rect 15653 12472 20000 12474
rect 15653 12416 15658 12472
rect 15714 12416 20000 12472
rect 15653 12414 20000 12416
rect 15653 12411 15719 12414
rect 19200 12384 20000 12414
rect 0 12202 800 12232
rect 3785 12202 3851 12205
rect 0 12200 3851 12202
rect 0 12144 3790 12200
rect 3846 12144 3851 12200
rect 0 12142 3851 12144
rect 0 12112 800 12142
rect 3785 12139 3851 12142
rect 19200 12066 20000 12096
rect 16254 12006 20000 12066
rect 3909 12000 4229 12001
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 11935 4229 11936
rect 9840 12000 10160 12001
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 11935 10160 11936
rect 15770 12000 16090 12001
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 15770 11935 16090 11936
rect 0 11794 800 11824
rect 3785 11794 3851 11797
rect 0 11792 3851 11794
rect 0 11736 3790 11792
rect 3846 11736 3851 11792
rect 0 11734 3851 11736
rect 0 11704 800 11734
rect 3785 11731 3851 11734
rect 13445 11794 13511 11797
rect 16254 11794 16314 12006
rect 19200 11976 20000 12006
rect 13445 11792 16314 11794
rect 13445 11736 13450 11792
rect 13506 11736 16314 11792
rect 13445 11734 16314 11736
rect 13445 11731 13511 11734
rect 17769 11658 17835 11661
rect 19200 11658 20000 11688
rect 17769 11656 20000 11658
rect 17769 11600 17774 11656
rect 17830 11600 20000 11656
rect 17769 11598 20000 11600
rect 17769 11595 17835 11598
rect 19200 11568 20000 11598
rect 6874 11456 7194 11457
rect 0 11386 800 11416
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7194 11456
rect 6874 11391 7194 11392
rect 12805 11456 13125 11457
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 11391 13125 11392
rect 2957 11386 3023 11389
rect 0 11384 3023 11386
rect 0 11328 2962 11384
rect 3018 11328 3023 11384
rect 0 11326 3023 11328
rect 0 11296 800 11326
rect 2957 11323 3023 11326
rect 16573 11250 16639 11253
rect 17401 11250 17467 11253
rect 19200 11250 20000 11280
rect 16573 11248 20000 11250
rect 16573 11192 16578 11248
rect 16634 11192 17406 11248
rect 17462 11192 20000 11248
rect 16573 11190 20000 11192
rect 16573 11187 16639 11190
rect 17401 11187 17467 11190
rect 19200 11160 20000 11190
rect 0 10978 800 11008
rect 3601 10978 3667 10981
rect 16389 10980 16455 10981
rect 16389 10978 16436 10980
rect 0 10976 3667 10978
rect 0 10920 3606 10976
rect 3662 10920 3667 10976
rect 0 10918 3667 10920
rect 16344 10976 16436 10978
rect 16344 10920 16394 10976
rect 16344 10918 16436 10920
rect 0 10888 800 10918
rect 3601 10915 3667 10918
rect 16389 10916 16436 10918
rect 16500 10916 16506 10980
rect 16389 10915 16455 10916
rect 3909 10912 4229 10913
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 10847 4229 10848
rect 9840 10912 10160 10913
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 10847 10160 10848
rect 15770 10912 16090 10913
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15770 10847 16090 10848
rect 16665 10842 16731 10845
rect 19200 10842 20000 10872
rect 16665 10840 20000 10842
rect 16665 10784 16670 10840
rect 16726 10784 20000 10840
rect 16665 10782 20000 10784
rect 16665 10779 16731 10782
rect 19200 10752 20000 10782
rect 9581 10706 9647 10709
rect 11421 10706 11487 10709
rect 15377 10708 15443 10709
rect 9581 10704 11487 10706
rect 9581 10648 9586 10704
rect 9642 10648 11426 10704
rect 11482 10648 11487 10704
rect 9581 10646 11487 10648
rect 9581 10643 9647 10646
rect 11421 10643 11487 10646
rect 15326 10644 15332 10708
rect 15396 10706 15443 10708
rect 15396 10704 15488 10706
rect 15438 10648 15488 10704
rect 15396 10646 15488 10648
rect 15396 10644 15443 10646
rect 15377 10643 15443 10644
rect 0 10570 800 10600
rect 2865 10570 2931 10573
rect 0 10568 2931 10570
rect 0 10512 2870 10568
rect 2926 10512 2931 10568
rect 0 10510 2931 10512
rect 0 10480 800 10510
rect 2865 10507 2931 10510
rect 12157 10570 12223 10573
rect 15653 10570 15719 10573
rect 12157 10568 15719 10570
rect 12157 10512 12162 10568
rect 12218 10512 15658 10568
rect 15714 10512 15719 10568
rect 12157 10510 15719 10512
rect 12157 10507 12223 10510
rect 15653 10507 15719 10510
rect 15377 10434 15443 10437
rect 19200 10434 20000 10464
rect 15377 10432 20000 10434
rect 15377 10376 15382 10432
rect 15438 10376 20000 10432
rect 15377 10374 20000 10376
rect 15377 10371 15443 10374
rect 6874 10368 7194 10369
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7194 10368
rect 6874 10303 7194 10304
rect 12805 10368 13125 10369
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 19200 10344 20000 10374
rect 12805 10303 13125 10304
rect 10041 10298 10107 10301
rect 11513 10298 11579 10301
rect 10041 10296 11579 10298
rect 10041 10240 10046 10296
rect 10102 10240 11518 10296
rect 11574 10240 11579 10296
rect 10041 10238 11579 10240
rect 10041 10235 10107 10238
rect 11513 10235 11579 10238
rect 0 10162 800 10192
rect 4061 10162 4127 10165
rect 0 10160 4127 10162
rect 0 10104 4066 10160
rect 4122 10104 4127 10160
rect 0 10102 4127 10104
rect 0 10072 800 10102
rect 4061 10099 4127 10102
rect 16389 10162 16455 10165
rect 16665 10162 16731 10165
rect 16389 10160 16731 10162
rect 16389 10104 16394 10160
rect 16450 10104 16670 10160
rect 16726 10104 16731 10160
rect 16389 10102 16731 10104
rect 16389 10099 16455 10102
rect 16665 10099 16731 10102
rect 1393 10026 1459 10029
rect 7557 10026 7623 10029
rect 1393 10024 7623 10026
rect 1393 9968 1398 10024
rect 1454 9968 7562 10024
rect 7618 9968 7623 10024
rect 1393 9966 7623 9968
rect 1393 9963 1459 9966
rect 7557 9963 7623 9966
rect 10593 10026 10659 10029
rect 16573 10026 16639 10029
rect 10593 10024 16639 10026
rect 10593 9968 10598 10024
rect 10654 9968 16578 10024
rect 16634 9968 16639 10024
rect 10593 9966 16639 9968
rect 10593 9963 10659 9966
rect 16573 9963 16639 9966
rect 11053 9890 11119 9893
rect 11605 9890 11671 9893
rect 11053 9888 11671 9890
rect 11053 9832 11058 9888
rect 11114 9832 11610 9888
rect 11666 9832 11671 9888
rect 11053 9830 11671 9832
rect 11053 9827 11119 9830
rect 11605 9827 11671 9830
rect 17125 9890 17191 9893
rect 19200 9890 20000 9920
rect 17125 9888 20000 9890
rect 17125 9832 17130 9888
rect 17186 9832 20000 9888
rect 17125 9830 20000 9832
rect 17125 9827 17191 9830
rect 3909 9824 4229 9825
rect 0 9754 800 9784
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 9759 4229 9760
rect 9840 9824 10160 9825
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 9759 10160 9760
rect 15770 9824 16090 9825
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 19200 9800 20000 9830
rect 15770 9759 16090 9760
rect 3509 9754 3575 9757
rect 0 9752 3575 9754
rect 0 9696 3514 9752
rect 3570 9696 3575 9752
rect 0 9694 3575 9696
rect 0 9664 800 9694
rect 3509 9691 3575 9694
rect 4429 9754 4495 9757
rect 5257 9754 5323 9757
rect 8569 9754 8635 9757
rect 4429 9752 8635 9754
rect 4429 9696 4434 9752
rect 4490 9696 5262 9752
rect 5318 9696 8574 9752
rect 8630 9696 8635 9752
rect 4429 9694 8635 9696
rect 4429 9691 4495 9694
rect 5257 9691 5323 9694
rect 8569 9691 8635 9694
rect 2681 9618 2747 9621
rect 3233 9618 3299 9621
rect 9581 9618 9647 9621
rect 2681 9616 9647 9618
rect 2681 9560 2686 9616
rect 2742 9560 3238 9616
rect 3294 9560 9586 9616
rect 9642 9560 9647 9616
rect 2681 9558 9647 9560
rect 2681 9555 2747 9558
rect 3233 9555 3299 9558
rect 9581 9555 9647 9558
rect 11513 9618 11579 9621
rect 15653 9618 15719 9621
rect 11513 9616 15719 9618
rect 11513 9560 11518 9616
rect 11574 9560 15658 9616
rect 15714 9560 15719 9616
rect 11513 9558 15719 9560
rect 11513 9555 11579 9558
rect 15653 9555 15719 9558
rect 4521 9482 4587 9485
rect 4705 9482 4771 9485
rect 9121 9482 9187 9485
rect 4521 9480 9187 9482
rect 4521 9424 4526 9480
rect 4582 9424 4710 9480
rect 4766 9424 9126 9480
rect 9182 9424 9187 9480
rect 4521 9422 9187 9424
rect 4521 9419 4587 9422
rect 4705 9419 4771 9422
rect 9121 9419 9187 9422
rect 10869 9482 10935 9485
rect 12801 9482 12867 9485
rect 10869 9480 12867 9482
rect 10869 9424 10874 9480
rect 10930 9424 12806 9480
rect 12862 9424 12867 9480
rect 10869 9422 12867 9424
rect 10869 9419 10935 9422
rect 12801 9419 12867 9422
rect 15285 9482 15351 9485
rect 15510 9482 15516 9484
rect 15285 9480 15516 9482
rect 15285 9424 15290 9480
rect 15346 9424 15516 9480
rect 15285 9422 15516 9424
rect 15285 9419 15351 9422
rect 15510 9420 15516 9422
rect 15580 9420 15586 9484
rect 18597 9482 18663 9485
rect 19200 9482 20000 9512
rect 18597 9480 20000 9482
rect 18597 9424 18602 9480
rect 18658 9424 20000 9480
rect 18597 9422 20000 9424
rect 18597 9419 18663 9422
rect 19200 9392 20000 9422
rect 0 9346 800 9376
rect 6177 9346 6243 9349
rect 0 9344 6243 9346
rect 0 9288 6182 9344
rect 6238 9288 6243 9344
rect 0 9286 6243 9288
rect 0 9256 800 9286
rect 6177 9283 6243 9286
rect 8518 9284 8524 9348
rect 8588 9346 8594 9348
rect 8845 9346 8911 9349
rect 8588 9344 8911 9346
rect 8588 9288 8850 9344
rect 8906 9288 8911 9344
rect 8588 9286 8911 9288
rect 8588 9284 8594 9286
rect 8845 9283 8911 9286
rect 6874 9280 7194 9281
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7194 9280
rect 6874 9215 7194 9216
rect 12805 9280 13125 9281
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 9215 13125 9216
rect 9489 9210 9555 9213
rect 7284 9208 9555 9210
rect 7284 9152 9494 9208
rect 9550 9152 9555 9208
rect 7284 9150 9555 9152
rect 3509 9074 3575 9077
rect 7284 9074 7344 9150
rect 9489 9147 9555 9150
rect 11973 9210 12039 9213
rect 11973 9208 12680 9210
rect 11973 9152 11978 9208
rect 12034 9152 12680 9208
rect 11973 9150 12680 9152
rect 11973 9147 12039 9150
rect 3509 9072 7344 9074
rect 3509 9016 3514 9072
rect 3570 9016 7344 9072
rect 3509 9014 7344 9016
rect 9029 9074 9095 9077
rect 12341 9074 12407 9077
rect 9029 9072 12407 9074
rect 9029 9016 9034 9072
rect 9090 9016 12346 9072
rect 12402 9016 12407 9072
rect 9029 9014 12407 9016
rect 12620 9074 12680 9150
rect 12985 9074 13051 9077
rect 12620 9072 13051 9074
rect 12620 9016 12990 9072
rect 13046 9016 13051 9072
rect 12620 9014 13051 9016
rect 3509 9011 3575 9014
rect 9029 9011 9095 9014
rect 12341 9011 12407 9014
rect 12985 9011 13051 9014
rect 17125 9074 17191 9077
rect 19200 9074 20000 9104
rect 17125 9072 20000 9074
rect 17125 9016 17130 9072
rect 17186 9016 20000 9072
rect 17125 9014 20000 9016
rect 17125 9011 17191 9014
rect 0 8938 800 8968
rect 3601 8938 3667 8941
rect 5073 8938 5139 8941
rect 9029 8938 9095 8941
rect 9581 8938 9647 8941
rect 0 8936 9647 8938
rect 0 8880 3606 8936
rect 3662 8880 5078 8936
rect 5134 8880 9034 8936
rect 9090 8880 9586 8936
rect 9642 8880 9647 8936
rect 0 8878 9647 8880
rect 12344 8938 12404 9011
rect 19200 8984 20000 9014
rect 12344 8878 16314 8938
rect 0 8848 800 8878
rect 3601 8875 3667 8878
rect 5073 8875 5139 8878
rect 9029 8875 9095 8878
rect 9581 8875 9647 8878
rect 10593 8802 10659 8805
rect 13077 8802 13143 8805
rect 10593 8800 13143 8802
rect 10593 8744 10598 8800
rect 10654 8744 13082 8800
rect 13138 8744 13143 8800
rect 10593 8742 13143 8744
rect 10593 8739 10659 8742
rect 13077 8739 13143 8742
rect 3909 8736 4229 8737
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 8671 4229 8672
rect 9840 8736 10160 8737
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 8671 10160 8672
rect 15770 8736 16090 8737
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 15770 8671 16090 8672
rect 16254 8666 16314 8878
rect 17033 8666 17099 8669
rect 19200 8666 20000 8696
rect 16254 8664 20000 8666
rect 16254 8608 17038 8664
rect 17094 8608 20000 8664
rect 16254 8606 20000 8608
rect 17033 8603 17099 8606
rect 19200 8576 20000 8606
rect 11053 8530 11119 8533
rect 17953 8530 18019 8533
rect 11053 8528 18019 8530
rect 11053 8472 11058 8528
rect 11114 8472 17958 8528
rect 18014 8472 18019 8528
rect 11053 8470 18019 8472
rect 11053 8467 11119 8470
rect 17953 8467 18019 8470
rect 0 8394 800 8424
rect 1393 8394 1459 8397
rect 0 8392 1459 8394
rect 0 8336 1398 8392
rect 1454 8336 1459 8392
rect 0 8334 1459 8336
rect 0 8304 800 8334
rect 1393 8331 1459 8334
rect 6085 8394 6151 8397
rect 8569 8394 8635 8397
rect 6085 8392 8635 8394
rect 6085 8336 6090 8392
rect 6146 8336 8574 8392
rect 8630 8336 8635 8392
rect 6085 8334 8635 8336
rect 6085 8331 6151 8334
rect 8569 8331 8635 8334
rect 10409 8394 10475 8397
rect 13721 8394 13787 8397
rect 10409 8392 13787 8394
rect 10409 8336 10414 8392
rect 10470 8336 13726 8392
rect 13782 8336 13787 8392
rect 10409 8334 13787 8336
rect 10409 8331 10475 8334
rect 13721 8331 13787 8334
rect 17585 8258 17651 8261
rect 19200 8258 20000 8288
rect 17585 8256 20000 8258
rect 17585 8200 17590 8256
rect 17646 8200 20000 8256
rect 17585 8198 20000 8200
rect 17585 8195 17651 8198
rect 6874 8192 7194 8193
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7194 8192
rect 6874 8127 7194 8128
rect 12805 8192 13125 8193
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 19200 8168 20000 8198
rect 12805 8127 13125 8128
rect 0 7986 800 8016
rect 1577 7986 1643 7989
rect 0 7984 1643 7986
rect 0 7928 1582 7984
rect 1638 7928 1643 7984
rect 0 7926 1643 7928
rect 0 7896 800 7926
rect 1577 7923 1643 7926
rect 7281 7986 7347 7989
rect 17309 7986 17375 7989
rect 17953 7986 18019 7989
rect 7281 7984 18019 7986
rect 7281 7928 7286 7984
rect 7342 7928 17314 7984
rect 17370 7928 17958 7984
rect 18014 7928 18019 7984
rect 7281 7926 18019 7928
rect 7281 7923 7347 7926
rect 17309 7923 17375 7926
rect 17953 7923 18019 7926
rect 3693 7850 3759 7853
rect 12617 7850 12683 7853
rect 3693 7848 12683 7850
rect 3693 7792 3698 7848
rect 3754 7792 12622 7848
rect 12678 7792 12683 7848
rect 3693 7790 12683 7792
rect 3693 7787 3759 7790
rect 12617 7787 12683 7790
rect 14733 7850 14799 7853
rect 16941 7850 17007 7853
rect 14733 7848 17007 7850
rect 14733 7792 14738 7848
rect 14794 7792 16946 7848
rect 17002 7792 17007 7848
rect 14733 7790 17007 7792
rect 14733 7787 14799 7790
rect 16941 7787 17007 7790
rect 18321 7850 18387 7853
rect 19200 7850 20000 7880
rect 18321 7848 20000 7850
rect 18321 7792 18326 7848
rect 18382 7792 20000 7848
rect 18321 7790 20000 7792
rect 18321 7787 18387 7790
rect 19200 7760 20000 7790
rect 3909 7648 4229 7649
rect 0 7578 800 7608
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 7583 4229 7584
rect 9840 7648 10160 7649
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 7583 10160 7584
rect 15770 7648 16090 7649
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 7583 16090 7584
rect 1761 7578 1827 7581
rect 0 7576 1827 7578
rect 0 7520 1766 7576
rect 1822 7520 1827 7576
rect 0 7518 1827 7520
rect 0 7488 800 7518
rect 1761 7515 1827 7518
rect 11881 7578 11947 7581
rect 12341 7578 12407 7581
rect 11881 7576 12407 7578
rect 11881 7520 11886 7576
rect 11942 7520 12346 7576
rect 12402 7520 12407 7576
rect 11881 7518 12407 7520
rect 11881 7515 11947 7518
rect 12341 7515 12407 7518
rect 2865 7442 2931 7445
rect 9029 7442 9095 7445
rect 2865 7440 9095 7442
rect 2865 7384 2870 7440
rect 2926 7384 9034 7440
rect 9090 7384 9095 7440
rect 2865 7382 9095 7384
rect 2865 7379 2931 7382
rect 9029 7379 9095 7382
rect 18045 7442 18111 7445
rect 19200 7442 20000 7472
rect 18045 7440 20000 7442
rect 18045 7384 18050 7440
rect 18106 7384 20000 7440
rect 18045 7382 20000 7384
rect 18045 7379 18111 7382
rect 19200 7352 20000 7382
rect 8753 7306 8819 7309
rect 17953 7306 18019 7309
rect 8753 7304 18019 7306
rect 8753 7248 8758 7304
rect 8814 7248 17958 7304
rect 18014 7248 18019 7304
rect 8753 7246 18019 7248
rect 8753 7243 8819 7246
rect 17953 7243 18019 7246
rect 0 7170 800 7200
rect 3509 7170 3575 7173
rect 0 7168 3575 7170
rect 0 7112 3514 7168
rect 3570 7112 3575 7168
rect 0 7110 3575 7112
rect 0 7080 800 7110
rect 3509 7107 3575 7110
rect 6874 7104 7194 7105
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7194 7104
rect 6874 7039 7194 7040
rect 12805 7104 13125 7105
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 7039 13125 7040
rect 16757 7034 16823 7037
rect 16254 7032 16823 7034
rect 16254 6976 16762 7032
rect 16818 6976 16823 7032
rect 16254 6974 16823 6976
rect 11145 6898 11211 6901
rect 15326 6898 15332 6900
rect 11145 6896 15332 6898
rect 11145 6840 11150 6896
rect 11206 6840 15332 6896
rect 11145 6838 15332 6840
rect 11145 6835 11211 6838
rect 15326 6836 15332 6838
rect 15396 6898 15402 6900
rect 16254 6898 16314 6974
rect 16757 6971 16823 6974
rect 18229 7034 18295 7037
rect 19200 7034 20000 7064
rect 18229 7032 20000 7034
rect 18229 6976 18234 7032
rect 18290 6976 20000 7032
rect 18229 6974 20000 6976
rect 18229 6971 18295 6974
rect 19200 6944 20000 6974
rect 16481 6900 16547 6901
rect 16430 6898 16436 6900
rect 15396 6838 16314 6898
rect 16390 6838 16436 6898
rect 16500 6896 16547 6900
rect 16542 6840 16547 6896
rect 15396 6836 15402 6838
rect 16430 6836 16436 6838
rect 16500 6836 16547 6840
rect 16481 6835 16547 6836
rect 0 6762 800 6792
rect 2957 6762 3023 6765
rect 0 6760 3023 6762
rect 0 6704 2962 6760
rect 3018 6704 3023 6760
rect 0 6702 3023 6704
rect 0 6672 800 6702
rect 2957 6699 3023 6702
rect 3509 6762 3575 6765
rect 4521 6762 4587 6765
rect 3509 6760 4587 6762
rect 3509 6704 3514 6760
rect 3570 6704 4526 6760
rect 4582 6704 4587 6760
rect 3509 6702 4587 6704
rect 3509 6699 3575 6702
rect 4521 6699 4587 6702
rect 10317 6762 10383 6765
rect 12709 6762 12775 6765
rect 10317 6760 12775 6762
rect 10317 6704 10322 6760
rect 10378 6704 12714 6760
rect 12770 6704 12775 6760
rect 10317 6702 12775 6704
rect 10317 6699 10383 6702
rect 12709 6699 12775 6702
rect 3909 6560 4229 6561
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 6495 4229 6496
rect 9840 6560 10160 6561
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 6495 10160 6496
rect 15770 6560 16090 6561
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 15770 6495 16090 6496
rect 17953 6490 18019 6493
rect 19200 6490 20000 6520
rect 17953 6488 20000 6490
rect 17953 6432 17958 6488
rect 18014 6432 20000 6488
rect 17953 6430 20000 6432
rect 17953 6427 18019 6430
rect 19200 6400 20000 6430
rect 0 6354 800 6384
rect 2405 6354 2471 6357
rect 0 6352 2471 6354
rect 0 6296 2410 6352
rect 2466 6296 2471 6352
rect 0 6294 2471 6296
rect 0 6264 800 6294
rect 2405 6291 2471 6294
rect 18137 6082 18203 6085
rect 19200 6082 20000 6112
rect 18137 6080 20000 6082
rect 18137 6024 18142 6080
rect 18198 6024 20000 6080
rect 18137 6022 20000 6024
rect 18137 6019 18203 6022
rect 6874 6016 7194 6017
rect 0 5946 800 5976
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7194 6016
rect 6874 5951 7194 5952
rect 12805 6016 13125 6017
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 19200 5992 20000 6022
rect 12805 5951 13125 5952
rect 1853 5946 1919 5949
rect 0 5944 1919 5946
rect 0 5888 1858 5944
rect 1914 5888 1919 5944
rect 0 5886 1919 5888
rect 0 5856 800 5886
rect 1853 5883 1919 5886
rect 12249 5810 12315 5813
rect 12709 5810 12775 5813
rect 12249 5808 12775 5810
rect 12249 5752 12254 5808
rect 12310 5752 12714 5808
rect 12770 5752 12775 5808
rect 12249 5750 12775 5752
rect 12249 5747 12315 5750
rect 12709 5747 12775 5750
rect 11237 5674 11303 5677
rect 16021 5674 16087 5677
rect 11237 5672 16087 5674
rect 11237 5616 11242 5672
rect 11298 5616 16026 5672
rect 16082 5616 16087 5672
rect 11237 5614 16087 5616
rect 11237 5611 11303 5614
rect 16021 5611 16087 5614
rect 18229 5674 18295 5677
rect 19200 5674 20000 5704
rect 18229 5672 20000 5674
rect 18229 5616 18234 5672
rect 18290 5616 20000 5672
rect 18229 5614 20000 5616
rect 18229 5611 18295 5614
rect 19200 5584 20000 5614
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 3909 5472 4229 5473
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 5407 4229 5408
rect 9840 5472 10160 5473
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 5407 10160 5408
rect 15770 5472 16090 5473
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 15770 5407 16090 5408
rect 18413 5266 18479 5269
rect 19200 5266 20000 5296
rect 18413 5264 20000 5266
rect 18413 5208 18418 5264
rect 18474 5208 20000 5264
rect 18413 5206 20000 5208
rect 18413 5203 18479 5206
rect 19200 5176 20000 5206
rect 0 5130 800 5160
rect 1577 5130 1643 5133
rect 0 5128 1643 5130
rect 0 5072 1582 5128
rect 1638 5072 1643 5128
rect 0 5070 1643 5072
rect 0 5040 800 5070
rect 1577 5067 1643 5070
rect 13721 4994 13787 4997
rect 16573 4994 16639 4997
rect 13721 4992 16639 4994
rect 13721 4936 13726 4992
rect 13782 4936 16578 4992
rect 16634 4936 16639 4992
rect 13721 4934 16639 4936
rect 13721 4931 13787 4934
rect 16573 4931 16639 4934
rect 6874 4928 7194 4929
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7194 4928
rect 6874 4863 7194 4864
rect 12805 4928 13125 4929
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 4863 13125 4864
rect 17861 4858 17927 4861
rect 19200 4858 20000 4888
rect 17861 4856 20000 4858
rect 17861 4800 17866 4856
rect 17922 4800 20000 4856
rect 17861 4798 20000 4800
rect 17861 4795 17927 4798
rect 19200 4768 20000 4798
rect 0 4722 800 4752
rect 2405 4722 2471 4725
rect 0 4720 2471 4722
rect 0 4664 2410 4720
rect 2466 4664 2471 4720
rect 0 4662 2471 4664
rect 0 4632 800 4662
rect 2405 4659 2471 4662
rect 18229 4450 18295 4453
rect 19200 4450 20000 4480
rect 18229 4448 20000 4450
rect 18229 4392 18234 4448
rect 18290 4392 20000 4448
rect 18229 4390 20000 4392
rect 18229 4387 18295 4390
rect 3909 4384 4229 4385
rect 0 4314 800 4344
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 4319 4229 4320
rect 9840 4384 10160 4385
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 4319 10160 4320
rect 15770 4384 16090 4385
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 19200 4360 20000 4390
rect 15770 4319 16090 4320
rect 1853 4314 1919 4317
rect 0 4312 1919 4314
rect 0 4256 1858 4312
rect 1914 4256 1919 4312
rect 0 4254 1919 4256
rect 0 4224 800 4254
rect 1853 4251 1919 4254
rect 11789 4042 11855 4045
rect 16297 4042 16363 4045
rect 11789 4040 16363 4042
rect 11789 3984 11794 4040
rect 11850 3984 16302 4040
rect 16358 3984 16363 4040
rect 11789 3982 16363 3984
rect 11789 3979 11855 3982
rect 16297 3979 16363 3982
rect 17861 4042 17927 4045
rect 19200 4042 20000 4072
rect 17861 4040 20000 4042
rect 17861 3984 17866 4040
rect 17922 3984 20000 4040
rect 17861 3982 20000 3984
rect 17861 3979 17927 3982
rect 19200 3952 20000 3982
rect 0 3906 800 3936
rect 2497 3906 2563 3909
rect 0 3904 2563 3906
rect 0 3848 2502 3904
rect 2558 3848 2563 3904
rect 0 3846 2563 3848
rect 0 3816 800 3846
rect 2497 3843 2563 3846
rect 6874 3840 7194 3841
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7194 3840
rect 6874 3775 7194 3776
rect 12805 3840 13125 3841
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 3775 13125 3776
rect 17585 3634 17651 3637
rect 19200 3634 20000 3664
rect 17585 3632 20000 3634
rect 17585 3576 17590 3632
rect 17646 3576 20000 3632
rect 17585 3574 20000 3576
rect 17585 3571 17651 3574
rect 19200 3544 20000 3574
rect 0 3498 800 3528
rect 1853 3498 1919 3501
rect 0 3496 1919 3498
rect 0 3440 1858 3496
rect 1914 3440 1919 3496
rect 0 3438 1919 3440
rect 0 3408 800 3438
rect 1853 3435 1919 3438
rect 3909 3296 4229 3297
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 3231 4229 3232
rect 9840 3296 10160 3297
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 3231 10160 3232
rect 15770 3296 16090 3297
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15770 3231 16090 3232
rect 0 3090 800 3120
rect 2405 3090 2471 3093
rect 0 3088 2471 3090
rect 0 3032 2410 3088
rect 2466 3032 2471 3088
rect 0 3030 2471 3032
rect 0 3000 800 3030
rect 2405 3027 2471 3030
rect 12249 3090 12315 3093
rect 12525 3090 12591 3093
rect 12249 3088 12591 3090
rect 12249 3032 12254 3088
rect 12310 3032 12530 3088
rect 12586 3032 12591 3088
rect 12249 3030 12591 3032
rect 12249 3027 12315 3030
rect 12525 3027 12591 3030
rect 18045 3090 18111 3093
rect 19200 3090 20000 3120
rect 18045 3088 20000 3090
rect 18045 3032 18050 3088
rect 18106 3032 20000 3088
rect 18045 3030 20000 3032
rect 18045 3027 18111 3030
rect 19200 3000 20000 3030
rect 6874 2752 7194 2753
rect 0 2682 800 2712
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7194 2752
rect 6874 2687 7194 2688
rect 12805 2752 13125 2753
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 12805 2687 13125 2688
rect 1853 2682 1919 2685
rect 0 2680 1919 2682
rect 0 2624 1858 2680
rect 1914 2624 1919 2680
rect 0 2622 1919 2624
rect 0 2592 800 2622
rect 1853 2619 1919 2622
rect 17585 2682 17651 2685
rect 19200 2682 20000 2712
rect 17585 2680 20000 2682
rect 17585 2624 17590 2680
rect 17646 2624 20000 2680
rect 17585 2622 20000 2624
rect 17585 2619 17651 2622
rect 19200 2592 20000 2622
rect 15510 2484 15516 2548
rect 15580 2546 15586 2548
rect 15837 2546 15903 2549
rect 15580 2544 15903 2546
rect 15580 2488 15842 2544
rect 15898 2488 15903 2544
rect 15580 2486 15903 2488
rect 15580 2484 15586 2486
rect 15837 2483 15903 2486
rect 0 2274 800 2304
rect 2957 2274 3023 2277
rect 0 2272 3023 2274
rect 0 2216 2962 2272
rect 3018 2216 3023 2272
rect 0 2214 3023 2216
rect 0 2184 800 2214
rect 2957 2211 3023 2214
rect 17309 2274 17375 2277
rect 19200 2274 20000 2304
rect 17309 2272 20000 2274
rect 17309 2216 17314 2272
rect 17370 2216 20000 2272
rect 17309 2214 20000 2216
rect 17309 2211 17375 2214
rect 3909 2208 4229 2209
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2143 4229 2144
rect 9840 2208 10160 2209
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2143 10160 2144
rect 15770 2208 16090 2209
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 19200 2184 20000 2214
rect 15770 2143 16090 2144
rect 0 1866 800 1896
rect 3325 1866 3391 1869
rect 0 1864 3391 1866
rect 0 1808 3330 1864
rect 3386 1808 3391 1864
rect 0 1806 3391 1808
rect 0 1776 800 1806
rect 3325 1803 3391 1806
rect 17585 1866 17651 1869
rect 19200 1866 20000 1896
rect 17585 1864 20000 1866
rect 17585 1808 17590 1864
rect 17646 1808 20000 1864
rect 17585 1806 20000 1808
rect 17585 1803 17651 1806
rect 19200 1776 20000 1806
rect 0 1458 800 1488
rect 2773 1458 2839 1461
rect 0 1456 2839 1458
rect 0 1400 2778 1456
rect 2834 1400 2839 1456
rect 0 1398 2839 1400
rect 0 1368 800 1398
rect 2773 1395 2839 1398
rect 18689 1458 18755 1461
rect 19200 1458 20000 1488
rect 18689 1456 20000 1458
rect 18689 1400 18694 1456
rect 18750 1400 20000 1456
rect 18689 1398 20000 1400
rect 18689 1395 18755 1398
rect 19200 1368 20000 1398
rect 0 1050 800 1080
rect 933 1050 999 1053
rect 0 1048 999 1050
rect 0 992 938 1048
rect 994 992 999 1048
rect 0 990 999 992
rect 0 960 800 990
rect 933 987 999 990
rect 17861 1050 17927 1053
rect 19200 1050 20000 1080
rect 17861 1048 20000 1050
rect 17861 992 17866 1048
rect 17922 992 20000 1048
rect 17861 990 20000 992
rect 17861 987 17927 990
rect 19200 960 20000 990
rect 0 642 800 672
rect 1209 642 1275 645
rect 0 640 1275 642
rect 0 584 1214 640
rect 1270 584 1275 640
rect 0 582 1275 584
rect 0 552 800 582
rect 1209 579 1275 582
rect 17677 642 17743 645
rect 19200 642 20000 672
rect 17677 640 20000 642
rect 17677 584 17682 640
rect 17738 584 20000 640
rect 17677 582 20000 584
rect 17677 579 17743 582
rect 19200 552 20000 582
rect 0 234 800 264
rect 3049 234 3115 237
rect 0 232 3115 234
rect 0 176 3054 232
rect 3110 176 3115 232
rect 0 174 3115 176
rect 0 144 800 174
rect 3049 171 3115 174
rect 18229 234 18295 237
rect 19200 234 20000 264
rect 18229 232 20000 234
rect 18229 176 18234 232
rect 18290 176 20000 232
rect 18229 174 20000 176
rect 18229 171 18295 174
rect 19200 144 20000 174
<< via3 >>
rect 6882 14716 6946 14720
rect 6882 14660 6886 14716
rect 6886 14660 6942 14716
rect 6942 14660 6946 14716
rect 6882 14656 6946 14660
rect 6962 14716 7026 14720
rect 6962 14660 6966 14716
rect 6966 14660 7022 14716
rect 7022 14660 7026 14716
rect 6962 14656 7026 14660
rect 7042 14716 7106 14720
rect 7042 14660 7046 14716
rect 7046 14660 7102 14716
rect 7102 14660 7106 14716
rect 7042 14656 7106 14660
rect 7122 14716 7186 14720
rect 7122 14660 7126 14716
rect 7126 14660 7182 14716
rect 7182 14660 7186 14716
rect 7122 14656 7186 14660
rect 12813 14716 12877 14720
rect 12813 14660 12817 14716
rect 12817 14660 12873 14716
rect 12873 14660 12877 14716
rect 12813 14656 12877 14660
rect 12893 14716 12957 14720
rect 12893 14660 12897 14716
rect 12897 14660 12953 14716
rect 12953 14660 12957 14716
rect 12893 14656 12957 14660
rect 12973 14716 13037 14720
rect 12973 14660 12977 14716
rect 12977 14660 13033 14716
rect 13033 14660 13037 14716
rect 12973 14656 13037 14660
rect 13053 14716 13117 14720
rect 13053 14660 13057 14716
rect 13057 14660 13113 14716
rect 13113 14660 13117 14716
rect 13053 14656 13117 14660
rect 8524 14452 8588 14516
rect 3917 14172 3981 14176
rect 3917 14116 3921 14172
rect 3921 14116 3977 14172
rect 3977 14116 3981 14172
rect 3917 14112 3981 14116
rect 3997 14172 4061 14176
rect 3997 14116 4001 14172
rect 4001 14116 4057 14172
rect 4057 14116 4061 14172
rect 3997 14112 4061 14116
rect 4077 14172 4141 14176
rect 4077 14116 4081 14172
rect 4081 14116 4137 14172
rect 4137 14116 4141 14172
rect 4077 14112 4141 14116
rect 4157 14172 4221 14176
rect 4157 14116 4161 14172
rect 4161 14116 4217 14172
rect 4217 14116 4221 14172
rect 4157 14112 4221 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 15778 14172 15842 14176
rect 15778 14116 15782 14172
rect 15782 14116 15838 14172
rect 15838 14116 15842 14172
rect 15778 14112 15842 14116
rect 15858 14172 15922 14176
rect 15858 14116 15862 14172
rect 15862 14116 15918 14172
rect 15918 14116 15922 14172
rect 15858 14112 15922 14116
rect 15938 14172 16002 14176
rect 15938 14116 15942 14172
rect 15942 14116 15998 14172
rect 15998 14116 16002 14172
rect 15938 14112 16002 14116
rect 16018 14172 16082 14176
rect 16018 14116 16022 14172
rect 16022 14116 16078 14172
rect 16078 14116 16082 14172
rect 16018 14112 16082 14116
rect 6882 13628 6946 13632
rect 6882 13572 6886 13628
rect 6886 13572 6942 13628
rect 6942 13572 6946 13628
rect 6882 13568 6946 13572
rect 6962 13628 7026 13632
rect 6962 13572 6966 13628
rect 6966 13572 7022 13628
rect 7022 13572 7026 13628
rect 6962 13568 7026 13572
rect 7042 13628 7106 13632
rect 7042 13572 7046 13628
rect 7046 13572 7102 13628
rect 7102 13572 7106 13628
rect 7042 13568 7106 13572
rect 7122 13628 7186 13632
rect 7122 13572 7126 13628
rect 7126 13572 7182 13628
rect 7182 13572 7186 13628
rect 7122 13568 7186 13572
rect 12813 13628 12877 13632
rect 12813 13572 12817 13628
rect 12817 13572 12873 13628
rect 12873 13572 12877 13628
rect 12813 13568 12877 13572
rect 12893 13628 12957 13632
rect 12893 13572 12897 13628
rect 12897 13572 12953 13628
rect 12953 13572 12957 13628
rect 12893 13568 12957 13572
rect 12973 13628 13037 13632
rect 12973 13572 12977 13628
rect 12977 13572 13033 13628
rect 13033 13572 13037 13628
rect 12973 13568 13037 13572
rect 13053 13628 13117 13632
rect 13053 13572 13057 13628
rect 13057 13572 13113 13628
rect 13113 13572 13117 13628
rect 13053 13568 13117 13572
rect 3917 13084 3981 13088
rect 3917 13028 3921 13084
rect 3921 13028 3977 13084
rect 3977 13028 3981 13084
rect 3917 13024 3981 13028
rect 3997 13084 4061 13088
rect 3997 13028 4001 13084
rect 4001 13028 4057 13084
rect 4057 13028 4061 13084
rect 3997 13024 4061 13028
rect 4077 13084 4141 13088
rect 4077 13028 4081 13084
rect 4081 13028 4137 13084
rect 4137 13028 4141 13084
rect 4077 13024 4141 13028
rect 4157 13084 4221 13088
rect 4157 13028 4161 13084
rect 4161 13028 4217 13084
rect 4217 13028 4221 13084
rect 4157 13024 4221 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 15778 13084 15842 13088
rect 15778 13028 15782 13084
rect 15782 13028 15838 13084
rect 15838 13028 15842 13084
rect 15778 13024 15842 13028
rect 15858 13084 15922 13088
rect 15858 13028 15862 13084
rect 15862 13028 15918 13084
rect 15918 13028 15922 13084
rect 15858 13024 15922 13028
rect 15938 13084 16002 13088
rect 15938 13028 15942 13084
rect 15942 13028 15998 13084
rect 15998 13028 16002 13084
rect 15938 13024 16002 13028
rect 16018 13084 16082 13088
rect 16018 13028 16022 13084
rect 16022 13028 16078 13084
rect 16078 13028 16082 13084
rect 16018 13024 16082 13028
rect 6882 12540 6946 12544
rect 6882 12484 6886 12540
rect 6886 12484 6942 12540
rect 6942 12484 6946 12540
rect 6882 12480 6946 12484
rect 6962 12540 7026 12544
rect 6962 12484 6966 12540
rect 6966 12484 7022 12540
rect 7022 12484 7026 12540
rect 6962 12480 7026 12484
rect 7042 12540 7106 12544
rect 7042 12484 7046 12540
rect 7046 12484 7102 12540
rect 7102 12484 7106 12540
rect 7042 12480 7106 12484
rect 7122 12540 7186 12544
rect 7122 12484 7126 12540
rect 7126 12484 7182 12540
rect 7182 12484 7186 12540
rect 7122 12480 7186 12484
rect 12813 12540 12877 12544
rect 12813 12484 12817 12540
rect 12817 12484 12873 12540
rect 12873 12484 12877 12540
rect 12813 12480 12877 12484
rect 12893 12540 12957 12544
rect 12893 12484 12897 12540
rect 12897 12484 12953 12540
rect 12953 12484 12957 12540
rect 12893 12480 12957 12484
rect 12973 12540 13037 12544
rect 12973 12484 12977 12540
rect 12977 12484 13033 12540
rect 13033 12484 13037 12540
rect 12973 12480 13037 12484
rect 13053 12540 13117 12544
rect 13053 12484 13057 12540
rect 13057 12484 13113 12540
rect 13113 12484 13117 12540
rect 13053 12480 13117 12484
rect 3917 11996 3981 12000
rect 3917 11940 3921 11996
rect 3921 11940 3977 11996
rect 3977 11940 3981 11996
rect 3917 11936 3981 11940
rect 3997 11996 4061 12000
rect 3997 11940 4001 11996
rect 4001 11940 4057 11996
rect 4057 11940 4061 11996
rect 3997 11936 4061 11940
rect 4077 11996 4141 12000
rect 4077 11940 4081 11996
rect 4081 11940 4137 11996
rect 4137 11940 4141 11996
rect 4077 11936 4141 11940
rect 4157 11996 4221 12000
rect 4157 11940 4161 11996
rect 4161 11940 4217 11996
rect 4217 11940 4221 11996
rect 4157 11936 4221 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 15778 11996 15842 12000
rect 15778 11940 15782 11996
rect 15782 11940 15838 11996
rect 15838 11940 15842 11996
rect 15778 11936 15842 11940
rect 15858 11996 15922 12000
rect 15858 11940 15862 11996
rect 15862 11940 15918 11996
rect 15918 11940 15922 11996
rect 15858 11936 15922 11940
rect 15938 11996 16002 12000
rect 15938 11940 15942 11996
rect 15942 11940 15998 11996
rect 15998 11940 16002 11996
rect 15938 11936 16002 11940
rect 16018 11996 16082 12000
rect 16018 11940 16022 11996
rect 16022 11940 16078 11996
rect 16078 11940 16082 11996
rect 16018 11936 16082 11940
rect 6882 11452 6946 11456
rect 6882 11396 6886 11452
rect 6886 11396 6942 11452
rect 6942 11396 6946 11452
rect 6882 11392 6946 11396
rect 6962 11452 7026 11456
rect 6962 11396 6966 11452
rect 6966 11396 7022 11452
rect 7022 11396 7026 11452
rect 6962 11392 7026 11396
rect 7042 11452 7106 11456
rect 7042 11396 7046 11452
rect 7046 11396 7102 11452
rect 7102 11396 7106 11452
rect 7042 11392 7106 11396
rect 7122 11452 7186 11456
rect 7122 11396 7126 11452
rect 7126 11396 7182 11452
rect 7182 11396 7186 11452
rect 7122 11392 7186 11396
rect 12813 11452 12877 11456
rect 12813 11396 12817 11452
rect 12817 11396 12873 11452
rect 12873 11396 12877 11452
rect 12813 11392 12877 11396
rect 12893 11452 12957 11456
rect 12893 11396 12897 11452
rect 12897 11396 12953 11452
rect 12953 11396 12957 11452
rect 12893 11392 12957 11396
rect 12973 11452 13037 11456
rect 12973 11396 12977 11452
rect 12977 11396 13033 11452
rect 13033 11396 13037 11452
rect 12973 11392 13037 11396
rect 13053 11452 13117 11456
rect 13053 11396 13057 11452
rect 13057 11396 13113 11452
rect 13113 11396 13117 11452
rect 13053 11392 13117 11396
rect 16436 10976 16500 10980
rect 16436 10920 16450 10976
rect 16450 10920 16500 10976
rect 16436 10916 16500 10920
rect 3917 10908 3981 10912
rect 3917 10852 3921 10908
rect 3921 10852 3977 10908
rect 3977 10852 3981 10908
rect 3917 10848 3981 10852
rect 3997 10908 4061 10912
rect 3997 10852 4001 10908
rect 4001 10852 4057 10908
rect 4057 10852 4061 10908
rect 3997 10848 4061 10852
rect 4077 10908 4141 10912
rect 4077 10852 4081 10908
rect 4081 10852 4137 10908
rect 4137 10852 4141 10908
rect 4077 10848 4141 10852
rect 4157 10908 4221 10912
rect 4157 10852 4161 10908
rect 4161 10852 4217 10908
rect 4217 10852 4221 10908
rect 4157 10848 4221 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 15778 10908 15842 10912
rect 15778 10852 15782 10908
rect 15782 10852 15838 10908
rect 15838 10852 15842 10908
rect 15778 10848 15842 10852
rect 15858 10908 15922 10912
rect 15858 10852 15862 10908
rect 15862 10852 15918 10908
rect 15918 10852 15922 10908
rect 15858 10848 15922 10852
rect 15938 10908 16002 10912
rect 15938 10852 15942 10908
rect 15942 10852 15998 10908
rect 15998 10852 16002 10908
rect 15938 10848 16002 10852
rect 16018 10908 16082 10912
rect 16018 10852 16022 10908
rect 16022 10852 16078 10908
rect 16078 10852 16082 10908
rect 16018 10848 16082 10852
rect 15332 10704 15396 10708
rect 15332 10648 15382 10704
rect 15382 10648 15396 10704
rect 15332 10644 15396 10648
rect 6882 10364 6946 10368
rect 6882 10308 6886 10364
rect 6886 10308 6942 10364
rect 6942 10308 6946 10364
rect 6882 10304 6946 10308
rect 6962 10364 7026 10368
rect 6962 10308 6966 10364
rect 6966 10308 7022 10364
rect 7022 10308 7026 10364
rect 6962 10304 7026 10308
rect 7042 10364 7106 10368
rect 7042 10308 7046 10364
rect 7046 10308 7102 10364
rect 7102 10308 7106 10364
rect 7042 10304 7106 10308
rect 7122 10364 7186 10368
rect 7122 10308 7126 10364
rect 7126 10308 7182 10364
rect 7182 10308 7186 10364
rect 7122 10304 7186 10308
rect 12813 10364 12877 10368
rect 12813 10308 12817 10364
rect 12817 10308 12873 10364
rect 12873 10308 12877 10364
rect 12813 10304 12877 10308
rect 12893 10364 12957 10368
rect 12893 10308 12897 10364
rect 12897 10308 12953 10364
rect 12953 10308 12957 10364
rect 12893 10304 12957 10308
rect 12973 10364 13037 10368
rect 12973 10308 12977 10364
rect 12977 10308 13033 10364
rect 13033 10308 13037 10364
rect 12973 10304 13037 10308
rect 13053 10364 13117 10368
rect 13053 10308 13057 10364
rect 13057 10308 13113 10364
rect 13113 10308 13117 10364
rect 13053 10304 13117 10308
rect 3917 9820 3981 9824
rect 3917 9764 3921 9820
rect 3921 9764 3977 9820
rect 3977 9764 3981 9820
rect 3917 9760 3981 9764
rect 3997 9820 4061 9824
rect 3997 9764 4001 9820
rect 4001 9764 4057 9820
rect 4057 9764 4061 9820
rect 3997 9760 4061 9764
rect 4077 9820 4141 9824
rect 4077 9764 4081 9820
rect 4081 9764 4137 9820
rect 4137 9764 4141 9820
rect 4077 9760 4141 9764
rect 4157 9820 4221 9824
rect 4157 9764 4161 9820
rect 4161 9764 4217 9820
rect 4217 9764 4221 9820
rect 4157 9760 4221 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 15778 9820 15842 9824
rect 15778 9764 15782 9820
rect 15782 9764 15838 9820
rect 15838 9764 15842 9820
rect 15778 9760 15842 9764
rect 15858 9820 15922 9824
rect 15858 9764 15862 9820
rect 15862 9764 15918 9820
rect 15918 9764 15922 9820
rect 15858 9760 15922 9764
rect 15938 9820 16002 9824
rect 15938 9764 15942 9820
rect 15942 9764 15998 9820
rect 15998 9764 16002 9820
rect 15938 9760 16002 9764
rect 16018 9820 16082 9824
rect 16018 9764 16022 9820
rect 16022 9764 16078 9820
rect 16078 9764 16082 9820
rect 16018 9760 16082 9764
rect 15516 9420 15580 9484
rect 8524 9284 8588 9348
rect 6882 9276 6946 9280
rect 6882 9220 6886 9276
rect 6886 9220 6942 9276
rect 6942 9220 6946 9276
rect 6882 9216 6946 9220
rect 6962 9276 7026 9280
rect 6962 9220 6966 9276
rect 6966 9220 7022 9276
rect 7022 9220 7026 9276
rect 6962 9216 7026 9220
rect 7042 9276 7106 9280
rect 7042 9220 7046 9276
rect 7046 9220 7102 9276
rect 7102 9220 7106 9276
rect 7042 9216 7106 9220
rect 7122 9276 7186 9280
rect 7122 9220 7126 9276
rect 7126 9220 7182 9276
rect 7182 9220 7186 9276
rect 7122 9216 7186 9220
rect 12813 9276 12877 9280
rect 12813 9220 12817 9276
rect 12817 9220 12873 9276
rect 12873 9220 12877 9276
rect 12813 9216 12877 9220
rect 12893 9276 12957 9280
rect 12893 9220 12897 9276
rect 12897 9220 12953 9276
rect 12953 9220 12957 9276
rect 12893 9216 12957 9220
rect 12973 9276 13037 9280
rect 12973 9220 12977 9276
rect 12977 9220 13033 9276
rect 13033 9220 13037 9276
rect 12973 9216 13037 9220
rect 13053 9276 13117 9280
rect 13053 9220 13057 9276
rect 13057 9220 13113 9276
rect 13113 9220 13117 9276
rect 13053 9216 13117 9220
rect 3917 8732 3981 8736
rect 3917 8676 3921 8732
rect 3921 8676 3977 8732
rect 3977 8676 3981 8732
rect 3917 8672 3981 8676
rect 3997 8732 4061 8736
rect 3997 8676 4001 8732
rect 4001 8676 4057 8732
rect 4057 8676 4061 8732
rect 3997 8672 4061 8676
rect 4077 8732 4141 8736
rect 4077 8676 4081 8732
rect 4081 8676 4137 8732
rect 4137 8676 4141 8732
rect 4077 8672 4141 8676
rect 4157 8732 4221 8736
rect 4157 8676 4161 8732
rect 4161 8676 4217 8732
rect 4217 8676 4221 8732
rect 4157 8672 4221 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 15778 8732 15842 8736
rect 15778 8676 15782 8732
rect 15782 8676 15838 8732
rect 15838 8676 15842 8732
rect 15778 8672 15842 8676
rect 15858 8732 15922 8736
rect 15858 8676 15862 8732
rect 15862 8676 15918 8732
rect 15918 8676 15922 8732
rect 15858 8672 15922 8676
rect 15938 8732 16002 8736
rect 15938 8676 15942 8732
rect 15942 8676 15998 8732
rect 15998 8676 16002 8732
rect 15938 8672 16002 8676
rect 16018 8732 16082 8736
rect 16018 8676 16022 8732
rect 16022 8676 16078 8732
rect 16078 8676 16082 8732
rect 16018 8672 16082 8676
rect 6882 8188 6946 8192
rect 6882 8132 6886 8188
rect 6886 8132 6942 8188
rect 6942 8132 6946 8188
rect 6882 8128 6946 8132
rect 6962 8188 7026 8192
rect 6962 8132 6966 8188
rect 6966 8132 7022 8188
rect 7022 8132 7026 8188
rect 6962 8128 7026 8132
rect 7042 8188 7106 8192
rect 7042 8132 7046 8188
rect 7046 8132 7102 8188
rect 7102 8132 7106 8188
rect 7042 8128 7106 8132
rect 7122 8188 7186 8192
rect 7122 8132 7126 8188
rect 7126 8132 7182 8188
rect 7182 8132 7186 8188
rect 7122 8128 7186 8132
rect 12813 8188 12877 8192
rect 12813 8132 12817 8188
rect 12817 8132 12873 8188
rect 12873 8132 12877 8188
rect 12813 8128 12877 8132
rect 12893 8188 12957 8192
rect 12893 8132 12897 8188
rect 12897 8132 12953 8188
rect 12953 8132 12957 8188
rect 12893 8128 12957 8132
rect 12973 8188 13037 8192
rect 12973 8132 12977 8188
rect 12977 8132 13033 8188
rect 13033 8132 13037 8188
rect 12973 8128 13037 8132
rect 13053 8188 13117 8192
rect 13053 8132 13057 8188
rect 13057 8132 13113 8188
rect 13113 8132 13117 8188
rect 13053 8128 13117 8132
rect 3917 7644 3981 7648
rect 3917 7588 3921 7644
rect 3921 7588 3977 7644
rect 3977 7588 3981 7644
rect 3917 7584 3981 7588
rect 3997 7644 4061 7648
rect 3997 7588 4001 7644
rect 4001 7588 4057 7644
rect 4057 7588 4061 7644
rect 3997 7584 4061 7588
rect 4077 7644 4141 7648
rect 4077 7588 4081 7644
rect 4081 7588 4137 7644
rect 4137 7588 4141 7644
rect 4077 7584 4141 7588
rect 4157 7644 4221 7648
rect 4157 7588 4161 7644
rect 4161 7588 4217 7644
rect 4217 7588 4221 7644
rect 4157 7584 4221 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 15778 7644 15842 7648
rect 15778 7588 15782 7644
rect 15782 7588 15838 7644
rect 15838 7588 15842 7644
rect 15778 7584 15842 7588
rect 15858 7644 15922 7648
rect 15858 7588 15862 7644
rect 15862 7588 15918 7644
rect 15918 7588 15922 7644
rect 15858 7584 15922 7588
rect 15938 7644 16002 7648
rect 15938 7588 15942 7644
rect 15942 7588 15998 7644
rect 15998 7588 16002 7644
rect 15938 7584 16002 7588
rect 16018 7644 16082 7648
rect 16018 7588 16022 7644
rect 16022 7588 16078 7644
rect 16078 7588 16082 7644
rect 16018 7584 16082 7588
rect 6882 7100 6946 7104
rect 6882 7044 6886 7100
rect 6886 7044 6942 7100
rect 6942 7044 6946 7100
rect 6882 7040 6946 7044
rect 6962 7100 7026 7104
rect 6962 7044 6966 7100
rect 6966 7044 7022 7100
rect 7022 7044 7026 7100
rect 6962 7040 7026 7044
rect 7042 7100 7106 7104
rect 7042 7044 7046 7100
rect 7046 7044 7102 7100
rect 7102 7044 7106 7100
rect 7042 7040 7106 7044
rect 7122 7100 7186 7104
rect 7122 7044 7126 7100
rect 7126 7044 7182 7100
rect 7182 7044 7186 7100
rect 7122 7040 7186 7044
rect 12813 7100 12877 7104
rect 12813 7044 12817 7100
rect 12817 7044 12873 7100
rect 12873 7044 12877 7100
rect 12813 7040 12877 7044
rect 12893 7100 12957 7104
rect 12893 7044 12897 7100
rect 12897 7044 12953 7100
rect 12953 7044 12957 7100
rect 12893 7040 12957 7044
rect 12973 7100 13037 7104
rect 12973 7044 12977 7100
rect 12977 7044 13033 7100
rect 13033 7044 13037 7100
rect 12973 7040 13037 7044
rect 13053 7100 13117 7104
rect 13053 7044 13057 7100
rect 13057 7044 13113 7100
rect 13113 7044 13117 7100
rect 13053 7040 13117 7044
rect 15332 6836 15396 6900
rect 16436 6896 16500 6900
rect 16436 6840 16486 6896
rect 16486 6840 16500 6896
rect 16436 6836 16500 6840
rect 3917 6556 3981 6560
rect 3917 6500 3921 6556
rect 3921 6500 3977 6556
rect 3977 6500 3981 6556
rect 3917 6496 3981 6500
rect 3997 6556 4061 6560
rect 3997 6500 4001 6556
rect 4001 6500 4057 6556
rect 4057 6500 4061 6556
rect 3997 6496 4061 6500
rect 4077 6556 4141 6560
rect 4077 6500 4081 6556
rect 4081 6500 4137 6556
rect 4137 6500 4141 6556
rect 4077 6496 4141 6500
rect 4157 6556 4221 6560
rect 4157 6500 4161 6556
rect 4161 6500 4217 6556
rect 4217 6500 4221 6556
rect 4157 6496 4221 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 15778 6556 15842 6560
rect 15778 6500 15782 6556
rect 15782 6500 15838 6556
rect 15838 6500 15842 6556
rect 15778 6496 15842 6500
rect 15858 6556 15922 6560
rect 15858 6500 15862 6556
rect 15862 6500 15918 6556
rect 15918 6500 15922 6556
rect 15858 6496 15922 6500
rect 15938 6556 16002 6560
rect 15938 6500 15942 6556
rect 15942 6500 15998 6556
rect 15998 6500 16002 6556
rect 15938 6496 16002 6500
rect 16018 6556 16082 6560
rect 16018 6500 16022 6556
rect 16022 6500 16078 6556
rect 16078 6500 16082 6556
rect 16018 6496 16082 6500
rect 6882 6012 6946 6016
rect 6882 5956 6886 6012
rect 6886 5956 6942 6012
rect 6942 5956 6946 6012
rect 6882 5952 6946 5956
rect 6962 6012 7026 6016
rect 6962 5956 6966 6012
rect 6966 5956 7022 6012
rect 7022 5956 7026 6012
rect 6962 5952 7026 5956
rect 7042 6012 7106 6016
rect 7042 5956 7046 6012
rect 7046 5956 7102 6012
rect 7102 5956 7106 6012
rect 7042 5952 7106 5956
rect 7122 6012 7186 6016
rect 7122 5956 7126 6012
rect 7126 5956 7182 6012
rect 7182 5956 7186 6012
rect 7122 5952 7186 5956
rect 12813 6012 12877 6016
rect 12813 5956 12817 6012
rect 12817 5956 12873 6012
rect 12873 5956 12877 6012
rect 12813 5952 12877 5956
rect 12893 6012 12957 6016
rect 12893 5956 12897 6012
rect 12897 5956 12953 6012
rect 12953 5956 12957 6012
rect 12893 5952 12957 5956
rect 12973 6012 13037 6016
rect 12973 5956 12977 6012
rect 12977 5956 13033 6012
rect 13033 5956 13037 6012
rect 12973 5952 13037 5956
rect 13053 6012 13117 6016
rect 13053 5956 13057 6012
rect 13057 5956 13113 6012
rect 13113 5956 13117 6012
rect 13053 5952 13117 5956
rect 3917 5468 3981 5472
rect 3917 5412 3921 5468
rect 3921 5412 3977 5468
rect 3977 5412 3981 5468
rect 3917 5408 3981 5412
rect 3997 5468 4061 5472
rect 3997 5412 4001 5468
rect 4001 5412 4057 5468
rect 4057 5412 4061 5468
rect 3997 5408 4061 5412
rect 4077 5468 4141 5472
rect 4077 5412 4081 5468
rect 4081 5412 4137 5468
rect 4137 5412 4141 5468
rect 4077 5408 4141 5412
rect 4157 5468 4221 5472
rect 4157 5412 4161 5468
rect 4161 5412 4217 5468
rect 4217 5412 4221 5468
rect 4157 5408 4221 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 15778 5468 15842 5472
rect 15778 5412 15782 5468
rect 15782 5412 15838 5468
rect 15838 5412 15842 5468
rect 15778 5408 15842 5412
rect 15858 5468 15922 5472
rect 15858 5412 15862 5468
rect 15862 5412 15918 5468
rect 15918 5412 15922 5468
rect 15858 5408 15922 5412
rect 15938 5468 16002 5472
rect 15938 5412 15942 5468
rect 15942 5412 15998 5468
rect 15998 5412 16002 5468
rect 15938 5408 16002 5412
rect 16018 5468 16082 5472
rect 16018 5412 16022 5468
rect 16022 5412 16078 5468
rect 16078 5412 16082 5468
rect 16018 5408 16082 5412
rect 6882 4924 6946 4928
rect 6882 4868 6886 4924
rect 6886 4868 6942 4924
rect 6942 4868 6946 4924
rect 6882 4864 6946 4868
rect 6962 4924 7026 4928
rect 6962 4868 6966 4924
rect 6966 4868 7022 4924
rect 7022 4868 7026 4924
rect 6962 4864 7026 4868
rect 7042 4924 7106 4928
rect 7042 4868 7046 4924
rect 7046 4868 7102 4924
rect 7102 4868 7106 4924
rect 7042 4864 7106 4868
rect 7122 4924 7186 4928
rect 7122 4868 7126 4924
rect 7126 4868 7182 4924
rect 7182 4868 7186 4924
rect 7122 4864 7186 4868
rect 12813 4924 12877 4928
rect 12813 4868 12817 4924
rect 12817 4868 12873 4924
rect 12873 4868 12877 4924
rect 12813 4864 12877 4868
rect 12893 4924 12957 4928
rect 12893 4868 12897 4924
rect 12897 4868 12953 4924
rect 12953 4868 12957 4924
rect 12893 4864 12957 4868
rect 12973 4924 13037 4928
rect 12973 4868 12977 4924
rect 12977 4868 13033 4924
rect 13033 4868 13037 4924
rect 12973 4864 13037 4868
rect 13053 4924 13117 4928
rect 13053 4868 13057 4924
rect 13057 4868 13113 4924
rect 13113 4868 13117 4924
rect 13053 4864 13117 4868
rect 3917 4380 3981 4384
rect 3917 4324 3921 4380
rect 3921 4324 3977 4380
rect 3977 4324 3981 4380
rect 3917 4320 3981 4324
rect 3997 4380 4061 4384
rect 3997 4324 4001 4380
rect 4001 4324 4057 4380
rect 4057 4324 4061 4380
rect 3997 4320 4061 4324
rect 4077 4380 4141 4384
rect 4077 4324 4081 4380
rect 4081 4324 4137 4380
rect 4137 4324 4141 4380
rect 4077 4320 4141 4324
rect 4157 4380 4221 4384
rect 4157 4324 4161 4380
rect 4161 4324 4217 4380
rect 4217 4324 4221 4380
rect 4157 4320 4221 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 15778 4380 15842 4384
rect 15778 4324 15782 4380
rect 15782 4324 15838 4380
rect 15838 4324 15842 4380
rect 15778 4320 15842 4324
rect 15858 4380 15922 4384
rect 15858 4324 15862 4380
rect 15862 4324 15918 4380
rect 15918 4324 15922 4380
rect 15858 4320 15922 4324
rect 15938 4380 16002 4384
rect 15938 4324 15942 4380
rect 15942 4324 15998 4380
rect 15998 4324 16002 4380
rect 15938 4320 16002 4324
rect 16018 4380 16082 4384
rect 16018 4324 16022 4380
rect 16022 4324 16078 4380
rect 16078 4324 16082 4380
rect 16018 4320 16082 4324
rect 6882 3836 6946 3840
rect 6882 3780 6886 3836
rect 6886 3780 6942 3836
rect 6942 3780 6946 3836
rect 6882 3776 6946 3780
rect 6962 3836 7026 3840
rect 6962 3780 6966 3836
rect 6966 3780 7022 3836
rect 7022 3780 7026 3836
rect 6962 3776 7026 3780
rect 7042 3836 7106 3840
rect 7042 3780 7046 3836
rect 7046 3780 7102 3836
rect 7102 3780 7106 3836
rect 7042 3776 7106 3780
rect 7122 3836 7186 3840
rect 7122 3780 7126 3836
rect 7126 3780 7182 3836
rect 7182 3780 7186 3836
rect 7122 3776 7186 3780
rect 12813 3836 12877 3840
rect 12813 3780 12817 3836
rect 12817 3780 12873 3836
rect 12873 3780 12877 3836
rect 12813 3776 12877 3780
rect 12893 3836 12957 3840
rect 12893 3780 12897 3836
rect 12897 3780 12953 3836
rect 12953 3780 12957 3836
rect 12893 3776 12957 3780
rect 12973 3836 13037 3840
rect 12973 3780 12977 3836
rect 12977 3780 13033 3836
rect 13033 3780 13037 3836
rect 12973 3776 13037 3780
rect 13053 3836 13117 3840
rect 13053 3780 13057 3836
rect 13057 3780 13113 3836
rect 13113 3780 13117 3836
rect 13053 3776 13117 3780
rect 3917 3292 3981 3296
rect 3917 3236 3921 3292
rect 3921 3236 3977 3292
rect 3977 3236 3981 3292
rect 3917 3232 3981 3236
rect 3997 3292 4061 3296
rect 3997 3236 4001 3292
rect 4001 3236 4057 3292
rect 4057 3236 4061 3292
rect 3997 3232 4061 3236
rect 4077 3292 4141 3296
rect 4077 3236 4081 3292
rect 4081 3236 4137 3292
rect 4137 3236 4141 3292
rect 4077 3232 4141 3236
rect 4157 3292 4221 3296
rect 4157 3236 4161 3292
rect 4161 3236 4217 3292
rect 4217 3236 4221 3292
rect 4157 3232 4221 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 15778 3292 15842 3296
rect 15778 3236 15782 3292
rect 15782 3236 15838 3292
rect 15838 3236 15842 3292
rect 15778 3232 15842 3236
rect 15858 3292 15922 3296
rect 15858 3236 15862 3292
rect 15862 3236 15918 3292
rect 15918 3236 15922 3292
rect 15858 3232 15922 3236
rect 15938 3292 16002 3296
rect 15938 3236 15942 3292
rect 15942 3236 15998 3292
rect 15998 3236 16002 3292
rect 15938 3232 16002 3236
rect 16018 3292 16082 3296
rect 16018 3236 16022 3292
rect 16022 3236 16078 3292
rect 16078 3236 16082 3292
rect 16018 3232 16082 3236
rect 6882 2748 6946 2752
rect 6882 2692 6886 2748
rect 6886 2692 6942 2748
rect 6942 2692 6946 2748
rect 6882 2688 6946 2692
rect 6962 2748 7026 2752
rect 6962 2692 6966 2748
rect 6966 2692 7022 2748
rect 7022 2692 7026 2748
rect 6962 2688 7026 2692
rect 7042 2748 7106 2752
rect 7042 2692 7046 2748
rect 7046 2692 7102 2748
rect 7102 2692 7106 2748
rect 7042 2688 7106 2692
rect 7122 2748 7186 2752
rect 7122 2692 7126 2748
rect 7126 2692 7182 2748
rect 7182 2692 7186 2748
rect 7122 2688 7186 2692
rect 12813 2748 12877 2752
rect 12813 2692 12817 2748
rect 12817 2692 12873 2748
rect 12873 2692 12877 2748
rect 12813 2688 12877 2692
rect 12893 2748 12957 2752
rect 12893 2692 12897 2748
rect 12897 2692 12953 2748
rect 12953 2692 12957 2748
rect 12893 2688 12957 2692
rect 12973 2748 13037 2752
rect 12973 2692 12977 2748
rect 12977 2692 13033 2748
rect 13033 2692 13037 2748
rect 12973 2688 13037 2692
rect 13053 2748 13117 2752
rect 13053 2692 13057 2748
rect 13057 2692 13113 2748
rect 13113 2692 13117 2748
rect 13053 2688 13117 2692
rect 15516 2484 15580 2548
rect 3917 2204 3981 2208
rect 3917 2148 3921 2204
rect 3921 2148 3977 2204
rect 3977 2148 3981 2204
rect 3917 2144 3981 2148
rect 3997 2204 4061 2208
rect 3997 2148 4001 2204
rect 4001 2148 4057 2204
rect 4057 2148 4061 2204
rect 3997 2144 4061 2148
rect 4077 2204 4141 2208
rect 4077 2148 4081 2204
rect 4081 2148 4137 2204
rect 4137 2148 4141 2204
rect 4077 2144 4141 2148
rect 4157 2204 4221 2208
rect 4157 2148 4161 2204
rect 4161 2148 4217 2204
rect 4217 2148 4221 2204
rect 4157 2144 4221 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 15778 2204 15842 2208
rect 15778 2148 15782 2204
rect 15782 2148 15838 2204
rect 15838 2148 15842 2204
rect 15778 2144 15842 2148
rect 15858 2204 15922 2208
rect 15858 2148 15862 2204
rect 15862 2148 15918 2204
rect 15918 2148 15922 2204
rect 15858 2144 15922 2148
rect 15938 2204 16002 2208
rect 15938 2148 15942 2204
rect 15942 2148 15998 2204
rect 15998 2148 16002 2204
rect 15938 2144 16002 2148
rect 16018 2204 16082 2208
rect 16018 2148 16022 2204
rect 16022 2148 16078 2204
rect 16078 2148 16082 2204
rect 16018 2144 16082 2148
<< metal4 >>
rect 3909 14176 4229 14736
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 13088 4229 14112
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 12000 4229 13024
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 10912 4229 11936
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 9824 4229 10848
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 8736 4229 9760
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 7648 4229 8672
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 6560 4229 7584
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 5472 4229 6496
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 4384 4229 5408
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 3296 4229 4320
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 2208 4229 3232
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2128 4229 2144
rect 6874 14720 7195 14736
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7195 14720
rect 6874 13632 7195 14656
rect 8523 14516 8589 14517
rect 8523 14452 8524 14516
rect 8588 14452 8589 14516
rect 8523 14451 8589 14452
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7195 13632
rect 6874 12544 7195 13568
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7195 12544
rect 6874 11456 7195 12480
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7195 11456
rect 6874 10368 7195 11392
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7195 10368
rect 6874 9280 7195 10304
rect 8526 9349 8586 14451
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 8523 9348 8589 9349
rect 8523 9284 8524 9348
rect 8588 9284 8589 9348
rect 8523 9283 8589 9284
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7195 9280
rect 6874 8192 7195 9216
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7195 8192
rect 6874 7104 7195 8128
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7195 7104
rect 6874 6016 7195 7040
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7195 6016
rect 6874 4928 7195 5952
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7195 4928
rect 6874 3840 7195 4864
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7195 3840
rect 6874 2752 7195 3776
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7195 2752
rect 6874 2128 7195 2688
rect 9840 8736 10160 9760
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 6560 10160 7584
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 2208 10160 3232
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12805 14720 13125 14736
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 13632 13125 14656
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 12544 13125 13568
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 11456 13125 12480
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 10368 13125 11392
rect 15770 14176 16090 14736
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 15770 13088 16090 14112
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 15770 12000 16090 13024
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 15770 10912 16090 11936
rect 16435 10980 16501 10981
rect 16435 10916 16436 10980
rect 16500 10916 16501 10980
rect 16435 10915 16501 10916
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15331 10708 15397 10709
rect 15331 10644 15332 10708
rect 15396 10644 15397 10708
rect 15331 10643 15397 10644
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 12805 9280 13125 10304
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 8192 13125 9216
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 12805 7104 13125 8128
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 6016 13125 7040
rect 15334 6901 15394 10643
rect 15770 9824 16090 10848
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 15515 9484 15581 9485
rect 15515 9420 15516 9484
rect 15580 9420 15581 9484
rect 15515 9419 15581 9420
rect 15331 6900 15397 6901
rect 15331 6836 15332 6900
rect 15396 6836 15397 6900
rect 15331 6835 15397 6836
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12805 4928 13125 5952
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 3840 13125 4864
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 2752 13125 3776
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 12805 2128 13125 2688
rect 15518 2549 15578 9419
rect 15770 8736 16090 9760
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 15770 7648 16090 8672
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 6560 16090 7584
rect 16438 6901 16498 10915
rect 16435 6900 16501 6901
rect 16435 6836 16436 6900
rect 16500 6836 16501 6900
rect 16435 6835 16501 6836
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 15770 5472 16090 6496
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 15770 4384 16090 5408
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 15770 3296 16090 4320
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15515 2548 15581 2549
rect 15515 2484 15516 2548
rect 15580 2484 15581 2548
rect 15515 2483 15581 2484
rect 15770 2208 16090 3232
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 15770 2128 16090 2144
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608763569
transform -1 0 18860 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608763569
transform 1 0 18216 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_168
timestamp 1608763569
transform 1 0 16560 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_180
timestamp 1608763569
transform 1 0 17664 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_22_187
timestamp 1608763569
transform 1 0 18308 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608763569
transform 1 0 15364 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_149
timestamp 1608763569
transform 1 0 14812 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_156
timestamp 1608763569
transform 1 0 15456 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_137
timestamp 1608763569
transform 1 0 13708 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608763569
transform 1 0 12512 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_106
timestamp 1608763569
transform 1 0 10856 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_118
timestamp 1608763569
transform 1 0 11960 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_125
timestamp 1608763569
transform 1 0 12604 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608763569
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_87
timestamp 1608763569
transform 1 0 9108 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_94
timestamp 1608763569
transform 1 0 9752 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_63
timestamp 1608763569
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_75
timestamp 1608763569
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608763569
transform 1 0 6808 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1608763569
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_56
timestamp 1608763569
transform 1 0 6256 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608763569
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_23
timestamp 1608763569
transform 1 0 3220 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1608763569
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1608763569
transform 1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608763569
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1608763569
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_11
timestamp 1608763569
transform 1 0 2116 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608763569
transform -1 0 18860 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608763569
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_174
timestamp 1608763569
transform 1 0 17112 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1608763569
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_184
timestamp 1608763569
transform 1 0 18032 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1608763569
transform 1 0 15088 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1608763569
transform 1 0 15640 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_149
timestamp 1608763569
transform 1 0 14812 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_156
timestamp 1608763569
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_162
timestamp 1608763569
transform 1 0 16008 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1608763569
transform 1 0 13616 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1608763569
transform 1 0 14444 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_135
timestamp 1608763569
transform 1 0 13524 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_140
timestamp 1608763569
transform 1 0 13984 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_144
timestamp 1608763569
transform 1 0 14352 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608763569
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_114
timestamp 1608763569
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1608763569
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_90
timestamp 1608763569
transform 1 0 9384 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_102
timestamp 1608763569
transform 1 0 10488 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_66
timestamp 1608763569
transform 1 0 7176 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_78
timestamp 1608763569
transform 1 0 8280 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1608763569
transform 1 0 5980 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1608763569
transform 1 0 6808 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608763569
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_52
timestamp 1608763569
transform 1 0 5888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1608763569
transform 1 0 6348 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1608763569
transform 1 0 3312 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_22
timestamp 1608763569
transform 1 0 3128 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_28
timestamp 1608763569
transform 1 0 3680 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_40
timestamp 1608763569
transform 1 0 4784 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1608763569
transform 1 0 1656 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1608763569
transform 1 0 2208 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1608763569
transform 1 0 2760 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608763569
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1608763569
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_10
timestamp 1608763569
transform 1 0 2024 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_16
timestamp 1608763569
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608763569
transform -1 0 18860 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608763569
transform -1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608763569
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_171
timestamp 1608763569
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_184
timestamp 1608763569
transform 1 0 18032 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1608763569
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608763569
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1608763569
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_159
timestamp 1608763569
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1608763569
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1608763569
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1608763569
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1608763569
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1608763569
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608763569
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1608763569
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1608763569
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1608763569
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1608763569
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608763569
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1608763569
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1608763569
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1608763569
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1608763569
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1608763569
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1608763569
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608763569
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_46
timestamp 1608763569
transform 1 0 5336 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_58
timestamp 1608763569
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1608763569
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1608763569
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1608763569
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1608763569
transform 1 0 3220 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1608763569
transform 1 0 4508 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608763569
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_21
timestamp 1608763569
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_32
timestamp 1608763569
transform 1 0 4048 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_36
timestamp 1608763569
transform 1 0 4416 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1608763569
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1608763569
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1608763569
transform 1 0 2208 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1608763569
transform 1 0 1840 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608763569
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608763569
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1608763569
transform 1 0 1380 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_11
timestamp 1608763569
transform 1 0 2116 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1608763569
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1608763569
transform 1 0 1748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_17
timestamp 1608763569
transform 1 0 2668 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608763569
transform -1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1608763569
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608763569
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1608763569
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1608763569
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1608763569
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1608763569
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1608763569
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1608763569
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608763569
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1608763569
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1608763569
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_70
timestamp 1608763569
transform 1 0 7544 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_82
timestamp 1608763569
transform 1 0 8648 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763569
transform 1 0 6072 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_52
timestamp 1608763569
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763569
transform 1 0 4416 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608763569
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1608763569
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_32
timestamp 1608763569
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _11_
timestamp 1608763569
transform 1 0 1840 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763569
transform 1 0 2300 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608763569
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1608763569
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp 1608763569
transform 1 0 1748 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_11
timestamp 1608763569
transform 1 0 2116 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608763569
transform -1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608763569
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_171
timestamp 1608763569
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_184
timestamp 1608763569
transform 1 0 18032 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_147
timestamp 1608763569
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_159
timestamp 1608763569
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1608763569
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608763569
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_115
timestamp 1608763569
transform 1 0 11684 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1608763569
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1608763569
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1608763569
transform 1 0 9752 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_84
timestamp 1608763569
transform 1 0 8832 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_92
timestamp 1608763569
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_103
timestamp 1608763569
transform 1 0 10580 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00
timestamp 1608763569
transform 1 0 7728 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_70
timestamp 1608763569
transform 1 0 7544 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1608763569
transform 1 0 5336 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608763569
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_42
timestamp 1608763569
transform 1 0 4968 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_55
timestamp 1608763569
transform 1 0 6164 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_62
timestamp 1608763569
transform 1 0 6808 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763569
transform 1 0 3496 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_21
timestamp 1608763569
transform 1 0 3036 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_25
timestamp 1608763569
transform 1 0 3404 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1608763569
transform 1 0 2208 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608763569
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1608763569
transform 1 0 1380 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_11
timestamp 1608763569
transform 1 0 2116 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608763569
transform -1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1608763569
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608763569
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1608763569
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1608763569
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1608763569
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_140
timestamp 1608763569
transform 1 0 13984 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763569
transform 1 0 12512 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1608763569
transform 1 0 11500 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_109
timestamp 1608763569
transform 1 0 11132 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_122
timestamp 1608763569
transform 1 0 12328 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763569
transform 1 0 9660 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608763569
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_89
timestamp 1608763569
transform 1 0 9292 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_77
timestamp 1608763569
transform 1 0 8188 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763569
transform 1 0 6716 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1608763569
transform 1 0 5612 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_47
timestamp 1608763569
transform 1 0 5428 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_58
timestamp 1608763569
transform 1 0 6440 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1608763569
transform 1 0 4600 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608763569
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_26
timestamp 1608763569
transform 1 0 3496 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1608763569
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_32
timestamp 1608763569
transform 1 0 4048 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_2_
timestamp 1608763569
transform 1 0 2668 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1608763569
transform 1 0 1656 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608763569
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1608763569
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_15
timestamp 1608763569
transform 1 0 2484 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608763569
transform -1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1608763569
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1608763569
transform 1 0 16928 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608763569
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_170
timestamp 1608763569
transform 1 0 16744 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1608763569
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_187
timestamp 1608763569
transform 1 0 18308 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1608763569
transform 1 0 15916 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_156
timestamp 1608763569
transform 1 0 15456 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_160
timestamp 1608763569
transform 1 0 15824 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763569
transform 1 0 13984 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_15_134
timestamp 1608763569
transform 1 0 13432 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1608763569
transform 1 0 12604 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608763569
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_117
timestamp 1608763569
transform 1 0 11868 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1608763569
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_123
timestamp 1608763569
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763569
transform 1 0 10396 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1608763569
transform 1 0 9384 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_85
timestamp 1608763569
transform 1 0 8924 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_89
timestamp 1608763569
transform 1 0 9292 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_99
timestamp 1608763569
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763569
transform 1 0 7452 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_68
timestamp 1608763569
transform 1 0 7360 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1608763569
transform 1 0 5336 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608763569
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_44
timestamp 1608763569
transform 1 0 5152 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_55
timestamp 1608763569
transform 1 0 6164 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_62
timestamp 1608763569
transform 1 0 6808 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1608763569
transform 1 0 4324 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_30
timestamp 1608763569
transform 1 0 3864 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_34
timestamp 1608763569
transform 1 0 4232 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763569
transform 1 0 2392 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1608763569
transform 1 0 1380 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608763569
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_12
timestamp 1608763569
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608763569
transform -1 0 18860 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608763569
transform -1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_188
timestamp 1608763569
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_188
timestamp 1608763569
transform 1 0 18400 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1608763569
transform 1 0 18032 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1608763569
transform 1 0 18032 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1608763569
transform 1 0 17388 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1608763569
transform 1 0 17020 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608763569
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_174
timestamp 1608763569
transform 1 0 17112 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1608763569
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_171
timestamp 1608763569
transform 1 0 16836 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_182
timestamp 1608763569
transform 1 0 17848 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763569
transform 1 0 15364 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1608763569
transform 1 0 16284 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1608763569
transform 1 0 15272 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608763569
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_152
timestamp 1608763569
transform 1 0 15088 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_163
timestamp 1608763569
transform 1 0 16100 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1608763569
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_154
timestamp 1608763569
transform 1 0 15272 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763569
transform 1 0 13524 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1608763569
transform 1 0 14260 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1608763569
transform 1 0 12880 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_127
timestamp 1608763569
transform 1 0 12788 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_137
timestamp 1608763569
transform 1 0 13708 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_131
timestamp 1608763569
transform 1 0 13156 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1608763569
transform 1 0 11592 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1608763569
transform 1 0 12328 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608763569
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_112
timestamp 1608763569
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_117
timestamp 1608763569
transform 1 0 11868 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1608763569
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_123
timestamp 1608763569
transform 1 0 12420 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_113
timestamp 1608763569
transform 1 0 11500 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_121
timestamp 1608763569
transform 1 0 12236 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1608763569
transform 1 0 8832 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1608763569
transform 1 0 10580 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1608763569
transform 1 0 10672 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1608763569
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608763569
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_93
timestamp 1608763569
transform 1 0 9660 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_101
timestamp 1608763569
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_86
timestamp 1608763569
transform 1 0 9016 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_102
timestamp 1608763569
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763569
transform 1 0 7544 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1608763569
transform 1 0 7820 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_71
timestamp 1608763569
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_82
timestamp 1608763569
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_64
timestamp 1608763569
transform 1 0 6992 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1608763569
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _12_
timestamp 1608763569
transform 1 0 6716 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608763569
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1608763569
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_59
timestamp 1608763569
transform 1 0 6532 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1608763569
transform 1 0 5704 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1608763569
transform 1 0 5704 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763569
transform 1 0 5060 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_47
timestamp 1608763569
transform 1 0 5428 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_46
timestamp 1608763569
transform 1 0 5336 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1608763569
transform 1 0 3864 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_1_
timestamp 1608763569
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763569
transform 1 0 4876 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608763569
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_25
timestamp 1608763569
transform 1 0 3404 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_29
timestamp 1608763569
transform 1 0 3772 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_39
timestamp 1608763569
transform 1 0 4692 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1608763569
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_41
timestamp 1608763569
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763569
transform 1 0 1932 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1608763569
transform 1 0 2944 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_18
timestamp 1608763569
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _31_
timestamp 1608763569
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1608763569
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1608763569
transform 1 0 1932 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608763569
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608763569
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1608763569
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_7
timestamp 1608763569
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608763569
transform -1 0 18860 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1608763569
transform 1 0 17848 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1608763569
transform 1 0 16744 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_168
timestamp 1608763569
transform 1 0 16560 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_179
timestamp 1608763569
transform 1 0 17572 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_186
timestamp 1608763569
transform 1 0 18216 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1608763569
transform 1 0 15732 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608763569
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1608763569
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_154
timestamp 1608763569
transform 1 0 15272 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_158
timestamp 1608763569
transform 1 0 15640 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1608763569
transform 1 0 12880 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_137
timestamp 1608763569
transform 1 0 13708 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763569
transform 1 0 10948 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763569
transform 1 0 12604 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_106
timestamp 1608763569
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_123
timestamp 1608763569
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1608763569
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608763569
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1608763569
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_102
timestamp 1608763569
transform 1 0 10488 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1608763569
transform 1 0 8556 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_78
timestamp 1608763569
transform 1 0 8280 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763569
transform 1 0 6808 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_12_50
timestamp 1608763569
transform 1 0 5704 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1608763569
transform 1 0 4876 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608763569
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_21
timestamp 1608763569
transform 1 0 3036 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1608763569
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_32
timestamp 1608763569
transform 1 0 4048 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_40
timestamp 1608763569
transform 1 0 4784 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763569
transform 1 0 1564 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608763569
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1608763569
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608763569
transform -1 0 18860 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_188
timestamp 1608763569
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1608763569
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1608763569
transform 1 0 16744 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608763569
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_179
timestamp 1608763569
transform 1 0 17572 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1608763569
transform 1 0 16100 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_161
timestamp 1608763569
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_166
timestamp 1608763569
transform 1 0 16376 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763569
transform 1 0 14444 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1608763569
transform 1 0 12880 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_127
timestamp 1608763569
transform 1 0 12788 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_137
timestamp 1608763569
transform 1 0 13708 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608763569
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_116
timestamp 1608763569
transform 1 0 11776 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_123
timestamp 1608763569
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763569
transform 1 0 10304 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1608763569
transform 1 0 7452 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763569
transform 1 0 8464 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_11_68
timestamp 1608763569
transform 1 0 7360 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_78
timestamp 1608763569
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1608763569
transform 1 0 5428 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608763569
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763569
transform 1 0 6440 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_43
timestamp 1608763569
transform 1 0 5060 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_56
timestamp 1608763569
transform 1 0 6256 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_62
timestamp 1608763569
transform 1 0 6808 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763569
transform 1 0 3588 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_25
timestamp 1608763569
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1608763569
transform 1 0 1656 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1608763569
transform 1 0 2576 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608763569
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1608763569
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_10
timestamp 1608763569
transform 1 0 2024 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608763569
transform -1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1608763569
transform 1 0 17940 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1608763569
transform 1 0 16928 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_170
timestamp 1608763569
transform 1 0 16744 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_181
timestamp 1608763569
transform 1 0 17756 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_187
timestamp 1608763569
transform 1 0 18308 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763569
transform 1 0 15272 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608763569
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_148
timestamp 1608763569
transform 1 0 14720 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1608763569
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_1_
timestamp 1608763569
transform 1 0 12880 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_2_
timestamp 1608763569
transform 1 0 13892 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_126
timestamp 1608763569
transform 1 0 12696 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_137
timestamp 1608763569
transform 1 0 13708 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1608763569
transform 1 0 11868 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763569
transform 1 0 11316 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_109
timestamp 1608763569
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_114
timestamp 1608763569
transform 1 0 11592 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763569
transform 1 0 9660 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608763569
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1608763569
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1608763569
transform 1 0 8556 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1608763569
transform 1 0 7636 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_10_64
timestamp 1608763569
transform 1 0 6992 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_70
timestamp 1608763569
transform 1 0 7544 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_80
timestamp 1608763569
transform 1 0 8464 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763569
transform 1 0 5520 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_46
timestamp 1608763569
transform 1 0 5336 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_1_
timestamp 1608763569
transform 1 0 4508 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608763569
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_25
timestamp 1608763569
transform 1 0 3404 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_32
timestamp 1608763569
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_36
timestamp 1608763569
transform 1 0 4416 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1608763569
transform 1 0 2576 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1608763569
transform 1 0 1564 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608763569
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1608763569
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_14
timestamp 1608763569
transform 1 0 2392 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608763569
transform -1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp 1608763569
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _15_
timestamp 1608763569
transform 1 0 17480 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1608763569
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1608763569
transform 1 0 16468 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608763569
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_176
timestamp 1608763569
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1608763569
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1608763569
transform 1 0 15456 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_153
timestamp 1608763569
transform 1 0 15180 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_165
timestamp 1608763569
transform 1 0 16284 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763569
transform 1 0 13708 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_132
timestamp 1608763569
transform 1 0 13248 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_136
timestamp 1608763569
transform 1 0 13616 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1608763569
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1608763569
transform 1 0 11316 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608763569
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_109
timestamp 1608763569
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1608763569
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1608763569
transform 1 0 10304 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_9_94
timestamp 1608763569
transform 1 0 9752 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763569
transform 1 0 8280 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1608763569
transform 1 0 7268 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_66
timestamp 1608763569
transform 1 0 7176 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_76
timestamp 1608763569
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1608763569
transform 1 0 5612 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608763569
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_47
timestamp 1608763569
transform 1 0 5428 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_58
timestamp 1608763569
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1608763569
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _10_
timestamp 1608763569
transform 1 0 3128 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_2_
timestamp 1608763569
transform 1 0 4600 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1608763569
transform 1 0 3588 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_25
timestamp 1608763569
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_36
timestamp 1608763569
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _30_
timestamp 1608763569
transform 1 0 1564 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1608763569
transform 1 0 2116 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608763569
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1608763569
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_9
timestamp 1608763569
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_20
timestamp 1608763569
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608763569
transform -1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1608763569
transform 1 0 17940 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1608763569
transform 1 0 16928 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_170
timestamp 1608763569
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_181
timestamp 1608763569
transform 1 0 17756 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_187
timestamp 1608763569
transform 1 0 18308 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763569
transform 1 0 15272 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608763569
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1608763569
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1608763569
transform 1 0 13064 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1608763569
transform 1 0 14168 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_128
timestamp 1608763569
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_139
timestamp 1608763569
transform 1 0 13892 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1608763569
transform 1 0 12052 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_115
timestamp 1608763569
transform 1 0 11684 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _13_
timestamp 1608763569
transform 1 0 9016 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763569
transform 1 0 10212 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608763569
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1608763569
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_89
timestamp 1608763569
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_93
timestamp 1608763569
transform 1 0 9660 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _09_
timestamp 1608763569
transform 1 0 7268 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1608763569
transform 1 0 8004 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_65
timestamp 1608763569
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_70
timestamp 1608763569
transform 1 0 7544 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_74
timestamp 1608763569
transform 1 0 7912 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1608763569
transform 1 0 6256 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_48
timestamp 1608763569
transform 1 0 5520 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _29_
timestamp 1608763569
transform 1 0 3312 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763569
transform 1 0 4048 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608763569
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_22
timestamp 1608763569
transform 1 0 3128 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_28
timestamp 1608763569
transform 1 0 3680 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _26_
timestamp 1608763569
transform 1 0 1656 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _27_
timestamp 1608763569
transform 1 0 2208 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _28_
timestamp 1608763569
transform 1 0 2760 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608763569
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1608763569
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_10
timestamp 1608763569
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_16
timestamp 1608763569
transform 1 0 2576 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608763569
transform -1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608763569
transform -1 0 18860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_188
timestamp 1608763569
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1608763569
transform 1 0 17848 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1608763569
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1608763569
transform 1 0 17388 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608763569
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_178
timestamp 1608763569
transform 1 0 17480 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_186
timestamp 1608763569
transform 1 0 18216 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1608763569
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_1_
timestamp 1608763569
transform 1 0 16652 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_167
timestamp 1608763569
transform 1 0 16468 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_172
timestamp 1608763569
transform 1 0 16928 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_176
timestamp 1608763569
transform 1 0 17296 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1608763569
transform 1 0 14628 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1608763569
transform 1 0 16100 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1608763569
transform 1 0 15640 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608763569
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1608763569
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_154
timestamp 1608763569
transform 1 0 15272 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_157
timestamp 1608763569
transform 1 0 15548 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763569
transform 1 0 12880 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763569
transform 1 0 14076 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_6_144
timestamp 1608763569
transform 1 0 14352 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_136
timestamp 1608763569
transform 1 0 13616 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_140
timestamp 1608763569
transform 1 0 13984 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _14_
timestamp 1608763569
transform 1 0 10856 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608763569
transform 1 0 12420 0 1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763569
transform 1 0 11132 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1608763569
transform 1 0 11316 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608763569
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_107
timestamp 1608763569
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_125
timestamp 1608763569
transform 1 0 12604 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_109
timestamp 1608763569
transform 1 0 11132 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1608763569
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763569
transform 1 0 9108 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1608763569
transform 1 0 10672 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1608763569
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608763569
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_86
timestamp 1608763569
transform 1 0 9016 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_102
timestamp 1608763569
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_84
timestamp 1608763569
transform 1 0 8832 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_103
timestamp 1608763569
transform 1 0 10580 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1608763569
transform 1 0 8004 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1608763569
transform 1 0 7084 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_6_74
timestamp 1608763569
transform 1 0 7912 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_71
timestamp 1608763569
transform 1 0 7636 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1608763569
transform 1 0 5520 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1608763569
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608763569
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763569
transform 1 0 6532 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_46
timestamp 1608763569
transform 1 0 5336 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_57
timestamp 1608763569
transform 1 0 6348 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_62
timestamp 1608763569
transform 1 0 6808 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_55
timestamp 1608763569
transform 1 0 6164 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1608763569
transform 1 0 4048 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763569
transform 1 0 4692 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1608763569
transform 1 0 4508 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608763569
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1608763569
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1608763569
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_36
timestamp 1608763569
transform 1 0 4416 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_30
timestamp 1608763569
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_36
timestamp 1608763569
transform 1 0 4416 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763569
transform 1 0 2392 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1608763569
transform 1 0 2944 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_18
timestamp 1608763569
transform 1 0 2760 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _24_
timestamp 1608763569
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _25_
timestamp 1608763569
transform 1 0 1656 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1608763569
transform 1 0 1932 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608763569
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608763569
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_7
timestamp 1608763569
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1608763569
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_10
timestamp 1608763569
transform 1 0 2024 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608763569
transform -1 0 18860 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1608763569
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1608763569
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1608763569
transform 1 0 16652 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608763569
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_167
timestamp 1608763569
transform 1 0 16468 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_178
timestamp 1608763569
transform 1 0 17480 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1608763569
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1608763569
transform 1 0 16192 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1608763569
transform 1 0 15180 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_151
timestamp 1608763569
transform 1 0 14996 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_162
timestamp 1608763569
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1608763569
transform 1 0 13800 0 1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_5_136
timestamp 1608763569
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1608763569
transform 1 0 11776 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608763569
transform 1 0 12420 0 1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1608763569
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_112
timestamp 1608763569
transform 1 0 11408 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1608763569
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763569
transform 1 0 9936 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_94
timestamp 1608763569
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1608763569
transform 1 0 6900 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763569
transform 1 0 8280 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_5_72
timestamp 1608763569
transform 1 0 7728 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763569
transform 1 0 5060 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1608763569
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1608763569
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_62
timestamp 1608763569
transform 1 0 6808 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1608763569
transform 1 0 4048 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1608763569
transform 1 0 3036 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_30
timestamp 1608763569
transform 1 0 3864 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_41
timestamp 1608763569
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763569
transform 1 0 1840 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608763569
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1608763569
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1608763569
transform 1 0 1748 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_14
timestamp 1608763569
transform 1 0 2392 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_20
timestamp 1608763569
transform 1 0 2944 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608763569
transform -1 0 18860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1608763569
transform 1 0 17848 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_2_
timestamp 1608763569
transform 1 0 16652 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_167
timestamp 1608763569
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_178
timestamp 1608763569
transform 1 0 17480 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_186
timestamp 1608763569
transform 1 0 18216 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1608763569
transform 1 0 14628 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1608763569
transform 1 0 15272 0 -1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1608763569
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1608763569
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1608763569
transform 1 0 12880 0 -1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_4_126
timestamp 1608763569
transform 1 0 12696 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_141
timestamp 1608763569
transform 1 0 14076 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1608763569
transform 1 0 11684 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1608763569
transform 1 0 12328 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_113
timestamp 1608763569
transform 1 0 11500 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_119
timestamp 1608763569
transform 1 0 12052 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763569
transform 1 0 10028 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1608763569
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1608763569
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_93
timestamp 1608763569
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1608763569
transform 1 0 8556 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_72
timestamp 1608763569
transform 1 0 7728 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_80
timestamp 1608763569
transform 1 0 8464 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763569
transform 1 0 6256 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_4_46
timestamp 1608763569
transform 1 0 5336 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_54
timestamp 1608763569
transform 1 0 6072 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1608763569
transform 1 0 4508 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763569
transform 1 0 3036 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1608763569
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1608763569
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1608763569
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_36
timestamp 1608763569
transform 1 0 4416 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _22_
timestamp 1608763569
transform 1 0 1656 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _23_
timestamp 1608763569
transform 1 0 2208 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608763569
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1608763569
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_10
timestamp 1608763569
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_16
timestamp 1608763569
transform 1 0 2576 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_20
timestamp 1608763569
transform 1 0 2944 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608763569
transform -1 0 18860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_188
timestamp 1608763569
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1608763569
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1608763569
transform 1 0 17388 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1608763569
transform 1 0 16928 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1608763569
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_170
timestamp 1608763569
transform 1 0 16744 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_175
timestamp 1608763569
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1608763569
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608763569
transform 1 0 15548 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_3_155
timestamp 1608763569
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1608763569
transform 1 0 13616 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1608763569
transform 1 0 13064 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1608763569
transform 1 0 14168 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_3_127
timestamp 1608763569
transform 1 0 12788 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_134
timestamp 1608763569
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_140
timestamp 1608763569
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1608763569
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1608763569
transform 1 0 11040 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1608763569
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608763569
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_106
timestamp 1608763569
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_117
timestamp 1608763569
transform 1 0 11868 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1608763569
transform 1 0 9384 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1608763569
transform 1 0 10028 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_88
timestamp 1608763569
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_94
timestamp 1608763569
transform 1 0 9752 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763569
transform 1 0 7728 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_70
timestamp 1608763569
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1608763569
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_48
timestamp 1608763569
transform 1 0 5520 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_60
timestamp 1608763569
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_62
timestamp 1608763569
transform 1 0 6808 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763569
transform 1 0 4048 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_3_29
timestamp 1608763569
transform 1 0 3772 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1608763569
transform 1 0 2300 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01
timestamp 1608763569
transform 1 0 1564 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608763569
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1608763569
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_11
timestamp 1608763569
transform 1 0 2116 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_17
timestamp 1608763569
transform 1 0 2668 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608763569
transform -1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1608763569
transform 1 0 17848 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1608763569
transform 1 0 17112 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_172
timestamp 1608763569
transform 1 0 16928 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_178
timestamp 1608763569
transform 1 0 17480 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_186
timestamp 1608763569
transform 1 0 18216 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1608763569
transform 1 0 14628 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1608763569
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608763569
transform 1 0 15732 0 -1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1608763569
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1608763569
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_157
timestamp 1608763569
transform 1 0 15548 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1608763569
transform 1 0 14076 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1608763569
transform 1 0 13616 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_140
timestamp 1608763569
transform 1 0 13984 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_145
timestamp 1608763569
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1608763569
transform 1 0 12420 0 -1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763569
transform 1 0 10764 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_121
timestamp 1608763569
transform 1 0 12236 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1608763569
transform 1 0 9752 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1608763569
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1608763569
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_93
timestamp 1608763569
transform 1 0 9660 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_103
timestamp 1608763569
transform 1 0 10580 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1608763569
transform 1 0 8556 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763569
transform 1 0 6900 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_79
timestamp 1608763569
transform 1 0 8372 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763569
transform 1 0 5244 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_2_44
timestamp 1608763569
transform 1 0 5152 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_61
timestamp 1608763569
transform 1 0 6716 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1608763569
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_22
timestamp 1608763569
transform 1 0 3128 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_30
timestamp 1608763569
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1608763569
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _20_
timestamp 1608763569
transform 1 0 1656 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1608763569
transform 1 0 2208 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1608763569
transform 1 0 2760 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608763569
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1608763569
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_10
timestamp 1608763569
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_16
timestamp 1608763569
transform 1 0 2576 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608763569
transform -1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608763569
transform -1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_188
timestamp 1608763569
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp 1608763569
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1608763569
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1608763569
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1608763569
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1608763569
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1608763569
transform 1 0 17664 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1608763569
transform 1 0 17388 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_178
timestamp 1608763569
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1608763569
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1608763569
transform 1 0 17112 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_173
timestamp 1608763569
transform 1 0 17020 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1608763569
transform 1 0 16928 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_176
timestamp 1608763569
transform 1 0 17296 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1608763569
transform 1 0 16652 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1608763569
transform 1 0 14904 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1608763569
transform 1 0 15456 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608763569
transform 1 0 15732 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1608763569
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_148
timestamp 1608763569
transform 1 0 14720 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1608763569
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_156
timestamp 1608763569
transform 1 0 15456 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1608763569
transform 1 0 14352 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608763569
transform 1 0 12880 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1608763569
transform 1 0 12972 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608763569
transform 1 0 14260 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_0_142
timestamp 1608763569
transform 1 0 14168 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_126
timestamp 1608763569
transform 1 0 12696 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_141
timestamp 1608763569
transform 1 0 14076 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1608763569
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1608763569
transform 1 0 11132 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1608763569
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1608763569
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_107
timestamp 1608763569
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1608763569
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1608763569
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_116
timestamp 1608763569
transform 1 0 11776 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1608763569
transform 1 0 9016 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1608763569
transform 1 0 9936 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1608763569
transform 1 0 9752 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608763569
transform 1 0 10580 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1608763569
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_84
timestamp 1608763569
transform 1 0 8832 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_90
timestamp 1608763569
transform 1 0 9384 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_94
timestamp 1608763569
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_100
timestamp 1608763569
transform 1 0 10304 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608763569
transform 1 0 8556 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1608763569
transform 1 0 7912 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1608763569
transform 1 0 7912 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1608763569
transform 1 0 8464 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78
timestamp 1608763569
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_78
timestamp 1608763569
transform 1 0 8280 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1608763569
transform 1 0 6900 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1608763569
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1608763569
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_72
timestamp 1608763569
transform 1 0 7728 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_44
timestamp 1608763569
transform 1 0 5152 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1608763569
transform 1 0 6256 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763569
transform 1 0 5980 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1608763569
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1608763569
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59
timestamp 1608763569
transform 1 0 6532 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1608763569
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_62
timestamp 1608763569
transform 1 0 6808 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1608763569
transform 1 0 5520 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46
timestamp 1608763569
transform 1 0 5336 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51
timestamp 1608763569
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1608763569
transform 1 0 3680 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763569
transform 1 0 3036 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763569
transform 1 0 4048 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46
timestamp 1608763569
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1608763569
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38
timestamp 1608763569
transform 1 0 4600 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_26
timestamp 1608763569
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_32
timestamp 1608763569
transform 1 0 4048 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763569
transform 1 0 2944 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19
timestamp 1608763569
transform 1 0 2852 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_16
timestamp 1608763569
transform 1 0 2576 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _19_
timestamp 1608763569
transform 1 0 2208 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763569
transform 1 0 2300 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11
timestamp 1608763569
transform 1 0 2116 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_10
timestamp 1608763569
transform 1 0 2024 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _18_
timestamp 1608763569
transform 1 0 1656 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763569
transform 1 0 1564 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608763569
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1608763569
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3
timestamp 1608763569
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp 1608763569
transform 1 0 1380 0 1 2720
box -38 -48 314 592
<< labels >>
rlabel metal2 s 7378 16200 7434 17000 4 IO_ISOL_N
port 1 nsew
rlabel metal2 s 5630 0 5686 800 4 SC_IN_BOT
port 2 nsew
rlabel metal2 s 6090 16200 6146 17000 4 SC_IN_TOP
port 3 nsew
rlabel metal2 s 6182 0 6238 800 4 SC_OUT_BOT
port 4 nsew
rlabel metal2 s 6734 16200 6790 17000 4 SC_OUT_TOP
port 5 nsew
rlabel metal2 s 202 0 258 800 4 bottom_grid_pin_0_
port 6 nsew
rlabel metal2 s 2686 0 2742 800 4 bottom_grid_pin_10_
port 7 nsew
rlabel metal2 s 3146 0 3202 800 4 bottom_grid_pin_12_
port 8 nsew
rlabel metal2 s 3606 0 3662 800 4 bottom_grid_pin_14_
port 9 nsew
rlabel metal2 s 4158 0 4214 800 4 bottom_grid_pin_16_
port 10 nsew
rlabel metal2 s 662 0 718 800 4 bottom_grid_pin_2_
port 11 nsew
rlabel metal2 s 1122 0 1178 800 4 bottom_grid_pin_4_
port 12 nsew
rlabel metal2 s 1674 0 1730 800 4 bottom_grid_pin_6_
port 13 nsew
rlabel metal2 s 2134 0 2190 800 4 bottom_grid_pin_8_
port 14 nsew
rlabel metal2 s 4618 0 4674 800 4 ccff_head
port 15 nsew
rlabel metal2 s 5170 0 5226 800 4 ccff_tail
port 16 nsew
rlabel metal3 s 0 8848 800 8968 4 chanx_left_in[0]
port 17 nsew
rlabel metal3 s 0 12928 800 13048 4 chanx_left_in[10]
port 18 nsew
rlabel metal3 s 0 13336 800 13456 4 chanx_left_in[11]
port 19 nsew
rlabel metal3 s 0 13744 800 13864 4 chanx_left_in[12]
port 20 nsew
rlabel metal3 s 0 14152 800 14272 4 chanx_left_in[13]
port 21 nsew
rlabel metal3 s 0 14560 800 14680 4 chanx_left_in[14]
port 22 nsew
rlabel metal3 s 0 14968 800 15088 4 chanx_left_in[15]
port 23 nsew
rlabel metal3 s 0 15376 800 15496 4 chanx_left_in[16]
port 24 nsew
rlabel metal3 s 0 15784 800 15904 4 chanx_left_in[17]
port 25 nsew
rlabel metal3 s 0 16192 800 16312 4 chanx_left_in[18]
port 26 nsew
rlabel metal3 s 0 16600 800 16720 4 chanx_left_in[19]
port 27 nsew
rlabel metal3 s 0 9256 800 9376 4 chanx_left_in[1]
port 28 nsew
rlabel metal3 s 0 9664 800 9784 4 chanx_left_in[2]
port 29 nsew
rlabel metal3 s 0 10072 800 10192 4 chanx_left_in[3]
port 30 nsew
rlabel metal3 s 0 10480 800 10600 4 chanx_left_in[4]
port 31 nsew
rlabel metal3 s 0 10888 800 11008 4 chanx_left_in[5]
port 32 nsew
rlabel metal3 s 0 11296 800 11416 4 chanx_left_in[6]
port 33 nsew
rlabel metal3 s 0 11704 800 11824 4 chanx_left_in[7]
port 34 nsew
rlabel metal3 s 0 12112 800 12232 4 chanx_left_in[8]
port 35 nsew
rlabel metal3 s 0 12520 800 12640 4 chanx_left_in[9]
port 36 nsew
rlabel metal3 s 0 552 800 672 4 chanx_left_out[0]
port 37 nsew
rlabel metal3 s 0 4632 800 4752 4 chanx_left_out[10]
port 38 nsew
rlabel metal3 s 0 5040 800 5160 4 chanx_left_out[11]
port 39 nsew
rlabel metal3 s 0 5448 800 5568 4 chanx_left_out[12]
port 40 nsew
rlabel metal3 s 0 5856 800 5976 4 chanx_left_out[13]
port 41 nsew
rlabel metal3 s 0 6264 800 6384 4 chanx_left_out[14]
port 42 nsew
rlabel metal3 s 0 6672 800 6792 4 chanx_left_out[15]
port 43 nsew
rlabel metal3 s 0 7080 800 7200 4 chanx_left_out[16]
port 44 nsew
rlabel metal3 s 0 7488 800 7608 4 chanx_left_out[17]
port 45 nsew
rlabel metal3 s 0 7896 800 8016 4 chanx_left_out[18]
port 46 nsew
rlabel metal3 s 0 8304 800 8424 4 chanx_left_out[19]
port 47 nsew
rlabel metal3 s 0 960 800 1080 4 chanx_left_out[1]
port 48 nsew
rlabel metal3 s 0 1368 800 1488 4 chanx_left_out[2]
port 49 nsew
rlabel metal3 s 0 1776 800 1896 4 chanx_left_out[3]
port 50 nsew
rlabel metal3 s 0 2184 800 2304 4 chanx_left_out[4]
port 51 nsew
rlabel metal3 s 0 2592 800 2712 4 chanx_left_out[5]
port 52 nsew
rlabel metal3 s 0 3000 800 3120 4 chanx_left_out[6]
port 53 nsew
rlabel metal3 s 0 3408 800 3528 4 chanx_left_out[7]
port 54 nsew
rlabel metal3 s 0 3816 800 3936 4 chanx_left_out[8]
port 55 nsew
rlabel metal3 s 0 4224 800 4344 4 chanx_left_out[9]
port 56 nsew
rlabel metal3 s 19200 8576 20000 8696 4 chanx_right_in[0]
port 57 nsew
rlabel metal3 s 19200 12792 20000 12912 4 chanx_right_in[10]
port 58 nsew
rlabel metal3 s 19200 13200 20000 13320 4 chanx_right_in[11]
port 59 nsew
rlabel metal3 s 19200 13744 20000 13864 4 chanx_right_in[12]
port 60 nsew
rlabel metal3 s 19200 14152 20000 14272 4 chanx_right_in[13]
port 61 nsew
rlabel metal3 s 19200 14560 20000 14680 4 chanx_right_in[14]
port 62 nsew
rlabel metal3 s 19200 14968 20000 15088 4 chanx_right_in[15]
port 63 nsew
rlabel metal3 s 19200 15376 20000 15496 4 chanx_right_in[16]
port 64 nsew
rlabel metal3 s 19200 15784 20000 15904 4 chanx_right_in[17]
port 65 nsew
rlabel metal3 s 19200 16192 20000 16312 4 chanx_right_in[18]
port 66 nsew
rlabel metal3 s 19200 16600 20000 16720 4 chanx_right_in[19]
port 67 nsew
rlabel metal3 s 19200 8984 20000 9104 4 chanx_right_in[1]
port 68 nsew
rlabel metal3 s 19200 9392 20000 9512 4 chanx_right_in[2]
port 69 nsew
rlabel metal3 s 19200 9800 20000 9920 4 chanx_right_in[3]
port 70 nsew
rlabel metal3 s 19200 10344 20000 10464 4 chanx_right_in[4]
port 71 nsew
rlabel metal3 s 19200 10752 20000 10872 4 chanx_right_in[5]
port 72 nsew
rlabel metal3 s 19200 11160 20000 11280 4 chanx_right_in[6]
port 73 nsew
rlabel metal3 s 19200 11568 20000 11688 4 chanx_right_in[7]
port 74 nsew
rlabel metal3 s 19200 11976 20000 12096 4 chanx_right_in[8]
port 75 nsew
rlabel metal3 s 19200 12384 20000 12504 4 chanx_right_in[9]
port 76 nsew
rlabel metal3 s 19200 144 20000 264 4 chanx_right_out[0]
port 77 nsew
rlabel metal3 s 19200 4360 20000 4480 4 chanx_right_out[10]
port 78 nsew
rlabel metal3 s 19200 4768 20000 4888 4 chanx_right_out[11]
port 79 nsew
rlabel metal3 s 19200 5176 20000 5296 4 chanx_right_out[12]
port 80 nsew
rlabel metal3 s 19200 5584 20000 5704 4 chanx_right_out[13]
port 81 nsew
rlabel metal3 s 19200 5992 20000 6112 4 chanx_right_out[14]
port 82 nsew
rlabel metal3 s 19200 6400 20000 6520 4 chanx_right_out[15]
port 83 nsew
rlabel metal3 s 19200 6944 20000 7064 4 chanx_right_out[16]
port 84 nsew
rlabel metal3 s 19200 7352 20000 7472 4 chanx_right_out[17]
port 85 nsew
rlabel metal3 s 19200 7760 20000 7880 4 chanx_right_out[18]
port 86 nsew
rlabel metal3 s 19200 8168 20000 8288 4 chanx_right_out[19]
port 87 nsew
rlabel metal3 s 19200 552 20000 672 4 chanx_right_out[1]
port 88 nsew
rlabel metal3 s 19200 960 20000 1080 4 chanx_right_out[2]
port 89 nsew
rlabel metal3 s 19200 1368 20000 1488 4 chanx_right_out[3]
port 90 nsew
rlabel metal3 s 19200 1776 20000 1896 4 chanx_right_out[4]
port 91 nsew
rlabel metal3 s 19200 2184 20000 2304 4 chanx_right_out[5]
port 92 nsew
rlabel metal3 s 19200 2592 20000 2712 4 chanx_right_out[6]
port 93 nsew
rlabel metal3 s 19200 3000 20000 3120 4 chanx_right_out[7]
port 94 nsew
rlabel metal3 s 19200 3544 20000 3664 4 chanx_right_out[8]
port 95 nsew
rlabel metal3 s 19200 3952 20000 4072 4 chanx_right_out[9]
port 96 nsew
rlabel metal2 s 6642 0 6698 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
port 97 nsew
rlabel metal2 s 7102 0 7158 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
port 98 nsew
rlabel metal2 s 7654 0 7710 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
port 99 nsew
rlabel metal2 s 8114 0 8170 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
port 100 nsew
rlabel metal2 s 8666 0 8722 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
port 101 nsew
rlabel metal2 s 9126 0 9182 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
port 102 nsew
rlabel metal2 s 9678 0 9734 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
port 103 nsew
rlabel metal2 s 10138 0 10194 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
port 104 nsew
rlabel metal2 s 10598 0 10654 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
port 105 nsew
rlabel metal2 s 11150 0 11206 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
port 106 nsew
rlabel metal2 s 11610 0 11666 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
port 107 nsew
rlabel metal2 s 12162 0 12218 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
port 108 nsew
rlabel metal2 s 12622 0 12678 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
port 109 nsew
rlabel metal2 s 13174 0 13230 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
port 110 nsew
rlabel metal2 s 13634 0 13690 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
port 111 nsew
rlabel metal2 s 14094 0 14150 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
port 112 nsew
rlabel metal2 s 14646 0 14702 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
port 113 nsew
rlabel metal2 s 15106 0 15162 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
port 114 nsew
rlabel metal2 s 15658 0 15714 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
port 115 nsew
rlabel metal2 s 16118 0 16174 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
port 116 nsew
rlabel metal2 s 16670 0 16726 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
port 117 nsew
rlabel metal2 s 17130 0 17186 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
port 118 nsew
rlabel metal2 s 17590 0 17646 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
port 119 nsew
rlabel metal2 s 18142 0 18198 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
port 120 nsew
rlabel metal2 s 18602 0 18658 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
port 121 nsew
rlabel metal2 s 19154 0 19210 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
port 122 nsew
rlabel metal2 s 19614 0 19670 800 4 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
port 123 nsew
rlabel metal2 s 8022 16200 8078 17000 4 prog_clk_0_N_in
port 124 nsew
rlabel metal3 s 0 144 800 264 4 prog_clk_0_W_out
port 125 nsew
rlabel metal2 s 8666 16200 8722 17000 4 top_width_0_height_0__pin_0_
port 126 nsew
rlabel metal2 s 11886 16200 11942 17000 4 top_width_0_height_0__pin_10_
port 127 nsew
rlabel metal2 s 14462 16200 14518 17000 4 top_width_0_height_0__pin_11_lower
port 128 nsew
rlabel metal2 s 3514 16200 3570 17000 4 top_width_0_height_0__pin_11_upper
port 129 nsew
rlabel metal2 s 12530 16200 12586 17000 4 top_width_0_height_0__pin_12_
port 130 nsew
rlabel metal2 s 15106 16200 15162 17000 4 top_width_0_height_0__pin_13_lower
port 131 nsew
rlabel metal2 s 4158 16200 4214 17000 4 top_width_0_height_0__pin_13_upper
port 132 nsew
rlabel metal2 s 13174 16200 13230 17000 4 top_width_0_height_0__pin_14_
port 133 nsew
rlabel metal2 s 15750 16200 15806 17000 4 top_width_0_height_0__pin_15_lower
port 134 nsew
rlabel metal2 s 4802 16200 4858 17000 4 top_width_0_height_0__pin_15_upper
port 135 nsew
rlabel metal2 s 13818 16200 13874 17000 4 top_width_0_height_0__pin_16_
port 136 nsew
rlabel metal2 s 16394 16200 16450 17000 4 top_width_0_height_0__pin_17_lower
port 137 nsew
rlabel metal2 s 5446 16200 5502 17000 4 top_width_0_height_0__pin_17_upper
port 138 nsew
rlabel metal2 s 17038 16200 17094 17000 4 top_width_0_height_0__pin_1_lower
port 139 nsew
rlabel metal2 s 294 16200 350 17000 4 top_width_0_height_0__pin_1_upper
port 140 nsew
rlabel metal2 s 9310 16200 9366 17000 4 top_width_0_height_0__pin_2_
port 141 nsew
rlabel metal2 s 17682 16200 17738 17000 4 top_width_0_height_0__pin_3_lower
port 142 nsew
rlabel metal2 s 938 16200 994 17000 4 top_width_0_height_0__pin_3_upper
port 143 nsew
rlabel metal2 s 9954 16200 10010 17000 4 top_width_0_height_0__pin_4_
port 144 nsew
rlabel metal2 s 18326 16200 18382 17000 4 top_width_0_height_0__pin_5_lower
port 145 nsew
rlabel metal2 s 1582 16200 1638 17000 4 top_width_0_height_0__pin_5_upper
port 146 nsew
rlabel metal2 s 10598 16200 10654 17000 4 top_width_0_height_0__pin_6_
port 147 nsew
rlabel metal2 s 18970 16200 19026 17000 4 top_width_0_height_0__pin_7_lower
port 148 nsew
rlabel metal2 s 2226 16200 2282 17000 4 top_width_0_height_0__pin_7_upper
port 149 nsew
rlabel metal2 s 11242 16200 11298 17000 4 top_width_0_height_0__pin_8_
port 150 nsew
rlabel metal2 s 19614 16200 19670 17000 4 top_width_0_height_0__pin_9_lower
port 151 nsew
rlabel metal2 s 2870 16200 2926 17000 4 top_width_0_height_0__pin_9_upper
port 152 nsew
rlabel metal4 s 3909 2128 4229 14736 4 VPWR
port 153 nsew
rlabel metal4 s 6875 2128 7195 14736 4 VGND
port 154 nsew
<< properties >>
string FIXED_BBOX 0 0 20000 17000
string GDS_FILE /ef/openfpga/openlane/runs/cbx_1__0_/results/magic/cbx_1__0_.gds
string GDS_END 872146
string GDS_START 98316
<< end >>
