* NGSPICE file created from sb_1__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_dfxbp_1 abstract view
.subckt scs8hd_dfxbp_1 CLK D Q QN vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_mux2_1 abstract view
.subckt scs8hd_mux2_1 A0 A1 S X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

.subckt sb_1__1_ bottom_left_grid_pin_34_ bottom_left_grid_pin_35_ bottom_left_grid_pin_36_
+ bottom_left_grid_pin_37_ bottom_left_grid_pin_38_ bottom_left_grid_pin_39_ bottom_left_grid_pin_40_
+ bottom_left_grid_pin_41_ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10]
+ chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15]
+ chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10]
+ chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15]
+ chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in[0] chanx_right_in[10]
+ chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15]
+ chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9]
+ chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13]
+ chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17]
+ chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12]
+ chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17]
+ chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17]
+ chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] left_top_grid_pin_42_ left_top_grid_pin_43_ left_top_grid_pin_44_
+ left_top_grid_pin_45_ left_top_grid_pin_46_ left_top_grid_pin_47_ left_top_grid_pin_48_
+ left_top_grid_pin_49_ prog_clk right_top_grid_pin_42_ right_top_grid_pin_43_ right_top_grid_pin_44_
+ right_top_grid_pin_45_ right_top_grid_pin_46_ right_top_grid_pin_47_ right_top_grid_pin_48_
+ right_top_grid_pin_49_ top_left_grid_pin_34_ top_left_grid_pin_35_ top_left_grid_pin_36_
+ top_left_grid_pin_37_ top_left_grid_pin_38_ top_left_grid_pin_39_ top_left_grid_pin_40_
+ top_left_grid_pin_41_ vpwr vgnd
XFILLER_7_7 vgnd vpwr scs8hd_decap_3
Xmem_right_track_2.scs8hd_dfxbp_1_3_ prog_clk mux_right_track_2.mux_l3_in_0_/S mux_right_track_2.mux_l4_in_0_/S
+ mem_right_track_2.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_0.mux_l2_in_3__A0 _029_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_7__S mux_top_track_4.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_25.scs8hd_buf_4_0_ mux_bottom_track_25.mux_l4_in_0_/X _103_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_13_111 vpwr vgnd scs8hd_fill_2
XFILLER_42_40 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_2__S mux_top_track_16.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_34 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.mux_l1_in_1_ chanx_right_in[11] chanx_right_in[4] mux_bottom_track_3.mux_l1_in_4_/S
+ mux_bottom_track_3.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_36_247 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l3_in_0__A0 mux_right_track_2.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l4_in_1__A1 mux_left_track_5.mux_l3_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l3_in_0__A1 mux_left_track_25.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_258 vpwr vgnd scs8hd_fill_2
XFILLER_27_236 vpwr vgnd scs8hd_fill_2
XFILLER_27_225 vgnd vpwr scs8hd_decap_4
XFILLER_6_118 vpwr vgnd scs8hd_fill_2
XFILLER_12_10 vpwr vgnd scs8hd_fill_2
XFILLER_12_32 vpwr vgnd scs8hd_fill_2
XFILLER_33_239 vgnd vpwr scs8hd_decap_3
XANTENNA__124__A chany_bottom_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_5_140 vpwr vgnd scs8hd_fill_2
XFILLER_5_173 vgnd vpwr scs8hd_decap_4
XFILLER_24_228 vpwr vgnd scs8hd_fill_2
XFILLER_24_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0__A1 chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_23_261 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.mux_l1_in_0__A0 top_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
XFILLER_15_217 vgnd vpwr scs8hd_fill_1
XFILLER_15_239 vpwr vgnd scs8hd_fill_2
X_131_ _131_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
X_062_ chanx_right_in[12] chanx_left_out[13] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_5.mux_l5_in_0__A1 mux_left_track_5.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_33.mux_l1_in_2__A1 chany_bottom_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_2_154 vpwr vgnd scs8hd_fill_2
XFILLER_2_110 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_3__S mux_bottom_track_3.mux_l1_in_4_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l3_in_0__S mux_bottom_track_1.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__119__A _119_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__D mux_bottom_track_5.mux_l2_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_2__A1 right_top_grid_pin_45_ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_1.mux_l2_in_0_/S mux_left_track_1.mux_l3_in_1_/S
+ mem_left_track_1.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_34_41 vpwr vgnd scs8hd_fill_2
XFILLER_11_220 vpwr vgnd scs8hd_fill_2
XFILLER_11_264 vpwr vgnd scs8hd_fill_2
X_114_ _114_/A chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
X_045_ _045_/HI _045_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_track_24.mux_l2_in_3__S mux_right_track_24.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_19 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_3.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_track_3.mux_l3_in_1_/S mux_bottom_track_3.mux_l4_in_0_/S
+ mem_bottom_track_3.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_25.mux_l3_in_0__S mux_bottom_track_25.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_0_ chany_top_in[17] chany_top_in[8] mux_bottom_track_17.mux_l1_in_0_/S
+ mux_bottom_track_17.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_33.mux_l2_in_1__A1 mux_left_track_33.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0__S mux_left_track_17.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_76 vpwr vgnd scs8hd_fill_2
XFILLER_20_32 vpwr vgnd scs8hd_fill_2
XFILLER_20_21 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_2__D mux_right_track_16.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_194 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_4__A1 chany_bottom_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_6_23 vpwr vgnd scs8hd_fill_2
XANTENNA__132__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l3_in_0__S mux_right_track_16.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
X_028_ _028_/HI _028_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_track_0.mux_l1_in_1__S mux_right_track_0.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_33.scs8hd_buf_4_0__A mux_left_track_33.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l2_in_1__A1 mux_right_track_2.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_33.scs8hd_buf_4_0_ mux_bottom_track_33.mux_l3_in_0_/X _099_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_25_175 vpwr vgnd scs8hd_fill_2
XFILLER_25_153 vgnd vpwr scs8hd_decap_3
XFILLER_31_53 vpwr vgnd scs8hd_fill_2
XFILLER_15_76 vpwr vgnd scs8hd_fill_2
XFILLER_15_98 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_1__A0 chanx_right_in[11] vgnd vpwr scs8hd_diode_2
XANTENNA__127__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_123 vgnd vpwr scs8hd_decap_3
XFILLER_31_101 vpwr vgnd scs8hd_fill_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_120 vpwr vgnd scs8hd_fill_2
XFILLER_16_142 vpwr vgnd scs8hd_fill_2
XFILLER_16_186 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_1__S mux_top_track_0.mux_l2_in_2_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_33.mux_l3_in_0__A1 mux_left_track_33.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_245 vgnd vpwr scs8hd_decap_8
XFILLER_22_145 vpwr vgnd scs8hd_fill_2
XFILLER_22_112 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l2_in_2__A0 left_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_2.mux_l2_in_0_/S mux_right_track_2.mux_l3_in_0_/S
+ mem_right_track_2.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_0.mux_l2_in_3__A1 chanx_left_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_26_97 vgnd vpwr scs8hd_decap_3
XFILLER_26_86 vgnd vpwr scs8hd_decap_4
XFILLER_42_63 vgnd vpwr scs8hd_decap_4
XFILLER_9_149 vpwr vgnd scs8hd_fill_2
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.mux_l1_in_0_ chany_top_in[13] chany_top_in[4] mux_bottom_track_3.mux_l1_in_4_/S
+ mux_bottom_track_3.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_36_226 vpwr vgnd scs8hd_fill_2
XFILLER_36_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l3_in_0__A1 mux_right_track_2.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_3__A0 bottom_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__D mux_top_track_8.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_160 vpwr vgnd scs8hd_fill_2
XFILLER_35_270 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_3.mux_l2_in_0__A0 mux_bottom_track_3.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_10_115 vpwr vgnd scs8hd_fill_2
XFILLER_12_77 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_37_30 vpwr vgnd scs8hd_fill_2
XFILLER_33_218 vpwr vgnd scs8hd_fill_2
XFILLER_18_215 vgnd vpwr scs8hd_decap_4
XFILLER_18_204 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_5.mux_l4_in_1__S mux_bottom_track_5.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_41_262 vgnd vpwr scs8hd_decap_12
XFILLER_41_251 vpwr vgnd scs8hd_fill_2
XFILLER_41_240 vpwr vgnd scs8hd_fill_2
XFILLER_26_270 vgnd vpwr scs8hd_decap_4
XFILLER_5_152 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l3_in_1__A0 mux_left_track_9.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_270 vpwr vgnd scs8hd_fill_2
XFILLER_32_251 vpwr vgnd scs8hd_fill_2
X_130_ chany_bottom_in[4] chany_top_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_23_240 vpwr vgnd scs8hd_fill_2
XFILLER_23_54 vgnd vpwr scs8hd_decap_4
XFILLER_23_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0__A1 top_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
X_061_ chanx_right_in[13] chanx_left_out[14] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_17.mux_l2_in_3__S mux_left_track_17.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_2__A0 chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_6__A0 left_top_grid_pin_48_ vgnd vpwr scs8hd_diode_2
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XANTENNA__135__A _135_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_56 vgnd vpwr scs8hd_decap_3
XFILLER_9_78 vpwr vgnd scs8hd_fill_2
XFILLER_14_251 vpwr vgnd scs8hd_fill_2
XFILLER_14_262 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_4__S mux_right_track_0.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_9.scs8hd_dfxbp_1_3_ prog_clk mux_left_track_9.mux_l3_in_1_/S mux_left_track_9.mux_l4_in_0_/S
+ mem_left_track_9.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_17.mux_l4_in_0__S mux_bottom_track_17.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_2__S mux_left_track_1.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
Xmem_left_track_1.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_1.mux_l1_in_0_/S mux_left_track_1.mux_l2_in_0_/S
+ mem_left_track_1.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_18_98 vpwr vgnd scs8hd_fill_2
XFILLER_34_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l4_in_0__A0 mux_left_track_9.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
X_113_ _113_/A chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_7_214 vgnd vpwr scs8hd_fill_1
XFILLER_11_232 vpwr vgnd scs8hd_fill_2
XFILLER_11_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_4.mux_l2_in_2__S mux_right_track_4.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_24.mux_l1_in_0__S mux_top_track_24.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
X_044_ _044_/HI _044_/LO vgnd vpwr scs8hd_conb_1
XFILLER_38_107 vgnd vpwr scs8hd_decap_3
XFILLER_15_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l3_in_0__S mux_left_track_5.mux_l3_in_3_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_3.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_3.mux_l2_in_3_/S mux_bottom_track_3.mux_l3_in_1_/S
+ mem_bottom_track_3.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XFILLER_37_162 vpwr vgnd scs8hd_fill_2
XFILLER_37_140 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.mux_l3_in_1__A0 mux_bottom_track_1.mux_l2_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__D mux_top_track_24.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l3_in_0__S mux_right_track_8.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_88 vpwr vgnd scs8hd_fill_2
XFILLER_4_228 vpwr vgnd scs8hd_fill_2
XFILLER_29_97 vpwr vgnd scs8hd_fill_2
XFILLER_29_53 vpwr vgnd scs8hd_fill_2
XFILLER_28_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l3_in_2__S mux_top_track_4.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_28_173 vpwr vgnd scs8hd_fill_2
XFILLER_19_184 vgnd vpwr scs8hd_decap_3
XFILLER_19_173 vgnd vpwr scs8hd_decap_4
XFILLER_34_176 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__D mux_bottom_track_25.mux_l2_in_3_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l4_in_0__S mux_top_track_8.mux_l4_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_40_124 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_25_187 vpwr vgnd scs8hd_fill_2
XFILLER_25_132 vpwr vgnd scs8hd_fill_2
XFILLER_15_11 vgnd vpwr scs8hd_decap_3
XFILLER_40_168 vpwr vgnd scs8hd_fill_2
XFILLER_40_146 vgnd vpwr scs8hd_decap_4
XFILLER_31_98 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__D mux_bottom_track_5.mux_l5_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_231 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_3_ _035_/HI chanx_left_in[16] mux_right_track_8.mux_l2_in_1_/S
+ mux_right_track_8.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_3.mux_l1_in_1__A1 chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_31_179 vpwr vgnd scs8hd_fill_2
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l4_in_0__A0 mux_bottom_track_1.mux_l3_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_224 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l2_in_3_ _036_/HI chanx_left_in[12] mux_top_track_0.mux_l2_in_2_/S
+ mux_top_track_0.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_22_157 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l2_in_2__A1 chany_bottom_in[16] vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_2.mux_l1_in_4_/S mux_right_track_2.mux_l2_in_0_/S
+ mem_right_track_2.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_13_157 vpwr vgnd scs8hd_fill_2
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_33.mux_l1_in_1__S mux_left_track_33.mux_l1_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_32.mux_l2_in_1__S mux_right_track_32.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_3__A1 bottom_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
XFILLER_8_150 vgnd vpwr scs8hd_fill_1
XFILLER_12_190 vpwr vgnd scs8hd_fill_2
XFILLER_42_208 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0__A1 mux_bottom_track_3.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_10_138 vpwr vgnd scs8hd_fill_2
XFILLER_12_23 vpwr vgnd scs8hd_fill_2
XFILLER_12_45 vpwr vgnd scs8hd_fill_2
XFILLER_37_75 vgnd vpwr scs8hd_fill_1
XFILLER_37_53 vpwr vgnd scs8hd_fill_2
XFILLER_18_238 vpwr vgnd scs8hd_fill_2
XFILLER_41_274 vgnd vpwr scs8hd_decap_3
Xmux_top_track_0.mux_l1_in_4_ chanx_left_in[0] chany_bottom_in[12] mux_top_track_0.mux_l1_in_1_/S
+ mux_top_track_0.mux_l1_in_4_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_4.mux_l2_in_5__S mux_right_track_4.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_197 vgnd vpwr scs8hd_fill_1
XFILLER_38_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l3_in_3__S mux_left_track_5.mux_l3_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_32_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l3_in_1__A1 mux_left_track_9.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_8.mux_l4_in_0_ mux_right_track_8.mux_l3_in_1_/X mux_right_track_8.mux_l3_in_0_/X
+ mux_right_track_8.mux_l4_in_0_/S mux_right_track_8.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_274 vgnd vpwr scs8hd_decap_3
XFILLER_23_77 vpwr vgnd scs8hd_fill_2
X_060_ chanx_right_in[14] chanx_left_out[15] vgnd vpwr scs8hd_buf_2
Xmux_top_track_0.mux_l4_in_0_ mux_top_track_0.mux_l3_in_1_/X mux_top_track_0.mux_l3_in_0_/X
+ mux_top_track_0.mux_l4_in_0_/S mux_top_track_0.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_3_3 vgnd vpwr scs8hd_decap_3
XFILLER_2_145 vpwr vgnd scs8hd_fill_2
XFILLER_2_134 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_2__A1 mux_bottom_track_1.mux_l1_in_4_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0__S mux_top_track_16.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_6__A1 left_top_grid_pin_47_ vgnd vpwr scs8hd_diode_2
XFILLER_9_35 vpwr vgnd scs8hd_fill_2
XFILLER_14_274 vgnd vpwr scs8hd_fill_1
XFILLER_36_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_4.mux_l2_in_2__A0 right_top_grid_pin_45_ vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_9.mux_l2_in_1_/S mux_left_track_9.mux_l3_in_1_/S
+ mem_left_track_9.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_20_255 vpwr vgnd scs8hd_fill_2
XANTENNA__061__A chanx_right_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_18_88 vpwr vgnd scs8hd_fill_2
XFILLER_18_77 vpwr vgnd scs8hd_fill_2
Xmem_left_track_1.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_33.mux_l3_in_0_/S mux_left_track_1.mux_l1_in_0_/S
+ mem_left_track_1.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_34_87 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l4_in_0__A1 mux_left_track_9.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
X_043_ _043_/HI _043_/LO vgnd vpwr scs8hd_conb_1
X_112_ chany_top_in[2] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_3__D mux_bottom_track_9.mux_l3_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_119 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l3_in_1_ mux_right_track_8.mux_l2_in_3_/X mux_right_track_8.mux_l2_in_2_/X
+ mux_right_track_8.mux_l3_in_0_/S mux_right_track_8.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmem_bottom_track_3.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_3.mux_l1_in_4_/S mux_bottom_track_3.mux_l2_in_3_/S
+ mem_bottom_track_3.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_6_270 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l3_in_1_ mux_top_track_0.mux_l2_in_3_/X mux_top_track_0.mux_l2_in_2_/X
+ mux_top_track_0.mux_l3_in_1_/S mux_top_track_0.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_1.mux_l3_in_1__A1 mux_bottom_track_1.mux_l2_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA__056__A chanx_right_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_4_207 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_4.mux_l3_in_1__A0 mux_right_track_4.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l2_in_1__S mux_bottom_track_3.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_6_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__D mux_right_track_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2__S mux_bottom_track_9.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_31_66 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.mux_l2_in_1__S mux_left_track_25.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_243 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_2_ chanx_left_in[6] chany_bottom_in[16] mux_right_track_8.mux_l2_in_1_/S
+ mux_right_track_8.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_16_166 vgnd vpwr scs8hd_fill_1
XFILLER_31_169 vgnd vpwr scs8hd_fill_1
XFILLER_31_114 vpwr vgnd scs8hd_fill_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l4_in_0__A1 mux_bottom_track_1.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_24.mux_l3_in_1__S mux_right_track_24.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_2_ chanx_left_in[2] mux_top_track_0.mux_l1_in_4_/X mux_top_track_0.mux_l2_in_2_/S
+ mux_top_track_0.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_39_236 vgnd vpwr scs8hd_decap_8
XFILLER_39_203 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l1_in_1__A0 top_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l4_in_0__A0 mux_right_track_4.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_right_track_2.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_0.mux_l4_in_0_/S mux_right_track_2.mux_l1_in_4_/S
+ mem_right_track_2.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_26_55 vpwr vgnd scs8hd_fill_2
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_42_98 vgnd vpwr scs8hd_decap_3
XFILLER_21_191 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_3__S mux_top_track_16.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_206 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.scs8hd_buf_4_0_ mux_bottom_track_5.mux_l5_in_0_/X _113_/A vgnd
+ vpwr scs8hd_buf_1
XANTENNA_mux_left_track_3.mux_l1_in_0__S mux_left_track_3.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_4__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA__064__A chanx_right_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_12_57 vgnd vpwr scs8hd_fill_1
XFILLER_41_220 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_0.mux_l1_in_3__A0 chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_3_ chany_bottom_in[2] chanx_right_in[12] mux_top_track_0.mux_l1_in_1_/S
+ mux_top_track_0.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_2__S mux_top_track_2.mux_l1_in_3_/S vgnd vpwr scs8hd_diode_2
XFILLER_5_132 vpwr vgnd scs8hd_fill_2
XFILLER_5_165 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l2_in_0__A0 mux_top_track_2.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_261 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_4_91 vgnd vpwr scs8hd_fill_1
XANTENNA__059__A _059_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_23 vpwr vgnd scs8hd_fill_2
XFILLER_2_102 vpwr vgnd scs8hd_fill_2
XFILLER_9_14 vpwr vgnd scs8hd_fill_2
XFILLER_29_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_4.mux_l2_in_2__A1 right_top_grid_pin_44_ vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_9.mux_l1_in_0_/S mux_left_track_9.mux_l2_in_1_/S
+ mem_left_track_9.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__D mux_right_track_2.mux_l1_in_4_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_267 vpwr vgnd scs8hd_fill_2
XFILLER_20_234 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_2__A0 chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_18_56 vpwr vgnd scs8hd_fill_2
XFILLER_18_23 vpwr vgnd scs8hd_fill_2
XFILLER_18_12 vpwr vgnd scs8hd_fill_2
XFILLER_34_22 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_042_ _042_/HI _042_/LO vgnd vpwr scs8hd_conb_1
X_111_ _111_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_7_227 vgnd vpwr scs8hd_decap_4
XFILLER_7_238 vgnd vpwr scs8hd_decap_4
XFILLER_11_256 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__D mux_top_track_16.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l3_in_0_ mux_right_track_8.mux_l2_in_1_/X mux_right_track_8.mux_l2_in_0_/X
+ mux_right_track_8.mux_l3_in_0_/S mux_right_track_8.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_bottom_track_3.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_1.mux_l4_in_0_/S mux_bottom_track_3.mux_l1_in_4_/S
+ mem_bottom_track_3.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_37_197 vpwr vgnd scs8hd_fill_2
XFILLER_37_175 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_1_/S mux_top_track_0.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__072__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l3_in_1__S mux_left_track_17.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l3_in_1__A1 mux_right_track_4.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_32.mux_l1_in_1__S mux_top_track_32.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l3_in_1__A0 mux_top_track_0.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_7 vgnd vpwr scs8hd_fill_1
XFILLER_3_274 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_3.mux_l1_in_4__A0 chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_10_90 vpwr vgnd scs8hd_fill_2
XFILLER_34_189 vpwr vgnd scs8hd_fill_2
XFILLER_34_145 vpwr vgnd scs8hd_fill_2
XFILLER_34_134 vgnd vpwr scs8hd_fill_1
XFILLER_19_142 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_2__S mux_right_track_0.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l1_in_3__S mux_left_track_3.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l3_in_0__S mux_left_track_1.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_1__A0 chanx_right_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_40_137 vpwr vgnd scs8hd_fill_2
XANTENNA__067__A _067_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_35 vpwr vgnd scs8hd_fill_2
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_33.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__D mux_left_track_25.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_200 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.mux_l2_in_1_ chany_bottom_in[6] mux_right_track_8.mux_l1_in_2_/X
+ mux_right_track_8.mux_l2_in_1_/S mux_right_track_8.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_4.mux_l3_in_0__S mux_right_track_4.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_148 vpwr vgnd scs8hd_fill_2
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_1_ mux_top_track_0.mux_l1_in_3_/X mux_top_track_0.mux_l1_in_2_/X
+ mux_top_track_0.mux_l2_in_2_/S mux_top_track_0.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_39_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_11_3 vgnd vpwr scs8hd_fill_1
XFILLER_22_137 vpwr vgnd scs8hd_fill_2
XFILLER_22_104 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l4_in_0__A1 mux_right_track_4.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_1__A1 top_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1__A0 chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_26_78 vpwr vgnd scs8hd_fill_2
XFILLER_26_23 vpwr vgnd scs8hd_fill_2
XFILLER_26_12 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_3__A0 _046_/HI vgnd vpwr scs8hd_diode_2
XFILLER_13_115 vpwr vgnd scs8hd_fill_2
XFILLER_42_11 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.scs8hd_buf_4_0_ mux_left_track_9.mux_l4_in_0_/X _071_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_21_170 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l4_in_0__A0 mux_top_track_0.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l4_in_0__S mux_top_track_4.mux_l4_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_13_126 vpwr vgnd scs8hd_fill_2
XFILLER_3_38 vgnd vpwr scs8hd_decap_4
XFILLER_29_270 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_5.mux_l3_in_0__A0 mux_bottom_track_5.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__D mux_right_track_2.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_35_240 vpwr vgnd scs8hd_fill_2
XFILLER_27_229 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.mux_l1_in_2_ chany_bottom_in[3] right_top_grid_pin_46_ mux_right_track_8.mux_l1_in_2_/S
+ mux_right_track_8.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__080__A chanx_left_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_37_11 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l1_in_3__A1 chanx_right_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_41_232 vgnd vpwr scs8hd_decap_8
XFILLER_41_210 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_2_ chanx_right_in[2] chanx_right_in[1] mux_top_track_0.mux_l1_in_1_/S
+ mux_top_track_0.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_5_111 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.scs8hd_buf_4_0_ mux_top_track_2.mux_l4_in_0_/X _134_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_top_track_2.mux_l2_in_0__A1 mux_top_track_2.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XFILLER_32_210 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0__A0 mux_left_track_1.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_254 vgnd vpwr scs8hd_decap_4
XANTENNA__075__A _075_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_169 vpwr vgnd scs8hd_fill_2
XFILLER_2_158 vpwr vgnd scs8hd_fill_2
XFILLER_2_114 vgnd vpwr scs8hd_fill_1
XFILLER_9_48 vpwr vgnd scs8hd_fill_2
XFILLER_14_243 vgnd vpwr scs8hd_fill_1
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_25.mux_l2_in_3_ _045_/HI chanx_left_in[19] mux_bottom_track_25.mux_l2_in_3_/S
+ mux_bottom_track_25.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_1_180 vgnd vpwr scs8hd_fill_1
Xmem_left_track_9.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_5.mux_l5_in_0_/S mux_left_track_9.mux_l1_in_0_/S
+ mem_left_track_9.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_0.mux_l2_in_2__A1 mux_top_track_0.mux_l1_in_4_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_46 vgnd vpwr scs8hd_fill_1
XFILLER_34_45 vpwr vgnd scs8hd_fill_2
X_110_ chany_top_in[4] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_11_224 vpwr vgnd scs8hd_fill_2
XFILLER_7_217 vgnd vpwr scs8hd_fill_1
XFILLER_11_268 vpwr vgnd scs8hd_fill_2
X_041_ _041_/HI _041_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_24.mux_l2_in_1__S mux_top_track_24.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l3_in_3__S mux_right_track_4.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_4.mux_l2_in_7_ _034_/HI chanx_left_in[14] mux_right_track_4.mux_l2_in_0_/S
+ mux_right_track_4.mux_l2_in_7_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_5.mux_l4_in_1__S mux_left_track_5.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_37_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_2__A0 chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_1_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_20_36 vpwr vgnd scs8hd_fill_2
XFILLER_20_25 vpwr vgnd scs8hd_fill_2
XFILLER_29_67 vpwr vgnd scs8hd_fill_2
XFILLER_29_34 vpwr vgnd scs8hd_fill_2
XFILLER_28_198 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_3_231 vgnd vpwr scs8hd_fill_1
XFILLER_6_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_4__A1 bottom_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_3_ _049_/HI chanx_left_in[16] mux_bottom_track_9.mux_l2_in_3_/S
+ mux_bottom_track_9.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_0.mux_l3_in_1__A1 mux_top_track_0.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_168 vpwr vgnd scs8hd_fill_2
XFILLER_34_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_3__D mux_right_track_4.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_25_113 vgnd vpwr scs8hd_decap_3
XFILLER_25_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_1__A1 chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_40_127 vgnd vpwr scs8hd_fill_1
XANTENNA__083__A _083_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_179 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_25.mux_l4_in_0_ mux_bottom_track_25.mux_l3_in_1_/X mux_bottom_track_25.mux_l3_in_0_/X
+ mux_bottom_track_25.mux_l4_in_0_/S mux_bottom_track_25.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XFILLER_31_57 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_0_ mux_right_track_8.mux_l1_in_1_/X mux_right_track_8.mux_l1_in_0_/X
+ mux_right_track_8.mux_l2_in_1_/S mux_right_track_8.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_124 vpwr vgnd scs8hd_fill_2
XFILLER_16_146 vpwr vgnd scs8hd_fill_2
XFILLER_16_157 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l2_in_1__A0 chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_0_ mux_top_track_0.mux_l1_in_1_/X mux_top_track_0.mux_l1_in_0_/X
+ mux_top_track_0.mux_l2_in_2_/S mux_top_track_0.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_22_149 vpwr vgnd scs8hd_fill_2
XFILLER_7_92 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l1_in_1__A1 chany_top_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_38_271 vgnd vpwr scs8hd_decap_4
XANTENNA__078__A chanx_left_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l2_in_3__A1 chanx_left_in[13] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l4_in_0__A1 mux_top_track_0.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_67 vgnd vpwr scs8hd_fill_1
XFILLER_42_23 vpwr vgnd scs8hd_fill_2
XFILLER_3_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l3_in_0__A1 mux_bottom_track_5.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_120 vgnd vpwr scs8hd_decap_3
XFILLER_8_142 vpwr vgnd scs8hd_fill_2
XFILLER_8_164 vpwr vgnd scs8hd_fill_2
XFILLER_35_230 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_25.mux_l3_in_1_ mux_bottom_track_25.mux_l2_in_3_/X mux_bottom_track_25.mux_l2_in_2_/X
+ mux_bottom_track_25.mux_l3_in_1_/S mux_bottom_track_25.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_mux2_1
Xmux_right_track_8.mux_l1_in_1_ right_top_grid_pin_42_ chany_top_in[16] mux_right_track_8.mux_l1_in_2_/S
+ mux_right_track_8.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_8.mux_l3_in_0__A0 mux_right_track_8.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_9.mux_l4_in_0_ mux_bottom_track_9.mux_l3_in_1_/X mux_bottom_track_9.mux_l3_in_0_/X
+ mux_bottom_track_9.mux_l4_in_0_/S mux_bottom_track_9.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_9.mux_l2_in_0__S mux_bottom_track_9.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_78 vpwr vgnd scs8hd_fill_2
XFILLER_18_219 vgnd vpwr scs8hd_fill_1
XFILLER_41_255 vgnd vpwr scs8hd_decap_4
XFILLER_26_274 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.mux_l1_in_1_ top_left_grid_pin_40_ top_left_grid_pin_38_ mux_top_track_0.mux_l1_in_1_/S
+ mux_top_track_0.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A0 chany_top_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_17_274 vgnd vpwr scs8hd_decap_3
XFILLER_32_255 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0__A1 mux_left_track_1.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1__S mux_bottom_track_17.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_5__A0 chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vpwr vgnd scs8hd_fill_2
XFILLER_4_82 vgnd vpwr scs8hd_decap_3
XFILLER_23_266 vpwr vgnd scs8hd_fill_2
XANTENNA__091__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_58 vgnd vpwr scs8hd_fill_1
XFILLER_0_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_14_211 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.mux_l3_in_1__S mux_top_track_16.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_266 vpwr vgnd scs8hd_fill_2
XFILLER_13_80 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_25.mux_l2_in_2_ chanx_left_in[18] chanx_left_in[9] mux_bottom_track_25.mux_l2_in_3_/S
+ mux_bottom_track_25.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_0__S mux_right_track_2.mux_l1_in_4_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_9.mux_l3_in_1_ mux_bottom_track_9.mux_l2_in_3_/X mux_bottom_track_9.mux_l2_in_2_/X
+ mux_bottom_track_9.mux_l3_in_1_/S mux_bottom_track_9.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_18_36 vpwr vgnd scs8hd_fill_2
XFILLER_34_79 vpwr vgnd scs8hd_fill_2
XANTENNA__086__A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_11_203 vpwr vgnd scs8hd_fill_2
XFILLER_11_236 vpwr vgnd scs8hd_fill_2
X_040_ _040_/HI _040_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_2.mux_l2_in_0__S mux_top_track_2.mux_l2_in_2_/S vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l2_in_6_ chanx_left_in[5] chany_bottom_in[14] mux_right_track_4.mux_l2_in_0_/S
+ mux_right_track_4.mux_l2_in_6_/X vgnd vpwr scs8hd_mux2_1
XFILLER_6_262 vpwr vgnd scs8hd_fill_2
XFILLER_34_3 vgnd vpwr scs8hd_decap_4
XFILLER_37_166 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_2__A1 right_top_grid_pin_46_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1__S mux_top_track_8.mux_l1_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_29_57 vpwr vgnd scs8hd_fill_2
XFILLER_28_111 vpwr vgnd scs8hd_fill_2
XFILLER_28_177 vpwr vgnd scs8hd_fill_2
XFILLER_28_144 vpwr vgnd scs8hd_fill_2
XFILLER_3_254 vpwr vgnd scs8hd_fill_2
XFILLER_3_210 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_2_ chanx_left_in[11] chanx_left_in[6] mux_bottom_track_9.mux_l2_in_3_/S
+ mux_bottom_track_9.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_70 vpwr vgnd scs8hd_fill_2
XFILLER_19_177 vgnd vpwr scs8hd_fill_1
XFILLER_19_155 vgnd vpwr scs8hd_decap_3
XFILLER_25_158 vpwr vgnd scs8hd_fill_2
XFILLER_25_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__D mux_right_track_24.mux_l2_in_2_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_191 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_3__S mux_bottom_track_9.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_4__A0 chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_213 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.scs8hd_dfxbp_1_3_ prog_clk mux_right_track_16.mux_l3_in_0_/S mux_right_track_16.mux_l4_in_0_/S
+ mem_right_track_16.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_31_128 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l2_in_1__A1 mux_right_track_8.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_91 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_1__A0 top_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_30_161 vpwr vgnd scs8hd_fill_2
XFILLER_30_150 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_7_60 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_1__A0 chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1__A0 right_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
XANTENNA__094__A _094_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_79 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A0 chany_top_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_8_154 vpwr vgnd scs8hd_fill_2
XFILLER_12_194 vpwr vgnd scs8hd_fill_2
XFILLER_16_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_2.mux_l1_in_3__S mux_right_track_2.mux_l1_in_4_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_187 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l3_in_0__S mux_right_track_0.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_3__A0 _038_/HI vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_25.mux_l3_in_0_ mux_bottom_track_25.mux_l2_in_1_/X mux_bottom_track_25.mux_l2_in_0_/X
+ mux_bottom_track_25.mux_l3_in_1_/S mux_bottom_track_25.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XANTENNA_mux_bottom_track_17.scs8hd_buf_4_0__A mux_bottom_track_17.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l2_in_1__S mux_left_track_3.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_0_ chany_top_in[6] chany_top_in[3] mux_right_track_8.mux_l1_in_2_/S
+ mux_right_track_8.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_12_27 vpwr vgnd scs8hd_fill_2
XFILLER_12_49 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__D mux_right_track_8.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l3_in_0__A1 mux_right_track_8.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA__089__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l3_in_0__A0 mux_top_track_4.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_ top_left_grid_pin_36_ top_left_grid_pin_34_ mux_top_track_0.mux_l1_in_1_/S
+ mux_top_track_0.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_2.mux_l2_in_3__S mux_top_track_2.mux_l2_in_2_/S vgnd vpwr scs8hd_diode_2
XFILLER_5_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_2__S mux_left_track_9.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l4_in_0__S mux_top_track_0.mux_l4_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A1 chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_32_234 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A0 mux_bottom_track_9.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0__A0 mux_right_track_16.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_5__A1 chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_23_201 vpwr vgnd scs8hd_fill_2
XFILLER_2_138 vpwr vgnd scs8hd_fill_2
XFILLER_2_149 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_25.mux_l2_in_1_ bottom_left_grid_pin_40_ mux_bottom_track_25.mux_l1_in_2_/X
+ mux_bottom_track_25.mux_l2_in_3_/S mux_bottom_track_25.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_mux2_1
XFILLER_1_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l1_in_0__A0 chany_top_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_20_204 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l3_in_0_ mux_bottom_track_9.mux_l2_in_1_/X mux_bottom_track_9.mux_l2_in_0_/X
+ mux_bottom_track_9.mux_l3_in_1_/S mux_bottom_track_9.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_58 vpwr vgnd scs8hd_fill_2
XFILLER_11_248 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.scs8hd_dfxbp_1_3_ prog_clk mux_left_track_17.mux_l3_in_1_/S mux_left_track_17.mux_l4_in_0_/S
+ mem_left_track_17.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_track_4.mux_l2_in_5_ chany_bottom_in[7] chany_bottom_in[5] mux_right_track_4.mux_l2_in_0_/S
+ mux_right_track_4.mux_l2_in_5_/X vgnd vpwr scs8hd_mux2_1
XFILLER_6_241 vgnd vpwr scs8hd_decap_4
XFILLER_6_274 vgnd vpwr scs8hd_fill_1
XFILLER_27_3 vgnd vpwr scs8hd_decap_4
X_099_ _099_/A chany_bottom_out[16] vgnd vpwr scs8hd_buf_2
XFILLER_37_101 vgnd vpwr scs8hd_decap_3
XFILLER_1_40 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l1_in_2__A0 chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l2_in_3_ _037_/HI chanx_left_in[17] mux_top_track_16.mux_l2_in_0_/S
+ mux_top_track_16.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_20_49 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_4__A0 bottom_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_25.mux_l1_in_2_ bottom_left_grid_pin_36_ chanx_right_in[18] mux_bottom_track_25.mux_l1_in_0_/S
+ mux_bottom_track_25.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__097__A chany_top_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_3_266 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_1_ bottom_left_grid_pin_38_ mux_bottom_track_9.mux_l1_in_2_/X
+ mux_bottom_track_9.mux_l2_in_3_/S mux_bottom_track_9.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_93 vgnd vpwr scs8hd_decap_3
XFILLER_34_137 vpwr vgnd scs8hd_fill_2
XFILLER_19_189 vpwr vgnd scs8hd_fill_2
XFILLER_19_123 vgnd vpwr scs8hd_decap_4
XFILLER_19_112 vpwr vgnd scs8hd_fill_2
XFILLER_35_90 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_24.mux_l1_in_1__A0 right_top_grid_pin_44_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l1_in_0__A0 chanx_right_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_31_26 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_16.mux_l2_in_0_/S mux_right_track_16.mux_l3_in_0_/S
+ mem_right_track_16.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_2.mux_l1_in_4__A1 chany_bottom_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_0_269 vpwr vgnd scs8hd_fill_2
XFILLER_0_258 vpwr vgnd scs8hd_fill_2
XFILLER_0_247 vgnd vpwr scs8hd_fill_1
XFILLER_0_203 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l1_in_4__A0 left_top_grid_pin_44_ vgnd vpwr scs8hd_diode_2
XFILLER_31_118 vpwr vgnd scs8hd_fill_2
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_4.mux_l4_in_1__S mux_right_track_4.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_1__A1 top_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
XFILLER_39_207 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l2_in_1__A0 mux_left_track_3.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1__A0 chanx_right_in[15] vgnd vpwr scs8hd_diode_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_2__D mux_bottom_track_33.mux_l2_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l3_in_3__A0 mux_bottom_track_5.mux_l2_in_7_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1__A1 chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_42_47 vgnd vpwr scs8hd_decap_12
XFILLER_42_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_1__A1 chany_top_in[17] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_2_ bottom_left_grid_pin_34_ chanx_right_in[16] mux_bottom_track_9.mux_l1_in_2_/S
+ mux_bottom_track_9.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_13_107 vpwr vgnd scs8hd_fill_2
XFILLER_21_195 vpwr vgnd scs8hd_fill_2
XFILLER_21_184 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A1 chany_top_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_29_240 vpwr vgnd scs8hd_fill_2
XFILLER_12_173 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l4_in_0_ mux_top_track_16.mux_l3_in_1_/X mux_top_track_16.mux_l3_in_0_/X
+ mux_top_track_16.mux_l4_in_0_/S mux_top_track_16.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_24.mux_l2_in_0__A0 mux_right_track_24.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_81 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_2.mux_l2_in_3__A1 chanx_left_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_35_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_254 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_3__A0 _050_/HI vgnd vpwr scs8hd_diode_2
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_26_254 vpwr vgnd scs8hd_fill_2
XFILLER_26_210 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l3_in_0__A1 mux_top_track_4.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l3_in_0__A0 mux_left_track_3.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_5.scs8hd_buf_4_0__A mux_bottom_track_5.mux_l5_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0__A0 mux_top_track_16.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_3.mux_l2_in_3_ _053_/HI left_top_grid_pin_49_ mux_left_track_3.mux_l2_in_2_/S
+ mux_left_track_3.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_5_136 vpwr vgnd scs8hd_fill_2
XFILLER_5_169 vpwr vgnd scs8hd_fill_2
XFILLER_17_221 vpwr vgnd scs8hd_fill_2
XFILLER_27_91 vpwr vgnd scs8hd_fill_2
XFILLER_17_254 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_2__S mux_bottom_track_1.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A1 mux_bottom_track_9.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_4.scs8hd_buf_4_0_ mux_right_track_4.mux_l5_in_0_/X _093_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_right_track_16.mux_l2_in_0__A1 mux_right_track_16.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l3_in_3_ mux_right_track_4.mux_l2_in_7_/X mux_right_track_4.mux_l2_in_6_/X
+ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l3_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_51 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__D mux_left_track_1.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_224 vpwr vgnd scs8hd_fill_2
XFILLER_23_27 vpwr vgnd scs8hd_fill_2
XFILLER_2_106 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l3_in_1_ mux_top_track_16.mux_l2_in_3_/X mux_top_track_16.mux_l2_in_2_/X
+ mux_top_track_16.mux_l3_in_0_/S mux_top_track_16.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_33.mux_l3_in_0__S ccff_tail vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0__S mux_bottom_track_5.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_18 vpwr vgnd scs8hd_fill_2
XFILLER_14_224 vpwr vgnd scs8hd_fill_2
XFILLER_14_235 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_25.mux_l2_in_0_ mux_bottom_track_25.mux_l1_in_1_/X mux_bottom_track_25.mux_l1_in_0_/X
+ mux_bottom_track_25.mux_l2_in_3_/S mux_bottom_track_25.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XFILLER_13_60 vgnd vpwr scs8hd_fill_1
XFILLER_1_172 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l1_in_0__A1 chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_20_238 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l2_in_7_ _048_/HI chanx_left_in[14] mux_bottom_track_5.mux_l2_in_1_/S
+ mux_bottom_track_5.mux_l2_in_7_/X vgnd vpwr scs8hd_mux2_1
XFILLER_9_261 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_25.mux_l1_in_2__S mux_bottom_track_25.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_18_27 vpwr vgnd scs8hd_fill_2
Xmux_left_track_3.mux_l1_in_4_ left_top_grid_pin_45_ left_top_grid_pin_43_ mux_left_track_3.mux_l1_in_0_/S
+ mux_left_track_3.mux_l1_in_4_/X vgnd vpwr scs8hd_mux2_1
Xmem_left_track_17.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_17.mux_l2_in_1_/S mux_left_track_17.mux_l3_in_1_/S
+ mem_left_track_17.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_24_70 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_32.mux_l1_in_1__A0 right_top_grid_pin_49_ vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l2_in_4_ right_top_grid_pin_49_ right_top_grid_pin_48_ mux_right_track_4.mux_l2_in_0_/S
+ mux_right_track_4.mux_l2_in_4_/X vgnd vpwr scs8hd_mux2_1
XFILLER_40_91 vgnd vpwr scs8hd_fill_1
X_098_ chany_top_in[16] chany_bottom_out[17] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_16.mux_l1_in_2__S mux_right_track_16.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l1_in_2__A1 chanx_right_in[13] vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l2_in_2_ chanx_left_in[8] chanx_left_in[7] mux_top_track_16.mux_l2_in_0_/S
+ mux_top_track_16.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
Xmux_left_track_3.mux_l4_in_0_ mux_left_track_3.mux_l3_in_1_/X mux_left_track_3.mux_l3_in_0_/X
+ mux_left_track_3.mux_l4_in_0_/S mux_left_track_3.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_20_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_4__A1 bottom_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XFILLER_28_135 vpwr vgnd scs8hd_fill_2
XFILLER_28_102 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_25.mux_l1_in_1_ chanx_right_in[9] chanx_right_in[0] mux_bottom_track_25.mux_l1_in_0_/S
+ mux_bottom_track_25.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_3_234 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_24.mux_l1_in_1__A0 chanx_right_in[18] vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l5_in_0_ mux_right_track_4.mux_l4_in_1_/X mux_right_track_4.mux_l4_in_0_/X
+ mux_right_track_4.mux_l5_in_0_/S mux_right_track_4.mux_l5_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_track_9.mux_l2_in_0_ mux_bottom_track_9.mux_l1_in_1_/X mux_bottom_track_9.mux_l1_in_0_/X
+ mux_bottom_track_9.mux_l2_in_3_/S mux_bottom_track_9.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_149 vpwr vgnd scs8hd_fill_2
XFILLER_19_92 vpwr vgnd scs8hd_fill_2
XFILLER_42_182 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_32.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_24.mux_l1_in_1__A1 chany_top_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_33_182 vgnd vpwr scs8hd_fill_1
XFILLER_33_160 vgnd vpwr scs8hd_decap_4
XFILLER_25_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_33.mux_l1_in_0__A1 chany_top_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_15_39 vgnd vpwr scs8hd_decap_3
Xmem_right_track_16.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_16.mux_l1_in_0_/S mux_right_track_16.mux_l2_in_0_/S
+ mem_right_track_16.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_1.mux_l1_in_4__A1 left_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_32.mux_l2_in_0__A0 mux_right_track_32.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_138 vpwr vgnd scs8hd_fill_2
XFILLER_24_182 vpwr vgnd scs8hd_fill_2
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A0 chany_top_in[12] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l2_in_1__A1 mux_left_track_3.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1__A1 chanx_right_in[8] vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.mux_l3_in_1_ mux_left_track_3.mux_l2_in_3_/X mux_left_track_3.mux_l2_in_2_/X
+ mux_left_track_3.mux_l3_in_1_/S mux_left_track_3.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_22_108 vpwr vgnd scs8hd_fill_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_5.mux_l3_in_3__A1 mux_bottom_track_5.mux_l2_in_6_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_193 vpwr vgnd scs8hd_fill_2
XFILLER_30_185 vpwr vgnd scs8hd_fill_2
XFILLER_38_241 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__D mux_left_track_3.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_26_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_24.mux_l2_in_0__A0 mux_top_track_24.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_59 vgnd vpwr scs8hd_decap_3
Xmux_right_track_4.mux_l4_in_1_ mux_right_track_4.mux_l3_in_3_/X mux_right_track_4.mux_l3_in_2_/X
+ mux_right_track_4.mux_l4_in_0_/S mux_right_track_4.mux_l4_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_21_174 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_1_ chanx_right_in[6] chanx_right_in[3] mux_bottom_track_9.mux_l1_in_2_/S
+ mux_bottom_track_9.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_13_119 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_5.mux_l2_in_3__S mux_bottom_track_5.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l4_in_0__S mux_bottom_track_3.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_93 vpwr vgnd scs8hd_fill_2
XFILLER_32_70 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l2_in_0__A1 mux_right_track_24.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1__A0 chanx_right_in[11] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_3__A1 left_top_grid_pin_48_ vgnd vpwr scs8hd_diode_2
XFILLER_35_266 vpwr vgnd scs8hd_fill_2
XFILLER_37_26 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l3_in_1__S mux_bottom_track_9.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_41_214 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_3.mux_l3_in_0__A1 mux_left_track_3.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_266 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.scs8hd_buf_4_0__A mux_top_track_0.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__D mux_bottom_track_9.mux_l4_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l4_in_0__S mux_left_track_25.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_115 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l2_in_0__A1 mux_top_track_16.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_3.mux_l2_in_2_ left_top_grid_pin_47_ mux_left_track_3.mux_l1_in_4_/X
+ mux_left_track_3.mux_l2_in_2_/S mux_left_track_3.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_5_148 vpwr vgnd scs8hd_fill_2
XFILLER_27_70 vgnd vpwr scs8hd_decap_4
XFILLER_17_211 vpwr vgnd scs8hd_fill_2
XFILLER_32_203 vgnd vpwr scs8hd_decap_4
XFILLER_17_266 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l3_in_2_ mux_right_track_4.mux_l2_in_5_/X mux_right_track_4.mux_l2_in_4_/X
+ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l3_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_236 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_2__S mux_bottom_track_17.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_top_track_4.scs8hd_dfxbp_1_4_ prog_clk mux_top_track_4.mux_l4_in_0_/S mux_top_track_4.mux_l5_in_0_/S
+ mem_top_track_4.scs8hd_dfxbp_1_4_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_23_258 vgnd vpwr scs8hd_fill_1
Xmux_top_track_16.mux_l3_in_0_ mux_top_track_16.mux_l2_in_1_/X mux_top_track_16.mux_l2_in_0_/X
+ mux_top_track_16.mux_l3_in_0_/S mux_top_track_16.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_17.mux_l2_in_2__A0 chanx_left_in[15] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0__A0 mux_top_track_8.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_203 vpwr vgnd scs8hd_fill_2
XFILLER_14_247 vpwr vgnd scs8hd_fill_2
XFILLER_14_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l2_in_1__S mux_right_track_2.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_5.mux_l2_in_6_ chanx_left_in[7] chanx_left_in[5] mux_bottom_track_5.mux_l2_in_1_/S
+ mux_bottom_track_5.mux_l2_in_6_/X vgnd vpwr scs8hd_mux2_1
XFILLER_9_273 vpwr vgnd scs8hd_fill_2
XFILLER_34_27 vpwr vgnd scs8hd_fill_2
Xmux_left_track_3.mux_l1_in_3_ chany_bottom_in[13] chany_bottom_in[4] mux_left_track_3.mux_l1_in_0_/S
+ mux_left_track_3.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
Xmem_right_track_0.scs8hd_dfxbp_1_3_ prog_clk mux_right_track_0.mux_l3_in_0_/S mux_right_track_0.mux_l4_in_0_/S
+ mem_right_track_0.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_32.mux_l1_in_1__A0 chanx_right_in[10] vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l2_in_3_ _030_/HI chanx_left_in[17] mux_right_track_16.mux_l2_in_0_/S
+ mux_right_track_16.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
Xmem_left_track_17.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_17.mux_l1_in_0_/S mux_left_track_17.mux_l2_in_1_/S
+ mem_left_track_17.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_8.mux_l1_in_2__S mux_right_track_8.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l3_in_1__S mux_top_track_2.mux_l3_in_1_/S vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l2_in_3_ right_top_grid_pin_47_ right_top_grid_pin_46_ mux_right_track_4.mux_l2_in_0_/S
+ mux_right_track_4.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_6_210 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_32.mux_l1_in_1__A1 right_top_grid_pin_45_ vgnd vpwr scs8hd_diode_2
XFILLER_41_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0__S mux_left_track_9.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
X_097_ chany_top_in[17] chany_bottom_out[18] vgnd vpwr scs8hd_buf_2
XFILLER_37_136 vgnd vpwr scs8hd_decap_4
XFILLER_37_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
XFILLER_1_75 vpwr vgnd scs8hd_fill_2
XFILLER_20_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l3_in_1__A0 mux_bottom_track_17.mux_l2_in_3_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l2_in_1_ chany_bottom_in[17] mux_top_track_16.mux_l1_in_2_/X
+ mux_top_track_16.mux_l2_in_0_/S mux_top_track_16.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_29_38 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l2_in_2__S mux_top_track_8.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__D mux_left_track_3.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_25.mux_l1_in_0_ chany_top_in[18] chany_top_in[9] mux_bottom_track_25.mux_l1_in_0_/S
+ mux_bottom_track_25.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_40 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_24.mux_l1_in_1__A1 chanx_right_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_19_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_6__S mux_bottom_track_5.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_10_84 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__D mux_top_track_24.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_161 vgnd vpwr scs8hd_decap_4
XFILLER_42_150 vpwr vgnd scs8hd_fill_2
XFILLER_34_117 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_4__A0 chanx_right_in[14] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_32.mux_l2_in_0__A0 mux_top_track_32.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_106 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1__A0 chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_18_191 vpwr vgnd scs8hd_fill_2
XFILLER_18_180 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_8.mux_l4_in_0_/S mux_right_track_16.mux_l1_in_0_/S
+ mem_right_track_16.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_0_227 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_3__D mux_bottom_track_17.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_32.mux_l2_in_0__A1 mux_right_track_32.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_128 vgnd vpwr scs8hd_fill_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A1 chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_21_83 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_2_ chany_bottom_in[8] chanx_right_in[17] mux_top_track_16.mux_l1_in_2_/S
+ mux_top_track_16.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_17.mux_l4_in_0__A0 mux_bottom_track_17.mux_l3_in_1_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_1_/S mux_left_track_3.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_30_142 vpwr vgnd scs8hd_fill_2
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_7_52 vpwr vgnd scs8hd_fill_2
XFILLER_7_96 vgnd vpwr scs8hd_fill_1
Xmux_right_track_16.mux_l4_in_0_ mux_right_track_16.mux_l3_in_1_/X mux_right_track_16.mux_l3_in_0_/X
+ mux_right_track_16.mux_l4_in_0_/S mux_right_track_16.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_38_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_33.mux_l1_in_0__S mux_bottom_track_33.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_24.mux_l2_in_0__A1 mux_top_track_24.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_33.scs8hd_dfxbp_1_1__D mux_left_track_33.mux_l1_in_3_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l4_in_0_ mux_right_track_4.mux_l3_in_1_/X mux_right_track_4.mux_l3_in_0_/X
+ mux_right_track_4.mux_l4_in_0_/S mux_right_track_4.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_21_153 vpwr vgnd scs8hd_fill_2
XFILLER_21_120 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_0_ chany_top_in[16] chany_top_in[6] mux_bottom_track_9.mux_l1_in_2_/S
+ mux_bottom_track_9.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_4.mux_l3_in_3__A0 mux_top_track_4.mux_l2_in_7_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1__A1 chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_8_146 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_32.mux_l3_in_0__S mux_top_track_32.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0__A0 mux_left_track_17.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_24.mux_l1_in_0__S mux_right_track_24.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_bottom_track_1.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_track_1.mux_l3_in_1_/S mux_bottom_track_1.mux_l4_in_0_/S
+ mem_bottom_track_1.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_9.mux_l2_in_3__A0 _049_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_3__A0 _030_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_2__A0 chanx_left_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_26_234 vgnd vpwr scs8hd_fill_1
Xmux_left_track_3.mux_l2_in_1_ mux_left_track_3.mux_l1_in_3_/X mux_left_track_3.mux_l1_in_2_/X
+ mux_left_track_3.mux_l2_in_2_/S mux_left_track_3.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_27_60 vgnd vpwr scs8hd_fill_1
XFILLER_17_234 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__D mux_top_track_0.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_270 vgnd vpwr scs8hd_decap_4
Xmux_right_track_16.mux_l3_in_1_ mux_right_track_16.mux_l2_in_3_/X mux_right_track_16.mux_l2_in_2_/X
+ mux_right_track_16.mux_l3_in_0_/S mux_right_track_16.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_9.mux_l2_in_3__S mux_left_track_9.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmem_right_track_24.scs8hd_dfxbp_1_3_ prog_clk mux_right_track_24.mux_l3_in_0_/S mux_right_track_24.mux_l4_in_0_/S
+ mem_right_track_24.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_4_182 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l3_in_1_ mux_right_track_4.mux_l2_in_3_/X mux_right_track_4.mux_l2_in_2_/X
+ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_97 vpwr vgnd scs8hd_fill_2
Xmem_top_track_4.scs8hd_dfxbp_1_3_ prog_clk mux_top_track_4.mux_l3_in_0_/S mux_top_track_4.mux_l4_in_0_/S
+ mem_top_track_4.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_31_270 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_3__D mux_left_track_5.mux_l3_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_2__A1 chanx_left_in[8] vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.scs8hd_buf_4_0_ mux_top_track_8.mux_l4_in_0_/X _131_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_top_track_8.mux_l2_in_0__A1 mux_top_track_8.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_270 vpwr vgnd scs8hd_fill_2
XFILLER_13_62 vgnd vpwr scs8hd_decap_3
XFILLER_13_84 vpwr vgnd scs8hd_fill_2
XFILLER_1_141 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l2_in_5_ bottom_left_grid_pin_41_ bottom_left_grid_pin_40_
+ mux_bottom_track_5.mux_l2_in_1_/S mux_bottom_track_5.mux_l2_in_5_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__100__A chany_top_in[14] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l3_in_1__A0 mux_bottom_track_25.mux_l2_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.mux_l1_in_2_ chany_bottom_in[0] chanx_right_in[13] mux_left_track_3.mux_l1_in_0_/S
+ mux_left_track_3.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_32.mux_l1_in_1__A1 chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_11_207 vpwr vgnd scs8hd_fill_2
Xmem_right_track_0.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_0.mux_l2_in_0_/S mux_right_track_0.mux_l3_in_0_/S
+ mem_right_track_0.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_5.mux_l2_in_7__A0 _048_/HI vgnd vpwr scs8hd_diode_2
Xmem_left_track_17.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_9.mux_l4_in_0_/S mux_left_track_17.mux_l1_in_0_/S
+ mem_left_track_17.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_track_16.mux_l2_in_2_ chanx_left_in[8] chany_bottom_in[17] mux_right_track_16.mux_l2_in_0_/S
+ mux_right_track_16.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_1_7 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_25.scs8hd_buf_4_0__A mux_bottom_track_25.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l2_in_2_ right_top_grid_pin_45_ right_top_grid_pin_44_ mux_right_track_4.mux_l2_in_0_/S
+ mux_right_track_4.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_5.mux_l2_in_2__A0 chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_10_273 vpwr vgnd scs8hd_fill_2
XFILLER_40_93 vpwr vgnd scs8hd_fill_2
X_096_ chany_top_in[18] chany_bottom_out[19] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0__S mux_bottom_track_1.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_6_266 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.mux_l1_in_1__A0 chanx_right_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_1_98 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_ mux_top_track_16.mux_l1_in_1_/X mux_top_track_16.mux_l1_in_0_/X
+ mux_top_track_16.mux_l2_in_0_/S mux_top_track_16.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_17.mux_l3_in_1__A1 mux_bottom_track_17.mux_l2_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_28 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_33.mux_l1_in_3__S mux_bottom_track_33.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_181 vpwr vgnd scs8hd_fill_2
XFILLER_28_148 vgnd vpwr scs8hd_decap_3
XFILLER_28_115 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_33.mux_l1_in_3__A0 _047_/HI vgnd vpwr scs8hd_diode_2
XFILLER_3_258 vpwr vgnd scs8hd_fill_2
XFILLER_3_214 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_25.mux_l4_in_0__A0 mux_bottom_track_25.mux_l3_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_10_74 vgnd vpwr scs8hd_fill_1
XFILLER_35_60 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_4.mux_l2_in_4__A1 chanx_right_in[7] vgnd vpwr scs8hd_diode_2
X_079_ _079_/A chanx_right_out[16] vgnd vpwr scs8hd_buf_2
XFILLER_25_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_32.mux_l2_in_0__A1 mux_top_track_32.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1__A1 chany_top_in[17] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__S mux_bottom_track_25.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l3_in_1__A0 mux_left_track_5.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_239 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0__S mux_left_track_17.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_195 vpwr vgnd scs8hd_fill_2
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_25.mux_l2_in_0__A0 mux_left_track_25.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_62 vpwr vgnd scs8hd_fill_2
XFILLER_21_51 vpwr vgnd scs8hd_fill_2
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_17.mux_l4_in_0__A1 mux_bottom_track_17.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_1_ chanx_right_in[15] chanx_right_in[8] mux_top_track_16.mux_l1_in_2_/S
+ mux_top_track_16.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_24.mux_l4_in_0__S mux_top_track_24.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__D mux_top_track_0.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0__S mux_right_track_16.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_165 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_24.mux_l2_in_3__A0 _032_/HI vgnd vpwr scs8hd_diode_2
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_162 vpwr vgnd scs8hd_fill_2
Xmem_left_track_25.scs8hd_dfxbp_1_3_ prog_clk mux_left_track_25.mux_l3_in_0_/S mux_left_track_25.mux_l4_in_0_/S
+ mem_left_track_25.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_132 vpwr vgnd scs8hd_fill_2
XFILLER_29_276 vgnd vpwr scs8hd_fill_1
XFILLER_29_254 vpwr vgnd scs8hd_fill_2
XFILLER_29_232 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l3_in_3__A1 mux_top_track_4.mux_l2_in_6_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_125 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_16.mux_l2_in_3__A0 _037_/HI vgnd vpwr scs8hd_diode_2
XFILLER_12_132 vpwr vgnd scs8hd_fill_2
XFILLER_32_83 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_0.mux_l1_in_1__S mux_top_track_0.mux_l1_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_12_198 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l2_in_0__A1 mux_left_track_17.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA__103__A _103_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_213 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l4_in_0__A0 mux_left_track_5.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_1.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_1.mux_l2_in_0_/S mux_bottom_track_1.mux_l3_in_1_/S
+ mem_bottom_track_1.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_9.mux_l2_in_3__A1 chanx_left_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.scs8hd_buf_4_0__A mux_top_track_8.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_3__A1 chanx_left_in[17] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l3_in_3_ mux_bottom_track_5.mux_l2_in_7_/X mux_bottom_track_5.mux_l2_in_6_/X
+ mux_bottom_track_5.mux_l3_in_2_/S mux_bottom_track_5.mux_l3_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_25.mux_l2_in_2__A1 chanx_left_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_26_224 vpwr vgnd scs8hd_fill_2
XFILLER_41_227 vgnd vpwr scs8hd_decap_3
Xmux_left_track_3.mux_l2_in_0_ mux_left_track_3.mux_l1_in_1_/X mux_left_track_3.mux_l1_in_0_/X
+ mux_left_track_3.mux_l2_in_2_/S mux_left_track_3.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_32_238 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l3_in_0_ mux_right_track_16.mux_l2_in_1_/X mux_right_track_16.mux_l2_in_0_/X
+ mux_right_track_16.mux_l3_in_0_/S mux_right_track_16.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_right_track_24.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_24.mux_l2_in_2_/S mux_right_track_24.mux_l3_in_0_/S
+ mem_right_track_24.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_4_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_3__S mux_bottom_track_1.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_87 vpwr vgnd scs8hd_fill_2
Xmem_top_track_4.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_4.mux_l2_in_0_/S mux_top_track_4.mux_l3_in_0_/S
+ mem_top_track_4.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_13_52 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_33.mux_l1_in_1__A0 chany_bottom_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l3_in_1__S mux_bottom_track_5.mux_l3_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_38_60 vpwr vgnd scs8hd_fill_2
XFILLER_1_197 vpwr vgnd scs8hd_fill_2
XFILLER_20_208 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_5.mux_l2_in_4_ bottom_left_grid_pin_39_ bottom_left_grid_pin_38_
+ mux_bottom_track_5.mux_l2_in_1_/S mux_bottom_track_5.mux_l2_in_4_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_25.mux_l3_in_1__A1 mux_bottom_track_25.mux_l2_in_2_/X vgnd
+ vpwr scs8hd_diode_2
Xmem_right_track_8.scs8hd_dfxbp_1_3_ prog_clk mux_right_track_8.mux_l3_in_0_/S mux_right_track_8.mux_l4_in_0_/S
+ mem_right_track_8.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_231 vgnd vpwr scs8hd_fill_1
XFILLER_9_242 vpwr vgnd scs8hd_fill_2
XFILLER_9_253 vpwr vgnd scs8hd_fill_2
XFILLER_34_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_25.mux_l2_in_3__S mux_bottom_track_25.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_3.mux_l1_in_1_ chanx_right_in[4] chany_top_in[19] mux_left_track_3.mux_l1_in_0_/S
+ mux_left_track_3.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmem_right_track_0.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_0.mux_l1_in_1_/S mux_right_track_0.mux_l2_in_0_/S
+ mem_right_track_0.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_5.mux_l2_in_7__A1 chanx_left_in[14] vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l2_in_1_ chany_bottom_in[8] mux_right_track_16.mux_l1_in_2_/X
+ mux_right_track_16.mux_l2_in_0_/S mux_right_track_16.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_1__A0 right_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l2_in_1_ right_top_grid_pin_43_ right_top_grid_pin_42_ mux_right_track_4.mux_l2_in_0_/S
+ mux_right_track_4.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_84 vpwr vgnd scs8hd_fill_2
XFILLER_24_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_2__A1 chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l5_in_0_ mux_bottom_track_5.mux_l4_in_1_/X mux_bottom_track_5.mux_l4_in_0_/X
+ mux_bottom_track_5.mux_l5_in_0_/S mux_bottom_track_5.mux_l5_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_241 vpwr vgnd scs8hd_fill_2
X_095_ _095_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_40_83 vpwr vgnd scs8hd_fill_2
XFILLER_27_7 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_3__D mux_top_track_2.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l1_in_1__A1 chany_top_in[18] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_3__S mux_right_track_16.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__111__A _111_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l3_in_0__S mux_bottom_track_17.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_33.mux_l2_in_0__A0 mux_left_track_33.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__D mux_bottom_track_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l1_in_3__A1 chanx_left_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2__S mux_left_track_1.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l4_in_0__A1 mux_bottom_track_25.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__D mux_left_track_9.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_19_138 vpwr vgnd scs8hd_fill_2
XFILLER_19_116 vgnd vpwr scs8hd_decap_4
XFILLER_19_105 vgnd vpwr scs8hd_decap_4
XFILLER_19_40 vpwr vgnd scs8hd_fill_2
XFILLER_42_196 vgnd vpwr scs8hd_decap_4
XFILLER_27_193 vpwr vgnd scs8hd_fill_2
X_078_ chanx_left_in[16] chanx_right_out[17] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_0.mux_l1_in_3__A0 chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__106__A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_4__S mux_top_track_0.mux_l1_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_2_270 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_0__S mux_left_track_5.mux_l2_in_7_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_2_ chany_bottom_in[1] right_top_grid_pin_47_ mux_right_track_16.mux_l1_in_0_/S
+ mux_right_track_16.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_2.mux_l2_in_0__A0 mux_right_track_2.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l3_in_1__A1 mux_left_track_5.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_4__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l4_in_1_ mux_bottom_track_5.mux_l3_in_3_/X mux_bottom_track_5.mux_l3_in_2_/X
+ mux_bottom_track_5.mux_l4_in_0_/S mux_bottom_track_5.mux_l4_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_24.mux_l2_in_3__A0 _039_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0__S mux_right_track_8.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_141 vpwr vgnd scs8hd_fill_2
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_25.mux_l2_in_0__A1 mux_left_track_25.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_2__S mux_top_track_4.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_ top_left_grid_pin_39_ top_left_grid_pin_35_ mux_top_track_16.mux_l1_in_2_/S
+ mux_top_track_16.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_2__D mux_left_track_17.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_24.mux_l2_in_3__A1 chanx_left_in[18] vgnd vpwr scs8hd_diode_2
XPHY_5 vgnd vpwr scs8hd_decap_3
Xmem_left_track_25.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_25.mux_l2_in_3_/S mux_left_track_25.mux_l3_in_0_/S
+ mem_left_track_25.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_7_21 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_32.scs8hd_dfxbp_1_2__D mux_right_track_32.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_65 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l3_in_0__S mux_top_track_8.mux_l3_in_1_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_2__A0 chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_29_266 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_track_9.mux_l3_in_1_/S mux_bottom_track_9.mux_l4_in_0_/S
+ mem_bottom_track_9.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_16.mux_l2_in_3__A1 chanx_left_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_32_40 vpwr vgnd scs8hd_fill_2
XFILLER_8_137 vgnd vpwr scs8hd_decap_3
XFILLER_12_177 vpwr vgnd scs8hd_fill_2
XFILLER_35_258 vpwr vgnd scs8hd_fill_2
XFILLER_35_236 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_1.mux_l1_in_0_/S mux_bottom_track_1.mux_l2_in_0_/S
+ mem_bottom_track_1.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_5.mux_l4_in_0__A1 mux_left_track_5.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_5.mux_l3_in_2_ mux_bottom_track_5.mux_l2_in_5_/X mux_bottom_track_5.mux_l2_in_4_/X
+ mux_bottom_track_5.mux_l3_in_2_/S mux_bottom_track_5.mux_l3_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_26_258 vpwr vgnd scs8hd_fill_2
XFILLER_17_203 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_3__A0 _042_/HI vgnd vpwr scs8hd_diode_2
XFILLER_27_40 vpwr vgnd scs8hd_fill_2
XFILLER_17_258 vgnd vpwr scs8hd_fill_1
Xmem_right_track_24.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_24.mux_l1_in_1_/S mux_right_track_24.mux_l2_in_2_/S
+ mem_right_track_24.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA__114__A _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_55 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__D mux_top_track_4.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_32.mux_l1_in_1__S mux_right_track_32.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmem_top_track_4.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_4.mux_l1_in_0_/S mux_top_track_4.mux_l2_in_0_/S
+ mem_top_track_4.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_31_261 vgnd vpwr scs8hd_fill_1
XFILLER_23_228 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l3_in_1__A0 mux_right_track_0.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__D mux_bottom_track_3.mux_l1_in_4_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_228 vpwr vgnd scs8hd_fill_2
XFILLER_14_239 vpwr vgnd scs8hd_fill_2
XFILLER_13_20 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_33.mux_l1_in_1__A1 chanx_right_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_1_176 vgnd vpwr scs8hd_decap_4
XFILLER_38_72 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_5.mux_l2_in_3_ bottom_left_grid_pin_37_ bottom_left_grid_pin_36_
+ mux_bottom_track_5.mux_l2_in_1_/S mux_bottom_track_5.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
Xmem_right_track_8.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_8.mux_l2_in_1_/S mux_right_track_8.mux_l3_in_0_/S
+ mem_right_track_8.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA__109__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_9_210 vpwr vgnd scs8hd_fill_2
XFILLER_13_261 vpwr vgnd scs8hd_fill_2
XFILLER_9_265 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_3__S mux_left_track_5.mux_l2_in_7_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_3.mux_l1_in_0_ chany_top_in[13] chany_top_in[4] mux_left_track_3.mux_l1_in_0_/S
+ mux_left_track_3.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_3.mux_l4_in_0__S mux_left_track_3.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_right_track_0.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_32.mux_l3_in_0_/S mux_right_track_0.mux_l1_in_1_/S
+ mem_right_track_0.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_39_180 vgnd vpwr scs8hd_fill_1
Xmux_right_track_16.mux_l2_in_0_ mux_right_track_16.mux_l1_in_1_/X mux_right_track_16.mux_l1_in_0_/X
+ mux_right_track_16.mux_l2_in_0_/S mux_right_track_16.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_4.mux_l2_in_0_ chany_top_in[14] mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_0_/S mux_right_track_4.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_1__A1 chany_top_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_24_74 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_8.mux_l2_in_3__S mux_right_track_8.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_5__S mux_top_track_4.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l4_in_0__A0 mux_right_track_0.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_202 vpwr vgnd scs8hd_fill_2
XFILLER_6_224 vpwr vgnd scs8hd_fill_2
XFILLER_10_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0__S mux_top_track_16.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
X_094_ _094_/A chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_37_106 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l3_in_1__S mux_left_track_9.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_7__A0 _041_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_33.mux_l2_in_0__A1 mux_left_track_33.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_194 vpwr vgnd scs8hd_fill_2
XFILLER_3_227 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.scs8hd_buf_4_0_ mux_bottom_track_1.mux_l4_in_0_/X _115_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_3_238 vgnd vpwr scs8hd_decap_4
XFILLER_10_65 vgnd vpwr scs8hd_decap_3
XFILLER_10_98 vpwr vgnd scs8hd_fill_2
XFILLER_42_120 vpwr vgnd scs8hd_fill_2
XFILLER_35_51 vgnd vpwr scs8hd_decap_3
XFILLER_35_95 vgnd vpwr scs8hd_decap_3
XFILLER_35_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_3__A1 right_top_grid_pin_48_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2__A0 chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__122__A chany_bottom_in[12] vgnd vpwr scs8hd_diode_2
X_077_ chanx_left_in[17] chanx_right_out[18] vgnd vpwr scs8hd_buf_2
XFILLER_32_6 vgnd vpwr scs8hd_decap_3
XFILLER_33_175 vgnd vpwr scs8hd_decap_4
XFILLER_33_153 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_2.mux_l2_in_0__A1 mux_right_track_2.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_1_ right_top_grid_pin_43_ chany_top_in[17] mux_right_track_16.mux_l1_in_0_/S
+ mux_right_track_16.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_0_208 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_5.mux_l4_in_0_ mux_bottom_track_5.mux_l3_in_1_/X mux_bottom_track_5.mux_l3_in_0_/X
+ mux_bottom_track_5.mux_l4_in_0_/S mux_bottom_track_5.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_24.mux_l2_in_3__A1 chanx_left_in[18] vgnd vpwr scs8hd_diode_2
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A0 chany_top_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_30_101 vpwr vgnd scs8hd_fill_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_3.mux_l1_in_1__S mux_bottom_track_3.mux_l1_in_4_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_131 vpwr vgnd scs8hd_fill_2
XFILLER_15_175 vpwr vgnd scs8hd_fill_2
Xmem_left_track_25.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_25.mux_l1_in_1_/S mux_left_track_25.mux_l2_in_3_/S
+ mem_left_track_25.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA__117__A chany_bottom_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_30_189 vpwr vgnd scs8hd_fill_2
XFILLER_15_197 vpwr vgnd scs8hd_fill_2
X_129_ chany_bottom_in[5] chany_top_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_17.mux_l2_in_3__A0 _051_/HI vgnd vpwr scs8hd_diode_2
XFILLER_7_99 vpwr vgnd scs8hd_fill_2
XFILLER_38_245 vgnd vpwr scs8hd_decap_8
XFILLER_42_19 vpwr vgnd scs8hd_fill_2
XFILLER_21_178 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_33.mux_l2_in_1__S mux_bottom_track_33.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_1__A0 chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_2__A1 mux_right_track_0.mux_l1_in_4_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__D mux_bottom_track_3.mux_l4_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_9.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_9.mux_l2_in_3_/S mux_bottom_track_9.mux_l3_in_1_/S
+ mem_bottom_track_9.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_16_64 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.mux_l1_in_1__S mux_left_track_25.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_96 vgnd vpwr scs8hd_decap_3
XFILLER_12_145 vpwr vgnd scs8hd_fill_2
XFILLER_16_97 vpwr vgnd scs8hd_fill_2
XFILLER_35_226 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_32.mux_l3_in_0_/S mux_bottom_track_1.mux_l1_in_0_/S
+ mem_bottom_track_1.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_24.mux_l2_in_1__S mux_right_track_24.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2__A0 bottom_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_6__S mux_left_track_5.mux_l2_in_7_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_5.mux_l3_in_1_ mux_bottom_track_5.mux_l2_in_3_/X mux_bottom_track_5.mux_l2_in_2_/X
+ mux_bottom_track_5.mux_l3_in_2_/S mux_bottom_track_5.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_7_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_5_119 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__D mux_right_track_8.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_3__A1 chanx_left_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_32_207 vgnd vpwr scs8hd_fill_1
XFILLER_27_74 vgnd vpwr scs8hd_fill_1
XFILLER_25_270 vpwr vgnd scs8hd_fill_2
Xmem_right_track_24.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_16.mux_l4_in_0_/S mux_right_track_24.mux_l1_in_1_/S
+ mem_right_track_24.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA__130__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_4_78 vpwr vgnd scs8hd_fill_2
XFILLER_4_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l3_in_0__A0 mux_left_track_9.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_4.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_2.mux_l4_in_0_/S mux_top_track_4.mux_l1_in_0_/S
+ mem_top_track_4.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_31_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l3_in_1__A1 mux_right_track_0.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_207 vgnd vpwr scs8hd_decap_4
XFILLER_13_43 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_1__A0 mux_bottom_track_1.mux_l1_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_3 vpwr vgnd scs8hd_fill_2
XFILLER_38_84 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l2_in_2_ bottom_left_grid_pin_35_ bottom_left_grid_pin_34_
+ mux_bottom_track_5.mux_l2_in_1_/S mux_bottom_track_5.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_5.mux_l2_in_5__A0 left_top_grid_pin_46_ vgnd vpwr scs8hd_diode_2
Xmem_right_track_8.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_8.mux_l1_in_2_/S mux_right_track_8.mux_l2_in_1_/S
+ mem_right_track_8.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_200 vgnd vpwr scs8hd_fill_1
XFILLER_13_273 vpwr vgnd scs8hd_fill_2
XANTENNA__125__A chany_bottom_in[9] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_24_97 vpwr vgnd scs8hd_fill_2
XFILLER_10_210 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l4_in_0__A1 mux_right_track_0.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
X_093_ _093_/A chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_6_247 vpwr vgnd scs8hd_fill_2
XFILLER_6_258 vpwr vgnd scs8hd_fill_2
XFILLER_10_265 vpwr vgnd scs8hd_fill_2
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
XFILLER_37_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_4__S mux_bottom_track_3.mux_l1_in_4_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_5.scs8hd_buf_4_0_ mux_left_track_5.mux_l5_in_0_/X _073_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_bottom_track_1.mux_l3_in_1__S mux_bottom_track_1.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_7__A1 chanx_left_in[15] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__D mux_top_track_4.mux_l5_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_129 vgnd vpwr scs8hd_decap_4
XFILLER_28_107 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l3_in_0__A0 mux_bottom_track_1.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_173 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_3__D mux_bottom_track_5.mux_l3_in_2_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_44 vpwr vgnd scs8hd_fill_2
XFILLER_19_53 vgnd vpwr scs8hd_decap_4
XFILLER_42_154 vgnd vpwr scs8hd_fill_1
XFILLER_27_162 vpwr vgnd scs8hd_fill_2
XFILLER_27_151 vpwr vgnd scs8hd_fill_2
XFILLER_19_75 vpwr vgnd scs8hd_fill_2
XFILLER_42_165 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_25.mux_l2_in_3__A0 _052_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2__A1 chanx_right_in[16] vgnd vpwr scs8hd_diode_2
X_076_ chanx_left_in[18] chanx_right_out[19] vgnd vpwr scs8hd_buf_2
XFILLER_18_140 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l1_in_0_ chany_top_in[8] chany_top_in[7] mux_right_track_16.mux_l1_in_0_/S
+ mux_right_track_16.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_33_187 vpwr vgnd scs8hd_fill_2
XFILLER_33_132 vpwr vgnd scs8hd_fill_2
XFILLER_18_173 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_25.mux_l3_in_1__S mux_bottom_track_25.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l1_in_0_ chany_top_in[5] chany_top_in[1] mux_right_track_4.mux_l1_in_0_/S
+ mux_right_track_4.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vpwr vgnd scs8hd_fill_2
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_17.mux_l2_in_1__S mux_left_track_17.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_3__D mux_right_track_16.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_87 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A1 chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_30_146 vpwr vgnd scs8hd_fill_2
XFILLER_30_124 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_7 vgnd vpwr scs8hd_decap_3
X_128_ chany_bottom_in[6] chany_top_out[7] vgnd vpwr scs8hd_buf_2
Xmem_left_track_25.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_17.mux_l4_in_0_/S mux_left_track_25.mux_l1_in_1_/S
+ mem_left_track_25.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_17.mux_l2_in_3__A1 left_top_grid_pin_47_ vgnd vpwr scs8hd_diode_2
XANTENNA__133__A _133_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l3_in_1__S mux_right_track_16.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_157 vpwr vgnd scs8hd_fill_2
XFILLER_7_56 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_33.scs8hd_buf_4_0__A mux_bottom_track_33.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
X_059_ _059_/A chanx_left_out[16] vgnd vpwr scs8hd_buf_2
XFILLER_38_224 vpwr vgnd scs8hd_fill_2
XFILLER_38_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.mux_l1_in_2__S mux_right_track_0.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_1__A1 mux_left_track_9.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0__S mux_left_track_1.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_9.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_9.mux_l1_in_2_/S mux_bottom_track_9.mux_l2_in_3_/S
+ mem_bottom_track_9.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_12_102 vpwr vgnd scs8hd_fill_2
XFILLER_16_10 vpwr vgnd scs8hd_fill_2
XFILLER_16_32 vpwr vgnd scs8hd_fill_2
XFILLER_16_87 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0__S mux_right_track_4.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_2__S mux_top_track_0.mux_l2_in_2_/S vgnd vpwr scs8hd_diode_2
XANTENNA__128__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2__A1 chanx_right_in[15] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ mux_bottom_track_5.mux_l3_in_2_/S mux_bottom_track_5.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_260 vpwr vgnd scs8hd_fill_2
XFILLER_27_53 vgnd vpwr scs8hd_decap_4
XFILLER_17_238 vgnd vpwr scs8hd_decap_4
XFILLER_17_216 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_4.mux_l3_in_0__S mux_top_track_4.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_40_274 vgnd vpwr scs8hd_fill_1
XFILLER_4_186 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l3_in_0__A1 mux_left_track_9.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_3__D mux_top_track_8.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__D mux_bottom_track_17.mux_l4_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_22_274 vgnd vpwr scs8hd_fill_1
XFILLER_1_123 vgnd vpwr scs8hd_decap_3
XFILLER_1_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_1__A1 mux_bottom_track_1.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_4__A0 chany_bottom_in[13] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l2_in_1_ chanx_right_in[14] chanx_right_in[7] mux_bottom_track_5.mux_l2_in_1_/S
+ mux_bottom_track_5.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmem_right_track_8.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_4.mux_l5_in_0_/S mux_right_track_8.mux_l1_in_2_/S
+ mem_right_track_8.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_5.mux_l2_in_5__A1 left_top_grid_pin_45_ vgnd vpwr scs8hd_diode_2
XFILLER_9_234 vpwr vgnd scs8hd_fill_2
XFILLER_13_252 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_4.mux_l2_in_1__A0 right_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
XFILLER_24_32 vgnd vpwr scs8hd_decap_4
XFILLER_40_97 vpwr vgnd scs8hd_fill_2
XFILLER_40_53 vpwr vgnd scs8hd_fill_2
X_092_ chanx_left_in[2] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_1_36 vpwr vgnd scs8hd_fill_2
XFILLER_5_270 vpwr vgnd scs8hd_fill_2
XFILLER_36_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.mux_l3_in_0__A1 mux_bottom_track_1.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_3__A0 _031_/HI vgnd vpwr scs8hd_diode_2
Xmem_right_track_32.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_32.mux_l2_in_0_/S mux_right_track_32.mux_l3_in_0_/S
+ mem_right_track_32.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_1.mux_l2_in_3__S mux_left_track_1.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_10_23 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_33.mux_l1_in_3_ _047_/HI chanx_left_in[10] mux_bottom_track_33.mux_l1_in_0_/S
+ mux_bottom_track_33.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_25.mux_l2_in_3__A1 left_top_grid_pin_48_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l3_in_0__A0 mux_right_track_4.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
X_075_ _075_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_24.mux_l1_in_1__S mux_top_track_24.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_3__S mux_right_track_4.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_7 vgnd vpwr scs8hd_fill_1
XFILLER_2_262 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l4_in_0__S mux_right_track_2.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_6 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_5.mux_l3_in_1__S mux_left_track_5.mux_l3_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_199 vpwr vgnd scs8hd_fill_2
XFILLER_21_55 vgnd vpwr scs8hd_decap_4
XFILLER_21_22 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__D mux_top_track_32.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l3_in_1__S mux_right_track_8.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l3_in_3__S mux_top_track_4.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.scs8hd_buf_4_0__A mux_left_track_5.mux_l5_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_111 vpwr vgnd scs8hd_fill_2
X_127_ _127_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
X_058_ chanx_right_in[16] chanx_left_out[17] vgnd vpwr scs8hd_buf_2
XFILLER_38_203 vgnd vpwr scs8hd_decap_4
XFILLER_21_136 vpwr vgnd scs8hd_fill_2
XFILLER_21_114 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_3__D mux_bottom_track_25.mux_l3_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0__A0 top_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_29_258 vpwr vgnd scs8hd_fill_2
XFILLER_29_236 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_5.mux_l5_in_0_/S mux_bottom_track_9.mux_l1_in_2_/S
+ mem_bottom_track_9.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_12_125 vgnd vpwr scs8hd_decap_4
XFILLER_16_55 vpwr vgnd scs8hd_fill_2
XFILLER_20_191 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__D mux_bottom_track_9.mux_l1_in_2_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_162 vpwr vgnd scs8hd_fill_2
XFILLER_26_228 vgnd vpwr scs8hd_decap_4
XFILLER_26_206 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_33.mux_l3_in_0_ mux_bottom_track_33.mux_l2_in_1_/X mux_bottom_track_33.mux_l2_in_0_/X
+ mux_bottom_track_33.mux_l3_in_0_/S mux_bottom_track_33.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XFILLER_34_272 vgnd vpwr scs8hd_decap_3
XFILLER_27_87 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_2__A0 chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_33.mux_l1_in_2__S mux_left_track_33.mux_l1_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_4_132 vpwr vgnd scs8hd_fill_2
XFILLER_4_110 vgnd vpwr scs8hd_decap_3
XFILLER_4_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__D mux_top_track_32.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_left_track_33.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_33.mux_l2_in_1_/S ccff_tail
+ mem_left_track_33.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_22_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0__S mux_bottom_track_9.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_56 vpwr vgnd scs8hd_fill_2
XFILLER_1_102 vpwr vgnd scs8hd_fill_2
XFILLER_13_67 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l1_in_4__A1 chany_bottom_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_38_64 vpwr vgnd scs8hd_fill_2
XFILLER_1_168 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l2_in_0_ chanx_right_in[5] mux_bottom_track_5.mux_l1_in_0_/X
+ mux_bottom_track_5.mux_l2_in_1_/S mux_bottom_track_5.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_13_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_6__S mux_right_track_4.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_33.mux_l2_in_1_ mux_bottom_track_33.mux_l1_in_3_/X mux_bottom_track_33.mux_l1_in_2_/X
+ mux_bottom_track_33.mux_l2_in_1_/S mux_bottom_track_33.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_mux2_1
XANTENNA_mux_right_track_4.mux_l2_in_1__A1 right_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_1__A0 mux_top_track_0.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_172 vpwr vgnd scs8hd_fill_2
XFILLER_40_32 vpwr vgnd scs8hd_fill_2
XFILLER_24_88 vpwr vgnd scs8hd_fill_2
XFILLER_24_66 vpwr vgnd scs8hd_fill_2
X_091_ _091_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_10_245 vpwr vgnd scs8hd_fill_2
XFILLER_40_87 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l2_in_1__S mux_top_track_16.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_131 vgnd vpwr scs8hd_fill_1
Xmem_right_track_32.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_32.mux_l1_in_0_/S mux_right_track_32.mux_l2_in_0_/S
+ mem_right_track_32.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_2.mux_l2_in_3__A1 chanx_left_in[13] vgnd vpwr scs8hd_diode_2
Xmux_top_track_24.mux_l2_in_3_ _039_/HI chanx_left_in[18] mux_top_track_24.mux_l2_in_2_/S
+ mux_top_track_24.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__062__A chanx_right_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_27_142 vpwr vgnd scs8hd_fill_2
XFILLER_19_109 vgnd vpwr scs8hd_fill_1
XFILLER_19_88 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_33.mux_l1_in_2_ chanx_left_in[0] bottom_left_grid_pin_41_ mux_bottom_track_33.mux_l1_in_0_/S
+ mux_bottom_track_33.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_42_178 vpwr vgnd scs8hd_fill_2
XFILLER_42_156 vgnd vpwr scs8hd_fill_1
XFILLER_42_134 vpwr vgnd scs8hd_fill_2
XFILLER_35_21 vpwr vgnd scs8hd_fill_2
XFILLER_27_197 vpwr vgnd scs8hd_fill_2
XFILLER_27_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l3_in_0__A1 mux_right_track_4.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0__S mux_top_track_2.mux_l1_in_3_/S vgnd vpwr scs8hd_diode_2
X_074_ _074_/A chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_0.mux_l3_in_0__A0 mux_top_track_0.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_274 vgnd vpwr scs8hd_fill_1
XFILLER_2_241 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_3__A0 bottom_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
XFILLER_33_112 vgnd vpwr scs8hd_decap_4
XFILLER_33_156 vpwr vgnd scs8hd_fill_2
XFILLER_2_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_5.mux_l2_in_0__A0 chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.scs8hd_buf_4_0__A mux_right_track_4.mux_l5_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA__057__A chanx_right_in[17] vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l2_in_3_ _051_/HI left_top_grid_pin_47_ mux_left_track_17.mux_l2_in_1_/S
+ mux_left_track_17.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_178 vpwr vgnd scs8hd_fill_2
XFILLER_24_145 vpwr vgnd scs8hd_fill_2
XFILLER_24_101 vpwr vgnd scs8hd_fill_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_34 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_3.mux_l2_in_2__S mux_bottom_track_3.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_25 vpwr vgnd scs8hd_fill_2
X_126_ chany_bottom_in[8] chany_top_out[9] vgnd vpwr scs8hd_buf_2
X_057_ chanx_right_in[17] chanx_left_out[18] vgnd vpwr scs8hd_buf_2
XFILLER_7_69 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_38_259 vgnd vpwr scs8hd_decap_12
XFILLER_30_6 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_3__D mux_right_track_0.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0__A1 top_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0__A0 chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_29_215 vpwr vgnd scs8hd_fill_2
XFILLER_16_23 vpwr vgnd scs8hd_fill_2
XFILLER_32_44 vgnd vpwr scs8hd_decap_3
XFILLER_32_11 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_3.mux_l2_in_2__A0 chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l2_in_2__S mux_left_track_25.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_88 vpwr vgnd scs8hd_fill_2
XFILLER_32_66 vpwr vgnd scs8hd_fill_2
XFILLER_20_170 vpwr vgnd scs8hd_fill_2
Xmux_top_track_24.mux_l4_in_0_ mux_top_track_24.mux_l3_in_1_/X mux_top_track_24.mux_l3_in_0_/X
+ mux_top_track_24.mux_l4_in_0_/S mux_top_track_24.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
X_109_ chany_top_in[5] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_19_270 vgnd vpwr scs8hd_decap_6
Xmux_left_track_9.mux_l2_in_3_ _028_/HI left_top_grid_pin_46_ mux_left_track_9.mux_l2_in_1_/S
+ mux_left_track_9.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_8_90 vpwr vgnd scs8hd_fill_2
XANTENNA__070__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_27_77 vgnd vpwr scs8hd_fill_1
XFILLER_27_66 vpwr vgnd scs8hd_fill_2
XFILLER_27_33 vgnd vpwr scs8hd_fill_1
XFILLER_17_207 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_2__A1 chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
Xmux_right_track_0.mux_l2_in_3_ _029_/HI chanx_left_in[12] mux_right_track_0.mux_l2_in_0_/S
+ mux_right_track_0.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_199 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l4_in_0_ mux_left_track_17.mux_l3_in_1_/X mux_left_track_17.mux_l3_in_0_/X
+ mux_left_track_17.mux_l4_in_0_/S mux_left_track_17.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_31_276 vgnd vpwr scs8hd_fill_1
XFILLER_31_254 vgnd vpwr scs8hd_decap_4
XFILLER_31_221 vpwr vgnd scs8hd_fill_2
XFILLER_16_251 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0__S mux_right_track_0.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l1_in_1__S mux_left_track_3.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l3_in_1__A0 mux_bottom_track_3.mux_l2_in_3_/X vgnd
+ vpwr scs8hd_diode_2
Xmem_left_track_33.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_33.mux_l1_in_3_/S mux_left_track_33.mux_l2_in_1_/S
+ mem_left_track_33.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_22_210 vpwr vgnd scs8hd_fill_2
XANTENNA__065__A chanx_right_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_114 vpwr vgnd scs8hd_fill_2
Xmux_top_track_24.mux_l3_in_1_ mux_top_track_24.mux_l2_in_3_/X mux_top_track_24.mux_l2_in_2_/X
+ mux_top_track_24.mux_l3_in_0_/S mux_top_track_24.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_38_32 vgnd vpwr scs8hd_decap_3
XFILLER_38_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l1_in_3__S mux_top_track_2.mux_l1_in_3_/S vgnd vpwr scs8hd_diode_2
XFILLER_9_214 vpwr vgnd scs8hd_fill_2
XFILLER_13_210 vgnd vpwr scs8hd_decap_4
XFILLER_13_265 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l3_in_0__S mux_top_track_0.mux_l3_in_1_/S vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_33.mux_l2_in_0_ mux_bottom_track_33.mux_l1_in_1_/X mux_bottom_track_33.mux_l1_in_0_/X
+ mux_bottom_track_33.mux_l2_in_1_/S mux_bottom_track_33.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XFILLER_9_269 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_1__A1 mux_top_track_0.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_80 vpwr vgnd scs8hd_fill_2
XFILLER_24_23 vpwr vgnd scs8hd_fill_2
XFILLER_24_12 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_4_ chany_bottom_in[15] chany_bottom_in[12] mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_4_/X vgnd vpwr scs8hd_mux2_1
Xmux_left_track_17.mux_l3_in_1_ mux_left_track_17.mux_l2_in_3_/X mux_left_track_17.mux_l2_in_2_/X
+ mux_left_track_17.mux_l3_in_1_/S mux_left_track_17.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
X_090_ chanx_left_in[4] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_6_206 vpwr vgnd scs8hd_fill_2
XFILLER_6_228 vpwr vgnd scs8hd_fill_2
XFILLER_10_202 vpwr vgnd scs8hd_fill_2
XFILLER_10_224 vpwr vgnd scs8hd_fill_2
XFILLER_10_257 vpwr vgnd scs8hd_fill_2
XFILLER_6_3 vgnd vpwr scs8hd_decap_3
Xmux_left_track_9.mux_l4_in_0_ mux_left_track_9.mux_l3_in_1_/X mux_left_track_9.mux_l3_in_0_/X
+ mux_left_track_9.mux_l4_in_0_/S mux_left_track_9.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_3.mux_l4_in_0__A0 mux_bottom_track_3.mux_l3_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_39_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l1_in_1__A0 right_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
XFILLER_36_198 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__D mux_right_track_2.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_right_track_32.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_24.mux_l4_in_0_/S mux_right_track_32.mux_l1_in_0_/S
+ mem_right_track_32.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_top_track_24.mux_l2_in_2_ chanx_left_in[9] chanx_left_in[3] mux_top_track_24.mux_l2_in_2_/S
+ mux_top_track_24.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_0.mux_l4_in_0_ mux_right_track_0.mux_l3_in_1_/X mux_right_track_0.mux_l3_in_0_/X
+ mux_right_track_0.mux_l4_in_0_/S mux_right_track_0.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_track_5.mux_l1_in_0_ chany_top_in[14] chany_top_in[5] mux_bottom_track_5.mux_l1_in_0_/S
+ mux_bottom_track_5.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_19_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.scs8hd_buf_4_0__A mux_bottom_track_3.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_33.mux_l1_in_1_ bottom_left_grid_pin_37_ chanx_right_in[19] mux_bottom_track_33.mux_l1_in_0_/S
+ mux_bottom_track_33.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_42_168 vgnd vpwr scs8hd_fill_1
XFILLER_42_146 vpwr vgnd scs8hd_fill_2
XFILLER_35_66 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_5.mux_l5_in_0__S mux_bottom_track_5.mux_l5_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_073_ _073_/A chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_0.mux_l3_in_0__A1 mux_top_track_0.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_3__A1 bottom_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
XFILLER_33_179 vgnd vpwr scs8hd_fill_1
XFILLER_18_187 vpwr vgnd scs8hd_fill_2
XFILLER_18_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_2__D mux_top_track_16.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l2_in_2_ left_top_grid_pin_43_ chany_bottom_in[17] mux_left_track_17.mux_l2_in_1_/S
+ mux_left_track_17.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_2_70 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0__A1 mux_bottom_track_5.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_24_124 vpwr vgnd scs8hd_fill_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_0.scs8hd_buf_4_0_ mux_right_track_0.mux_l4_in_0_/X _095_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA__073__A _073_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l3_in_1_ mux_left_track_9.mux_l2_in_3_/X mux_left_track_9.mux_l2_in_2_/X
+ mux_left_track_9.mux_l3_in_1_/S mux_left_track_9.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_15_135 vpwr vgnd scs8hd_fill_2
X_125_ chany_bottom_in[9] chany_top_out[10] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_8.mux_l2_in_0__A0 mux_right_track_8.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_48 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_32.mux_l1_in_2__S mux_top_track_32.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
X_056_ chanx_right_in[18] chanx_left_out[19] vgnd vpwr scs8hd_buf_2
XFILLER_23_6 vpwr vgnd scs8hd_fill_2
XFILLER_21_149 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l3_in_1_ mux_right_track_0.mux_l2_in_3_/X mux_right_track_0.mux_l2_in_2_/X
+ mux_right_track_0.mux_l3_in_0_/S mux_right_track_0.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_0.mux_l2_in_3__S mux_right_track_0.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0__A1 chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l1_in_4__S mux_left_track_3.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_260 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l3_in_1__S mux_left_track_1.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA__068__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_16_68 vpwr vgnd scs8hd_fill_2
XFILLER_32_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_2__A1 mux_bottom_track_3.mux_l1_in_4_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_2__D mux_left_track_25.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l3_in_1__S mux_right_track_4.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
X_108_ chany_top_in[6] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_7_120 vpwr vgnd scs8hd_fill_2
XFILLER_7_153 vgnd vpwr scs8hd_decap_3
XFILLER_7_175 vpwr vgnd scs8hd_fill_2
XFILLER_7_197 vpwr vgnd scs8hd_fill_2
XFILLER_21_3 vpwr vgnd scs8hd_fill_2
X_039_ _039_/HI _039_/LO vgnd vpwr scs8hd_conb_1
Xmux_left_track_9.mux_l2_in_2_ left_top_grid_pin_42_ chany_bottom_in[16] mux_left_track_9.mux_l2_in_1_/S
+ mux_left_track_9.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_40_200 vpwr vgnd scs8hd_fill_2
XFILLER_25_274 vgnd vpwr scs8hd_decap_3
XFILLER_25_241 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_4.mux_l4_in_1__S mux_top_track_4.mux_l4_in_0_/S vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l2_in_2_ chanx_left_in[2] mux_right_track_0.mux_l1_in_4_/X
+ mux_right_track_0.mux_l2_in_0_/S mux_right_track_0.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_27 vpwr vgnd scs8hd_fill_2
XFILLER_4_145 vpwr vgnd scs8hd_fill_2
XFILLER_16_241 vgnd vpwr scs8hd_decap_4
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_266 vpwr vgnd scs8hd_fill_2
XFILLER_31_200 vpwr vgnd scs8hd_fill_2
XFILLER_16_263 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l3_in_1__A1 mux_bottom_track_3.mux_l2_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_4__A0 right_top_grid_pin_49_ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__D mux_right_track_4.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_left_track_33.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_25.mux_l4_in_0_/S mux_left_track_33.mux_l1_in_3_/S
+ mem_left_track_33.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_22_222 vgnd vpwr scs8hd_decap_4
XFILLER_22_266 vpwr vgnd scs8hd_fill_2
XFILLER_13_47 vgnd vpwr scs8hd_decap_3
XANTENNA__081__A chanx_left_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_8_7 vgnd vpwr scs8hd_decap_4
Xmux_top_track_24.mux_l3_in_0_ mux_top_track_24.mux_l2_in_1_/X mux_top_track_24.mux_l2_in_0_/X
+ mux_top_track_24.mux_l3_in_0_/S mux_top_track_24.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_38_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA__076__A chanx_left_in[18] vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_3_ chany_bottom_in[2] right_top_grid_pin_48_ mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
Xmux_left_track_17.mux_l3_in_0_ mux_left_track_17.mux_l2_in_1_/X mux_left_track_17.mux_l2_in_0_/X
+ mux_left_track_17.mux_l3_in_1_/S mux_left_track_17.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_2.mux_l2_in_3_ _038_/HI chanx_left_in[19] mux_top_track_2.mux_l2_in_2_/S
+ mux_top_track_2.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_269 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_33.mux_l2_in_0__S mux_left_track_33.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_24.mux_l2_in_3_ _032_/HI chanx_left_in[18] mux_right_track_24.mux_l2_in_2_/S
+ mux_right_track_24.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_5.mux_l1_in_0__S mux_bottom_track_5.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l4_in_0__A1 mux_bottom_track_3.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l3_in_3__A0 mux_right_track_4.mux_l2_in_7_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_1__A1 chany_top_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_32.mux_l3_in_0__S mux_right_track_32.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_177 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_17.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_track_17.mux_l3_in_0_/S
+ mux_bottom_track_17.mux_l4_in_0_/S mem_bottom_track_17.scs8hd_dfxbp_1_3_/QN vgnd
+ vpwr scs8hd_dfxbp_1
Xmux_top_track_24.mux_l2_in_1_ chany_bottom_in[18] mux_top_track_24.mux_l1_in_2_/X
+ mux_top_track_24.mux_l2_in_2_/S mux_top_track_24.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_42_103 vpwr vgnd scs8hd_fill_2
XFILLER_35_56 vpwr vgnd scs8hd_fill_2
XFILLER_35_34 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_33.mux_l1_in_0_ chanx_right_in[10] chany_top_in[10] mux_bottom_track_33.mux_l1_in_0_/S
+ mux_bottom_track_33.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
X_072_ chanx_right_in[2] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_24.mux_l2_in_2__S mux_top_track_24.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_136 vpwr vgnd scs8hd_fill_2
XFILLER_18_177 vgnd vpwr scs8hd_fill_1
XFILLER_18_144 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l2_in_1_ chany_bottom_in[8] mux_left_track_17.mux_l1_in_2_/X
+ mux_left_track_17.mux_l2_in_1_/S mux_left_track_17.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_2.mux_l1_in_4_ chanx_left_in[4] chany_bottom_in[13] mux_top_track_2.mux_l1_in_3_/S
+ mux_top_track_2.mux_l1_in_4_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_158 vgnd vpwr scs8hd_fill_1
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_9.mux_l3_in_0_ mux_left_track_9.mux_l2_in_1_/X mux_left_track_9.mux_l2_in_0_/X
+ mux_left_track_9.mux_l3_in_1_/S mux_left_track_9.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_2.mux_l1_in_3__A0 chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_21_14 vpwr vgnd scs8hd_fill_2
XFILLER_30_128 vgnd vpwr scs8hd_decap_3
XFILLER_15_158 vpwr vgnd scs8hd_fill_2
X_124_ chany_bottom_in[10] chany_top_out[11] vgnd vpwr scs8hd_buf_2
X_055_ _055_/HI _055_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_track_8.mux_l2_in_0__A1 mux_right_track_8.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_91 vpwr vgnd scs8hd_fill_2
Xmux_top_track_24.mux_l1_in_2_ chany_bottom_in[9] chanx_right_in[19] mux_top_track_24.mux_l1_in_1_/S
+ mux_top_track_24.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_4.mux_l2_in_0__A0 top_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
XFILLER_38_228 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_0_/S mux_right_track_0.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_16_6 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.mux_l4_in_0_ mux_top_track_2.mux_l3_in_1_/X mux_top_track_2.mux_l3_in_0_/X
+ mux_top_track_2.mux_l4_in_0_/S mux_top_track_2.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_14_180 vgnd vpwr scs8hd_decap_4
Xmux_right_track_24.mux_l4_in_0_ mux_right_track_24.mux_l3_in_1_/X mux_right_track_24.mux_l3_in_0_/X
+ mux_right_track_24.mux_l4_in_0_/S mux_right_track_24.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_4__D mux_right_track_4.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A0 chany_top_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_37_272 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l1_in_0__A0 chany_top_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__084__A chanx_left_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_35_209 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_2_ chany_bottom_in[7] chanx_right_in[17] mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
X_038_ _038_/HI _038_/LO vgnd vpwr scs8hd_conb_1
XFILLER_11_172 vgnd vpwr scs8hd_decap_4
X_107_ _107_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_14_3 vgnd vpwr scs8hd_decap_4
XFILLER_34_264 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_2.mux_l2_in_2__A0 chanx_left_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_19_261 vgnd vpwr scs8hd_fill_1
Xmux_left_track_9.mux_l2_in_1_ chany_bottom_in[6] mux_left_track_9.mux_l1_in_2_/X
+ mux_left_track_9.mux_l2_in_1_/S mux_left_track_9.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_8_81 vpwr vgnd scs8hd_fill_2
XANTENNA__079__A _079_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_57 vgnd vpwr scs8hd_fill_1
Xmux_right_track_0.mux_l2_in_1_ mux_right_track_0.mux_l1_in_3_/X mux_right_track_0.mux_l1_in_2_/X
+ mux_right_track_0.mux_l2_in_0_/S mux_right_track_0.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_3.mux_l3_in_0__S mux_bottom_track_3.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.mux_l3_in_1_ mux_top_track_2.mux_l2_in_3_/X mux_top_track_2.mux_l2_in_2_/X
+ mux_top_track_2.mux_l3_in_1_/S mux_top_track_2.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_24.mux_l3_in_1_ mux_right_track_24.mux_l2_in_3_/X mux_right_track_24.mux_l2_in_2_/X
+ mux_right_track_24.mux_l3_in_0_/S mux_right_track_24.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_4__A1 right_top_grid_pin_48_ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__D mux_right_track_16.mux_l4_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_1__S mux_bottom_track_9.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_38_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.mux_l3_in_0__S mux_left_track_25.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l3_in_1__A0 mux_top_track_2.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_227 vgnd vpwr scs8hd_decap_4
XFILLER_9_238 vpwr vgnd scs8hd_fill_2
XFILLER_9_249 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_2_ chany_bottom_in[3] chanx_right_in[16] mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_0_182 vpwr vgnd scs8hd_fill_2
Xmem_left_track_5.scs8hd_dfxbp_1_4_ prog_clk mux_left_track_5.mux_l4_in_0_/S mux_left_track_5.mux_l5_in_0_/S
+ mem_left_track_5.scs8hd_dfxbp_1_4_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_24.mux_l4_in_0__S mux_right_track_24.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2__S mux_bottom_track_17.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_142 vgnd vpwr scs8hd_decap_4
Xmux_right_track_0.mux_l1_in_2_ right_top_grid_pin_46_ right_top_grid_pin_44_ mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_58 vpwr vgnd scs8hd_fill_2
XFILLER_24_36 vgnd vpwr scs8hd_fill_1
XFILLER_40_79 vpwr vgnd scs8hd_fill_2
XFILLER_40_57 vgnd vpwr scs8hd_decap_3
Xmux_top_track_2.mux_l2_in_2_ chanx_left_in[13] mux_top_track_2.mux_l1_in_4_/X mux_top_track_2.mux_l2_in_2_/S
+ mux_top_track_2.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__092__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
Xmux_right_track_24.mux_l2_in_2_ chanx_left_in[9] chany_bottom_in[18] mux_right_track_24.mux_l2_in_2_/S
+ mux_right_track_24.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_4.mux_l3_in_3__A1 mux_right_track_4.mux_l2_in_6_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_80 vgnd vpwr scs8hd_decap_4
XFILLER_14_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_33.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_1__S mux_right_track_2.mux_l1_in_4_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_274 vgnd vpwr scs8hd_decap_3
XFILLER_36_134 vgnd vpwr scs8hd_fill_1
XFILLER_36_101 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_17.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_17.mux_l2_in_2_/S
+ mux_bottom_track_17.mux_l3_in_0_/S mem_bottom_track_17.scs8hd_dfxbp_1_2_/QN vgnd
+ vpwr scs8hd_dfxbp_1
Xmux_top_track_24.mux_l2_in_0_ mux_top_track_24.mux_l1_in_1_/X mux_top_track_24.mux_l1_in_0_/X
+ mux_top_track_24.mux_l2_in_2_/S mux_top_track_24.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_3.mux_l1_in_1__A0 chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l4_in_0__A0 mux_top_track_2.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_19_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_3__A0 bottom_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
XANTENNA__087__A _087_/A vgnd vpwr scs8hd_diode_2
X_071_ _071_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_2.mux_l2_in_1__S mux_top_track_2.mux_l2_in_2_/S vgnd vpwr scs8hd_diode_2
XFILLER_2_266 vpwr vgnd scs8hd_fill_2
XFILLER_2_211 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0__S mux_left_track_9.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_top_track_2.scs8hd_dfxbp_1_3_ prog_clk mux_top_track_2.mux_l3_in_1_/S mux_top_track_2.mux_l4_in_0_/S
+ mem_top_track_2.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_left_track_17.mux_l2_in_0_ mux_left_track_17.mux_l1_in_1_/X mux_left_track_17.mux_l1_in_0_/X
+ mux_left_track_17.mux_l2_in_1_/S mux_left_track_17.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_24.mux_l1_in_0__A0 chany_top_in[11] vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.mux_l1_in_3_ chany_bottom_in[4] chanx_right_in[13] mux_top_track_2.mux_l1_in_3_/S
+ mux_top_track_2.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_8.mux_l1_in_2__S mux_top_track_8.mux_l1_in_1_/S vgnd vpwr scs8hd_diode_2
Xmux_left_track_5.mux_l2_in_7_ _055_/HI left_top_grid_pin_49_ mux_left_track_5.mux_l2_in_7_/S
+ mux_left_track_5.mux_l2_in_7_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_2.mux_l1_in_3__A1 chanx_right_in[13] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_3__A0 chany_bottom_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_15_115 vpwr vgnd scs8hd_fill_2
XFILLER_15_126 vgnd vpwr scs8hd_decap_3
X_054_ _054_/HI _054_/LO vgnd vpwr scs8hd_conb_1
X_123_ _123_/A chany_top_out[12] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_3.mux_l2_in_0__A0 mux_left_track_3.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_0__A1 mux_top_track_4.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_4.scs8hd_buf_4_0_ mux_top_track_4.mux_l5_in_0_/X _133_/A vgnd vpwr
+ scs8hd_buf_1
Xmux_top_track_24.mux_l1_in_1_ chanx_right_in[18] chanx_right_in[9] mux_top_track_24.mux_l1_in_1_/S
+ mux_top_track_24.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_16.mux_l1_in_0__A0 top_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l3_in_2__A0 mux_bottom_track_5.mux_l2_in_5_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A1 chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0__A1 chany_top_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_3__D mux_right_track_24.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_129 vgnd vpwr scs8hd_fill_1
XFILLER_16_59 vgnd vpwr scs8hd_decap_3
XFILLER_32_36 vpwr vgnd scs8hd_fill_2
XFILLER_20_140 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_3_ _043_/HI chanx_left_in[12] mux_bottom_track_1.mux_l2_in_0_/S
+ mux_bottom_track_1.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_11_151 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_1_ chanx_right_in[8] chany_top_in[17] mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
X_106_ chany_top_in[8] chany_bottom_out[9] vgnd vpwr scs8hd_buf_2
X_037_ _037_/HI _037_/LO vgnd vpwr scs8hd_conb_1
XFILLER_19_240 vpwr vgnd scs8hd_fill_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XFILLER_34_243 vpwr vgnd scs8hd_fill_2
XFILLER_34_210 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_2__A0 left_top_grid_pin_46_ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l2_in_0_ mux_left_track_9.mux_l1_in_1_/X mux_left_track_9.mux_l1_in_0_/X
+ mux_left_track_9.mux_l2_in_1_/S mux_left_track_9.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_2.mux_l2_in_2__A1 mux_top_track_2.mux_l1_in_4_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_93 vpwr vgnd scs8hd_fill_2
XFILLER_27_36 vpwr vgnd scs8hd_fill_2
XFILLER_25_232 vgnd vpwr scs8hd_decap_3
XFILLER_40_224 vpwr vgnd scs8hd_fill_2
XFILLER_40_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.mux_l4_in_0__S mux_left_track_17.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_254 vpwr vgnd scs8hd_fill_2
XANTENNA__095__A _095_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_0_/S mux_right_track_0.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_158 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_5.mux_l4_in_1__A0 mux_bottom_track_5.mux_l3_in_3_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_1_/S mux_top_track_2.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_24.mux_l3_in_0_ mux_right_track_24.mux_l2_in_1_/X mux_right_track_24.mux_l2_in_0_/X
+ mux_right_track_24.mux_l3_in_0_/S mux_right_track_24.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_32.mux_l2_in_0__S mux_top_track_32.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_2.mux_l1_in_4__S mux_right_track_2.mux_l1_in_4_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l3_in_1__S mux_right_track_0.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l2_in_2__S mux_left_track_3.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_16 vpwr vgnd scs8hd_fill_2
XFILLER_1_106 vpwr vgnd scs8hd_fill_2
XFILLER_38_68 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__D mux_right_track_8.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_128 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_4_ chanx_left_in[1] bottom_left_grid_pin_40_ mux_bottom_track_1.mux_l1_in_0_/S
+ mux_bottom_track_1.mux_l1_in_4_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_4__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l3_in_1__A1 mux_top_track_2.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_235 vpwr vgnd scs8hd_fill_2
XFILLER_13_257 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l3_in_1__A0 mux_left_track_1.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_ chanx_right_in[6] chany_top_in[16] mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmem_left_track_5.scs8hd_dfxbp_1_3_ prog_clk mux_left_track_5.mux_l3_in_3_/S mux_left_track_5.mux_l4_in_0_/S
+ mem_left_track_5.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__D mux_bottom_track_25.mux_l4_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_5_94 vpwr vgnd scs8hd_fill_2
XFILLER_39_176 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_5.mux_l5_in_0__A0 mux_bottom_track_5.mux_l4_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_36 vpwr vgnd scs8hd_fill_2
XFILLER_40_25 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_1_ right_top_grid_pin_42_ chany_top_in[19] mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_track_1.mux_l4_in_0_ mux_bottom_track_1.mux_l3_in_1_/X mux_bottom_track_1.mux_l3_in_0_/X
+ mux_bottom_track_1.mux_l4_in_0_/S mux_bottom_track_1.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_2.mux_l2_in_1_ mux_top_track_2.mux_l1_in_3_/X mux_top_track_2.mux_l1_in_2_/X
+ mux_top_track_2.mux_l2_in_2_/S mux_top_track_2.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_right_track_24.mux_l2_in_1_ chany_bottom_in[9] mux_right_track_24.mux_l1_in_2_/X
+ mux_right_track_24.mux_l2_in_2_/S mux_right_track_24.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_1_19 vpwr vgnd scs8hd_fill_2
XFILLER_5_231 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_32.mux_l1_in_0__A0 chany_top_in[15] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_17.mux_l1_in_0_/S
+ mux_bottom_track_17.mux_l2_in_2_/S mem_bottom_track_17.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_3.mux_l1_in_1__A1 chany_top_in[19] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l4_in_0__A1 mux_top_track_2.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l4_in_0__A0 mux_left_track_1.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_3__A1 bottom_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
XFILLER_42_138 vpwr vgnd scs8hd_fill_2
XFILLER_42_116 vpwr vgnd scs8hd_fill_2
XFILLER_27_179 vpwr vgnd scs8hd_fill_2
XFILLER_27_146 vgnd vpwr scs8hd_decap_3
X_070_ chanx_right_in[4] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_4_3 vgnd vpwr scs8hd_decap_4
XFILLER_2_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_24.mux_l1_in_0__A0 top_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
XFILLER_18_113 vpwr vgnd scs8hd_fill_2
XFILLER_41_193 vpwr vgnd scs8hd_fill_2
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_33_149 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l2_in_3__A0 _035_/HI vgnd vpwr scs8hd_diode_2
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l1_in_0__S mux_bottom_track_1.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_top_track_2.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_2.mux_l2_in_2_/S mux_top_track_2.mux_l3_in_1_/S
+ mem_top_track_2.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_24.mux_l1_in_0__A1 chany_top_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_2_84 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.mux_l3_in_1_ mux_bottom_track_1.mux_l2_in_3_/X mux_bottom_track_1.mux_l2_in_2_/X
+ mux_bottom_track_1.mux_l3_in_1_/S mux_bottom_track_1.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_149 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.mux_l1_in_2_ chanx_right_in[4] chanx_right_in[3] mux_top_track_2.mux_l1_in_3_/S
+ mux_top_track_2.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_32_182 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_32.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_21_38 vpwr vgnd scs8hd_fill_2
Xmux_right_track_24.mux_l1_in_2_ chany_bottom_in[0] right_top_grid_pin_48_ mux_right_track_24.mux_l1_in_1_/S
+ mux_right_track_24.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__D mux_bottom_track_33.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_5.mux_l2_in_6_ left_top_grid_pin_48_ left_top_grid_pin_47_ mux_left_track_5.mux_l2_in_7_/S
+ mux_left_track_5.mux_l2_in_6_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_1.mux_l1_in_3__A1 chany_bottom_in[12] vgnd vpwr scs8hd_diode_2
XANTENNA__098__A chany_top_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_23_193 vpwr vgnd scs8hd_fill_2
X_122_ chany_bottom_in[12] chany_top_out[13] vgnd vpwr scs8hd_buf_2
X_053_ _053_/HI _053_/LO vgnd vpwr scs8hd_conb_1
XFILLER_11_60 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_3.mux_l2_in_0__A1 mux_left_track_3.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0__A1 top_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
Xmux_top_track_24.mux_l1_in_0_ top_left_grid_pin_40_ top_left_grid_pin_36_ mux_top_track_24.mux_l1_in_1_/S
+ mux_top_track_24.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_5.mux_l3_in_2__A1 mux_bottom_track_5.mux_l2_in_4_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_219 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__S mux_bottom_track_25.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_27 vpwr vgnd scs8hd_fill_2
XFILLER_20_174 vpwr vgnd scs8hd_fill_2
XFILLER_20_152 vgnd vpwr scs8hd_fill_1
XFILLER_28_274 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.mux_l2_in_2_ chanx_left_in[2] mux_bottom_track_1.mux_l1_in_4_/X
+ mux_bottom_track_1.mux_l2_in_0_/S mux_bottom_track_1.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_7_112 vpwr vgnd scs8hd_fill_2
XFILLER_7_123 vgnd vpwr scs8hd_decap_4
X_105_ chany_top_in[9] chany_bottom_out[10] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_24.mux_l3_in_0__S mux_top_track_24.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_0_ chany_top_in[8] chany_top_in[7] mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
X_036_ _036_/HI _036_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2__A0 bottom_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0__A0 top_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0__S mux_right_track_16.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_2__A1 mux_left_track_1.mux_l1_in_4_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l5_in_0__S mux_left_track_5.mux_l5_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_50 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_7__A0 _034_/HI vgnd vpwr scs8hd_diode_2
XFILLER_25_266 vpwr vgnd scs8hd_fill_2
XFILLER_40_258 vgnd vpwr scs8hd_decap_12
XFILLER_40_236 vgnd vpwr scs8hd_decap_12
XFILLER_4_115 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l4_in_1__A1 mux_bottom_track_5.mux_l3_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_258 vgnd vpwr scs8hd_fill_1
XFILLER_31_236 vpwr vgnd scs8hd_fill_2
XFILLER_31_225 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_16_211 vgnd vpwr scs8hd_fill_1
XFILLER_17_81 vpwr vgnd scs8hd_fill_2
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_91 vpwr vgnd scs8hd_fill_2
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_3_ bottom_left_grid_pin_38_ bottom_left_grid_pin_36_
+ mux_bottom_track_1.mux_l1_in_0_/S mux_bottom_track_1.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_17.mux_l2_in_1__A0 bottom_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
XFILLER_13_214 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l3_in_1__A1 mux_left_track_1.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_269 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_0_ chany_top_in[11] chany_top_in[6] mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
Xmem_left_track_5.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_5.mux_l2_in_7_/S mux_left_track_5.mux_l3_in_3_/S
+ mem_left_track_5.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_1.mux_l1_in_3__S mux_bottom_track_1.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_62 vgnd vpwr scs8hd_decap_3
XFILLER_8_273 vpwr vgnd scs8hd_fill_2
XFILLER_5_84 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_3__D mux_left_track_1.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_0_ chany_top_in[12] chany_top_in[2] mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l5_in_0__A1 mux_bottom_track_5.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_15 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.mux_l2_in_0_ mux_top_track_2.mux_l1_in_1_/X mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_2_/S mux_top_track_2.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_32.mux_l1_in_0__A0 top_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
XFILLER_10_206 vpwr vgnd scs8hd_fill_2
XFILLER_10_228 vpwr vgnd scs8hd_fill_2
Xmux_right_track_24.mux_l2_in_0_ mux_right_track_24.mux_l1_in_1_/X mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_2_/S mux_right_track_24.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_5.mux_l2_in_1__S mux_bottom_track_5.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_210 vpwr vgnd scs8hd_fill_2
XFILLER_5_254 vpwr vgnd scs8hd_fill_2
XFILLER_14_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_32.mux_l1_in_0__A1 chany_top_in[10] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_9.mux_l4_in_0_/S
+ mux_bottom_track_17.mux_l1_in_0_/S mem_bottom_track_17.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_17.mux_l3_in_0__A0 mux_bottom_track_17.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l4_in_0__A1 mux_left_track_1.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_158 vpwr vgnd scs8hd_fill_2
XFILLER_27_114 vpwr vgnd scs8hd_fill_2
XFILLER_2_224 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_24.mux_l1_in_0__A1 top_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
XFILLER_18_158 vgnd vpwr scs8hd_decap_4
XFILLER_18_136 vpwr vgnd scs8hd_fill_2
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XFILLER_25_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_3__A1 chanx_left_in[16] vgnd vpwr scs8hd_diode_2
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_top_track_2.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_2.mux_l1_in_3_/S mux_top_track_2.mux_l2_in_2_/S
+ mem_top_track_2.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_4.mux_l2_in_3__A0 chanx_right_in[5] vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.mux_l1_in_1_ top_left_grid_pin_41_ top_left_grid_pin_39_ mux_top_track_2.mux_l1_in_3_/S
+ mux_top_track_2.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ mux_bottom_track_1.mux_l3_in_1_/S mux_bottom_track_1.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_2_74 vgnd vpwr scs8hd_decap_4
XFILLER_2_41 vgnd vpwr scs8hd_decap_3
Xmux_right_track_24.mux_l1_in_1_ right_top_grid_pin_44_ chany_top_in[18] mux_right_track_24.mux_l1_in_1_/S
+ mux_right_track_24.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_24_128 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0__S mux_bottom_track_17.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0__A0 chany_top_in[8] vgnd vpwr scs8hd_diode_2
Xmux_left_track_5.mux_l2_in_5_ left_top_grid_pin_46_ left_top_grid_pin_45_ mux_left_track_5.mux_l2_in_7_/S
+ mux_left_track_5.mux_l2_in_5_/X vgnd vpwr scs8hd_mux2_1
X_121_ chany_bottom_in[13] chany_top_out[14] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_25.mux_l1_in_2__A0 bottom_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
X_052_ _052_/HI _052_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_16.mux_l4_in_0__S mux_top_track_16.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_209 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l1_in_0__S mux_left_track_5.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_253 vpwr vgnd scs8hd_fill_2
XFILLER_37_242 vpwr vgnd scs8hd_fill_2
XFILLER_37_231 vgnd vpwr scs8hd_fill_1
XFILLER_32_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0__S mux_right_track_8.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_25.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_track_25.mux_l3_in_1_/S
+ mux_bottom_track_25.mux_l4_in_0_/S mem_bottom_track_25.scs8hd_dfxbp_1_3_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_4.mux_l3_in_2__A0 mux_top_track_4.mux_l2_in_5_/X vgnd vpwr
+ scs8hd_diode_2
X_035_ _035_/HI _035_/LO vgnd vpwr scs8hd_conb_1
XFILLER_22_93 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_1_ mux_bottom_track_1.mux_l1_in_3_/X mux_bottom_track_1.mux_l1_in_2_/X
+ mux_bottom_track_1.mux_l2_in_0_/S mux_bottom_track_1.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
XFILLER_11_120 vpwr vgnd scs8hd_fill_2
X_104_ chany_top_in[10] chany_bottom_out[11] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2__A1 chanx_right_in[17] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0__A1 top_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_2__A0 chanx_left_in[11] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_2__A0 chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_6_190 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_4.mux_l2_in_7__A1 chanx_left_in[14] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_1__A0 bottom_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
XFILLER_40_204 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__D mux_left_track_3.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0__S mux_top_track_8.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_40_248 vgnd vpwr scs8hd_decap_6
XFILLER_4_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_4__S mux_bottom_track_5.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_204 vpwr vgnd scs8hd_fill_2
XFILLER_16_267 vgnd vpwr scs8hd_decap_8
XFILLER_3_193 vpwr vgnd scs8hd_fill_2
XFILLER_3_160 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l4_in_1__A0 mux_top_track_4.mux_l3_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_38_37 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_2_ bottom_left_grid_pin_34_ chanx_right_in[15] mux_bottom_track_1.mux_l1_in_0_/S
+ mux_bottom_track_1.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_17.mux_l2_in_1__A1 mux_bottom_track_17.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__D mux_bottom_track_17.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_248 vpwr vgnd scs8hd_fill_2
XFILLER_21_270 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l3_in_1__A0 mux_bottom_track_9.mux_l2_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_196 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l3_in_1__A0 mux_right_track_16.mux_l2_in_3_/X vgnd
+ vpwr scs8hd_diode_2
Xmem_left_track_5.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_5.mux_l1_in_0_/S mux_left_track_5.mux_l2_in_7_/S
+ mem_left_track_5.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_25.mux_l3_in_0__A0 mux_bottom_track_25.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_241 vgnd vpwr scs8hd_decap_4
XFILLER_12_270 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.scs8hd_buf_4_0__A mux_top_track_16.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_3__S mux_bottom_track_17.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_49 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l1_in_4__A0 left_top_grid_pin_45_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_32.mux_l1_in_0__A1 top_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
XFILLER_6_8 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_5.mux_l2_in_6__A0 chanx_left_in[7] vgnd vpwr scs8hd_diode_2
Xmux_left_track_5.mux_l3_in_3_ mux_left_track_5.mux_l2_in_7_/X mux_left_track_5.mux_l2_in_6_/X
+ mux_left_track_5.mux_l3_in_3_/S mux_left_track_5.mux_l3_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_14_50 vpwr vgnd scs8hd_fill_2
XFILLER_30_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_1__A0 chanx_right_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_5_200 vgnd vpwr scs8hd_fill_1
XFILLER_5_266 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l5_in_0__A0 mux_top_track_4.mux_l4_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l1_in_0__A0 chany_top_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_36_148 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l2_in_2__S mux_right_track_2.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l3_in_0__A1 mux_bottom_track_17.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l3_in_0__S mux_left_track_3.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_38 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_33.mux_l1_in_2__A0 chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l4_in_0__A0 mux_bottom_track_9.mux_l3_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l4_in_0__A0 mux_right_track_16.mux_l3_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_203 vpwr vgnd scs8hd_fill_2
XFILLER_2_258 vpwr vgnd scs8hd_fill_2
XFILLER_41_140 vpwr vgnd scs8hd_fill_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XFILLER_33_118 vpwr vgnd scs8hd_fill_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_26_192 vgnd vpwr scs8hd_decap_3
XFILLER_18_148 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_9.mux_l2_in_1__S mux_left_track_9.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_2.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_0.mux_l4_in_0_/S mux_top_track_2.mux_l1_in_3_/S
+ mem_top_track_2.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_3.mux_l2_in_3__A0 _053_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_3__A1 top_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.mux_l1_in_0_ top_left_grid_pin_37_ top_left_grid_pin_35_ mux_top_track_2.mux_l1_in_3_/S
+ mux_top_track_2.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_17.mux_l1_in_0__A1 chany_top_in[7] vgnd vpwr scs8hd_diode_2
Xmux_right_track_24.mux_l1_in_0_ chany_top_in[11] chany_top_in[9] mux_right_track_24.mux_l1_in_1_/S
+ mux_right_track_24.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_left_track_5.mux_l2_in_4_ left_top_grid_pin_44_ left_top_grid_pin_43_ mux_left_track_5.mux_l2_in_7_/S
+ mux_left_track_5.mux_l2_in_4_/X vgnd vpwr scs8hd_mux2_1
XFILLER_21_18 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__D mux_left_track_5.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l3_in_0__A0 mux_left_track_5.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_3__S mux_top_track_8.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
X_120_ chany_bottom_in[14] chany_top_out[15] vgnd vpwr scs8hd_buf_2
X_051_ _051_/HI _051_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_track_25.mux_l1_in_2__A1 chanx_right_in[18] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_2__D mux_top_track_24.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_7__S mux_bottom_track_5.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_51 vpwr vgnd scs8hd_fill_2
XFILLER_11_62 vpwr vgnd scs8hd_fill_2
XFILLER_11_95 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.scs8hd_buf_4_0__A mux_right_track_16.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_24.mux_l2_in_2__A0 chanx_left_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_14_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_33.mux_l2_in_1__A0 mux_bottom_track_33.mux_l1_in_3_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_5.mux_l5_in_0_ mux_left_track_5.mux_l4_in_1_/X mux_left_track_5.mux_l4_in_0_/X
+ mux_left_track_5.mux_l5_in_0_/S mux_left_track_5.mux_l5_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_37_276 vgnd vpwr scs8hd_fill_1
XFILLER_37_210 vpwr vgnd scs8hd_fill_2
XFILLER_20_187 vpwr vgnd scs8hd_fill_2
XFILLER_20_154 vgnd vpwr scs8hd_decap_4
XFILLER_28_254 vpwr vgnd scs8hd_fill_2
XFILLER_28_210 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l3_in_2__A1 mux_top_track_4.mux_l2_in_4_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_25.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_25.mux_l2_in_3_/S
+ mux_bottom_track_25.mux_l3_in_1_/S mem_bottom_track_25.scs8hd_dfxbp_1_2_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.mux_l2_in_2__A0 chanx_left_in[8] vgnd vpwr scs8hd_diode_2
X_034_ _034_/HI _034_/LO vgnd vpwr scs8hd_conb_1
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_0_/S mux_bottom_track_1.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_7_158 vpwr vgnd scs8hd_fill_2
X_103_ _103_/A chany_bottom_out[12] vgnd vpwr scs8hd_buf_2
XFILLER_11_176 vgnd vpwr scs8hd_fill_1
XFILLER_19_276 vgnd vpwr scs8hd_fill_1
XFILLER_19_254 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l2_in_2__A1 chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_14_7 vgnd vpwr scs8hd_fill_1
XFILLER_8_41 vgnd vpwr scs8hd_decap_3
XFILLER_8_63 vgnd vpwr scs8hd_decap_3
XFILLER_8_85 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_16.mux_l2_in_2__A1 chany_bottom_in[17] vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.scs8hd_buf_4_0_ mux_left_track_1.mux_l4_in_0_/X _075_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_bottom_track_25.mux_l2_in_1__A1 mux_bottom_track_25.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l1_in_1__S mux_bottom_track_33.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_33.scs8hd_dfxbp_1_2__D mux_left_track_33.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_128 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_24.mux_l3_in_1__A0 mux_right_track_24.mux_l2_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l3_in_0__A0 mux_bottom_track_33.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_224 vpwr vgnd scs8hd_fill_2
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_5.mux_l4_in_1_ mux_left_track_5.mux_l3_in_3_/X mux_left_track_5.mux_l3_in_2_/X
+ mux_left_track_5.mux_l4_in_0_/S mux_left_track_5.mux_l4_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_24.mux_l1_in_1__S mux_right_track_24.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_249 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l4_in_1__A1 mux_top_track_4.mux_l3_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l3_in_1__A0 mux_top_track_16.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_1_ chanx_right_in[12] chanx_right_in[2] mux_bottom_track_1.mux_l1_in_0_/S
+ mux_bottom_track_1.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_13_227 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l3_in_1__A1 mux_bottom_track_9.mux_l2_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_33.mux_l1_in_0__A0 chany_top_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l3_in_1__A1 mux_right_track_16.mux_l2_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__D mux_top_track_0.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XFILLER_0_175 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_4.mux_l5_in_0__S mux_right_track_4.mux_l5_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_5.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_3.mux_l4_in_0_/S mux_left_track_5.mux_l1_in_0_/S
+ mem_left_track_5.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_25.mux_l3_in_0__A1 mux_bottom_track_25.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_253 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_32.mux_l1_in_3__A0 _033_/HI vgnd vpwr scs8hd_diode_2
XFILLER_5_42 vpwr vgnd scs8hd_fill_2
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_39_146 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_24.mux_l4_in_0__A0 mux_right_track_24.mux_l3_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l1_in_4__A1 left_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_4__D mux_left_track_5.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_6__A1 chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0__A0 chany_top_in[4] vgnd vpwr scs8hd_diode_2
Xmux_left_track_5.mux_l3_in_2_ mux_left_track_5.mux_l2_in_5_/X mux_left_track_5.mux_l2_in_4_/X
+ mux_left_track_5.mux_l3_in_3_/S mux_left_track_5.mux_l3_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_38_190 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_5.mux_l2_in_1__A1 chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_14_84 vgnd vpwr scs8hd_fill_1
XFILLER_5_234 vpwr vgnd scs8hd_fill_2
XFILLER_39_70 vgnd vpwr scs8hd_decap_4
XFILLER_36_127 vgnd vpwr scs8hd_decap_4
XFILLER_36_105 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_16.mux_l4_in_0__A0 mux_top_track_16.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA__101__A chany_top_in[13] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l5_in_0__A1 mux_top_track_4.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l1_in_0__A1 chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_35_160 vgnd vpwr scs8hd_decap_4
XFILLER_35_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_33.mux_l1_in_2__A1 bottom_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l4_in_0__A1 mux_bottom_track_9.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l4_in_0__A1 mux_right_track_16.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_83 vgnd vpwr scs8hd_decap_3
XFILLER_41_163 vgnd vpwr scs8hd_fill_1
XPHY_72 vgnd vpwr scs8hd_decap_3
XFILLER_33_108 vpwr vgnd scs8hd_fill_2
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_26_171 vpwr vgnd scs8hd_fill_2
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_2__A0 right_top_grid_pin_46_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l2_in_3__A1 left_top_grid_pin_49_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_1__S mux_bottom_track_1.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_10 vpwr vgnd scs8hd_fill_2
XFILLER_1_270 vpwr vgnd scs8hd_fill_2
XFILLER_32_163 vgnd vpwr scs8hd_decap_3
Xmux_left_track_5.mux_l2_in_3_ left_top_grid_pin_42_ chany_bottom_in[14] mux_left_track_5.mux_l2_in_7_/S
+ mux_left_track_5.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_5.mux_l3_in_0__A1 mux_left_track_5.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_24.mux_l2_in_2__A0 chanx_left_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_23_152 vpwr vgnd scs8hd_fill_2
XFILLER_15_119 vgnd vpwr scs8hd_decap_3
X_050_ _050_/HI _050_/LO vgnd vpwr scs8hd_conb_1
XFILLER_11_30 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_24.mux_l2_in_2__A1 chany_bottom_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_14_163 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_33.mux_l2_in_1__A1 mux_bottom_track_33.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_35_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_1__S mux_bottom_track_25.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_28_266 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_0.mux_l2_in_1__A0 mux_right_track_0.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_25.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_25.mux_l1_in_0_/S
+ mux_bottom_track_25.mux_l2_in_3_/S mem_bottom_track_25.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_17.mux_l1_in_1__S mux_left_track_17.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_155 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_2__A1 chanx_left_in[7] vgnd vpwr scs8hd_diode_2
X_033_ _033_/HI _033_/LO vgnd vpwr scs8hd_conb_1
XFILLER_22_84 vpwr vgnd scs8hd_fill_2
X_102_ chany_top_in[12] chany_bottom_out[13] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__D mux_top_track_2.mux_l1_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_247 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_1__S mux_right_track_16.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_19_266 vpwr vgnd scs8hd_fill_2
XFILLER_19_233 vgnd vpwr scs8hd_fill_1
XFILLER_8_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_24.mux_l3_in_1__A0 mux_top_track_24.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_170 vgnd vpwr scs8hd_fill_1
XFILLER_27_29 vgnd vpwr scs8hd_decap_4
XFILLER_25_214 vgnd vpwr scs8hd_decap_3
XFILLER_40_228 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l1_in_0__S mux_left_track_1.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__D mux_right_track_32.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_24.mux_l3_in_1__A1 mux_right_track_24.mux_l2_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_2__A0 chanx_left_in[11] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l3_in_0__A1 mux_bottom_track_33.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_31_217 vpwr vgnd scs8hd_fill_2
XFILLER_16_203 vpwr vgnd scs8hd_fill_2
XFILLER_16_247 vpwr vgnd scs8hd_fill_2
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_5.mux_l4_in_0_ mux_left_track_5.mux_l3_in_1_/X mux_left_track_5.mux_l3_in_0_/X
+ mux_left_track_5.mux_l4_in_0_/S mux_left_track_5.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_4.mux_l1_in_0__S mux_right_track_4.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_173 vgnd vpwr scs8hd_decap_4
XANTENNA__104__A chany_top_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2__S mux_top_track_0.mux_l1_in_1_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l3_in_0__A0 mux_right_track_0.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_228 vpwr vgnd scs8hd_fill_2
XFILLER_22_206 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_0_ chany_top_in[12] chany_top_in[2] mux_bottom_track_1.mux_l1_in_0_/S
+ mux_bottom_track_1.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_16.mux_l3_in_1__A1 mux_top_track_16.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_13_217 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_32.mux_l1_in_3__A0 _040_/HI vgnd vpwr scs8hd_diode_2
XFILLER_13_239 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_4.mux_l2_in_0__S mux_top_track_4.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_33.mux_l1_in_0__A1 chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_28_50 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.scs8hd_buf_4_0__A mux_left_track_3.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_24.mux_l4_in_0__A0 mux_top_track_24.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__D mux_left_track_9.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_32.mux_l1_in_3__A1 chanx_left_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_8_265 vpwr vgnd scs8hd_fill_2
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XFILLER_12_250 vpwr vgnd scs8hd_fill_2
XFILLER_39_114 vpwr vgnd scs8hd_fill_2
XFILLER_39_103 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_32.scs8hd_dfxbp_1_0__D mux_right_track_24.mux_l4_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_98 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_24.mux_l4_in_0__A1 mux_right_track_24.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l3_in_1__A0 mux_top_track_8.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l1_in_0__A1 chany_top_in[0] vgnd vpwr scs8hd_diode_2
Xmux_left_track_5.mux_l3_in_1_ mux_left_track_5.mux_l2_in_3_/X mux_left_track_5.mux_l2_in_2_/X
+ mux_left_track_5.mux_l3_in_3_/S mux_left_track_5.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_30_40 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_5.mux_l3_in_2__S mux_bottom_track_5.mux_l3_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_41 vgnd vpwr scs8hd_decap_3
XFILLER_14_63 vgnd vpwr scs8hd_decap_4
XFILLER_30_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l4_in_0__A1 mux_top_track_16.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_6__A0 chanx_left_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_19_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l4_in_0__S mux_bottom_track_9.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_7 vgnd vpwr scs8hd_fill_1
XPHY_84 vgnd vpwr scs8hd_decap_3
XFILLER_41_197 vpwr vgnd scs8hd_fill_2
XFILLER_41_175 vpwr vgnd scs8hd_fill_2
XFILLER_41_153 vgnd vpwr scs8hd_decap_4
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_40 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_1__A0 chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XPHY_40 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_72 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_2__A1 right_top_grid_pin_44_ vgnd vpwr scs8hd_diode_2
XFILLER_37_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__D mux_top_track_2.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA__112__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l4_in_0__A0 mux_top_track_8.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_88 vgnd vpwr scs8hd_fill_1
XFILLER_32_186 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l3_in_1__S mux_bottom_track_17.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_5.mux_l2_in_2_ chany_bottom_in[5] chany_bottom_in[1] mux_left_track_5.mux_l2_in_7_/S
+ mux_left_track_5.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
Xmux_left_track_25.mux_l2_in_3_ _052_/HI left_top_grid_pin_48_ mux_left_track_25.mux_l2_in_3_/S
+ mux_left_track_25.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_3__D mux_bottom_track_1.mux_l3_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_24.mux_l2_in_2__A1 chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_3__S mux_left_track_1.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_197 vpwr vgnd scs8hd_fill_2
XFILLER_23_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__D mux_left_track_9.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_131 vgnd vpwr scs8hd_decap_3
XANTENNA__107__A _107_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_186 vpwr vgnd scs8hd_fill_2
XFILLER_14_197 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l2_in_2__A0 left_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l3_in_0__S mux_right_track_2.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_234 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_1__S mux_left_track_5.mux_l2_in_7_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_123 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_1__A1 mux_right_track_0.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0__A0 mux_left_track_9.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_234 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_25.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_17.mux_l4_in_0_/S
+ mux_bottom_track_25.mux_l1_in_0_/S mem_bottom_track_25.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_8.mux_l2_in_1__S mux_right_track_8.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_116 vpwr vgnd scs8hd_fill_2
XFILLER_7_127 vgnd vpwr scs8hd_fill_1
X_101_ chany_top_in[13] chany_bottom_out[14] vgnd vpwr scs8hd_buf_2
XFILLER_11_112 vpwr vgnd scs8hd_fill_2
XFILLER_11_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_4.mux_l2_in_3__S mux_top_track_4.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l4_in_0__S mux_top_track_2.mux_l4_in_0_/S vgnd vpwr scs8hd_diode_2
X_032_ _032_/HI _032_/LO vgnd vpwr scs8hd_conb_1
XFILLER_7_149 vpwr vgnd scs8hd_fill_2
XFILLER_19_212 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_3__D mux_left_track_17.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1__A0 chanx_right_in[12] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_24.mux_l3_in_1__A1 mux_top_track_24.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_237 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l3_in_1__S mux_top_track_8.mux_l3_in_1_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_2__A1 chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l3_in_1__A0 mux_left_track_17.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_259 vpwr vgnd scs8hd_fill_2
XFILLER_17_41 vpwr vgnd scs8hd_fill_2
XFILLER_17_85 vpwr vgnd scs8hd_fill_2
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_95 vpwr vgnd scs8hd_fill_2
XFILLER_33_62 vgnd vpwr scs8hd_decap_4
XFILLER_3_152 vpwr vgnd scs8hd_fill_2
Xmux_left_track_25.mux_l4_in_0_ mux_left_track_25.mux_l3_in_1_/X mux_left_track_25.mux_l3_in_0_/X
+ mux_left_track_25.mux_l4_in_0_/S mux_left_track_25.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__120__A chany_bottom_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_12_6 vpwr vgnd scs8hd_fill_2
XFILLER_30_251 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l3_in_0__A1 mux_right_track_0.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_218 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.scs8hd_buf_4_0__A mux_right_track_2.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_32.mux_l1_in_3__A1 chanx_left_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0__A0 mux_bottom_track_1.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_24.mux_l4_in_0__A1 mux_top_track_24.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_84 vpwr vgnd scs8hd_fill_2
XFILLER_28_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_4__A0 left_top_grid_pin_44_ vgnd vpwr scs8hd_diode_2
XFILLER_12_262 vpwr vgnd scs8hd_fill_2
XANTENNA__115__A _115_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_3__D mux_top_track_4.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_32.mux_l1_in_2__S mux_right_track_32.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_88 vgnd vpwr scs8hd_fill_1
XFILLER_10_3 vgnd vpwr scs8hd_decap_4
XFILLER_40_19 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l4_in_0__A0 mux_left_track_17.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l3_in_1__A1 mux_top_track_8.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_3_/S mux_left_track_5.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__D mux_bottom_track_3.mux_l2_in_3_/S
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_25.mux_l3_in_1_ mux_left_track_25.mux_l2_in_3_/X mux_left_track_25.mux_l2_in_2_/X
+ mux_left_track_25.mux_l3_in_0_/S mux_left_track_25.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_5_214 vpwr vgnd scs8hd_fill_2
XFILLER_5_258 vpwr vgnd scs8hd_fill_2
XFILLER_14_97 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_29_192 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_6__A1 chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_4__S mux_left_track_5.mux_l2_in_7_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_4
XFILLER_35_151 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_5.mux_l3_in_3__A0 mux_left_track_5.mux_l2_in_7_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_228 vpwr vgnd scs8hd_fill_2
XFILLER_26_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_6__S mux_top_track_4.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.mux_l2_in_2__A0 left_top_grid_pin_44_ vgnd vpwr scs8hd_diode_2
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XFILLER_26_184 vpwr vgnd scs8hd_fill_2
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_25_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_1__A1 chany_top_in[16] vgnd vpwr scs8hd_diode_2
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_16.mux_l1_in_1__S mux_top_track_16.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_62 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l4_in_0__A1 mux_top_track_8.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_78 vgnd vpwr scs8hd_fill_1
XFILLER_2_23 vpwr vgnd scs8hd_fill_2
XFILLER_32_121 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l2_in_1_ chanx_right_in[14] chanx_right_in[5] mux_left_track_5.mux_l2_in_7_/S
+ mux_left_track_5.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_left_track_25.mux_l2_in_2_ left_top_grid_pin_44_ chany_bottom_in[18] mux_left_track_25.mux_l2_in_3_/S
+ mux_left_track_25.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_24.scs8hd_buf_4_0__A mux_top_track_24.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_84 vpwr vgnd scs8hd_fill_2
XFILLER_36_73 vpwr vgnd scs8hd_fill_2
XFILLER_14_143 vpwr vgnd scs8hd_fill_2
XANTENNA__123__A _123_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_2__A1 chany_bottom_in[17] vgnd vpwr scs8hd_diode_2
Xmux_top_track_32.mux_l1_in_3_ _040_/HI chanx_left_in[10] mux_top_track_32.mux_l1_in_0_/S
+ mux_top_track_32.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_20_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.mux_l3_in_1__A0 mux_left_track_25.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0__A1 mux_left_track_9.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_224 vpwr vgnd scs8hd_fill_2
X_031_ _031_/HI _031_/LO vgnd vpwr scs8hd_conb_1
XFILLER_22_53 vpwr vgnd scs8hd_fill_2
X_100_ chany_top_in[14] chany_bottom_out[15] vgnd vpwr scs8hd_buf_2
XFILLER_11_168 vpwr vgnd scs8hd_fill_2
XFILLER_11_179 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.scs8hd_buf_4_0_ mux_top_track_16.mux_l4_in_0_/X _127_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_bottom_track_3.mux_l1_in_2__S mux_bottom_track_3.mux_l1_in_4_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__118__A chany_bottom_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1__A1 chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_8_11 vgnd vpwr scs8hd_fill_1
XFILLER_6_194 vgnd vpwr scs8hd_fill_1
XFILLER_10_190 vpwr vgnd scs8hd_fill_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.scs8hd_buf_4_0__A mux_bottom_track_1.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l3_in_1__A1 mux_left_track_17.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__D mux_bottom_track_5.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_25.mux_l1_in_2__S mux_left_track_25.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_33.mux_l1_in_3__A0 _054_/HI vgnd vpwr scs8hd_diode_2
XFILLER_3_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.mux_l4_in_0__A0 mux_left_track_25.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_24.mux_l2_in_2__S mux_right_track_24.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_7__S mux_left_track_5.mux_l2_in_7_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_24.scs8hd_buf_4_0__A mux_right_track_24.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_274 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__D mux_right_track_16.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0__A1 mux_bottom_track_1.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_32.mux_l3_in_0_ mux_top_track_32.mux_l2_in_1_/X mux_top_track_32.mux_l2_in_0_/X
+ mux_top_track_32.mux_l3_in_0_/S mux_top_track_32.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_3__A0 chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_4__A1 left_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
XFILLER_12_274 vgnd vpwr scs8hd_fill_1
XFILLER_5_67 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_33.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_33.mux_l2_in_1_/S
+ mux_bottom_track_33.mux_l3_in_0_/S mem_bottom_track_33.scs8hd_dfxbp_1_2_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA__131__A _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0__A0 chany_top_in[14] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0__S mux_right_track_0.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_3_ _042_/HI chanx_left_in[16] mux_top_track_8.mux_l2_in_1_/S
+ mux_top_track_8.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_17.mux_l4_in_0__A1 mux_left_track_17.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_193 vgnd vpwr scs8hd_fill_1
XFILLER_14_10 vpwr vgnd scs8hd_fill_2
XFILLER_14_87 vpwr vgnd scs8hd_fill_2
Xmux_left_track_25.mux_l3_in_0_ mux_left_track_25.mux_l2_in_1_/X mux_left_track_25.mux_l2_in_0_/X
+ mux_left_track_25.mux_l3_in_0_/S mux_left_track_25.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_30_97 vpwr vgnd scs8hd_fill_2
XFILLER_39_95 vpwr vgnd scs8hd_fill_2
XFILLER_39_40 vpwr vgnd scs8hd_fill_2
XFILLER_29_171 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0__S mux_top_track_0.mux_l2_in_2_/S vgnd vpwr scs8hd_diode_2
XANTENNA__126__A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_4_270 vpwr vgnd scs8hd_fill_2
Xmux_top_track_32.mux_l2_in_1_ mux_top_track_32.mux_l1_in_3_/X mux_top_track_32.mux_l1_in_2_/X
+ mux_top_track_32.mux_l2_in_1_/S mux_top_track_32.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_2.mux_l2_in_2__A0 chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_2_207 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_5.mux_l3_in_3__A1 mux_left_track_5.mux_l2_in_6_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_41_30 vpwr vgnd scs8hd_fill_2
XPHY_75 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_25.mux_l2_in_2__A1 chany_bottom_in[18] vgnd vpwr scs8hd_diode_2
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_41_85 vpwr vgnd scs8hd_fill_2
XFILLER_2_46 vgnd vpwr scs8hd_decap_3
XFILLER_32_199 vpwr vgnd scs8hd_fill_2
XFILLER_17_152 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__D mux_top_track_8.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_5.mux_l2_in_0_ chany_top_in[15] mux_left_track_5.mux_l1_in_0_/X mux_left_track_5.mux_l2_in_7_/S
+ mux_left_track_5.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_left_track_25.mux_l2_in_1_ chany_bottom_in[11] mux_left_track_25.mux_l1_in_2_/X
+ mux_left_track_25.mux_l2_in_3_/S mux_left_track_25.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_111 vpwr vgnd scs8hd_fill_2
XFILLER_23_100 vpwr vgnd scs8hd_fill_2
Xmux_top_track_24.scs8hd_buf_4_0_ mux_top_track_24.mux_l4_in_0_/X _123_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_4__D mux_bottom_track_5.mux_l4_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_6 vpwr vgnd scs8hd_fill_2
XFILLER_11_55 vgnd vpwr scs8hd_decap_3
XFILLER_11_66 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_5.mux_l4_in_0__S mux_bottom_track_5.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l4_in_0_ mux_top_track_8.mux_l3_in_1_/X mux_top_track_8.mux_l3_in_0_/X
+ mux_top_track_8.mux_l4_in_0_/S mux_top_track_8.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_42_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l3_in_1__A0 mux_right_track_2.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_32.mux_l1_in_2_ chanx_left_in[1] chany_bottom_in[10] mux_top_track_32.mux_l1_in_0_/S
+ mux_top_track_32.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_37_214 vpwr vgnd scs8hd_fill_2
XFILLER_20_158 vgnd vpwr scs8hd_fill_1
XFILLER_20_136 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.scs8hd_dfxbp_1_3_ prog_clk mux_top_track_16.mux_l3_in_0_/S mux_top_track_16.mux_l4_in_0_/S
+ mem_top_track_16.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_170 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_25.mux_l3_in_1__A1 mux_left_track_25.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_258 vpwr vgnd scs8hd_fill_2
X_030_ _030_/HI _030_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_17.mux_l2_in_2__S mux_left_track_17.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_65 vpwr vgnd scs8hd_fill_2
XFILLER_22_32 vpwr vgnd scs8hd_fill_2
XFILLER_22_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_34_206 vpwr vgnd scs8hd_fill_2
XFILLER_19_258 vgnd vpwr scs8hd_fill_1
XFILLER_19_236 vpwr vgnd scs8hd_fill_2
XFILLER_8_23 vpwr vgnd scs8hd_fill_2
XANTENNA__134__A _134_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_25.mux_l1_in_2_ chany_bottom_in[9] chanx_right_in[18] mux_left_track_25.mux_l1_in_1_/S
+ mux_left_track_25.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_33_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l1_in_3__S mux_right_track_0.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_209 vpwr vgnd scs8hd_fill_2
XFILLER_33_272 vgnd vpwr scs8hd_decap_4
Xmux_top_track_8.mux_l3_in_1_ mux_top_track_8.mux_l2_in_3_/X mux_top_track_8.mux_l2_in_2_/X
+ mux_top_track_8.mux_l3_in_1_/S mux_top_track_8.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_1.mux_l2_in_1__S mux_left_track_1.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1__A0 top_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
XFILLER_16_228 vpwr vgnd scs8hd_fill_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l4_in_0__A0 mux_right_track_2.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_33.mux_l1_in_3__A1 left_top_grid_pin_49_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_1__S mux_right_track_4.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_3__S mux_top_track_0.mux_l2_in_2_/S vgnd vpwr scs8hd_diode_2
XANTENNA__129__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l4_in_0__A1 mux_left_track_25.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.scs8hd_buf_4_0_ mux_bottom_track_3.mux_l4_in_0_/X _114_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_0_90 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_0_113 vgnd vpwr scs8hd_decap_4
XFILLER_0_179 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_4.mux_l3_in_1__S mux_top_track_4.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_3__A1 right_top_grid_pin_49_ vgnd vpwr scs8hd_diode_2
XFILLER_8_224 vpwr vgnd scs8hd_fill_2
XFILLER_5_46 vpwr vgnd scs8hd_fill_2
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_33.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_33.mux_l1_in_0_/S
+ mux_bottom_track_33.mux_l2_in_1_/S mem_bottom_track_33.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
Xmux_top_track_8.mux_l2_in_2_ chanx_left_in[11] chanx_left_in[6] mux_top_track_8.mux_l2_in_1_/S
+ mux_top_track_8.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_4.mux_l2_in_0__A1 mux_right_track_4.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0__A0 mux_top_track_0.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__D mux_bottom_track_25.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_65 vgnd vpwr scs8hd_decap_4
XFILLER_5_227 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A0 chany_top_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_5_238 vgnd vpwr scs8hd_decap_4
XFILLER_35_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l2_in_2__A1 mux_right_track_2.mux_l1_in_4_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_32.mux_l2_in_0_ mux_top_track_32.mux_l1_in_1_/X mux_top_track_32.mux_l1_in_0_/X
+ mux_top_track_32.mux_l2_in_1_/S mux_top_track_32.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_32.scs8hd_buf_4_0_ mux_top_track_32.mux_l3_in_0_/X _119_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_18_109 vpwr vgnd scs8hd_fill_2
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_33.mux_l1_in_0__S mux_left_track_33.mux_l1_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_274 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_3.mux_l1_in_2__A0 bottom_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XFILLER_32_145 vpwr vgnd scs8hd_fill_2
XFILLER_32_101 vgnd vpwr scs8hd_decap_3
XFILLER_17_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_32.mux_l2_in_0__S mux_right_track_32.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ mux_left_track_25.mux_l2_in_3_/S mux_left_track_25.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_123 vgnd vpwr scs8hd_decap_3
Xmux_right_track_32.mux_l1_in_3_ _033_/HI chanx_left_in[10] mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_9.mux_l2_in_3__A0 _028_/HI vgnd vpwr scs8hd_diode_2
XFILLER_11_34 vpwr vgnd scs8hd_fill_2
XFILLER_36_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_4__S mux_right_track_4.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_24.mux_l1_in_2__S mux_top_track_24.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l3_in_1__A1 mux_right_track_2.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_6 vpwr vgnd scs8hd_fill_2
Xmux_top_track_32.mux_l1_in_1_ chanx_right_in[10] chanx_right_in[0] mux_top_track_32.mux_l1_in_0_/S
+ mux_top_track_32.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_1.mux_l1_in_4__A0 chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l3_in_2__S mux_left_track_5.mux_l3_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_148 vpwr vgnd scs8hd_fill_2
XFILLER_9_193 vgnd vpwr scs8hd_decap_4
Xmem_top_track_16.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_16.mux_l2_in_0_/S mux_top_track_16.mux_l3_in_0_/S
+ mem_top_track_16.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_2__D mux_top_track_32.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l2_in_1__A0 mux_bottom_track_3.mux_l1_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_88 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l1_in_0_ chany_top_in[14] chany_top_in[5] mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_27_270 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_9.mux_l4_in_0__S mux_left_track_9.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_46 vpwr vgnd scs8hd_fill_2
XFILLER_8_68 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.scs8hd_buf_4_0__A mux_bottom_track_9.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_25.mux_l1_in_1_ chanx_right_in[9] chany_top_in[18] mux_left_track_25.mux_l1_in_1_/S
+ mux_left_track_25.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
X_089_ chanx_left_in[5] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_6_163 vgnd vpwr scs8hd_decap_4
Xmux_top_track_8.mux_l3_in_0_ mux_top_track_8.mux_l2_in_1_/X mux_top_track_8.mux_l2_in_0_/X
+ mux_top_track_8.mux_l3_in_1_/S mux_top_track_8.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__060__A chanx_right_in[14] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1__A1 top_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XFILLER_16_207 vgnd vpwr scs8hd_decap_4
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_2.mux_l4_in_0__A1 mux_right_track_2.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_251 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__D mux_bottom_track_9.mux_l2_in_3_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_3__A0 _043_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_7__A0 _055_/HI vgnd vpwr scs8hd_diode_2
XFILLER_30_210 vpwr vgnd scs8hd_fill_2
Xmux_right_track_32.mux_l3_in_0_ mux_right_track_32.mux_l2_in_1_/X mux_right_track_32.mux_l2_in_0_/X
+ mux_right_track_32.mux_l3_in_0_/S mux_right_track_32.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_top_track_0.scs8hd_dfxbp_1_3_ prog_clk mux_top_track_0.mux_l3_in_1_/S mux_top_track_0.mux_l4_in_0_/S
+ mem_top_track_0.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_3.mux_l3_in_0__A0 mux_bottom_track_3.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_254 vgnd vpwr scs8hd_decap_3
XFILLER_28_54 vpwr vgnd scs8hd_fill_2
XFILLER_28_32 vgnd vpwr scs8hd_decap_3
XFILLER_28_10 vpwr vgnd scs8hd_fill_2
XFILLER_0_125 vgnd vpwr scs8hd_decap_3
XFILLER_0_147 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_33.mux_l1_in_3__S mux_left_track_33.mux_l1_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_210 vpwr vgnd scs8hd_fill_2
Xmem_right_track_4.scs8hd_dfxbp_1_4_ prog_clk mux_right_track_4.mux_l4_in_0_/S mux_right_track_4.mux_l5_in_0_/S
+ mem_right_track_4.scs8hd_dfxbp_1_4_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_3.mux_l2_in_0__S mux_bottom_track_3.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_247 vpwr vgnd scs8hd_fill_2
XFILLER_8_269 vpwr vgnd scs8hd_fill_2
XFILLER_12_254 vpwr vgnd scs8hd_fill_2
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_33.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_25.mux_l4_in_0_/S
+ mux_bottom_track_33.mux_l1_in_0_/S mem_bottom_track_33.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_39_118 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l2_in_1_ chany_bottom_in[16] mux_top_track_8.mux_l1_in_2_/X mux_top_track_8.mux_l2_in_1_/S
+ mux_top_track_8.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_0.scs8hd_buf_4_0_ mux_top_track_0.mux_l4_in_0_/X _135_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__D mux_right_track_0.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0__A1 mux_top_track_0.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l3_in_0__S mux_bottom_track_33.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_38_162 vgnd vpwr scs8hd_decap_3
XFILLER_38_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1__S mux_bottom_track_9.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_11 vgnd vpwr scs8hd_decap_3
XFILLER_14_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.mux_l2_in_0__S mux_left_track_25.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_88 vpwr vgnd scs8hd_fill_2
Xmux_right_track_32.mux_l2_in_1_ mux_right_track_32.mux_l1_in_3_/X mux_right_track_32.mux_l1_in_2_/X
+ mux_right_track_32.mux_l2_in_0_/S mux_right_track_32.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A1 chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_39_53 vpwr vgnd scs8hd_fill_2
XFILLER_29_184 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_4.mux_l2_in_7__S mux_right_track_4.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_24.mux_l3_in_0__S mux_right_track_24.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0__A0 chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_6_90 vpwr vgnd scs8hd_fill_2
XFILLER_41_179 vpwr vgnd scs8hd_fill_2
XFILLER_41_102 vgnd vpwr scs8hd_decap_4
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_154 vpwr vgnd scs8hd_fill_2
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
Xmux_top_track_8.mux_l1_in_2_ chany_bottom_in[6] chanx_right_in[16] mux_top_track_8.mux_l1_in_1_/S
+ mux_top_track_8.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_3.mux_l1_in_2__A1 chanx_right_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_1_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_2__S mux_top_track_16.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_32_113 vpwr vgnd scs8hd_fill_2
XFILLER_32_168 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_23_179 vpwr vgnd scs8hd_fill_2
XFILLER_23_146 vgnd vpwr scs8hd_decap_4
XFILLER_23_135 vpwr vgnd scs8hd_fill_2
Xmux_right_track_32.mux_l1_in_2_ chany_bottom_in[19] chany_bottom_in[10] mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__063__A _063_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_13 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_3__A1 left_top_grid_pin_46_ vgnd vpwr scs8hd_diode_2
XFILLER_36_54 vpwr vgnd scs8hd_fill_2
XFILLER_36_32 vpwr vgnd scs8hd_fill_2
XFILLER_36_21 vgnd vpwr scs8hd_decap_4
XFILLER_14_113 vpwr vgnd scs8hd_fill_2
XFILLER_22_190 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_2.mux_l1_in_1__S mux_top_track_2.mux_l1_in_3_/S vgnd vpwr scs8hd_diode_2
Xmem_left_track_3.scs8hd_dfxbp_1_3_ prog_clk mux_left_track_3.mux_l3_in_1_/S mux_left_track_3.mux_l4_in_0_/S
+ mem_left_track_3.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_37_238 vpwr vgnd scs8hd_fill_2
XFILLER_37_227 vgnd vpwr scs8hd_decap_4
Xmux_top_track_32.mux_l1_in_0_ top_left_grid_pin_41_ top_left_grid_pin_37_ mux_top_track_32.mux_l1_in_0_/S
+ mux_top_track_32.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_37_249 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_4__A1 bottom_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_16.mux_l1_in_2_/S mux_top_track_16.mux_l2_in_0_/S
+ mem_top_track_16.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_36_260 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_5.scs8hd_dfxbp_1_4_ prog_clk mux_bottom_track_5.mux_l4_in_0_/S mux_bottom_track_5.mux_l5_in_0_/S
+ mem_bottom_track_5.scs8hd_dfxbp_1_4_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA__058__A chanx_right_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_22_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_1__A1 mux_bottom_track_3.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_116 vpwr vgnd scs8hd_fill_2
XFILLER_42_252 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_34_219 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_3.mux_l2_in_3__S mux_bottom_track_3.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.scs8hd_buf_4_0__A mux_top_track_4.mux_l5_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_25.mux_l1_in_0_ chany_top_in[9] chany_top_in[3] mux_left_track_25.mux_l1_in_1_/S
+ mux_left_track_25.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
X_088_ chanx_left_in[6] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_1.mux_l4_in_0__S mux_bottom_track_1.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_6_197 vgnd vpwr scs8hd_fill_1
XFILLER_25_219 vpwr vgnd scs8hd_fill_2
XFILLER_19_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__D mux_right_track_0.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l2_in_7_ _041_/HI chanx_left_in[15] mux_top_track_4.mux_l2_in_0_/S
+ mux_top_track_4.mux_l2_in_7_/X vgnd vpwr scs8hd_mux2_1
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_263 vpwr vgnd scs8hd_fill_2
XFILLER_17_45 vpwr vgnd scs8hd_fill_2
XFILLER_17_89 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_25.mux_l2_in_3__S mux_left_track_25.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_22 vpwr vgnd scs8hd_fill_2
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_156 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_3__A1 chanx_left_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_3_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_32.scs8hd_buf_4_0__A mux_top_track_32.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_7__A1 left_top_grid_pin_49_ vgnd vpwr scs8hd_diode_2
XFILLER_30_255 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_0.mux_l2_in_2_/S mux_top_track_0.mux_l3_in_1_/S
+ mem_top_track_0.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_15_263 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__D mux_top_track_8.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l3_in_0__A1 mux_bottom_track_3.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_3__A0 right_top_grid_pin_47_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l4_in_0__S mux_bottom_track_25.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_266 vpwr vgnd scs8hd_fill_2
XFILLER_21_222 vpwr vgnd scs8hd_fill_2
XANTENNA__071__A _071_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l3_in_0__S mux_left_track_17.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_88 vpwr vgnd scs8hd_fill_2
Xmem_right_track_4.scs8hd_dfxbp_1_3_ prog_clk mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l4_in_0_/S
+ mem_right_track_4.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_5_15 vpwr vgnd scs8hd_fill_2
XFILLER_8_204 vpwr vgnd scs8hd_fill_2
XFILLER_8_259 vpwr vgnd scs8hd_fill_2
XFILLER_12_266 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_32.mux_l1_in_0__S mux_top_track_32.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l4_in_0__S mux_right_track_16.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_ mux_top_track_8.mux_l1_in_1_/X mux_top_track_8.mux_l1_in_0_/X
+ mux_top_track_8.mux_l2_in_1_/S mux_top_track_8.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_0.mux_l2_in_1__S mux_right_track_0.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_270 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l1_in_2__S mux_left_track_3.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA__066__A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_30_23 vpwr vgnd scs8hd_fill_2
XFILLER_14_46 vpwr vgnd scs8hd_fill_2
Xmux_right_track_32.mux_l2_in_0_ mux_right_track_32.mux_l1_in_1_/X mux_right_track_32.mux_l1_in_0_/X
+ mux_right_track_32.mux_l2_in_0_/S mux_right_track_32.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__D mux_left_track_17.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l3_in_2__A0 mux_right_track_4.mux_l2_in_5_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_4__S mux_top_track_2.mux_l1_in_3_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l3_in_1__S mux_top_track_0.mux_l3_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_4_251 vgnd vpwr scs8hd_decap_3
XFILLER_4_262 vpwr vgnd scs8hd_fill_2
XFILLER_35_111 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0__A1 chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A0 top_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XFILLER_26_144 vpwr vgnd scs8hd_fill_2
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_136 vpwr vgnd scs8hd_fill_2
XFILLER_41_114 vpwr vgnd scs8hd_fill_2
XFILLER_41_11 vpwr vgnd scs8hd_fill_2
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_26_188 vpwr vgnd scs8hd_fill_2
XFILLER_25_89 vpwr vgnd scs8hd_fill_2
XFILLER_25_23 vpwr vgnd scs8hd_fill_2
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_32.scs8hd_buf_4_0__A mux_right_track_32.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_210 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_1_ chanx_right_in[11] chanx_right_in[6] mux_top_track_8.mux_l1_in_1_/S
+ mux_top_track_8.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_2_27 vpwr vgnd scs8hd_fill_2
XFILLER_1_254 vpwr vgnd scs8hd_fill_2
XFILLER_32_125 vgnd vpwr scs8hd_fill_1
Xmux_left_track_17.scs8hd_buf_4_0_ mux_left_track_17.mux_l4_in_0_/X _067_/A vgnd vpwr
+ scs8hd_buf_1
Xmux_right_track_32.mux_l1_in_1_ right_top_grid_pin_49_ right_top_grid_pin_45_ mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_3__D mux_right_track_2.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_47 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l4_in_1__A0 mux_right_track_4.mux_l3_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_2__A0 chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_36_88 vpwr vgnd scs8hd_fill_2
XFILLER_14_147 vpwr vgnd scs8hd_fill_2
XFILLER_14_169 vpwr vgnd scs8hd_fill_2
Xmem_left_track_3.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_3.mux_l2_in_2_/S mux_left_track_3.mux_l3_in_1_/S
+ mem_left_track_3.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_20_106 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_8.mux_l4_in_0_/S mux_top_track_16.mux_l1_in_2_/S
+ mem_top_track_16.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_3__D mux_top_track_16.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_81 vpwr vgnd scs8hd_fill_2
XFILLER_36_272 vgnd vpwr scs8hd_decap_3
XFILLER_28_228 vgnd vpwr scs8hd_decap_4
XFILLER_28_206 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_5.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_track_5.mux_l3_in_2_/S mux_bottom_track_5.mux_l4_in_0_/S
+ mem_bottom_track_5.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_22_57 vpwr vgnd scs8hd_fill_2
XFILLER_11_128 vpwr vgnd scs8hd_fill_2
XANTENNA__074__A _074_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_6 vpwr vgnd scs8hd_fill_2
XFILLER_19_217 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_0.mux_l1_in_4__A0 chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_42_264 vgnd vpwr scs8hd_decap_12
X_087_ _087_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_10_150 vgnd vpwr scs8hd_fill_1
XFILLER_10_194 vpwr vgnd scs8hd_fill_2
XFILLER_12_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_32.mux_l1_in_3__S mux_top_track_32.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_1__A0 mux_top_track_2.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_264 vpwr vgnd scs8hd_fill_2
XFILLER_33_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l5_in_0__A0 mux_right_track_4.mux_l4_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_4.mux_l2_in_6_ chanx_left_in[14] chanx_left_in[5] mux_top_track_4.mux_l2_in_0_/S
+ mux_top_track_4.mux_l2_in_6_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__069__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_top_track_8.scs8hd_dfxbp_1_3_ prog_clk mux_top_track_8.mux_l3_in_1_/S mux_top_track_8.mux_l4_in_0_/S
+ mem_top_track_8.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_3__D mux_left_track_25.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_135 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l3_in_2__S mux_right_track_4.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_24.mux_l2_in_0__S mux_top_track_24.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_0.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_0.mux_l1_in_1_/S mux_top_track_0.mux_l2_in_2_/S
+ mem_top_track_0.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_15_231 vpwr vgnd scs8hd_fill_2
XFILLER_15_275 vpwr vgnd scs8hd_fill_2
XFILLER_31_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l4_in_0__S mux_left_track_5.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_3__A1 right_top_grid_pin_46_ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_0_82 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_3__A0 _036_/HI vgnd vpwr scs8hd_diode_2
XFILLER_28_67 vgnd vpwr scs8hd_decap_4
XFILLER_28_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l4_in_0__S mux_right_track_8.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_24.scs8hd_dfxbp_1_3_ prog_clk mux_top_track_24.mux_l3_in_0_/S mux_top_track_24.mux_l4_in_0_/S
+ mem_top_track_24.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
Xmem_right_track_4.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_4.mux_l2_in_0_/S mux_right_track_4.mux_l3_in_0_/S
+ mem_right_track_4.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_2.mux_l3_in_0__A0 mux_top_track_2.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_186 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__D mux_right_track_4.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_3_ _050_/HI left_top_grid_pin_48_ mux_left_track_1.mux_l2_in_0_/S
+ mux_left_track_1.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_14_69 vpwr vgnd scs8hd_fill_2
XANTENNA__082__A chanx_left_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_39_99 vpwr vgnd scs8hd_fill_2
XFILLER_39_66 vpwr vgnd scs8hd_fill_2
Xmux_left_track_25.scs8hd_buf_4_0_ mux_left_track_25.mux_l4_in_0_/X _063_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_29_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l3_in_2__A1 mux_right_track_4.mux_l2_in_4_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_241 vgnd vpwr scs8hd_decap_4
XFILLER_4_274 vgnd vpwr scs8hd_fill_1
XFILLER_35_156 vpwr vgnd scs8hd_fill_2
XFILLER_35_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_3.mux_l1_in_0__A0 chany_top_in[13] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A1 top_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_4__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_33.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_2__A0 bottom_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XANTENNA__077__A chanx_left_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_26_167 vpwr vgnd scs8hd_fill_2
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_4
XFILLER_41_34 vgnd vpwr scs8hd_decap_3
XFILLER_41_23 vgnd vpwr scs8hd_decap_4
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XFILLER_41_89 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_0_ top_left_grid_pin_38_ top_left_grid_pin_34_ mux_top_track_8.mux_l1_in_1_/S
+ mux_top_track_8.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_9_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_33.mux_l2_in_1__S mux_left_track_33.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_1_266 vpwr vgnd scs8hd_fill_2
XFILLER_17_123 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l1_in_4_ left_top_grid_pin_44_ left_top_grid_pin_42_ mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_4_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_104 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_right_track_32.mux_l1_in_0_ chany_top_in[15] chany_top_in[10] mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_115 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_2.mux_l1_in_2__A1 chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l4_in_1__A1 mux_right_track_4.mux_l3_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2__A0 chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_36_67 vgnd vpwr scs8hd_decap_4
XFILLER_36_45 vpwr vgnd scs8hd_fill_2
XFILLER_14_126 vgnd vpwr scs8hd_decap_3
Xmem_left_track_3.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_3.mux_l1_in_0_/S mux_left_track_3.mux_l2_in_2_/S
+ mem_left_track_3.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_left_track_1.mux_l4_in_0_ mux_left_track_1.mux_l3_in_1_/X mux_left_track_1.mux_l3_in_0_/X
+ mux_left_track_1.mux_l4_in_0_/S mux_left_track_1.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_24.mux_l2_in_3__S mux_top_track_24.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l3_in_1__A0 mux_bottom_track_5.mux_l2_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_170 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0__S mux_bottom_track_17.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_bottom_track_5.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_5.mux_l2_in_1_/S mux_bottom_track_5.mux_l3_in_2_/S
+ mem_bottom_track_5.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_22_69 vgnd vpwr scs8hd_decap_4
XANTENNA__090__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_27_240 vpwr vgnd scs8hd_fill_2
XFILLER_19_229 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l1_in_4__A1 chany_bottom_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_42_276 vgnd vpwr scs8hd_fill_1
XFILLER_8_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l3_in_0__S mux_top_track_16.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
X_086_ chanx_left_in[8] chanx_right_out[9] vgnd vpwr scs8hd_buf_2
XFILLER_6_122 vpwr vgnd scs8hd_fill_2
XFILLER_10_173 vpwr vgnd scs8hd_fill_2
XFILLER_26_6 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l2_in_1__A0 mux_left_track_1.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_1__A1 mux_top_track_2.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_251 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l5_in_0__A1 mux_right_track_4.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_276 vgnd vpwr scs8hd_fill_1
Xmux_top_track_4.mux_l2_in_5_ chany_bottom_in[14] chany_bottom_in[5] mux_top_track_4.mux_l2_in_0_/S
+ mux_top_track_4.mux_l2_in_5_/X vgnd vpwr scs8hd_mux2_1
Xmem_top_track_8.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_8.mux_l2_in_1_/S mux_top_track_8.mux_l3_in_1_/S
+ mem_top_track_8.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_17_14 vpwr vgnd scs8hd_fill_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_68 vpwr vgnd scs8hd_fill_2
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_57 vpwr vgnd scs8hd_fill_2
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.mux_l3_in_1_ mux_left_track_1.mux_l2_in_3_/X mux_left_track_1.mux_l2_in_2_/X
+ mux_left_track_1.mux_l3_in_1_/S mux_left_track_1.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__085__A chanx_left_in[9] vgnd vpwr scs8hd_diode_2
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XFILLER_24_210 vpwr vgnd scs8hd_fill_2
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XFILLER_3_103 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_5.mux_l4_in_0__A0 mux_bottom_track_5.mux_l3_in_1_/X vgnd
+ vpwr scs8hd_diode_2
Xmem_top_track_0.scs8hd_dfxbp_1_0_ prog_clk ccff_head mux_top_track_0.mux_l1_in_1_/S
+ mem_top_track_0.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_15_210 vgnd vpwr scs8hd_decap_4
XFILLER_15_243 vgnd vpwr scs8hd_fill_1
XFILLER_30_224 vgnd vpwr scs8hd_decap_3
XFILLER_30_202 vpwr vgnd scs8hd_fill_2
X_069_ chanx_right_in[5] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_21_235 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_left_track_33.scs8hd_buf_4_0_ mux_left_track_33.mux_l3_in_0_/X _059_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_top_track_0.mux_l2_in_3__A1 chanx_left_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_0_117 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_8.mux_l1_in_0__S mux_top_track_8.mux_l1_in_1_/S vgnd vpwr scs8hd_diode_2
Xmem_top_track_24.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_24.mux_l2_in_2_/S mux_top_track_24.mux_l3_in_0_/S
+ mem_top_track_24.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
Xmem_right_track_4.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_4.mux_l1_in_0_/S mux_right_track_4.mux_l2_in_0_/S
+ mem_right_track_4.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_8_228 vpwr vgnd scs8hd_fill_2
XFILLER_12_224 vpwr vgnd scs8hd_fill_2
XFILLER_12_235 vpwr vgnd scs8hd_fill_2
XFILLER_12_246 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l3_in_0__A0 mux_left_track_1.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l3_in_0__A1 mux_top_track_2.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l3_in_1__S mux_bottom_track_3.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_10_9 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_right_track_2.scs8hd_buf_4_0_ mux_right_track_2.mux_l4_in_0_/X _094_/A vgnd vpwr
+ scs8hd_buf_1
Xmux_left_track_1.mux_l2_in_2_ left_top_grid_pin_46_ mux_left_track_1.mux_l1_in_4_/X
+ mux_left_track_1.mux_l2_in_0_/S mux_left_track_1.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__D mux_right_track_24.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_30_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_2__S mux_bottom_track_9.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_23 vpwr vgnd scs8hd_fill_2
XFILLER_29_143 vgnd vpwr scs8hd_decap_3
XFILLER_29_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.mux_l3_in_1__S mux_left_track_25.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_80 vpwr vgnd scs8hd_fill_2
XFILLER_35_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l1_in_0__A1 chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_6_82 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_2__A1 bottom_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_25_36 vpwr vgnd scs8hd_fill_2
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XFILLER_41_68 vpwr vgnd scs8hd_fill_2
XFILLER_41_46 vgnd vpwr scs8hd_decap_12
XANTENNA__093__A _093_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_2__A0 chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_17_179 vpwr vgnd scs8hd_fill_2
XFILLER_15_80 vgnd vpwr scs8hd_decap_3
Xmux_left_track_1.mux_l1_in_3_ chany_bottom_in[19] chany_bottom_in[12] mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_2__S mux_right_track_2.mux_l1_in_4_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l2_in_0__S mux_left_track_3.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_190 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l2_in_3_ _031_/HI chanx_left_in[13] mux_right_track_2.mux_l2_in_0_/S
+ mux_right_track_2.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_17.scs8hd_buf_4_0__A mux_left_track_17.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__D mux_right_track_4.mux_l5_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__088__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l3_in_3_ mux_top_track_4.mux_l2_in_7_/X mux_top_track_4.mux_l2_in_6_/X
+ mux_top_track_4.mux_l3_in_0_/S mux_top_track_4.mux_l3_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_1.mux_l1_in_2__A1 chanx_right_in[12] vgnd vpwr scs8hd_diode_2
Xmem_left_track_3.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_1.mux_l4_in_0_/S mux_left_track_3.mux_l1_in_0_/S
+ mem_left_track_3.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_right_track_32.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_2__S mux_top_track_2.mux_l2_in_2_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1__S mux_left_track_9.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_119 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l3_in_1__A1 mux_bottom_track_5.mux_l2_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_153 vpwr vgnd scs8hd_fill_2
XFILLER_9_175 vpwr vgnd scs8hd_fill_2
XFILLER_13_193 vpwr vgnd scs8hd_fill_2
XFILLER_9_197 vgnd vpwr scs8hd_fill_1
XFILLER_36_230 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_5.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_5.mux_l1_in_0_/S mux_bottom_track_5.mux_l2_in_1_/S
+ mem_bottom_track_5.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_11_108 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l3_in_1__A0 mux_right_track_8.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_200 vgnd vpwr scs8hd_fill_1
XFILLER_42_222 vpwr vgnd scs8hd_fill_2
X_085_ chanx_left_in[9] chanx_right_out[10] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1__A0 chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_6_112 vgnd vpwr scs8hd_decap_4
XFILLER_6_145 vpwr vgnd scs8hd_fill_2
XFILLER_6_167 vgnd vpwr scs8hd_fill_1
XFILLER_12_81 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l1_in_4_ chany_bottom_in[13] chany_bottom_in[11] mux_right_track_2.mux_l1_in_4_/S
+ mux_right_track_2.mux_l1_in_4_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_1.mux_l2_in_1__A1 mux_left_track_1.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_263 vpwr vgnd scs8hd_fill_2
Xmux_top_track_4.mux_l2_in_4_ chanx_right_in[14] chanx_right_in[7] mux_top_track_4.mux_l2_in_0_/S
+ mux_top_track_4.mux_l2_in_4_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_4.mux_l2_in_6__A0 chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_8.mux_l1_in_1_/S mux_top_track_8.mux_l2_in_1_/S
+ mem_top_track_8.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_1_/S mux_left_track_1.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_255 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l4_in_0__A1 mux_bottom_track_5.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_2.mux_l4_in_0_ mux_right_track_2.mux_l3_in_1_/X mux_right_track_2.mux_l3_in_0_/X
+ mux_right_track_2.mux_l4_in_0_/S mux_right_track_2.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
X_068_ chanx_right_in[6] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_2_192 vpwr vgnd scs8hd_fill_2
Xmux_top_track_4.mux_l5_in_0_ mux_top_track_4.mux_l4_in_1_/X mux_top_track_4.mux_l4_in_0_/X
+ mux_top_track_4.mux_l5_in_0_/S mux_top_track_4.mux_l5_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_17_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l4_in_0__A0 mux_right_track_8.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_82 vgnd vpwr scs8hd_decap_4
XANTENNA__096__A chany_top_in[18] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0__A0 mux_bottom_track_17.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
Xmem_top_track_24.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_24.mux_l1_in_1_/S mux_top_track_24.mux_l2_in_2_/S
+ mem_top_track_24.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmem_right_track_4.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_2.mux_l4_in_0_/S mux_right_track_4.mux_l1_in_0_/S
+ mem_right_track_4.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_12_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l3_in_0__A1 mux_left_track_1.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_9.scs8hd_buf_4_0_ mux_bottom_track_9.mux_l4_in_0_/X _111_/A vgnd
+ vpwr scs8hd_buf_1
XANTENNA_mux_top_track_32.mux_l2_in_1__S mux_top_track_32.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_16.scs8hd_buf_4_0_ mux_right_track_16.mux_l4_in_0_/X _087_/A vgnd
+ vpwr scs8hd_buf_1
Xmux_left_track_1.mux_l2_in_1_ mux_left_track_1.mux_l1_in_3_/X mux_left_track_1.mux_l1_in_2_/X
+ mux_left_track_1.mux_l2_in_0_/S mux_left_track_1.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_38_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l2_in_3__S mux_left_track_3.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l4_in_0__S mux_left_track_1.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_3__D mux_right_track_8.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_57 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l3_in_1_ mux_right_track_2.mux_l2_in_3_/X mux_right_track_2.mux_l2_in_2_/X
+ mux_right_track_2.mux_l3_in_0_/S mux_right_track_2.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_29_188 vpwr vgnd scs8hd_fill_2
Xmux_top_track_4.mux_l4_in_1_ mux_top_track_4.mux_l3_in_3_/X mux_top_track_4.mux_l3_in_2_/X
+ mux_top_track_4.mux_l4_in_0_/S mux_top_track_4.mux_l4_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_4.mux_l4_in_0__S mux_right_track_4.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__D mux_bottom_track_33.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_106 vgnd vpwr scs8hd_fill_1
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_26_136 vpwr vgnd scs8hd_fill_2
XFILLER_26_125 vpwr vgnd scs8hd_fill_2
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XFILLER_41_58 vgnd vpwr scs8hd_fill_1
XFILLER_1_235 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l5_in_0__S mux_top_track_4.mux_l5_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_17_114 vgnd vpwr scs8hd_decap_3
XFILLER_40_183 vpwr vgnd scs8hd_fill_2
XFILLER_40_172 vpwr vgnd scs8hd_fill_2
XFILLER_40_150 vgnd vpwr scs8hd_fill_1
XFILLER_32_117 vpwr vgnd scs8hd_fill_2
XFILLER_25_191 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_2__A1 chany_bottom_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_2__A0 top_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_2_ chany_bottom_in[2] chanx_right_in[12] mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_139 vpwr vgnd scs8hd_fill_2
XFILLER_31_161 vpwr vgnd scs8hd_fill_2
XFILLER_11_17 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l2_in_2_ chanx_left_in[4] mux_right_track_2.mux_l1_in_4_/X
+ mux_right_track_2.mux_l2_in_0_/S mux_right_track_2.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2__A0 bottom_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l3_in_2_ mux_top_track_4.mux_l2_in_5_/X mux_top_track_4.mux_l2_in_4_/X
+ mux_top_track_4.mux_l3_in_0_/S mux_top_track_4.mux_l3_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_16.mux_l1_in_2__A0 chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_22_194 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.scs8hd_buf_4_0__A mux_left_track_1.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_1__A0 chanx_right_in[9] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1__S mux_bottom_track_1.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_132 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_5.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_3.mux_l4_in_0_/S mux_bottom_track_5.mux_l1_in_0_/S
+ mem_bottom_track_5.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__D mux_left_track_1.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l3_in_1__A1 mux_right_track_8.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA__099__A _099_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_234 vgnd vpwr scs8hd_decap_12
XFILLER_42_212 vgnd vpwr scs8hd_decap_4
XFILLER_27_220 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_4.mux_l3_in_1__A0 mux_top_track_4.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_142 vpwr vgnd scs8hd_fill_2
X_084_ chanx_left_in[10] chanx_right_out[11] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1__A1 chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_19_7 vgnd vpwr scs8hd_fill_1
Xmux_right_track_2.mux_l1_in_3_ chany_bottom_in[4] right_top_grid_pin_49_ mux_right_track_2.mux_l1_in_4_/S
+ mux_right_track_2.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_9.mux_l2_in_1__A0 bottom_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_1__A0 chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l2_in_3_ chanx_right_in[5] top_left_grid_pin_41_ mux_top_track_4.mux_l2_in_0_/S
+ mux_top_track_4.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_4.mux_l2_in_6__A1 chany_bottom_in[14] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_1__S mux_bottom_track_25.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__A0 mux_bottom_track_25.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_top_track_8.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_4.mux_l5_in_0_/S mux_top_track_8.mux_l1_in_1_/S
+ mem_top_track_8.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_33_26 vpwr vgnd scs8hd_fill_2
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_267 vgnd vpwr scs8hd_decap_8
Xmux_right_track_24.scs8hd_buf_4_0_ mux_right_track_24.mux_l4_in_0_/X _083_/A vgnd
+ vpwr scs8hd_buf_1
XANTENNA_mux_top_track_24.mux_l3_in_1__S mux_top_track_24.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_245 vpwr vgnd scs8hd_fill_2
XFILLER_15_267 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_16.mux_l1_in_1__S mux_right_track_16.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
X_067_ _067_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_8.mux_l4_in_0__A1 mux_right_track_8.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_259 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_4.mux_l4_in_0__A0 mux_top_track_4.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_37 vpwr vgnd scs8hd_fill_2
Xmem_top_track_24.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_16.mux_l4_in_0_/S mux_top_track_24.mux_l1_in_1_/S
+ mem_top_track_24.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_17.mux_l2_in_0__A1 mux_bottom_track_17.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_19 vpwr vgnd scs8hd_fill_2
XFILLER_8_208 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l3_in_0__A0 mux_bottom_track_9.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l3_in_0__A0 mux_right_track_16.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_91 vgnd vpwr scs8hd_fill_1
X_119_ _119_/A chany_top_out[16] vgnd vpwr scs8hd_buf_2
XFILLER_7_274 vgnd vpwr scs8hd_decap_3
XFILLER_38_123 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_0_/S mux_left_track_1.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l1_in_3__A0 chany_bottom_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_30_27 vpwr vgnd scs8hd_fill_2
XFILLER_39_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_5__A0 bottom_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_0_/S mux_right_track_2.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_29_101 vpwr vgnd scs8hd_fill_2
Xmux_top_track_4.mux_l4_in_0_ mux_top_track_4.mux_l3_in_1_/X mux_top_track_4.mux_l3_in_0_/X
+ mux_top_track_4.mux_l4_in_0_/S mux_top_track_4.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_4.mux_l1_in_0__S mux_top_track_4.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_0__A0 chany_top_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_4_211 vgnd vpwr scs8hd_fill_1
XFILLER_4_266 vpwr vgnd scs8hd_fill_2
XFILLER_29_80 vpwr vgnd scs8hd_fill_2
XFILLER_35_115 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_4__S mux_bottom_track_1.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_6_40 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l1_in_2__A0 chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_41_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__D mux_left_track_1.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_26_148 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_33.mux_l1_in_1__A0 bottom_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XFILLER_1_258 vpwr vgnd scs8hd_fill_2
XFILLER_1_214 vpwr vgnd scs8hd_fill_2
XFILLER_17_148 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_2__S mux_bottom_track_5.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_1_ chanx_right_in[2] chany_top_in[12] mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_31_70 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_4.mux_l2_in_2__A1 top_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l2_in_2__A0 left_top_grid_pin_47_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2__A0 chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_31_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.scs8hd_buf_4_0__A mux_right_track_0.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_31_184 vgnd vpwr scs8hd_decap_4
Xmux_right_track_2.mux_l2_in_1_ mux_right_track_2.mux_l1_in_3_/X mux_right_track_2.mux_l1_in_2_/X
+ mux_right_track_2.mux_l2_in_0_/S mux_right_track_2.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2__A1 chanx_right_in[16] vgnd vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l3_in_1_ mux_top_track_4.mux_l2_in_3_/X mux_top_track_4.mux_l2_in_2_/X
+ mux_top_track_4.mux_l3_in_0_/S mux_top_track_4.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_9.mux_l3_in_0__S mux_bottom_track_9.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2__A1 right_top_grid_pin_47_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_1__A1 chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l2_in_1__A0 chany_bottom_in[9] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l2_in_0__A0 mux_bottom_track_33.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_166 vpwr vgnd scs8hd_fill_2
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
XFILLER_36_243 vpwr vgnd scs8hd_fill_2
XFILLER_36_210 vpwr vgnd scs8hd_fill_2
XFILLER_3_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_1__S mux_bottom_track_17.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_32.scs8hd_buf_4_0_ mux_right_track_32.mux_l3_in_0_/X _079_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_42_246 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l3_in_1__A0 mux_left_track_3.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_276 vgnd vpwr scs8hd_fill_1
XFILLER_27_254 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l3_in_1__A1 mux_top_track_4.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_1__A0 chany_bottom_in[17] vgnd vpwr scs8hd_diode_2
X_083_ _083_/A chanx_right_out[12] vgnd vpwr scs8hd_buf_2
Xmux_right_track_2.mux_l1_in_2_ right_top_grid_pin_47_ right_top_grid_pin_45_ mux_right_track_2.mux_l1_in_4_/S
+ mux_right_track_2.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_210 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l2_in_0__S mux_right_track_2.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_268 vpwr vgnd scs8hd_fill_2
XFILLER_33_235 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_1__A1 mux_bottom_track_9.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l2_in_2_ top_left_grid_pin_40_ top_left_grid_pin_39_ mux_top_track_4.mux_l2_in_0_/S
+ mux_top_track_4.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
Xmux_left_track_33.mux_l1_in_3_ _054_/HI left_top_grid_pin_49_ mux_left_track_33.mux_l1_in_3_/S
+ mux_left_track_33.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_16.mux_l2_in_1__A1 mux_right_track_16.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__A1 mux_bottom_track_25.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_224 vpwr vgnd scs8hd_fill_2
XFILLER_33_49 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l3_in_0__A0 mux_right_track_24.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_139 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_1__S mux_right_track_8.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l3_in_0__S mux_top_track_2.mux_l3_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_15_235 vpwr vgnd scs8hd_fill_2
X_135_ _135_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
X_066_ chanx_right_in[8] chanx_left_out[9] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_17.mux_l2_in_3_ _044_/HI chanx_left_in[17] mux_bottom_track_17.mux_l2_in_2_/S
+ mux_bottom_track_17.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_24_6 vgnd vpwr scs8hd_decap_4
XFILLER_0_86 vgnd vpwr scs8hd_decap_4
XFILLER_9_62 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_4.mux_l4_in_0__A1 mux_top_track_4.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l4_in_0__A0 mux_left_track_3.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l3_in_0__A0 mux_top_track_16.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_3__D mux_left_track_3.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_1__S mux_top_track_8.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_20_271 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l3_in_0__A1 mux_bottom_track_9.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__D mux_top_track_16.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_5__S mux_bottom_track_5.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l3_in_0__A1 mux_right_track_16.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_93 vgnd vpwr scs8hd_decap_3
XFILLER_18_60 vpwr vgnd scs8hd_fill_2
XFILLER_7_231 vgnd vpwr scs8hd_fill_1
XFILLER_11_260 vpwr vgnd scs8hd_fill_2
X_118_ chany_bottom_in[16] chany_top_out[17] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_32.mux_l1_in_2__A0 chany_bottom_in[19] vgnd vpwr scs8hd_diode_2
X_049_ _049_/HI _049_/LO vgnd vpwr scs8hd_conb_1
XFILLER_38_102 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_3.mux_l1_in_3__A1 chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_39_15 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_5__A1 bottom_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
XFILLER_29_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_2__D mux_bottom_track_17.mux_l2_in_2_/S
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_33.mux_l3_in_0_ mux_left_track_33.mux_l2_in_1_/X mux_left_track_33.mux_l2_in_0_/X
+ ccff_tail mux_left_track_33.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_5.mux_l2_in_0__A1 mux_left_track_5.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_24.mux_l1_in_2__A0 chany_bottom_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_28_190 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_33.mux_l1_in_1__A1 chanx_right_in[19] vgnd vpwr scs8hd_diode_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_24.mux_l1_in_2__A1 right_top_grid_pin_48_ vgnd vpwr scs8hd_diode_2
XFILLER_41_27 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_33.scs8hd_dfxbp_1_0__D mux_left_track_25.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_193 vpwr vgnd scs8hd_fill_2
XPHY_39 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_3.mux_l2_in_3_ _046_/HI chanx_left_in[13] mux_bottom_track_3.mux_l2_in_3_/S
+ mux_bottom_track_3.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_track_17.mux_l4_in_0_ mux_bottom_track_17.mux_l3_in_1_/X mux_bottom_track_17.mux_l3_in_0_/X
+ mux_bottom_track_17.mux_l4_in_0_/S mux_bottom_track_17.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XANTENNA_mux_right_track_32.mux_l2_in_1__A0 mux_right_track_32.mux_l1_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_163 vgnd vpwr scs8hd_decap_3
XFILLER_40_141 vgnd vpwr scs8hd_decap_3
Xmux_left_track_1.mux_l1_in_0_ chany_top_in[2] chany_top_in[0] mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_0.mux_l1_in_1__A0 right_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
XFILLER_15_94 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l2_in_2__A1 mux_left_track_3.mux_l1_in_4_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_32.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_32.mux_l2_in_1_/S mux_top_track_32.mux_l3_in_0_/S
+ mem_top_track_32.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_2.mux_l2_in_3__S mux_right_track_2.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2__A1 chanx_right_in[17] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l4_in_0__S mux_right_track_0.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_119 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.scs8hd_buf_4_0__A mux_left_track_9.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_0_/S mux_right_track_2.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_3.mux_l3_in_1__S mux_left_track_3.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_0_/S mux_top_track_4.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_left_track_33.mux_l2_in_1_ mux_left_track_33.mux_l1_in_3_/X mux_left_track_33.mux_l1_in_2_/X
+ mux_left_track_33.mux_l2_in_1_/S mux_left_track_33.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_39_263 vgnd vpwr scs8hd_decap_12
XFILLER_36_49 vgnd vpwr scs8hd_decap_3
XFILLER_36_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_24.mux_l2_in_1__A0 chany_bottom_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_22_163 vpwr vgnd scs8hd_fill_2
XFILLER_22_141 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_2__S mux_left_track_9.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_93 vpwr vgnd scs8hd_fill_2
XFILLER_26_82 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l2_in_1__A1 mux_right_track_24.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__D ccff_head vgnd vpwr scs8hd_diode_2
XFILLER_9_101 vpwr vgnd scs8hd_fill_2
XFILLER_13_130 vpwr vgnd scs8hd_fill_2
XFILLER_13_174 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l1_in_2__A0 chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l2_in_0__A1 mux_bottom_track_33.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l1_in_4_ chanx_left_in[3] bottom_left_grid_pin_41_ mux_bottom_track_3.mux_l1_in_4_/S
+ mux_bottom_track_3.mux_l1_in_4_/X vgnd vpwr scs8hd_mux2_1
XFILLER_3_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l3_in_1_ mux_bottom_track_17.mux_l2_in_3_/X mux_bottom_track_17.mux_l2_in_2_/X
+ mux_bottom_track_17.mux_l3_in_0_/S mux_bottom_track_17.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_mux2_1
XANTENNA_mux_right_track_32.mux_l3_in_0__A0 mux_right_track_32.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__D mux_left_track_5.mux_l2_in_7_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0__A0 mux_right_track_0.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_203 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_3.mux_l3_in_1__A1 mux_left_track_3.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_266 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_1__A1 mux_top_track_16.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
X_082_ chanx_left_in[12] chanx_right_out[13] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_10_111 vpwr vgnd scs8hd_fill_2
XFILLER_10_177 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_3__D mux_top_track_24.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_2.mux_l1_in_1_ right_top_grid_pin_43_ chany_top_in[13] mux_right_track_2.mux_l1_in_4_/S
+ mux_right_track_2.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_33_214 vpwr vgnd scs8hd_fill_2
XFILLER_18_255 vpwr vgnd scs8hd_fill_2
XFILLER_18_222 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_3.mux_l4_in_0_ mux_bottom_track_3.mux_l3_in_1_/X mux_bottom_track_3.mux_l3_in_0_/X
+ mux_bottom_track_3.mux_l4_in_0_/S mux_bottom_track_3.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_24.mux_l3_in_0__A0 mux_top_track_24.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_4.mux_l2_in_1_ top_left_grid_pin_38_ top_left_grid_pin_37_ mux_top_track_4.mux_l2_in_0_/S
+ mux_top_track_4.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_left_track_33.mux_l1_in_2_ left_top_grid_pin_45_ chany_bottom_in[15] mux_left_track_33.mux_l1_in_3_/S
+ mux_left_track_33.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_17_18 vpwr vgnd scs8hd_fill_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_24.mux_l3_in_0__A1 mux_right_track_24.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_1__A0 chany_bottom_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_3__A0 _044_/HI vgnd vpwr scs8hd_diode_2
XFILLER_15_214 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_25.scs8hd_buf_4_0__A mux_left_track_25.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_206 vpwr vgnd scs8hd_fill_2
XFILLER_23_50 vpwr vgnd scs8hd_fill_2
X_134_ _134_/A chany_top_out[1] vgnd vpwr scs8hd_buf_2
X_065_ chanx_right_in[9] chanx_left_out[10] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_17.mux_l2_in_2_ chanx_left_in[15] chanx_left_in[8] mux_bottom_track_17.mux_l2_in_2_/S
+ mux_bottom_track_17.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_2_173 vpwr vgnd scs8hd_fill_2
XFILLER_0_10 vpwr vgnd scs8hd_fill_2
XFILLER_0_32 vgnd vpwr scs8hd_decap_3
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XFILLER_21_239 vgnd vpwr scs8hd_decap_3
XFILLER_9_52 vpwr vgnd scs8hd_fill_2
XFILLER_9_74 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l4_in_0__A1 mux_left_track_3.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l1_in_2__S mux_bottom_track_33.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l3_in_0__A1 mux_top_track_16.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_206 vpwr vgnd scs8hd_fill_2
XFILLER_12_228 vpwr vgnd scs8hd_fill_2
XFILLER_12_239 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_32.mux_l1_in_2__A0 chanx_left_in[1] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l3_in_1_ mux_bottom_track_3.mux_l2_in_3_/X mux_bottom_track_3.mux_l2_in_2_/X
+ mux_bottom_track_3.mux_l3_in_1_/S mux_bottom_track_3.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_117_ chany_bottom_in[17] chany_top_out[18] vgnd vpwr scs8hd_buf_2
XFILLER_34_93 vgnd vpwr scs8hd_fill_1
XFILLER_7_210 vgnd vpwr scs8hd_decap_4
XFILLER_7_254 vpwr vgnd scs8hd_fill_2
XFILLER_11_272 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_32.mux_l1_in_2__A1 chany_bottom_in[10] vgnd vpwr scs8hd_diode_2
X_048_ _048_/HI _048_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_track_24.mux_l1_in_2__S mux_right_track_24.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_38_158 vpwr vgnd scs8hd_fill_2
XFILLER_38_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l3_in_0__A0 mux_top_track_8.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_136 vpwr vgnd scs8hd_fill_2
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_20_84 vpwr vgnd scs8hd_fill_2
XFILLER_4_224 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_24.mux_l1_in_2__A1 chanx_right_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_35_128 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_3__D mux_top_track_0.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_5__A0 chany_bottom_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_6_86 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_32.mux_l2_in_1__A0 mux_top_track_32.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_109 vgnd vpwr scs8hd_fill_1
XFILLER_19_180 vgnd vpwr scs8hd_decap_3
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_34_172 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_2__A0 chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l2_in_2_ chanx_left_in[4] mux_bottom_track_3.mux_l1_in_4_/X
+ mux_bottom_track_3.mux_l2_in_3_/S mux_bottom_track_3.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_1_227 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_32.mux_l2_in_1__A1 mux_right_track_32.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_120 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.scs8hd_buf_4_0__A mux_right_track_8.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_62 vgnd vpwr scs8hd_decap_3
XFILLER_31_94 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l1_in_1__A1 chany_top_in[19] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0__A0 chany_top_in[11] vgnd vpwr scs8hd_diode_2
Xmem_top_track_32.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_32.mux_l1_in_0_/S mux_top_track_32.mux_l2_in_1_/S
+ mem_top_track_32.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_0.mux_l1_in_0__S mux_top_track_0.mux_l1_in_1_/S vgnd vpwr scs8hd_diode_2
XANTENNA__102__A chany_top_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_16_150 vgnd vpwr scs8hd_decap_3
XFILLER_31_175 vpwr vgnd scs8hd_fill_2
XFILLER_39_275 vpwr vgnd scs8hd_fill_2
XFILLER_39_220 vpwr vgnd scs8hd_fill_2
Xmux_left_track_33.mux_l2_in_0_ mux_left_track_33.mux_l1_in_1_/X mux_left_track_33.mux_l1_in_0_/X
+ mux_left_track_33.mux_l2_in_1_/S mux_left_track_33.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_36_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_24.mux_l2_in_1__A1 mux_top_track_24.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_109 vpwr vgnd scs8hd_fill_2
XFILLER_22_186 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_32.mux_l3_in_0__A0 mux_top_track_32.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_153 vpwr vgnd scs8hd_fill_2
XFILLER_13_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l2_in_1__A0 chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_2__S mux_bottom_track_1.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2__A1 chanx_right_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_98 vgnd vpwr scs8hd_decap_3
XFILLER_3_21 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.mux_l1_in_3_ bottom_left_grid_pin_39_ bottom_left_grid_pin_37_
+ mux_bottom_track_3.mux_l1_in_4_/S mux_bottom_track_3.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_track_17.mux_l3_in_0_ mux_bottom_track_17.mux_l2_in_1_/X mux_bottom_track_17.mux_l2_in_0_/X
+ mux_bottom_track_17.mux_l3_in_0_/S mux_bottom_track_17.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XANTENNA_mux_right_track_32.mux_l3_in_0__A1 mux_right_track_32.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_3__A0 _045_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0__A1 mux_right_track_0.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_226 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_081_ chanx_left_in[13] chanx_right_out[14] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_5.mux_l3_in_0__S mux_bottom_track_5.mux_l3_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_6_149 vpwr vgnd scs8hd_fill_2
XFILLER_12_85 vgnd vpwr scs8hd_decap_3
XFILLER_12_96 vgnd vpwr scs8hd_decap_4
Xmux_right_track_2.mux_l1_in_0_ chany_top_in[4] chany_top_in[0] mux_right_track_2.mux_l1_in_4_/S
+ mux_right_track_2.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_37_71 vgnd vpwr scs8hd_decap_4
XFILLER_18_267 vgnd vpwr scs8hd_decap_8
XFILLER_18_234 vpwr vgnd scs8hd_fill_2
Xmux_left_track_33.mux_l1_in_1_ chany_bottom_in[10] chanx_right_in[10] mux_left_track_33.mux_l1_in_3_/S
+ mux_left_track_33.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A0 chany_top_in[12] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_24.mux_l3_in_0__A1 mux_top_track_24.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_4.mux_l2_in_0_ top_left_grid_pin_36_ mux_top_track_4.mux_l1_in_0_/X
+ mux_top_track_4.mux_l2_in_0_/S mux_top_track_4.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_5_193 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_25.mux_l2_in_2__S mux_bottom_track_25.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_33_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l3_in_0__A0 mux_left_track_17.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2__S mux_left_track_17.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_3__A1 chanx_left_in[17] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_1__A1 mux_top_track_8.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_259 vpwr vgnd scs8hd_fill_2
X_133_ _133_/A chany_top_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_30_229 vgnd vpwr scs8hd_decap_3
XFILLER_23_270 vpwr vgnd scs8hd_fill_2
XFILLER_23_73 vpwr vgnd scs8hd_fill_2
XFILLER_23_62 vpwr vgnd scs8hd_fill_2
X_064_ chanx_right_in[10] chanx_left_out[11] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__D mux_top_track_2.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_1_ bottom_left_grid_pin_39_ mux_bottom_track_17.mux_l1_in_2_/X
+ mux_bottom_track_17.mux_l2_in_2_/S mux_bottom_track_17.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_mux2_1
XANTENNA__110__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_2__S mux_right_track_16.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_218 vpwr vgnd scs8hd_fill_2
XFILLER_9_31 vpwr vgnd scs8hd_fill_2
XFILLER_14_270 vgnd vpwr scs8hd_decap_4
XFILLER_9_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__D mux_bottom_track_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_251 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_32.mux_l1_in_2__A1 chany_bottom_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1__S mux_left_track_1.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__D mux_left_track_5.mux_l5_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ mux_bottom_track_3.mux_l3_in_1_/S mux_bottom_track_3.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_18_40 vgnd vpwr scs8hd_decap_4
XFILLER_18_84 vpwr vgnd scs8hd_fill_2
XFILLER_18_73 vpwr vgnd scs8hd_fill_2
X_116_ chany_bottom_in[18] chany_top_out[19] vgnd vpwr scs8hd_buf_2
XFILLER_34_83 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_3__A0 left_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
XANTENNA__105__A chany_top_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_7_266 vpwr vgnd scs8hd_fill_2
XFILLER_11_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_3__S mux_top_track_0.mux_l1_in_1_/S vgnd vpwr scs8hd_diode_2
X_047_ _047_/HI _047_/LO vgnd vpwr scs8hd_conb_1
XFILLER_38_148 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_25.mux_l1_in_2__A0 chany_bottom_in[9] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l3_in_0__A1 mux_top_track_8.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_148 vpwr vgnd scs8hd_fill_2
XFILLER_37_170 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_17.mux_l1_in_2_ bottom_left_grid_pin_35_ chanx_right_in[17] mux_bottom_track_17.mux_l1_in_0_/S
+ mux_bottom_track_17.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_203 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_1__S mux_top_track_4.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.scs8hd_buf_4_0_ mux_right_track_8.mux_l4_in_0_/X _091_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_4_247 vpwr vgnd scs8hd_fill_2
XFILLER_4_258 vpwr vgnd scs8hd_fill_2
XFILLER_35_107 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__D mux_left_track_17.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_5__A1 chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_32.scs8hd_dfxbp_1_1__D mux_right_track_32.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_32.mux_l2_in_1__A1 mux_top_track_32.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_19 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.mux_l2_in_1_ mux_bottom_track_3.mux_l1_in_3_/X mux_bottom_track_3.mux_l1_in_2_/X
+ mux_bottom_track_3.mux_l2_in_3_/S mux_bottom_track_3.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_19 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_17.mux_l1_in_2__A1 chanx_right_in[17] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l3_in_2__A0 mux_left_track_5.mux_l2_in_5_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_239 vgnd vpwr scs8hd_decap_3
XFILLER_25_162 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l3_in_3__S mux_bottom_track_5.mux_l3_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_187 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.mux_l2_in_1__A0 chany_bottom_in[11] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0__A1 chany_top_in[6] vgnd vpwr scs8hd_diode_2
Xmem_top_track_32.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_24.mux_l4_in_0_/S mux_top_track_32.mux_l1_in_0_/S
+ mem_top_track_32.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_16_162 vpwr vgnd scs8hd_fill_2
XFILLER_31_165 vgnd vpwr scs8hd_decap_4
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_3.scs8hd_buf_4_0_ mux_left_track_3.mux_l4_in_0_/X _074_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_39_232 vpwr vgnd scs8hd_fill_2
XFILLER_26_51 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_32.mux_l3_in_0__A1 mux_top_track_32.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_83 vgnd vpwr scs8hd_decap_8
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XFILLER_9_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l2_in_1__A1 mux_left_track_17.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__D mux_top_track_4.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA__113__A _113_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l1_in_2_ bottom_left_grid_pin_35_ chanx_right_in[13] mux_bottom_track_3.mux_l1_in_4_/S
+ mux_bottom_track_3.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_32.mux_l1_in_0__S mux_right_track_32.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l4_in_1__A0 mux_left_track_5.mux_l3_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_191 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.mux_l3_in_0__A0 mux_left_track_25.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_3__A1 chanx_left_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_42_216 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__D mux_bottom_track_1.mux_l4_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_4__S mux_left_track_1.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_080_ chanx_left_in[14] chanx_right_out[15] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_3__D mux_left_track_9.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_10_146 vgnd vpwr scs8hd_decap_4
XFILLER_5_3 vgnd vpwr scs8hd_decap_3
XFILLER_12_53 vpwr vgnd scs8hd_fill_2
Xmux_left_track_33.mux_l1_in_0_ chany_top_in[10] chany_top_in[1] mux_left_track_33.mux_l1_in_3_/S
+ mux_left_track_33.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_2.mux_l3_in_1__S mux_right_track_2.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA__108__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A1 chany_top_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.scs8hd_buf_4_0_ mux_bottom_track_17.mux_l4_in_0_/X _107_/A vgnd
+ vpwr scs8hd_buf_1
XANTENNA_mux_left_track_5.mux_l2_in_2__S mux_left_track_5.mux_l2_in_7_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_109 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_4.mux_l1_in_0__A0 chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l3_in_0__A1 mux_left_track_17.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_2__S mux_right_track_8.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_4__S mux_top_track_4.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_15_227 vpwr vgnd scs8hd_fill_2
XFILLER_15_249 vgnd vpwr scs8hd_decap_4
X_132_ chany_bottom_in[2] chany_top_out[3] vgnd vpwr scs8hd_buf_2
X_063_ _063_/A chanx_left_out[12] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_17.mux_l2_in_0_ mux_bottom_track_17.mux_l1_in_1_/X mux_bottom_track_17.mux_l1_in_0_/X
+ mux_bottom_track_17.mux_l2_in_2_/S mux_bottom_track_17.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XANTENNA_mux_left_track_33.mux_l1_in_2__A0 left_top_grid_pin_45_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l5_in_0__A0 mux_left_track_5.mux_l4_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_186 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l3_in_0__S mux_left_track_9.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_23 vgnd vpwr scs8hd_decap_4
XFILLER_20_263 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l1_in_2__A0 right_top_grid_pin_47_ vgnd vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l1_in_0_ top_left_grid_pin_35_ top_left_grid_pin_34_ mux_top_track_4.mux_l1_in_0_/S
+ mux_top_track_4.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_62 vpwr vgnd scs8hd_fill_2
Xmem_left_track_1.scs8hd_dfxbp_1_3_ prog_clk mux_left_track_1.mux_l3_in_1_/S mux_left_track_1.mux_l4_in_0_/S
+ mem_left_track_1.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_5.mux_l2_in_3__A1 chany_bottom_in[14] vgnd vpwr scs8hd_diode_2
X_046_ _046_/HI _046_/LO vgnd vpwr scs8hd_conb_1
XFILLER_7_234 vpwr vgnd scs8hd_fill_2
X_115_ _115_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_11_252 vpwr vgnd scs8hd_fill_2
XANTENNA__121__A chany_bottom_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_22_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.mux_l1_in_2__A1 chanx_right_in[18] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_33.mux_l2_in_1__A0 mux_left_track_33.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_193 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_1_ chanx_right_in[8] chanx_right_in[1] mux_bottom_track_17.mux_l1_in_0_/S
+ mux_bottom_track_17.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_2.scs8hd_buf_4_0__A mux_top_track_2.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_62 vgnd vpwr scs8hd_decap_3
XFILLER_20_53 vpwr vgnd scs8hd_fill_2
XFILLER_35_119 vgnd vpwr scs8hd_decap_3
XFILLER_29_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__S mux_bottom_track_3.mux_l1_in_4_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__116__A chany_bottom_in[18] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_4__A0 chany_bottom_in[15] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_4__D mux_top_track_4.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
X_029_ _029_/HI _029_/LO vgnd vpwr scs8hd_conb_1
XFILLER_3_270 vpwr vgnd scs8hd_fill_2
XFILLER_6_44 vpwr vgnd scs8hd_fill_2
XFILLER_6_55 vpwr vgnd scs8hd_fill_2
XFILLER_26_119 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_32.mux_l1_in_3__S mux_right_track_32.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_3 vpwr vgnd scs8hd_fill_2
XFILLER_34_163 vgnd vpwr scs8hd_decap_3
XFILLER_34_130 vgnd vpwr scs8hd_decap_4
XFILLER_19_160 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_3_/S mux_bottom_track_3.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_41_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l2_in_1__A0 mux_right_track_2.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l2_in_0__S mux_bottom_track_33.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l3_in_2__A1 mux_left_track_5.mux_l2_in_4_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_3__D mux_bottom_track_3.mux_l3_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_119 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_25.mux_l2_in_1__A1 mux_left_track_25.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l1_in_0__S mux_left_track_25.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
XFILLER_31_30 vpwr vgnd scs8hd_fill_2
XFILLER_0_273 vpwr vgnd scs8hd_fill_2
XFILLER_0_262 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_33.mux_l3_in_0__A0 mux_left_track_33.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_188 vgnd vpwr scs8hd_fill_1
XFILLER_31_144 vpwr vgnd scs8hd_fill_2
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_24.mux_l2_in_0__S mux_right_track_24.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_5__S mux_left_track_5.mux_l2_in_7_/S vgnd vpwr
+ scs8hd_diode_2
.ends

