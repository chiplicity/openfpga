VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__0_
  CLASS BLOCK ;
  FOREIGN sb_0__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 120.000 BY 120.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 3.440 120.000 4.040 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 10.240 120.000 10.840 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 17.040 120.000 17.640 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 2.400 3.360 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 2.400 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 2.400 ;
    END
  END address[5]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 24.520 120.000 25.120 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 2.400 8.800 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 31.320 120.000 31.920 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 38.120 120.000 38.720 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 2.400 14.920 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 2.400 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 2.400 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 45.600 120.000 46.200 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 52.400 120.000 53.000 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 2.400 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.070 117.600 6.350 120.000 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 2.400 21.040 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 2.400 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 2.400 27.160 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 2.400 33.280 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 2.400 38.720 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 2.400 44.840 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.030 117.600 18.310 120.000 ;
    END
  END chanx_right_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 59.200 120.000 59.800 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 66.680 120.000 67.280 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 73.480 120.000 74.080 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 2.400 50.960 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 2.400 57.080 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 2.400 63.200 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.990 117.600 30.270 120.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 2.400 68.640 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 2.400 74.760 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.950 117.600 42.230 120.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 53.910 117.600 54.190 120.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.870 117.600 66.150 120.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.830 117.600 78.110 120.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 2.400 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 80.280 120.000 80.880 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 2.400 80.880 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 2.400 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 2.400 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 2.400 ;
    END
  END enable
  PIN right_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 2.400 87.000 ;
    END
  END right_bottom_grid_pin_11_
  PIN right_bottom_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 101.360 120.000 101.960 ;
    END
  END right_bottom_grid_pin_13_
  PIN right_bottom_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 2.400 ;
    END
  END right_bottom_grid_pin_15_
  PIN right_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.790 117.600 90.070 120.000 ;
    END
  END right_bottom_grid_pin_1_
  PIN right_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 2.400 ;
    END
  END right_bottom_grid_pin_3_
  PIN right_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 87.760 120.000 88.360 ;
    END
  END right_bottom_grid_pin_5_
  PIN right_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 2.400 ;
    END
  END right_bottom_grid_pin_7_
  PIN right_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 94.560 120.000 95.160 ;
    END
  END right_bottom_grid_pin_9_
  PIN right_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 2.400 93.120 ;
    END
  END right_top_grid_pin_10_
  PIN top_left_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 2.400 110.800 ;
    END
  END top_left_grid_pin_11_
  PIN top_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 2.400 116.920 ;
    END
  END top_left_grid_pin_13_
  PIN top_left_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 113.710 117.600 113.990 120.000 ;
    END
  END top_left_grid_pin_15_
  PIN top_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 2.400 98.560 ;
    END
  END top_left_grid_pin_1_
  PIN top_left_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 2.400 ;
    END
  END top_left_grid_pin_3_
  PIN top_left_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 2.400 104.680 ;
    END
  END top_left_grid_pin_5_
  PIN top_left_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 101.750 117.600 102.030 120.000 ;
    END
  END top_left_grid_pin_7_
  PIN top_left_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 108.840 120.000 109.440 ;
    END
  END top_left_grid_pin_9_
  PIN top_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 115.640 120.000 116.240 ;
    END
  END top_right_grid_pin_11_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 24.720 10.640 26.320 109.040 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 44.720 10.640 46.320 109.040 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 114.080 108.885 ;
      LAYER met1 ;
        RECT 0.070 10.640 118.150 109.040 ;
      LAYER met2 ;
        RECT 0.090 117.320 5.790 118.050 ;
        RECT 6.630 117.320 17.750 118.050 ;
        RECT 18.590 117.320 29.710 118.050 ;
        RECT 30.550 117.320 41.670 118.050 ;
        RECT 42.510 117.320 53.630 118.050 ;
        RECT 54.470 117.320 65.590 118.050 ;
        RECT 66.430 117.320 77.550 118.050 ;
        RECT 78.390 117.320 89.510 118.050 ;
        RECT 90.350 117.320 101.470 118.050 ;
        RECT 102.310 117.320 113.430 118.050 ;
        RECT 114.270 117.320 118.130 118.050 ;
        RECT 0.090 2.680 118.130 117.320 ;
        RECT 0.090 0.270 3.490 2.680 ;
        RECT 4.330 0.270 11.310 2.680 ;
        RECT 12.150 0.270 19.130 2.680 ;
        RECT 19.970 0.270 27.410 2.680 ;
        RECT 28.250 0.270 35.230 2.680 ;
        RECT 36.070 0.270 43.510 2.680 ;
        RECT 44.350 0.270 51.330 2.680 ;
        RECT 52.170 0.270 59.150 2.680 ;
        RECT 59.990 0.270 67.430 2.680 ;
        RECT 68.270 0.270 75.250 2.680 ;
        RECT 76.090 0.270 83.530 2.680 ;
        RECT 84.370 0.270 91.350 2.680 ;
        RECT 92.190 0.270 99.170 2.680 ;
        RECT 100.010 0.270 107.450 2.680 ;
        RECT 108.290 0.270 115.270 2.680 ;
        RECT 116.110 0.270 118.130 2.680 ;
      LAYER met3 ;
        RECT 2.800 115.920 117.200 116.320 ;
        RECT 0.270 115.240 117.200 115.920 ;
        RECT 0.270 111.200 118.370 115.240 ;
        RECT 2.800 109.840 118.370 111.200 ;
        RECT 2.800 109.800 117.200 109.840 ;
        RECT 0.270 108.440 117.200 109.800 ;
        RECT 0.270 105.080 118.370 108.440 ;
        RECT 2.800 103.680 118.370 105.080 ;
        RECT 0.270 102.360 118.370 103.680 ;
        RECT 0.270 100.960 117.200 102.360 ;
        RECT 0.270 98.960 118.370 100.960 ;
        RECT 2.800 97.560 118.370 98.960 ;
        RECT 0.270 95.560 118.370 97.560 ;
        RECT 0.270 94.160 117.200 95.560 ;
        RECT 0.270 93.520 118.370 94.160 ;
        RECT 2.800 92.120 118.370 93.520 ;
        RECT 0.270 88.760 118.370 92.120 ;
        RECT 0.270 87.400 117.200 88.760 ;
        RECT 2.800 87.360 117.200 87.400 ;
        RECT 2.800 86.000 118.370 87.360 ;
        RECT 0.270 81.280 118.370 86.000 ;
        RECT 2.800 79.880 117.200 81.280 ;
        RECT 0.270 75.160 118.370 79.880 ;
        RECT 2.800 74.480 118.370 75.160 ;
        RECT 2.800 73.760 117.200 74.480 ;
        RECT 0.270 73.080 117.200 73.760 ;
        RECT 0.270 69.040 118.370 73.080 ;
        RECT 2.800 67.680 118.370 69.040 ;
        RECT 2.800 67.640 117.200 67.680 ;
        RECT 0.270 66.280 117.200 67.640 ;
        RECT 0.270 63.600 118.370 66.280 ;
        RECT 2.800 62.200 118.370 63.600 ;
        RECT 0.270 60.200 118.370 62.200 ;
        RECT 0.270 58.800 117.200 60.200 ;
        RECT 0.270 57.480 118.370 58.800 ;
        RECT 2.800 56.080 118.370 57.480 ;
        RECT 0.270 53.400 118.370 56.080 ;
        RECT 0.270 52.000 117.200 53.400 ;
        RECT 0.270 51.360 118.370 52.000 ;
        RECT 2.800 49.960 118.370 51.360 ;
        RECT 0.270 46.600 118.370 49.960 ;
        RECT 0.270 45.240 117.200 46.600 ;
        RECT 2.800 45.200 117.200 45.240 ;
        RECT 2.800 43.840 118.370 45.200 ;
        RECT 0.270 39.120 118.370 43.840 ;
        RECT 2.800 37.720 117.200 39.120 ;
        RECT 0.270 33.680 118.370 37.720 ;
        RECT 2.800 32.320 118.370 33.680 ;
        RECT 2.800 32.280 117.200 32.320 ;
        RECT 0.270 30.920 117.200 32.280 ;
        RECT 0.270 27.560 118.370 30.920 ;
        RECT 2.800 26.160 118.370 27.560 ;
        RECT 0.270 25.520 118.370 26.160 ;
        RECT 0.270 24.120 117.200 25.520 ;
        RECT 0.270 21.440 118.370 24.120 ;
        RECT 2.800 20.040 118.370 21.440 ;
        RECT 0.270 18.040 118.370 20.040 ;
        RECT 0.270 16.640 117.200 18.040 ;
        RECT 0.270 15.320 118.370 16.640 ;
        RECT 2.800 13.920 118.370 15.320 ;
        RECT 0.270 11.240 118.370 13.920 ;
        RECT 0.270 9.840 117.200 11.240 ;
        RECT 0.270 9.200 118.370 9.840 ;
        RECT 2.800 7.800 118.370 9.200 ;
        RECT 0.270 4.440 118.370 7.800 ;
        RECT 0.270 3.760 117.200 4.440 ;
        RECT 2.800 3.360 117.200 3.760 ;
      LAYER met4 ;
        RECT 0.295 10.640 24.320 109.040 ;
        RECT 26.720 10.640 44.320 109.040 ;
        RECT 46.720 10.640 106.320 109.040 ;
  END
END sb_0__0_
END LIBRARY

