VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cby_0__1_
  CLASS BLOCK ;
  FOREIGN cby_0__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 200.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 8.200 80.000 8.800 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 2.400 7.440 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 24.520 80.000 25.120 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 197.600 3.130 200.000 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.370 197.600 8.650 200.000 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 197.600 14.170 200.000 ;
    END
  END address[6]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 41.520 80.000 42.120 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 2.400 21.720 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.870 197.600 20.150 200.000 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 2.400 36.000 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.390 197.600 25.670 200.000 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 57.840 80.000 58.440 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.370 197.600 31.650 200.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 74.840 80.000 75.440 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 36.890 197.600 37.170 200.000 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 2.400 50.280 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 2.400 64.560 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 91.160 80.000 91.760 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 2.400 78.840 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 108.160 80.000 108.760 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 124.480 80.000 125.080 ;
    END
  END chany_bottom_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 141.480 80.000 142.080 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 2.400 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 2.400 93.120 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 2.400 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 157.800 80.000 158.400 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 174.800 80.000 175.400 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 2.400 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.870 197.600 43.150 200.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 2.400 107.400 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 2.400 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 48.390 197.600 48.670 200.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 2.400 121.680 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 2.400 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 53.910 197.600 54.190 200.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.890 197.600 60.170 200.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.410 197.600 65.690 200.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 2.400 135.960 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 2.400 150.240 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 2.400 ;
    END
  END enable
  PIN left_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 2.400 ;
    END
  END left_grid_pin_0_
  PIN left_grid_pin_10_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 2.400 ;
    END
  END left_grid_pin_10_
  PIN left_grid_pin_12_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 2.400 178.800 ;
    END
  END left_grid_pin_12_
  PIN left_grid_pin_14_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 2.400 ;
    END
  END left_grid_pin_14_
  PIN left_grid_pin_2_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 191.120 80.000 191.720 ;
    END
  END left_grid_pin_2_
  PIN left_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 2.400 164.520 ;
    END
  END left_grid_pin_4_
  PIN left_grid_pin_6_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 2.400 ;
    END
  END left_grid_pin_6_
  PIN left_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.390 197.600 71.670 200.000 ;
    END
  END left_grid_pin_8_
  PIN right_grid_pin_3_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.910 197.600 77.190 200.000 ;
    END
  END right_grid_pin_3_
  PIN right_grid_pin_7_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 2.400 193.080 ;
    END
  END right_grid_pin_7_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 18.055 10.640 19.655 187.920 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 31.385 10.640 32.985 187.920 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 74.060 187.765 ;
      LAYER met1 ;
        RECT 0.530 10.640 77.670 198.180 ;
      LAYER met2 ;
        RECT 0.550 197.320 2.570 198.290 ;
        RECT 3.410 197.320 8.090 198.290 ;
        RECT 8.930 197.320 13.610 198.290 ;
        RECT 14.450 197.320 19.590 198.290 ;
        RECT 20.430 197.320 25.110 198.290 ;
        RECT 25.950 197.320 31.090 198.290 ;
        RECT 31.930 197.320 36.610 198.290 ;
        RECT 37.450 197.320 42.590 198.290 ;
        RECT 43.430 197.320 48.110 198.290 ;
        RECT 48.950 197.320 53.630 198.290 ;
        RECT 54.470 197.320 59.610 198.290 ;
        RECT 60.450 197.320 65.130 198.290 ;
        RECT 65.970 197.320 71.110 198.290 ;
        RECT 71.950 197.320 76.630 198.290 ;
        RECT 77.470 197.320 77.650 198.290 ;
        RECT 0.550 2.680 77.650 197.320 ;
        RECT 0.550 0.270 2.110 2.680 ;
        RECT 2.950 0.270 7.170 2.680 ;
        RECT 8.010 0.270 12.690 2.680 ;
        RECT 13.530 0.270 17.750 2.680 ;
        RECT 18.590 0.270 23.270 2.680 ;
        RECT 24.110 0.270 28.790 2.680 ;
        RECT 29.630 0.270 33.850 2.680 ;
        RECT 34.690 0.270 39.370 2.680 ;
        RECT 40.210 0.270 44.430 2.680 ;
        RECT 45.270 0.270 49.950 2.680 ;
        RECT 50.790 0.270 55.470 2.680 ;
        RECT 56.310 0.270 60.530 2.680 ;
        RECT 61.370 0.270 66.050 2.680 ;
        RECT 66.890 0.270 71.110 2.680 ;
        RECT 71.950 0.270 76.630 2.680 ;
        RECT 77.470 0.270 77.650 2.680 ;
      LAYER met3 ;
        RECT 2.800 192.120 77.890 192.480 ;
        RECT 2.800 192.080 77.200 192.120 ;
        RECT 0.310 190.720 77.200 192.080 ;
        RECT 0.310 179.200 77.890 190.720 ;
        RECT 2.800 177.800 77.890 179.200 ;
        RECT 0.310 175.800 77.890 177.800 ;
        RECT 0.310 174.400 77.200 175.800 ;
        RECT 0.310 164.920 77.890 174.400 ;
        RECT 2.800 163.520 77.890 164.920 ;
        RECT 0.310 158.800 77.890 163.520 ;
        RECT 0.310 157.400 77.200 158.800 ;
        RECT 0.310 150.640 77.890 157.400 ;
        RECT 2.800 149.240 77.890 150.640 ;
        RECT 0.310 142.480 77.890 149.240 ;
        RECT 0.310 141.080 77.200 142.480 ;
        RECT 0.310 136.360 77.890 141.080 ;
        RECT 2.800 134.960 77.890 136.360 ;
        RECT 0.310 125.480 77.890 134.960 ;
        RECT 0.310 124.080 77.200 125.480 ;
        RECT 0.310 122.080 77.890 124.080 ;
        RECT 2.800 120.680 77.890 122.080 ;
        RECT 0.310 109.160 77.890 120.680 ;
        RECT 0.310 107.800 77.200 109.160 ;
        RECT 2.800 107.760 77.200 107.800 ;
        RECT 2.800 106.400 77.890 107.760 ;
        RECT 0.310 93.520 77.890 106.400 ;
        RECT 2.800 92.160 77.890 93.520 ;
        RECT 2.800 92.120 77.200 92.160 ;
        RECT 0.310 90.760 77.200 92.120 ;
        RECT 0.310 79.240 77.890 90.760 ;
        RECT 2.800 77.840 77.890 79.240 ;
        RECT 0.310 75.840 77.890 77.840 ;
        RECT 0.310 74.440 77.200 75.840 ;
        RECT 0.310 64.960 77.890 74.440 ;
        RECT 2.800 63.560 77.890 64.960 ;
        RECT 0.310 58.840 77.890 63.560 ;
        RECT 0.310 57.440 77.200 58.840 ;
        RECT 0.310 50.680 77.890 57.440 ;
        RECT 2.800 49.280 77.890 50.680 ;
        RECT 0.310 42.520 77.890 49.280 ;
        RECT 0.310 41.120 77.200 42.520 ;
        RECT 0.310 36.400 77.890 41.120 ;
        RECT 2.800 35.000 77.890 36.400 ;
        RECT 0.310 25.520 77.890 35.000 ;
        RECT 0.310 24.120 77.200 25.520 ;
        RECT 0.310 22.120 77.890 24.120 ;
        RECT 2.800 20.720 77.890 22.120 ;
        RECT 0.310 9.200 77.890 20.720 ;
        RECT 0.310 8.335 77.200 9.200 ;
      LAYER met4 ;
        RECT 15.935 10.640 17.655 187.920 ;
        RECT 20.055 10.640 30.985 187.920 ;
        RECT 33.385 10.640 72.985 187.920 ;
  END
END cby_0__1_
END LIBRARY

