magic
tech EFS8A
magscale 1 2
timestamp 1602529802
<< locali >>
rect 15243 23137 15370 23171
rect 24627 20961 24662 20995
rect 7147 15997 7182 16031
rect 24501 14943 24535 14977
rect 24501 14909 24615 14943
rect 6463 14569 6469 14603
rect 6463 14501 6497 14569
rect 24627 14433 24662 14467
rect 7935 13481 7941 13515
rect 11615 13481 11621 13515
rect 7935 13413 7969 13481
rect 11615 13413 11649 13481
rect 4439 12393 4445 12427
rect 4439 12325 4473 12393
rect 15663 10217 15669 10251
rect 15663 10149 15697 10217
rect 17359 10081 17394 10115
rect 2599 9129 2605 9163
rect 5635 9129 5641 9163
rect 2599 9061 2633 9129
rect 5635 9061 5669 9129
rect 19487 8585 19625 8619
rect 12811 6103 12845 6171
rect 12811 6069 12817 6103
rect 23063 5729 23098 5763
rect 13093 5015 13127 5321
rect 3007 4641 3042 4675
rect 13369 4471 13403 4777
rect 16589 4131 16623 4233
rect 13921 3927 13955 4097
rect 1547 3689 1685 3723
rect 20855 3553 20982 3587
rect 4307 3485 4537 3519
rect 9131 2839 9165 2907
rect 9131 2805 9137 2839
rect 1547 2397 1685 2431
rect 4077 2363 4111 2465
rect 6101 2295 6135 2601
rect 13461 2295 13495 2397
<< viali >>
rect 6009 24293 6043 24327
rect 5917 24157 5951 24191
rect 6561 24157 6595 24191
rect 5273 23817 5307 23851
rect 9137 23817 9171 23851
rect 16221 23817 16255 23851
rect 18521 23817 18555 23851
rect 20637 23817 20671 23851
rect 25145 23817 25179 23851
rect 4951 23749 4985 23783
rect 6193 23749 6227 23783
rect 19993 23749 20027 23783
rect 1444 23613 1478 23647
rect 1869 23613 1903 23647
rect 4880 23613 4914 23647
rect 8652 23613 8686 23647
rect 13620 23613 13654 23647
rect 14013 23613 14047 23647
rect 16037 23613 16071 23647
rect 16589 23613 16623 23647
rect 18337 23613 18371 23647
rect 18889 23613 18923 23647
rect 19508 23613 19542 23647
rect 20453 23613 20487 23647
rect 24660 23613 24694 23647
rect 1547 23545 1581 23579
rect 21005 23545 21039 23579
rect 5917 23477 5951 23511
rect 7021 23477 7055 23511
rect 8723 23477 8757 23511
rect 13691 23477 13725 23511
rect 19579 23477 19613 23511
rect 24731 23477 24765 23511
rect 11069 23273 11103 23307
rect 15439 23273 15473 23307
rect 6469 23205 6503 23239
rect 8033 23205 8067 23239
rect 1444 23137 1478 23171
rect 5340 23137 5374 23171
rect 10885 23137 10919 23171
rect 15209 23137 15243 23171
rect 6377 23069 6411 23103
rect 7021 23069 7055 23103
rect 7941 23069 7975 23103
rect 8217 23069 8251 23103
rect 1547 22933 1581 22967
rect 5411 22933 5445 22967
rect 1593 22729 1627 22763
rect 5365 22729 5399 22763
rect 5917 22729 5951 22763
rect 8585 22729 8619 22763
rect 7297 22593 7331 22627
rect 7941 22593 7975 22627
rect 9229 22593 9263 22627
rect 8804 22525 8838 22559
rect 8907 22525 8941 22559
rect 7113 22457 7147 22491
rect 7389 22457 7423 22491
rect 6285 22389 6319 22423
rect 8217 22389 8251 22423
rect 10977 22389 11011 22423
rect 15301 22389 15335 22423
rect 6101 22185 6135 22219
rect 7205 22185 7239 22219
rect 11483 22185 11517 22219
rect 7389 22117 7423 22151
rect 6009 22049 6043 22083
rect 7481 22049 7515 22083
rect 11412 22049 11446 22083
rect 13804 22049 13838 22083
rect 12541 21845 12575 21879
rect 13875 21845 13909 21879
rect 11805 21641 11839 21675
rect 13829 21641 13863 21675
rect 12541 21505 12575 21539
rect 12817 21505 12851 21539
rect 1444 21437 1478 21471
rect 1869 21437 1903 21471
rect 10701 21437 10735 21471
rect 11437 21437 11471 21471
rect 12173 21437 12207 21471
rect 1547 21369 1581 21403
rect 11529 21369 11563 21403
rect 12633 21369 12667 21403
rect 5825 21301 5859 21335
rect 7389 21301 7423 21335
rect 11437 21029 11471 21063
rect 12909 21029 12943 21063
rect 13001 21029 13035 21063
rect 24593 20961 24627 20995
rect 11345 20893 11379 20927
rect 11805 20893 11839 20927
rect 13185 20893 13219 20927
rect 12725 20757 12759 20791
rect 24731 20757 24765 20791
rect 11253 20553 11287 20587
rect 11805 20553 11839 20587
rect 24685 20553 24719 20587
rect 11345 20417 11379 20451
rect 12725 20417 12759 20451
rect 13001 20417 13035 20451
rect 12817 20281 12851 20315
rect 12173 20213 12207 20247
rect 13645 20213 13679 20247
rect 13369 20009 13403 20043
rect 13093 19941 13127 19975
rect 12449 19873 12483 19907
rect 12633 19125 12667 19159
rect 11529 17833 11563 17867
rect 24777 17833 24811 17867
rect 11345 17697 11379 17731
rect 24593 17697 24627 17731
rect 11437 16949 11471 16983
rect 24593 16949 24627 16983
rect 6412 16609 6446 16643
rect 8217 16609 8251 16643
rect 7573 16541 7607 16575
rect 6515 16405 6549 16439
rect 6377 16201 6411 16235
rect 25145 16201 25179 16235
rect 8769 16133 8803 16167
rect 8217 16065 8251 16099
rect 7113 15997 7147 16031
rect 24660 15997 24694 16031
rect 7251 15929 7285 15963
rect 7665 15929 7699 15963
rect 8033 15929 8067 15963
rect 8309 15929 8343 15963
rect 24731 15861 24765 15895
rect 7573 15589 7607 15623
rect 6101 15521 6135 15555
rect 6561 15453 6595 15487
rect 7481 15453 7515 15487
rect 7941 15453 7975 15487
rect 7205 15317 7239 15351
rect 8493 15317 8527 15351
rect 6101 15113 6135 15147
rect 7481 15113 7515 15147
rect 14197 15113 14231 15147
rect 24777 15113 24811 15147
rect 8309 15045 8343 15079
rect 8677 14977 8711 15011
rect 24501 14977 24535 15011
rect 25145 14977 25179 15011
rect 5708 14909 5742 14943
rect 9137 14909 9171 14943
rect 9321 14909 9355 14943
rect 14013 14909 14047 14943
rect 7757 14841 7791 14875
rect 7858 14841 7892 14875
rect 9229 14841 9263 14875
rect 5779 14773 5813 14807
rect 6469 14773 6503 14807
rect 7021 14773 7055 14807
rect 14657 14773 14691 14807
rect 6469 14569 6503 14603
rect 9781 14569 9815 14603
rect 5089 14501 5123 14535
rect 8033 14501 8067 14535
rect 1409 14433 1443 14467
rect 9689 14433 9723 14467
rect 10149 14433 10183 14467
rect 24593 14433 24627 14467
rect 6101 14365 6135 14399
rect 7941 14365 7975 14399
rect 8309 14365 8343 14399
rect 1593 14297 1627 14331
rect 7021 14297 7055 14331
rect 7757 14297 7791 14331
rect 24731 14229 24765 14263
rect 2421 14025 2455 14059
rect 7113 14025 7147 14059
rect 8493 14025 8527 14059
rect 11437 14025 11471 14059
rect 24685 14025 24719 14059
rect 7573 13889 7607 13923
rect 8769 13889 8803 13923
rect 14749 13889 14783 13923
rect 1409 13821 1443 13855
rect 1961 13821 1995 13855
rect 3065 13821 3099 13855
rect 5089 13821 5123 13855
rect 5365 13821 5399 13855
rect 5733 13821 5767 13855
rect 9356 13821 9390 13855
rect 10517 13821 10551 13855
rect 12484 13821 12518 13855
rect 12909 13821 12943 13855
rect 2973 13753 3007 13787
rect 7389 13753 7423 13787
rect 7894 13753 7928 13787
rect 9781 13753 9815 13787
rect 10838 13753 10872 13787
rect 14841 13753 14875 13787
rect 15393 13753 15427 13787
rect 1593 13685 1627 13719
rect 2789 13685 2823 13719
rect 5273 13685 5307 13719
rect 6193 13685 6227 13719
rect 6561 13685 6595 13719
rect 9137 13685 9171 13719
rect 9459 13685 9493 13719
rect 10333 13685 10367 13719
rect 12587 13685 12621 13719
rect 14473 13685 14507 13719
rect 1547 13481 1581 13515
rect 6469 13481 6503 13515
rect 7481 13481 7515 13515
rect 7941 13481 7975 13515
rect 8493 13481 8527 13515
rect 9781 13481 9815 13515
rect 11621 13481 11655 13515
rect 12173 13481 12207 13515
rect 14749 13481 14783 13515
rect 2605 13413 2639 13447
rect 5911 13413 5945 13447
rect 14381 13413 14415 13447
rect 15485 13413 15519 13447
rect 1476 13345 1510 13379
rect 9689 13345 9723 13379
rect 10149 13345 10183 13379
rect 13737 13345 13771 13379
rect 2513 13277 2547 13311
rect 2881 13277 2915 13311
rect 4077 13277 4111 13311
rect 5549 13277 5583 13311
rect 7573 13277 7607 13311
rect 11253 13277 11287 13311
rect 15393 13277 15427 13311
rect 2237 13209 2271 13243
rect 15945 13209 15979 13243
rect 1961 13141 1995 13175
rect 5273 13141 5307 13175
rect 9321 13141 9355 13175
rect 10701 13141 10735 13175
rect 7849 12937 7883 12971
rect 8309 12937 8343 12971
rect 12587 12937 12621 12971
rect 13645 12937 13679 12971
rect 15025 12937 15059 12971
rect 15301 12937 15335 12971
rect 15761 12937 15795 12971
rect 15991 12937 16025 12971
rect 4261 12869 4295 12903
rect 4721 12869 4755 12903
rect 8953 12869 8987 12903
rect 11805 12869 11839 12903
rect 13921 12869 13955 12903
rect 2513 12801 2547 12835
rect 2789 12801 2823 12835
rect 5733 12801 5767 12835
rect 6653 12801 6687 12835
rect 9597 12801 9631 12835
rect 10517 12801 10551 12835
rect 1685 12733 1719 12767
rect 2421 12733 2455 12767
rect 3341 12733 3375 12767
rect 5365 12733 5399 12767
rect 5641 12733 5675 12767
rect 7113 12733 7147 12767
rect 7297 12733 7331 12767
rect 8769 12733 8803 12767
rect 9229 12733 9263 12767
rect 9781 12733 9815 12767
rect 10241 12733 10275 12767
rect 11161 12733 11195 12767
rect 12484 12733 12518 12767
rect 13277 12733 13311 12767
rect 14105 12733 14139 12767
rect 15920 12733 15954 12767
rect 16313 12733 16347 12767
rect 3249 12665 3283 12699
rect 3662 12665 3696 12699
rect 10793 12665 10827 12699
rect 11345 12665 11379 12699
rect 14426 12665 14460 12699
rect 5089 12597 5123 12631
rect 6193 12597 6227 12631
rect 6929 12597 6963 12631
rect 12265 12597 12299 12631
rect 2329 12393 2363 12427
rect 4445 12393 4479 12427
rect 4997 12393 5031 12427
rect 5549 12393 5583 12427
rect 9045 12393 9079 12427
rect 11069 12393 11103 12427
rect 24777 12393 24811 12427
rect 2605 12325 2639 12359
rect 3525 12325 3559 12359
rect 6561 12325 6595 12359
rect 10701 12325 10735 12359
rect 11345 12325 11379 12359
rect 3157 12257 3191 12291
rect 6009 12257 6043 12291
rect 6377 12257 6411 12291
rect 8125 12257 8159 12291
rect 8309 12257 8343 12291
rect 9965 12257 9999 12291
rect 10425 12257 10459 12291
rect 11621 12257 11655 12291
rect 14172 12257 14206 12291
rect 15393 12257 15427 12291
rect 24593 12257 24627 12291
rect 2513 12189 2547 12223
rect 4077 12189 4111 12223
rect 8401 12189 8435 12223
rect 11529 12189 11563 12223
rect 13093 12189 13127 12223
rect 9413 12121 9447 12155
rect 1685 12053 1719 12087
rect 3893 12053 3927 12087
rect 6929 12053 6963 12087
rect 14243 12053 14277 12087
rect 15577 12053 15611 12087
rect 2881 11849 2915 11883
rect 8677 11849 8711 11883
rect 11621 11849 11655 11883
rect 14197 11849 14231 11883
rect 15393 11849 15427 11883
rect 11253 11781 11287 11815
rect 16497 11781 16531 11815
rect 2513 11713 2547 11747
rect 3065 11713 3099 11747
rect 4905 11713 4939 11747
rect 5917 11713 5951 11747
rect 7757 11713 7791 11747
rect 9137 11713 9171 11747
rect 10517 11713 10551 11747
rect 12449 11713 12483 11747
rect 15577 11713 15611 11747
rect 16037 11713 16071 11747
rect 1685 11645 1719 11679
rect 1961 11645 1995 11679
rect 3709 11645 3743 11679
rect 12265 11645 12299 11679
rect 12541 11645 12575 11679
rect 23740 11645 23774 11679
rect 2145 11577 2179 11611
rect 3157 11577 3191 11611
rect 4629 11577 4663 11611
rect 4721 11577 4755 11611
rect 7389 11577 7423 11611
rect 7481 11577 7515 11611
rect 9229 11577 9263 11611
rect 9781 11577 9815 11611
rect 10701 11577 10735 11611
rect 10793 11577 10827 11611
rect 15669 11577 15703 11611
rect 24593 11577 24627 11611
rect 4169 11509 4203 11543
rect 6285 11509 6319 11543
rect 7205 11509 7239 11543
rect 8309 11509 8343 11543
rect 10149 11509 10183 11543
rect 14473 11509 14507 11543
rect 15025 11509 15059 11543
rect 23811 11509 23845 11543
rect 24225 11509 24259 11543
rect 2329 11305 2363 11339
rect 3893 11305 3927 11339
rect 5365 11305 5399 11339
rect 7389 11305 7423 11339
rect 9137 11305 9171 11339
rect 9965 11305 9999 11339
rect 5089 11237 5123 11271
rect 6101 11237 6135 11271
rect 8217 11237 8251 11271
rect 10425 11237 10459 11271
rect 10977 11237 11011 11271
rect 15393 11237 15427 11271
rect 15485 11237 15519 11271
rect 16037 11237 16071 11271
rect 16957 11237 16991 11271
rect 17049 11237 17083 11271
rect 1476 11169 1510 11203
rect 2697 11169 2731 11203
rect 2881 11169 2915 11203
rect 4537 11169 4571 11203
rect 11897 11169 11931 11203
rect 13645 11169 13679 11203
rect 1961 11101 1995 11135
rect 3157 11101 3191 11135
rect 6009 11101 6043 11135
rect 6285 11101 6319 11135
rect 8125 11101 8159 11135
rect 8769 11101 8803 11135
rect 10333 11101 10367 11135
rect 12541 11101 12575 11135
rect 13369 11101 13403 11135
rect 17233 11101 17267 11135
rect 1547 11033 1581 11067
rect 3433 10965 3467 10999
rect 7849 10965 7883 10999
rect 16497 10965 16531 10999
rect 2697 10761 2731 10795
rect 4537 10761 4571 10795
rect 6009 10761 6043 10795
rect 7849 10761 7883 10795
rect 9229 10761 9263 10795
rect 11253 10761 11287 10795
rect 11897 10761 11931 10795
rect 13645 10761 13679 10795
rect 14381 10761 14415 10795
rect 15393 10761 15427 10795
rect 15669 10761 15703 10795
rect 24777 10761 24811 10795
rect 9597 10693 9631 10727
rect 10977 10693 11011 10727
rect 1685 10625 1719 10659
rect 3341 10625 3375 10659
rect 3617 10625 3651 10659
rect 6285 10625 6319 10659
rect 7113 10625 7147 10659
rect 8309 10625 8343 10659
rect 12725 10625 12759 10659
rect 14473 10625 14507 10659
rect 16497 10625 16531 10659
rect 17141 10625 17175 10659
rect 10057 10557 10091 10591
rect 18153 10557 18187 10591
rect 24593 10557 24627 10591
rect 25145 10557 25179 10591
rect 1777 10489 1811 10523
rect 2329 10489 2363 10523
rect 4721 10489 4755 10523
rect 4813 10489 4847 10523
rect 5365 10489 5399 10523
rect 8217 10489 8251 10523
rect 8671 10489 8705 10523
rect 10378 10489 10412 10523
rect 12817 10489 12851 10523
rect 13369 10489 13403 10523
rect 14794 10489 14828 10523
rect 16589 10489 16623 10523
rect 18061 10489 18095 10523
rect 2973 10421 3007 10455
rect 4169 10421 4203 10455
rect 9873 10421 9907 10455
rect 12265 10421 12299 10455
rect 16313 10421 16347 10455
rect 17417 10421 17451 10455
rect 17785 10421 17819 10455
rect 5273 10217 5307 10251
rect 8401 10217 8435 10251
rect 9965 10217 9999 10251
rect 10701 10217 10735 10251
rect 12725 10217 12759 10251
rect 15025 10217 15059 10251
rect 15669 10217 15703 10251
rect 17463 10217 17497 10251
rect 23719 10217 23753 10251
rect 2605 10149 2639 10183
rect 3433 10149 3467 10183
rect 4439 10149 4473 10183
rect 7205 10149 7239 10183
rect 7757 10149 7791 10183
rect 11253 10149 11287 10183
rect 13185 10149 13219 10183
rect 13737 10149 13771 10183
rect 16957 10149 16991 10183
rect 18429 10149 18463 10183
rect 18521 10149 18555 10183
rect 4997 10081 5031 10115
rect 8585 10081 8619 10115
rect 9873 10081 9907 10115
rect 10149 10081 10183 10115
rect 11621 10081 11655 10115
rect 17325 10081 17359 10115
rect 23648 10081 23682 10115
rect 1409 10013 1443 10047
rect 2513 10013 2547 10047
rect 3157 10013 3191 10047
rect 4077 10013 4111 10047
rect 7113 10013 7147 10047
rect 13093 10013 13127 10047
rect 15301 10013 15335 10047
rect 19073 10013 19107 10047
rect 16221 9945 16255 9979
rect 1869 9877 1903 9911
rect 2329 9877 2363 9911
rect 3801 9877 3835 9911
rect 6929 9877 6963 9911
rect 8769 9877 8803 9911
rect 14565 9877 14599 9911
rect 1547 9673 1581 9707
rect 7757 9673 7791 9707
rect 8125 9673 8159 9707
rect 11621 9673 11655 9707
rect 13369 9673 13403 9707
rect 13645 9673 13679 9707
rect 15393 9673 15427 9707
rect 17877 9673 17911 9707
rect 23857 9673 23891 9707
rect 4629 9605 4663 9639
rect 6653 9605 6687 9639
rect 8493 9605 8527 9639
rect 9413 9605 9447 9639
rect 12173 9605 12207 9639
rect 19165 9605 19199 9639
rect 4077 9537 4111 9571
rect 4997 9537 5031 9571
rect 14749 9537 14783 9571
rect 18613 9537 18647 9571
rect 19533 9537 19567 9571
rect 1476 9469 1510 9503
rect 1869 9469 1903 9503
rect 2329 9469 2363 9503
rect 2789 9469 2823 9503
rect 5800 9469 5834 9503
rect 6837 9469 6871 9503
rect 8577 9469 8611 9503
rect 9689 9469 9723 9503
rect 12449 9469 12483 9503
rect 14197 9469 14231 9503
rect 14657 9469 14691 9503
rect 16037 9469 16071 9503
rect 16221 9469 16255 9503
rect 3157 9401 3191 9435
rect 3433 9401 3467 9435
rect 4169 9401 4203 9435
rect 6285 9401 6319 9435
rect 7199 9401 7233 9435
rect 9137 9401 9171 9435
rect 9597 9401 9631 9435
rect 12770 9401 12804 9435
rect 16773 9401 16807 9435
rect 18705 9401 18739 9435
rect 3801 9333 3835 9367
rect 5365 9333 5399 9367
rect 5871 9333 5905 9367
rect 8769 9333 8803 9367
rect 10701 9333 10735 9367
rect 11161 9333 11195 9367
rect 14013 9333 14047 9367
rect 15853 9333 15887 9367
rect 17325 9333 17359 9367
rect 18429 9333 18463 9367
rect 2605 9129 2639 9163
rect 3157 9129 3191 9163
rect 5089 9129 5123 9163
rect 5641 9129 5675 9163
rect 6469 9129 6503 9163
rect 13553 9129 13587 9163
rect 15117 9129 15151 9163
rect 16497 9129 16531 9163
rect 18889 9129 18923 9163
rect 6837 9061 6871 9095
rect 7113 9061 7147 9095
rect 7205 9061 7239 9095
rect 11069 9061 11103 9095
rect 12541 9061 12575 9095
rect 12633 9061 12667 9095
rect 13185 9061 13219 9095
rect 15622 9061 15656 9095
rect 4077 8993 4111 9027
rect 5273 8993 5307 9027
rect 8585 8993 8619 9027
rect 9873 8993 9907 9027
rect 17141 8993 17175 9027
rect 18705 8993 18739 9027
rect 2237 8925 2271 8959
rect 7389 8925 7423 8959
rect 8125 8925 8159 8959
rect 10977 8925 11011 8959
rect 11621 8925 11655 8959
rect 15301 8925 15335 8959
rect 17049 8925 17083 8959
rect 10333 8857 10367 8891
rect 1593 8789 1627 8823
rect 2053 8789 2087 8823
rect 3525 8789 3559 8823
rect 3801 8789 3835 8823
rect 4261 8789 4295 8823
rect 4537 8789 4571 8823
rect 6193 8789 6227 8823
rect 8401 8789 8435 8823
rect 8769 8789 8803 8823
rect 10057 8789 10091 8823
rect 10701 8789 10735 8823
rect 12265 8789 12299 8823
rect 14197 8789 14231 8823
rect 16221 8789 16255 8823
rect 18337 8789 18371 8823
rect 4261 8585 4295 8619
rect 5089 8585 5123 8619
rect 6193 8585 6227 8619
rect 7113 8585 7147 8619
rect 8585 8585 8619 8619
rect 9781 8585 9815 8619
rect 10793 8585 10827 8619
rect 11069 8585 11103 8619
rect 12265 8585 12299 8619
rect 12633 8585 12667 8619
rect 14657 8585 14691 8619
rect 17141 8585 17175 8619
rect 18613 8585 18647 8619
rect 19625 8585 19659 8619
rect 3801 8517 3835 8551
rect 6653 8517 6687 8551
rect 7757 8517 7791 8551
rect 7941 8517 7975 8551
rect 16681 8517 16715 8551
rect 2697 8449 2731 8483
rect 5273 8449 5307 8483
rect 5917 8449 5951 8483
rect 7849 8449 7883 8483
rect 13185 8449 13219 8483
rect 14105 8449 14139 8483
rect 15761 8449 15795 8483
rect 18061 8449 18095 8483
rect 1685 8381 1719 8415
rect 3157 8381 3191 8415
rect 3525 8381 3559 8415
rect 3709 8381 3743 8415
rect 7628 8381 7662 8415
rect 8953 8381 8987 8415
rect 9873 8381 9907 8415
rect 13645 8381 13679 8415
rect 13921 8381 13955 8415
rect 19416 8381 19450 8415
rect 1501 8313 1535 8347
rect 5365 8313 5399 8347
rect 7481 8313 7515 8347
rect 9413 8313 9447 8347
rect 10194 8313 10228 8347
rect 15025 8313 15059 8347
rect 15853 8313 15887 8347
rect 16405 8313 16439 8347
rect 1777 8245 1811 8279
rect 2421 8245 2455 8279
rect 4629 8245 4663 8279
rect 11437 8245 11471 8279
rect 15301 8245 15335 8279
rect 19901 8245 19935 8279
rect 3341 8041 3375 8075
rect 4353 8041 4387 8075
rect 5549 8041 5583 8075
rect 10793 8041 10827 8075
rect 12173 8041 12207 8075
rect 17141 8041 17175 8075
rect 1863 7973 1897 8007
rect 8309 7973 8343 8007
rect 10425 7973 10459 8007
rect 14289 7973 14323 8007
rect 15622 7973 15656 8007
rect 4169 7905 4203 7939
rect 4629 7905 4663 7939
rect 4905 7905 4939 7939
rect 6193 7905 6227 7939
rect 7573 7905 7607 7939
rect 9965 7905 9999 7939
rect 10149 7905 10183 7939
rect 11069 7905 11103 7939
rect 11989 7905 12023 7939
rect 12357 7905 12391 7939
rect 13461 7905 13495 7939
rect 13645 7905 13679 7939
rect 14013 7905 14047 7939
rect 15301 7905 15335 7939
rect 17141 7905 17175 7939
rect 17509 7905 17543 7939
rect 1501 7837 1535 7871
rect 3709 7837 3743 7871
rect 7941 7837 7975 7871
rect 7738 7769 7772 7803
rect 16221 7769 16255 7803
rect 2421 7701 2455 7735
rect 2973 7701 3007 7735
rect 5917 7701 5951 7735
rect 6285 7701 6319 7735
rect 7113 7701 7147 7735
rect 7481 7701 7515 7735
rect 7849 7701 7883 7735
rect 8585 7701 8619 7735
rect 8953 7701 8987 7735
rect 9413 7701 9447 7735
rect 4445 7497 4479 7531
rect 7665 7497 7699 7531
rect 8677 7497 8711 7531
rect 9762 7497 9796 7531
rect 10241 7497 10275 7531
rect 11989 7497 12023 7531
rect 14289 7497 14323 7531
rect 14933 7497 14967 7531
rect 15485 7497 15519 7531
rect 17049 7497 17083 7531
rect 17509 7497 17543 7531
rect 25145 7497 25179 7531
rect 1869 7429 1903 7463
rect 8309 7429 8343 7463
rect 9873 7429 9907 7463
rect 17785 7429 17819 7463
rect 8401 7361 8435 7395
rect 9965 7361 9999 7395
rect 10609 7361 10643 7395
rect 14013 7361 14047 7395
rect 16405 7361 16439 7395
rect 1685 7293 1719 7327
rect 2513 7293 2547 7327
rect 2973 7293 3007 7327
rect 3525 7293 3559 7327
rect 3709 7293 3743 7327
rect 5089 7293 5123 7327
rect 5825 7293 5859 7327
rect 6837 7293 6871 7327
rect 8180 7293 8214 7327
rect 12633 7293 12667 7327
rect 13093 7293 13127 7327
rect 15092 7293 15126 7327
rect 18153 7293 18187 7327
rect 24660 7293 24694 7327
rect 4169 7225 4203 7259
rect 6561 7225 6595 7259
rect 8033 7225 8067 7259
rect 9597 7225 9631 7259
rect 10977 7225 11011 7259
rect 13369 7225 13403 7259
rect 13461 7225 13495 7259
rect 16129 7225 16163 7259
rect 16221 7225 16255 7259
rect 18061 7225 18095 7259
rect 2145 7157 2179 7191
rect 2789 7157 2823 7191
rect 5457 7157 5491 7191
rect 6193 7157 6227 7191
rect 7021 7157 7055 7191
rect 9137 7157 9171 7191
rect 9413 7157 9447 7191
rect 11345 7157 11379 7191
rect 15163 7157 15197 7191
rect 15945 7157 15979 7191
rect 24731 7157 24765 7191
rect 2789 6953 2823 6987
rect 3157 6953 3191 6987
rect 3801 6953 3835 6987
rect 9781 6953 9815 6987
rect 13185 6953 13219 6987
rect 13461 6953 13495 6987
rect 15117 6953 15151 6987
rect 16313 6953 16347 6987
rect 18521 6953 18555 6987
rect 3525 6885 3559 6919
rect 6469 6885 6503 6919
rect 8769 6885 8803 6919
rect 11069 6885 11103 6919
rect 12627 6885 12661 6919
rect 15485 6885 15519 6919
rect 2053 6817 2087 6851
rect 2973 6817 3007 6851
rect 4077 6817 4111 6851
rect 4629 6817 4663 6851
rect 8033 6817 8067 6851
rect 8180 6817 8214 6851
rect 9689 6817 9723 6851
rect 10149 6817 10183 6851
rect 11253 6817 11287 6851
rect 16865 6817 16899 6851
rect 18429 6817 18463 6851
rect 18889 6817 18923 6851
rect 23765 6817 23799 6851
rect 4445 6749 4479 6783
rect 6377 6749 6411 6783
rect 6837 6749 6871 6783
rect 8401 6749 8435 6783
rect 11713 6749 11747 6783
rect 12265 6749 12299 6783
rect 14197 6749 14231 6783
rect 15393 6749 15427 6783
rect 15669 6749 15703 6783
rect 17233 6749 17267 6783
rect 17601 6749 17635 6783
rect 18153 6749 18187 6783
rect 6009 6681 6043 6715
rect 6745 6681 6779 6715
rect 7113 6681 7147 6715
rect 13829 6681 13863 6715
rect 1685 6613 1719 6647
rect 5273 6613 5307 6647
rect 5549 6613 5583 6647
rect 6634 6613 6668 6647
rect 7665 6613 7699 6647
rect 8309 6613 8343 6647
rect 9045 6613 9079 6647
rect 9413 6613 9447 6647
rect 10701 6613 10735 6647
rect 11437 6613 11471 6647
rect 16773 6613 16807 6647
rect 17003 6613 17037 6647
rect 17141 6613 17175 6647
rect 23949 6613 23983 6647
rect 5346 6409 5380 6443
rect 5825 6409 5859 6443
rect 6561 6409 6595 6443
rect 7573 6409 7607 6443
rect 7849 6409 7883 6443
rect 8309 6409 8343 6443
rect 9137 6409 9171 6443
rect 9873 6409 9907 6443
rect 10701 6409 10735 6443
rect 12265 6409 12299 6443
rect 14565 6409 14599 6443
rect 16681 6409 16715 6443
rect 17233 6409 17267 6443
rect 19073 6409 19107 6443
rect 23949 6409 23983 6443
rect 25145 6409 25179 6443
rect 5457 6341 5491 6375
rect 8171 6341 8205 6375
rect 11345 6341 11379 6375
rect 2237 6273 2271 6307
rect 5549 6273 5583 6307
rect 8401 6273 8435 6307
rect 9413 6273 9447 6307
rect 9965 6273 9999 6307
rect 15025 6273 15059 6307
rect 18521 6273 18555 6307
rect 24225 6273 24259 6307
rect 2973 6205 3007 6239
rect 3249 6205 3283 6239
rect 3709 6205 3743 6239
rect 3893 6205 3927 6239
rect 6837 6205 6871 6239
rect 9597 6205 9631 6239
rect 9744 6205 9778 6239
rect 11161 6205 11195 6239
rect 11621 6205 11655 6239
rect 12449 6205 12483 6239
rect 13645 6205 13679 6239
rect 16824 6205 16858 6239
rect 18061 6205 18095 6239
rect 18613 6205 18647 6239
rect 19441 6205 19475 6239
rect 1593 6137 1627 6171
rect 1685 6137 1719 6171
rect 5089 6137 5123 6171
rect 5181 6137 5215 6171
rect 8033 6137 8067 6171
rect 8769 6137 8803 6171
rect 10977 6137 11011 6171
rect 14841 6137 14875 6171
rect 15346 6137 15380 6171
rect 16911 6137 16945 6171
rect 24317 6137 24351 6171
rect 24869 6137 24903 6171
rect 2605 6069 2639 6103
rect 4169 6069 4203 6103
rect 4537 6069 4571 6103
rect 7021 6069 7055 6103
rect 10241 6069 10275 6103
rect 12817 6069 12851 6103
rect 13369 6069 13403 6103
rect 14013 6069 14047 6103
rect 15945 6069 15979 6103
rect 16221 6069 16255 6103
rect 17785 6069 17819 6103
rect 23397 6069 23431 6103
rect 1869 5865 1903 5899
rect 2237 5865 2271 5899
rect 3893 5865 3927 5899
rect 5825 5865 5859 5899
rect 7297 5865 7331 5899
rect 11161 5865 11195 5899
rect 12541 5865 12575 5899
rect 15117 5865 15151 5899
rect 15945 5865 15979 5899
rect 2605 5797 2639 5831
rect 4398 5797 4432 5831
rect 9505 5797 9539 5831
rect 12173 5797 12207 5831
rect 12817 5797 12851 5831
rect 16681 5797 16715 5831
rect 18245 5797 18279 5831
rect 24225 5797 24259 5831
rect 1409 5729 1443 5763
rect 4997 5729 5031 5763
rect 6377 5729 6411 5763
rect 6745 5729 6779 5763
rect 7849 5729 7883 5763
rect 7996 5729 8030 5763
rect 9689 5729 9723 5763
rect 9836 5729 9870 5763
rect 11713 5729 11747 5763
rect 11897 5729 11931 5763
rect 13921 5729 13955 5763
rect 14105 5729 14139 5763
rect 14749 5729 14783 5763
rect 15393 5729 15427 5763
rect 17509 5729 17543 5763
rect 23029 5729 23063 5763
rect 2513 5661 2547 5695
rect 3157 5661 3191 5695
rect 4077 5661 4111 5695
rect 6837 5661 6871 5695
rect 8217 5661 8251 5695
rect 8953 5661 8987 5695
rect 10057 5661 10091 5695
rect 14381 5661 14415 5695
rect 16589 5661 16623 5695
rect 18153 5661 18187 5695
rect 18429 5661 18463 5695
rect 24133 5661 24167 5695
rect 1593 5593 1627 5627
rect 6101 5593 6135 5627
rect 10885 5593 10919 5627
rect 15577 5593 15611 5627
rect 17141 5593 17175 5627
rect 24685 5593 24719 5627
rect 3433 5525 3467 5559
rect 5365 5525 5399 5559
rect 7757 5525 7791 5559
rect 8125 5525 8159 5559
rect 8493 5525 8527 5559
rect 9965 5525 9999 5559
rect 10149 5525 10183 5559
rect 13553 5525 13587 5559
rect 23167 5525 23201 5559
rect 1685 5321 1719 5355
rect 9229 5321 9263 5355
rect 9689 5321 9723 5355
rect 12633 5321 12667 5355
rect 13093 5321 13127 5355
rect 16957 5321 16991 5355
rect 17509 5321 17543 5355
rect 23121 5321 23155 5355
rect 24685 5321 24719 5355
rect 25053 5321 25087 5355
rect 25375 5321 25409 5355
rect 4997 5253 5031 5287
rect 5917 5253 5951 5287
rect 6285 5253 6319 5287
rect 7987 5253 8021 5287
rect 8125 5253 8159 5287
rect 11897 5253 11931 5287
rect 12955 5253 12989 5287
rect 3065 5185 3099 5219
rect 8217 5185 8251 5219
rect 2421 5117 2455 5151
rect 4537 5117 4571 5151
rect 5733 5117 5767 5151
rect 6837 5117 6871 5151
rect 7849 5117 7883 5151
rect 9413 5117 9447 5151
rect 9597 5117 9631 5151
rect 10241 5117 10275 5151
rect 10885 5117 10919 5151
rect 11253 5117 11287 5151
rect 12173 5117 12207 5151
rect 12852 5117 12886 5151
rect 4629 5049 4663 5083
rect 5641 5049 5675 5083
rect 7297 5049 7331 5083
rect 7665 5049 7699 5083
rect 8585 5049 8619 5083
rect 11529 5049 11563 5083
rect 16313 5253 16347 5287
rect 23397 5185 23431 5219
rect 13277 5117 13311 5151
rect 13829 5117 13863 5151
rect 14289 5117 14323 5151
rect 14565 5117 14599 5151
rect 15209 5117 15243 5151
rect 15393 5117 15427 5151
rect 18061 5117 18095 5151
rect 18705 5117 18739 5151
rect 23765 5117 23799 5151
rect 25304 5117 25338 5151
rect 13645 5049 13679 5083
rect 14841 5049 14875 5083
rect 15714 5049 15748 5083
rect 19625 5049 19659 5083
rect 2145 4981 2179 5015
rect 3709 4981 3743 5015
rect 6561 4981 6595 5015
rect 7021 4981 7055 5015
rect 8953 4981 8987 5015
rect 10701 4981 10735 5015
rect 13093 4981 13127 5015
rect 16681 4981 16715 5015
rect 17785 4981 17819 5015
rect 22293 4981 22327 5015
rect 23949 4981 23983 5015
rect 25789 4981 25823 5015
rect 2513 4777 2547 4811
rect 2881 4777 2915 4811
rect 5733 4777 5767 4811
rect 7389 4777 7423 4811
rect 8493 4777 8527 4811
rect 9965 4777 9999 4811
rect 13093 4777 13127 4811
rect 13369 4777 13403 4811
rect 15117 4777 15151 4811
rect 16957 4777 16991 4811
rect 1409 4709 1443 4743
rect 3111 4709 3145 4743
rect 4537 4709 4571 4743
rect 7665 4709 7699 4743
rect 9229 4709 9263 4743
rect 10879 4709 10913 4743
rect 11805 4709 11839 4743
rect 1777 4641 1811 4675
rect 2973 4641 3007 4675
rect 6193 4641 6227 4675
rect 6469 4641 6503 4675
rect 8217 4641 8251 4675
rect 11437 4641 11471 4675
rect 12684 4641 12718 4675
rect 4445 4573 4479 4607
rect 4721 4573 4755 4607
rect 6653 4573 6687 4607
rect 7573 4573 7607 4607
rect 10517 4573 10551 4607
rect 12081 4573 12115 4607
rect 12771 4573 12805 4607
rect 8861 4505 8895 4539
rect 10241 4505 10275 4539
rect 12449 4505 12483 4539
rect 15714 4709 15748 4743
rect 17141 4709 17175 4743
rect 22569 4709 22603 4743
rect 24133 4709 24167 4743
rect 13829 4641 13863 4675
rect 14105 4641 14139 4675
rect 14657 4641 14691 4675
rect 17233 4641 17267 4675
rect 18797 4641 18831 4675
rect 14197 4573 14231 4607
rect 15393 4573 15427 4607
rect 18705 4573 18739 4607
rect 22477 4573 22511 4607
rect 22753 4573 22787 4607
rect 24041 4573 24075 4607
rect 24317 4573 24351 4607
rect 3709 4437 3743 4471
rect 5457 4437 5491 4471
rect 6929 4437 6963 4471
rect 13369 4437 13403 4471
rect 13461 4437 13495 4471
rect 16313 4437 16347 4471
rect 18245 4437 18279 4471
rect 1869 4233 1903 4267
rect 2973 4233 3007 4267
rect 3525 4233 3559 4267
rect 3755 4233 3789 4267
rect 3893 4233 3927 4267
rect 4261 4233 4295 4267
rect 4629 4233 4663 4267
rect 16589 4233 16623 4267
rect 16865 4233 16899 4267
rect 21557 4233 21591 4267
rect 23949 4233 23983 4267
rect 6193 4165 6227 4199
rect 7389 4165 7423 4199
rect 8677 4165 8711 4199
rect 9735 4165 9769 4199
rect 19073 4165 19107 4199
rect 23489 4165 23523 4199
rect 3985 4097 4019 4131
rect 12541 4097 12575 4131
rect 13921 4097 13955 4131
rect 14013 4097 14047 4131
rect 14841 4097 14875 4131
rect 15393 4097 15427 4131
rect 16497 4097 16531 4131
rect 16589 4097 16623 4131
rect 22109 4097 22143 4131
rect 22753 4097 22787 4131
rect 24501 4097 24535 4131
rect 1777 4029 1811 4063
rect 2513 4029 2547 4063
rect 3617 4029 3651 4063
rect 5089 4029 5123 4063
rect 5273 4029 5307 4063
rect 5641 4029 5675 4063
rect 7481 4029 7515 4063
rect 9505 4029 9539 4063
rect 9664 4029 9698 4063
rect 10425 4029 10459 4063
rect 10609 4029 10643 4063
rect 11529 4029 11563 4063
rect 1685 3961 1719 3995
rect 5917 3961 5951 3995
rect 7822 3961 7856 3995
rect 10149 3961 10183 3995
rect 10930 3961 10964 3995
rect 12265 3961 12299 3995
rect 12633 3961 12667 3995
rect 13185 3961 13219 3995
rect 14197 4029 14231 4063
rect 14749 4029 14783 4063
rect 17141 4029 17175 4063
rect 17877 4029 17911 4063
rect 18153 4029 18187 4063
rect 20704 4029 20738 4063
rect 21097 4029 21131 4063
rect 15853 3961 15887 3995
rect 15945 3961 15979 3995
rect 18061 3961 18095 3995
rect 21925 3961 21959 3995
rect 22201 3961 22235 3995
rect 24225 3961 24259 3995
rect 24317 3961 24351 3995
rect 6561 3893 6595 3927
rect 8401 3893 8435 3927
rect 9045 3893 9079 3927
rect 11805 3893 11839 3927
rect 13737 3893 13771 3927
rect 13921 3893 13955 3927
rect 19625 3893 19659 3927
rect 20775 3893 20809 3927
rect 23029 3893 23063 3927
rect 1685 3689 1719 3723
rect 3617 3689 3651 3723
rect 6285 3689 6319 3723
rect 7941 3689 7975 3723
rect 9321 3689 9355 3723
rect 10885 3689 10919 3723
rect 14473 3689 14507 3723
rect 14841 3689 14875 3723
rect 16589 3689 16623 3723
rect 22109 3689 22143 3723
rect 24225 3689 24259 3723
rect 24915 3689 24949 3723
rect 2421 3621 2455 3655
rect 3157 3621 3191 3655
rect 5365 3621 5399 3655
rect 6561 3621 6595 3655
rect 7066 3621 7100 3655
rect 10609 3621 10643 3655
rect 11253 3621 11287 3655
rect 12034 3621 12068 3655
rect 13645 3621 13679 3655
rect 15622 3621 15656 3655
rect 17233 3621 17267 3655
rect 18429 3621 18463 3655
rect 18797 3621 18831 3655
rect 22201 3621 22235 3655
rect 1476 3553 1510 3587
rect 4236 3553 4270 3587
rect 7665 3553 7699 3587
rect 8309 3553 8343 3587
rect 9873 3553 9907 3587
rect 10333 3553 10367 3587
rect 13277 3553 13311 3587
rect 16221 3553 16255 3587
rect 20821 3553 20855 3587
rect 22569 3553 22603 3587
rect 23800 3553 23834 3587
rect 24593 3553 24627 3587
rect 24844 3553 24878 3587
rect 2789 3485 2823 3519
rect 4537 3485 4571 3519
rect 5273 3485 5307 3519
rect 5917 3485 5951 3519
rect 6745 3485 6779 3519
rect 8493 3485 8527 3519
rect 11713 3485 11747 3519
rect 13553 3485 13587 3519
rect 13829 3485 13863 3519
rect 15301 3485 15335 3519
rect 17141 3485 17175 3519
rect 17785 3485 17819 3519
rect 18705 3485 18739 3519
rect 18981 3485 19015 3519
rect 2697 3417 2731 3451
rect 8953 3417 8987 3451
rect 12909 3417 12943 3451
rect 1869 3349 1903 3383
rect 2237 3349 2271 3383
rect 2586 3349 2620 3383
rect 4629 3349 4663 3383
rect 4997 3349 5031 3383
rect 12633 3349 12667 3383
rect 16865 3349 16899 3383
rect 21051 3349 21085 3383
rect 23903 3349 23937 3383
rect 1961 3145 1995 3179
rect 3065 3145 3099 3179
rect 3433 3145 3467 3179
rect 5089 3145 5123 3179
rect 5457 3145 5491 3179
rect 5825 3145 5859 3179
rect 6285 3145 6319 3179
rect 7113 3145 7147 3179
rect 9689 3145 9723 3179
rect 9965 3145 9999 3179
rect 10333 3145 10367 3179
rect 11713 3145 11747 3179
rect 13553 3145 13587 3179
rect 14105 3145 14139 3179
rect 17325 3145 17359 3179
rect 17877 3145 17911 3179
rect 19073 3145 19107 3179
rect 23029 3145 23063 3179
rect 23489 3145 23523 3179
rect 24869 3145 24903 3179
rect 5346 3077 5380 3111
rect 14381 3077 14415 3111
rect 19901 3077 19935 3111
rect 5549 3009 5583 3043
rect 7297 3009 7331 3043
rect 8309 3009 8343 3043
rect 8769 3009 8803 3043
rect 10885 3009 10919 3043
rect 13185 3009 13219 3043
rect 14565 3009 14599 3043
rect 16681 3009 16715 3043
rect 18153 3009 18187 3043
rect 18429 3009 18463 3043
rect 21649 3009 21683 3043
rect 22661 3009 22695 3043
rect 2697 2941 2731 2975
rect 4169 2941 4203 2975
rect 5181 2941 5215 2975
rect 6561 2941 6595 2975
rect 19717 2941 19751 2975
rect 21224 2941 21258 2975
rect 22268 2941 22302 2975
rect 24133 2941 24167 2975
rect 24276 2941 24310 2975
rect 2789 2873 2823 2907
rect 4353 2873 4387 2907
rect 7389 2873 7423 2907
rect 7941 2873 7975 2907
rect 10609 2873 10643 2907
rect 10701 2873 10735 2907
rect 12541 2873 12575 2907
rect 12633 2873 12667 2907
rect 14886 2873 14920 2907
rect 15761 2873 15795 2907
rect 16405 2873 16439 2907
rect 16497 2873 16531 2907
rect 18245 2873 18279 2907
rect 24363 2873 24397 2907
rect 4721 2805 4755 2839
rect 8677 2805 8711 2839
rect 9137 2805 9171 2839
rect 12265 2805 12299 2839
rect 15485 2805 15519 2839
rect 16221 2805 16255 2839
rect 19441 2805 19475 2839
rect 20913 2805 20947 2839
rect 21327 2805 21361 2839
rect 22339 2805 22373 2839
rect 1869 2601 1903 2635
rect 4399 2601 4433 2635
rect 5089 2601 5123 2635
rect 5917 2601 5951 2635
rect 6101 2601 6135 2635
rect 6377 2601 6411 2635
rect 7251 2601 7285 2635
rect 9137 2601 9171 2635
rect 10793 2601 10827 2635
rect 11161 2601 11195 2635
rect 11621 2601 11655 2635
rect 11989 2601 12023 2635
rect 14841 2601 14875 2635
rect 18153 2601 18187 2635
rect 20545 2601 20579 2635
rect 23397 2601 23431 2635
rect 2237 2533 2271 2567
rect 5273 2533 5307 2567
rect 1476 2465 1510 2499
rect 3065 2465 3099 2499
rect 3157 2465 3191 2499
rect 4077 2465 4111 2499
rect 4328 2465 4362 2499
rect 4813 2465 4847 2499
rect 1685 2397 1719 2431
rect 5641 2397 5675 2431
rect 3433 2329 3467 2363
rect 4077 2329 4111 2363
rect 7941 2533 7975 2567
rect 8217 2533 8251 2567
rect 8309 2533 8343 2567
rect 9505 2533 9539 2567
rect 9965 2533 9999 2567
rect 10517 2533 10551 2567
rect 12817 2533 12851 2567
rect 13369 2533 13403 2567
rect 15301 2533 15335 2567
rect 15669 2533 15703 2567
rect 16221 2533 16255 2567
rect 16957 2533 16991 2567
rect 18337 2533 18371 2567
rect 7180 2465 7214 2499
rect 8861 2465 8895 2499
rect 11437 2465 11471 2499
rect 14197 2465 14231 2499
rect 17049 2465 17083 2499
rect 17785 2465 17819 2499
rect 18429 2465 18463 2499
rect 19901 2465 19935 2499
rect 21224 2465 21258 2499
rect 21649 2465 21683 2499
rect 22753 2465 22787 2499
rect 6653 2397 6687 2431
rect 9873 2397 9907 2431
rect 12725 2397 12759 2431
rect 13461 2397 13495 2431
rect 15566 2397 15600 2431
rect 16497 2397 16531 2431
rect 19717 2397 19751 2431
rect 14013 2329 14047 2363
rect 14381 2329 14415 2363
rect 17233 2329 17267 2363
rect 20085 2329 20119 2363
rect 22937 2329 22971 2363
rect 3893 2261 3927 2295
rect 5411 2261 5445 2295
rect 5549 2261 5583 2295
rect 6101 2261 6135 2295
rect 7665 2261 7699 2295
rect 12449 2261 12483 2295
rect 13461 2261 13495 2295
rect 13737 2261 13771 2295
rect 19349 2261 19383 2295
rect 21327 2261 21361 2295
<< metal1 >>
rect 14 27480 20 27532
rect 72 27520 78 27532
rect 1026 27520 1032 27532
rect 72 27492 1032 27520
rect 72 27480 78 27492
rect 1026 27480 1032 27492
rect 1084 27480 1090 27532
rect 3142 27480 3148 27532
rect 3200 27520 3206 27532
rect 3970 27520 3976 27532
rect 3200 27492 3976 27520
rect 3200 27480 3206 27492
rect 3970 27480 3976 27492
rect 4028 27480 4034 27532
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 5997 24327 6055 24333
rect 5997 24293 6009 24327
rect 6043 24324 6055 24327
rect 6086 24324 6092 24336
rect 6043 24296 6092 24324
rect 6043 24293 6055 24296
rect 5997 24287 6055 24293
rect 6086 24284 6092 24296
rect 6144 24284 6150 24336
rect 5905 24191 5963 24197
rect 5905 24157 5917 24191
rect 5951 24188 5963 24191
rect 5994 24188 6000 24200
rect 5951 24160 6000 24188
rect 5951 24157 5963 24160
rect 5905 24151 5963 24157
rect 5994 24148 6000 24160
rect 6052 24148 6058 24200
rect 6549 24191 6607 24197
rect 6549 24157 6561 24191
rect 6595 24188 6607 24191
rect 6638 24188 6644 24200
rect 6595 24160 6644 24188
rect 6595 24157 6607 24160
rect 6549 24151 6607 24157
rect 6638 24148 6644 24160
rect 6696 24148 6702 24200
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 5258 23848 5264 23860
rect 5219 23820 5264 23848
rect 5258 23808 5264 23820
rect 5316 23808 5322 23860
rect 9125 23851 9183 23857
rect 9125 23817 9137 23851
rect 9171 23848 9183 23851
rect 9582 23848 9588 23860
rect 9171 23820 9588 23848
rect 9171 23817 9183 23820
rect 9125 23811 9183 23817
rect 4939 23783 4997 23789
rect 4939 23749 4951 23783
rect 4985 23780 4997 23783
rect 5994 23780 6000 23792
rect 4985 23752 6000 23780
rect 4985 23749 4997 23752
rect 4939 23743 4997 23749
rect 5994 23740 6000 23752
rect 6052 23780 6058 23792
rect 6181 23783 6239 23789
rect 6181 23780 6193 23783
rect 6052 23752 6193 23780
rect 6052 23740 6058 23752
rect 6181 23749 6193 23752
rect 6227 23749 6239 23783
rect 6181 23743 6239 23749
rect 1026 23604 1032 23656
rect 1084 23644 1090 23656
rect 1432 23647 1490 23653
rect 1432 23644 1444 23647
rect 1084 23616 1444 23644
rect 1084 23604 1090 23616
rect 1432 23613 1444 23616
rect 1478 23644 1490 23647
rect 1857 23647 1915 23653
rect 1857 23644 1869 23647
rect 1478 23616 1869 23644
rect 1478 23613 1490 23616
rect 1432 23607 1490 23613
rect 1857 23613 1869 23616
rect 1903 23613 1915 23647
rect 1857 23607 1915 23613
rect 4868 23647 4926 23653
rect 4868 23613 4880 23647
rect 4914 23644 4926 23647
rect 5258 23644 5264 23656
rect 4914 23616 5264 23644
rect 4914 23613 4926 23616
rect 4868 23607 4926 23613
rect 5258 23604 5264 23616
rect 5316 23604 5322 23656
rect 8640 23647 8698 23653
rect 8640 23613 8652 23647
rect 8686 23644 8698 23647
rect 9140 23644 9168 23811
rect 9582 23808 9588 23820
rect 9640 23808 9646 23860
rect 16209 23851 16267 23857
rect 16209 23817 16221 23851
rect 16255 23848 16267 23851
rect 18230 23848 18236 23860
rect 16255 23820 18236 23848
rect 16255 23817 16267 23820
rect 16209 23811 16267 23817
rect 18230 23808 18236 23820
rect 18288 23808 18294 23860
rect 18509 23851 18567 23857
rect 18509 23817 18521 23851
rect 18555 23848 18567 23851
rect 20346 23848 20352 23860
rect 18555 23820 20352 23848
rect 18555 23817 18567 23820
rect 18509 23811 18567 23817
rect 20346 23808 20352 23820
rect 20404 23808 20410 23860
rect 20625 23851 20683 23857
rect 20625 23817 20637 23851
rect 20671 23848 20683 23851
rect 22462 23848 22468 23860
rect 20671 23820 22468 23848
rect 20671 23817 20683 23820
rect 20625 23811 20683 23817
rect 22462 23808 22468 23820
rect 22520 23808 22526 23860
rect 25130 23848 25136 23860
rect 25091 23820 25136 23848
rect 25130 23808 25136 23820
rect 25188 23808 25194 23860
rect 19981 23783 20039 23789
rect 19981 23749 19993 23783
rect 20027 23780 20039 23783
rect 24670 23780 24676 23792
rect 20027 23752 24676 23780
rect 20027 23749 20039 23752
rect 19981 23743 20039 23749
rect 8686 23616 9168 23644
rect 13608 23647 13666 23653
rect 8686 23613 8698 23616
rect 8640 23607 8698 23613
rect 13608 23613 13620 23647
rect 13654 23644 13666 23647
rect 13906 23644 13912 23656
rect 13654 23616 13912 23644
rect 13654 23613 13666 23616
rect 13608 23607 13666 23613
rect 13906 23604 13912 23616
rect 13964 23644 13970 23656
rect 14001 23647 14059 23653
rect 14001 23644 14013 23647
rect 13964 23616 14013 23644
rect 13964 23604 13970 23616
rect 14001 23613 14013 23616
rect 14047 23613 14059 23647
rect 16022 23644 16028 23656
rect 15935 23616 16028 23644
rect 14001 23607 14059 23613
rect 16022 23604 16028 23616
rect 16080 23644 16086 23656
rect 16577 23647 16635 23653
rect 16577 23644 16589 23647
rect 16080 23616 16589 23644
rect 16080 23604 16086 23616
rect 16577 23613 16589 23616
rect 16623 23613 16635 23647
rect 18322 23644 18328 23656
rect 18235 23616 18328 23644
rect 16577 23607 16635 23613
rect 18322 23604 18328 23616
rect 18380 23644 18386 23656
rect 18877 23647 18935 23653
rect 18877 23644 18889 23647
rect 18380 23616 18889 23644
rect 18380 23604 18386 23616
rect 18877 23613 18889 23616
rect 18923 23613 18935 23647
rect 18877 23607 18935 23613
rect 19496 23647 19554 23653
rect 19496 23613 19508 23647
rect 19542 23644 19554 23647
rect 19996 23644 20024 23743
rect 24670 23740 24676 23752
rect 24728 23740 24734 23792
rect 19542 23616 20024 23644
rect 20441 23647 20499 23653
rect 19542 23613 19554 23616
rect 19496 23607 19554 23613
rect 20441 23613 20453 23647
rect 20487 23613 20499 23647
rect 20441 23607 20499 23613
rect 24648 23647 24706 23653
rect 24648 23613 24660 23647
rect 24694 23644 24706 23647
rect 25130 23644 25136 23656
rect 24694 23616 25136 23644
rect 24694 23613 24706 23616
rect 24648 23607 24706 23613
rect 1535 23579 1593 23585
rect 1535 23545 1547 23579
rect 1581 23576 1593 23579
rect 3786 23576 3792 23588
rect 1581 23548 3792 23576
rect 1581 23545 1593 23548
rect 1535 23539 1593 23545
rect 3786 23536 3792 23548
rect 3844 23536 3850 23588
rect 19334 23536 19340 23588
rect 19392 23576 19398 23588
rect 20456 23576 20484 23607
rect 25130 23604 25136 23616
rect 25188 23604 25194 23656
rect 20993 23579 21051 23585
rect 20993 23576 21005 23579
rect 19392 23548 21005 23576
rect 19392 23536 19398 23548
rect 20993 23545 21005 23548
rect 21039 23545 21051 23579
rect 20993 23539 21051 23545
rect 5905 23511 5963 23517
rect 5905 23477 5917 23511
rect 5951 23508 5963 23511
rect 6086 23508 6092 23520
rect 5951 23480 6092 23508
rect 5951 23477 5963 23480
rect 5905 23471 5963 23477
rect 6086 23468 6092 23480
rect 6144 23468 6150 23520
rect 7006 23508 7012 23520
rect 6967 23480 7012 23508
rect 7006 23468 7012 23480
rect 7064 23468 7070 23520
rect 8110 23468 8116 23520
rect 8168 23508 8174 23520
rect 8711 23511 8769 23517
rect 8711 23508 8723 23511
rect 8168 23480 8723 23508
rect 8168 23468 8174 23480
rect 8711 23477 8723 23480
rect 8757 23477 8769 23511
rect 8711 23471 8769 23477
rect 13679 23511 13737 23517
rect 13679 23477 13691 23511
rect 13725 23508 13737 23511
rect 13814 23508 13820 23520
rect 13725 23480 13820 23508
rect 13725 23477 13737 23480
rect 13679 23471 13737 23477
rect 13814 23468 13820 23480
rect 13872 23468 13878 23520
rect 19426 23468 19432 23520
rect 19484 23508 19490 23520
rect 19567 23511 19625 23517
rect 19567 23508 19579 23511
rect 19484 23480 19579 23508
rect 19484 23468 19490 23480
rect 19567 23477 19579 23480
rect 19613 23477 19625 23511
rect 19567 23471 19625 23477
rect 22738 23468 22744 23520
rect 22796 23508 22802 23520
rect 24719 23511 24777 23517
rect 24719 23508 24731 23511
rect 22796 23480 24731 23508
rect 22796 23468 22802 23480
rect 24719 23477 24731 23480
rect 24765 23477 24777 23511
rect 24719 23471 24777 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 7466 23304 7472 23316
rect 6104 23276 7472 23304
rect 106 23128 112 23180
rect 164 23168 170 23180
rect 1432 23171 1490 23177
rect 1432 23168 1444 23171
rect 164 23140 1444 23168
rect 164 23128 170 23140
rect 1432 23137 1444 23140
rect 1478 23168 1490 23171
rect 1578 23168 1584 23180
rect 1478 23140 1584 23168
rect 1478 23137 1490 23140
rect 1432 23131 1490 23137
rect 1578 23128 1584 23140
rect 1636 23128 1642 23180
rect 5350 23177 5356 23180
rect 5328 23171 5356 23177
rect 5328 23168 5340 23171
rect 5263 23140 5340 23168
rect 5328 23137 5340 23140
rect 5408 23168 5414 23180
rect 6104 23168 6132 23276
rect 7466 23264 7472 23276
rect 7524 23264 7530 23316
rect 11057 23307 11115 23313
rect 11057 23273 11069 23307
rect 11103 23304 11115 23307
rect 11698 23304 11704 23316
rect 11103 23276 11704 23304
rect 11103 23273 11115 23276
rect 11057 23267 11115 23273
rect 11698 23264 11704 23276
rect 11756 23264 11762 23316
rect 15427 23307 15485 23313
rect 15427 23273 15439 23307
rect 15473 23304 15485 23307
rect 16022 23304 16028 23316
rect 15473 23276 16028 23304
rect 15473 23273 15485 23276
rect 15427 23267 15485 23273
rect 16022 23264 16028 23276
rect 16080 23264 16086 23316
rect 6454 23236 6460 23248
rect 6415 23208 6460 23236
rect 6454 23196 6460 23208
rect 6512 23196 6518 23248
rect 8018 23236 8024 23248
rect 7979 23208 8024 23236
rect 8018 23196 8024 23208
rect 8076 23196 8082 23248
rect 5408 23140 6132 23168
rect 10873 23171 10931 23177
rect 5328 23131 5356 23137
rect 5350 23128 5356 23131
rect 5408 23128 5414 23140
rect 10873 23137 10885 23171
rect 10919 23168 10931 23171
rect 11054 23168 11060 23180
rect 10919 23140 11060 23168
rect 10919 23137 10931 23140
rect 10873 23131 10931 23137
rect 11054 23128 11060 23140
rect 11112 23128 11118 23180
rect 15197 23171 15255 23177
rect 15197 23137 15209 23171
rect 15243 23168 15255 23171
rect 15286 23168 15292 23180
rect 15243 23140 15292 23168
rect 15243 23137 15255 23140
rect 15197 23131 15255 23137
rect 15286 23128 15292 23140
rect 15344 23128 15350 23180
rect 6365 23103 6423 23109
rect 6365 23100 6377 23103
rect 5552 23072 6377 23100
rect 5552 22976 5580 23072
rect 6365 23069 6377 23072
rect 6411 23069 6423 23103
rect 6365 23063 6423 23069
rect 6638 23060 6644 23112
rect 6696 23100 6702 23112
rect 7009 23103 7067 23109
rect 7009 23100 7021 23103
rect 6696 23072 7021 23100
rect 6696 23060 6702 23072
rect 7009 23069 7021 23072
rect 7055 23100 7067 23103
rect 7926 23100 7932 23112
rect 7055 23072 7932 23100
rect 7055 23069 7067 23072
rect 7009 23063 7067 23069
rect 7926 23060 7932 23072
rect 7984 23060 7990 23112
rect 8202 23100 8208 23112
rect 8163 23072 8208 23100
rect 8202 23060 8208 23072
rect 8260 23060 8266 23112
rect 1535 22967 1593 22973
rect 1535 22933 1547 22967
rect 1581 22964 1593 22967
rect 2498 22964 2504 22976
rect 1581 22936 2504 22964
rect 1581 22933 1593 22936
rect 1535 22927 1593 22933
rect 2498 22924 2504 22936
rect 2556 22924 2562 22976
rect 5399 22967 5457 22973
rect 5399 22933 5411 22967
rect 5445 22964 5457 22967
rect 5534 22964 5540 22976
rect 5445 22936 5540 22964
rect 5445 22933 5457 22936
rect 5399 22927 5457 22933
rect 5534 22924 5540 22936
rect 5592 22924 5598 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1578 22760 1584 22772
rect 1539 22732 1584 22760
rect 1578 22720 1584 22732
rect 1636 22720 1642 22772
rect 5350 22760 5356 22772
rect 5311 22732 5356 22760
rect 5350 22720 5356 22732
rect 5408 22720 5414 22772
rect 5534 22720 5540 22772
rect 5592 22760 5598 22772
rect 5905 22763 5963 22769
rect 5905 22760 5917 22763
rect 5592 22732 5917 22760
rect 5592 22720 5598 22732
rect 5905 22729 5917 22732
rect 5951 22729 5963 22763
rect 5905 22723 5963 22729
rect 7926 22720 7932 22772
rect 7984 22760 7990 22772
rect 8573 22763 8631 22769
rect 8573 22760 8585 22763
rect 7984 22732 8585 22760
rect 7984 22720 7990 22732
rect 8573 22729 8585 22732
rect 8619 22729 8631 22763
rect 8573 22723 8631 22729
rect 7006 22584 7012 22636
rect 7064 22624 7070 22636
rect 7285 22627 7343 22633
rect 7285 22624 7297 22627
rect 7064 22596 7297 22624
rect 7064 22584 7070 22596
rect 7285 22593 7297 22596
rect 7331 22593 7343 22627
rect 7285 22587 7343 22593
rect 7929 22627 7987 22633
rect 7929 22593 7941 22627
rect 7975 22624 7987 22627
rect 8202 22624 8208 22636
rect 7975 22596 8208 22624
rect 7975 22593 7987 22596
rect 7929 22587 7987 22593
rect 8202 22584 8208 22596
rect 8260 22584 8266 22636
rect 9217 22627 9275 22633
rect 9217 22624 9229 22627
rect 8807 22596 9229 22624
rect 8220 22556 8248 22584
rect 8807 22565 8835 22596
rect 9217 22593 9229 22596
rect 9263 22593 9275 22627
rect 9217 22587 9275 22593
rect 8792 22559 8850 22565
rect 8792 22556 8804 22559
rect 8220 22528 8804 22556
rect 8792 22525 8804 22528
rect 8838 22525 8850 22559
rect 8792 22519 8850 22525
rect 8895 22559 8953 22565
rect 8895 22525 8907 22559
rect 8941 22556 8953 22559
rect 10870 22556 10876 22568
rect 8941 22528 10876 22556
rect 8941 22525 8953 22528
rect 8895 22519 8953 22525
rect 10870 22516 10876 22528
rect 10928 22516 10934 22568
rect 7101 22491 7159 22497
rect 7101 22457 7113 22491
rect 7147 22488 7159 22491
rect 7374 22488 7380 22500
rect 7147 22460 7380 22488
rect 7147 22457 7159 22460
rect 7101 22451 7159 22457
rect 7374 22448 7380 22460
rect 7432 22448 7438 22500
rect 5994 22380 6000 22432
rect 6052 22420 6058 22432
rect 6273 22423 6331 22429
rect 6273 22420 6285 22423
rect 6052 22392 6285 22420
rect 6052 22380 6058 22392
rect 6273 22389 6285 22392
rect 6319 22420 6331 22423
rect 6454 22420 6460 22432
rect 6319 22392 6460 22420
rect 6319 22389 6331 22392
rect 6273 22383 6331 22389
rect 6454 22380 6460 22392
rect 6512 22380 6518 22432
rect 8018 22380 8024 22432
rect 8076 22420 8082 22432
rect 8202 22420 8208 22432
rect 8076 22392 8208 22420
rect 8076 22380 8082 22392
rect 8202 22380 8208 22392
rect 8260 22380 8266 22432
rect 10962 22420 10968 22432
rect 10923 22392 10968 22420
rect 10962 22380 10968 22392
rect 11020 22380 11026 22432
rect 13998 22380 14004 22432
rect 14056 22420 14062 22432
rect 15286 22420 15292 22432
rect 14056 22392 15292 22420
rect 14056 22380 14062 22392
rect 15286 22380 15292 22392
rect 15344 22380 15350 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 6086 22216 6092 22228
rect 6047 22188 6092 22216
rect 6086 22176 6092 22188
rect 6144 22176 6150 22228
rect 7006 22176 7012 22228
rect 7064 22216 7070 22228
rect 7193 22219 7251 22225
rect 7193 22216 7205 22219
rect 7064 22188 7205 22216
rect 7064 22176 7070 22188
rect 7193 22185 7205 22188
rect 7239 22185 7251 22219
rect 7193 22179 7251 22185
rect 10962 22176 10968 22228
rect 11020 22216 11026 22228
rect 11471 22219 11529 22225
rect 11471 22216 11483 22219
rect 11020 22188 11483 22216
rect 11020 22176 11026 22188
rect 11471 22185 11483 22188
rect 11517 22185 11529 22219
rect 11471 22179 11529 22185
rect 7374 22148 7380 22160
rect 7335 22120 7380 22148
rect 7374 22108 7380 22120
rect 7432 22108 7438 22160
rect 5994 22080 6000 22092
rect 5955 22052 6000 22080
rect 5994 22040 6000 22052
rect 6052 22040 6058 22092
rect 7469 22083 7527 22089
rect 7469 22049 7481 22083
rect 7515 22080 7527 22083
rect 8202 22080 8208 22092
rect 7515 22052 8208 22080
rect 7515 22049 7527 22052
rect 7469 22043 7527 22049
rect 7374 21972 7380 22024
rect 7432 22012 7438 22024
rect 7484 22012 7512 22043
rect 8202 22040 8208 22052
rect 8260 22040 8266 22092
rect 11400 22083 11458 22089
rect 11400 22049 11412 22083
rect 11446 22080 11458 22083
rect 11790 22080 11796 22092
rect 11446 22052 11796 22080
rect 11446 22049 11458 22052
rect 11400 22043 11458 22049
rect 11790 22040 11796 22052
rect 11848 22040 11854 22092
rect 13792 22083 13850 22089
rect 13792 22049 13804 22083
rect 13838 22080 13850 22083
rect 13906 22080 13912 22092
rect 13838 22052 13912 22080
rect 13838 22049 13850 22052
rect 13792 22043 13850 22049
rect 13906 22040 13912 22052
rect 13964 22040 13970 22092
rect 7432 21984 7512 22012
rect 7432 21972 7438 21984
rect 12526 21876 12532 21888
rect 12487 21848 12532 21876
rect 12526 21836 12532 21848
rect 12584 21836 12590 21888
rect 12894 21836 12900 21888
rect 12952 21876 12958 21888
rect 13863 21879 13921 21885
rect 13863 21876 13875 21879
rect 12952 21848 13875 21876
rect 12952 21836 12958 21848
rect 13863 21845 13875 21848
rect 13909 21845 13921 21879
rect 13863 21839 13921 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 11790 21672 11796 21684
rect 11751 21644 11796 21672
rect 11790 21632 11796 21644
rect 11848 21632 11854 21684
rect 13817 21675 13875 21681
rect 13817 21641 13829 21675
rect 13863 21672 13875 21675
rect 13906 21672 13912 21684
rect 13863 21644 13912 21672
rect 13863 21641 13875 21644
rect 13817 21635 13875 21641
rect 13906 21632 13912 21644
rect 13964 21672 13970 21684
rect 15746 21672 15752 21684
rect 13964 21644 15752 21672
rect 13964 21632 13970 21644
rect 15746 21632 15752 21644
rect 15804 21632 15810 21684
rect 11808 21604 11836 21632
rect 11808 21576 12848 21604
rect 12526 21536 12532 21548
rect 12487 21508 12532 21536
rect 12526 21496 12532 21508
rect 12584 21496 12590 21548
rect 12820 21545 12848 21576
rect 12805 21539 12863 21545
rect 12805 21505 12817 21539
rect 12851 21505 12863 21539
rect 12805 21499 12863 21505
rect 1210 21428 1216 21480
rect 1268 21468 1274 21480
rect 1432 21471 1490 21477
rect 1432 21468 1444 21471
rect 1268 21440 1444 21468
rect 1268 21428 1274 21440
rect 1432 21437 1444 21440
rect 1478 21468 1490 21471
rect 1857 21471 1915 21477
rect 1857 21468 1869 21471
rect 1478 21440 1869 21468
rect 1478 21437 1490 21440
rect 1432 21431 1490 21437
rect 1857 21437 1869 21440
rect 1903 21437 1915 21471
rect 1857 21431 1915 21437
rect 10689 21471 10747 21477
rect 10689 21437 10701 21471
rect 10735 21468 10747 21471
rect 11422 21468 11428 21480
rect 10735 21440 11428 21468
rect 10735 21437 10747 21440
rect 10689 21431 10747 21437
rect 11422 21428 11428 21440
rect 11480 21468 11486 21480
rect 12161 21471 12219 21477
rect 12161 21468 12173 21471
rect 11480 21440 12173 21468
rect 11480 21428 11486 21440
rect 12161 21437 12173 21440
rect 12207 21437 12219 21471
rect 12161 21431 12219 21437
rect 1535 21403 1593 21409
rect 1535 21369 1547 21403
rect 1581 21400 1593 21403
rect 11514 21400 11520 21412
rect 1581 21372 7604 21400
rect 11475 21372 11520 21400
rect 1581 21369 1593 21372
rect 1535 21363 1593 21369
rect 5074 21292 5080 21344
rect 5132 21332 5138 21344
rect 5813 21335 5871 21341
rect 5813 21332 5825 21335
rect 5132 21304 5825 21332
rect 5132 21292 5138 21304
rect 5813 21301 5825 21304
rect 5859 21332 5871 21335
rect 5994 21332 6000 21344
rect 5859 21304 6000 21332
rect 5859 21301 5871 21304
rect 5813 21295 5871 21301
rect 5994 21292 6000 21304
rect 6052 21292 6058 21344
rect 7374 21332 7380 21344
rect 7335 21304 7380 21332
rect 7374 21292 7380 21304
rect 7432 21292 7438 21344
rect 7576 21332 7604 21372
rect 11514 21360 11520 21372
rect 11572 21360 11578 21412
rect 12176 21400 12204 21431
rect 12621 21403 12679 21409
rect 12621 21400 12633 21403
rect 12176 21372 12633 21400
rect 12621 21369 12633 21372
rect 12667 21369 12679 21403
rect 12621 21363 12679 21369
rect 11698 21332 11704 21344
rect 7576 21304 11704 21332
rect 11698 21292 11704 21304
rect 11756 21292 11762 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 11425 21063 11483 21069
rect 11425 21029 11437 21063
rect 11471 21060 11483 21063
rect 11514 21060 11520 21072
rect 11471 21032 11520 21060
rect 11471 21029 11483 21032
rect 11425 21023 11483 21029
rect 11514 21020 11520 21032
rect 11572 21020 11578 21072
rect 12894 21060 12900 21072
rect 12855 21032 12900 21060
rect 12894 21020 12900 21032
rect 12952 21020 12958 21072
rect 12989 21063 13047 21069
rect 12989 21029 13001 21063
rect 13035 21060 13047 21063
rect 13078 21060 13084 21072
rect 13035 21032 13084 21060
rect 13035 21029 13047 21032
rect 12989 21023 13047 21029
rect 13078 21020 13084 21032
rect 13136 21020 13142 21072
rect 24581 20995 24639 21001
rect 24581 20961 24593 20995
rect 24627 20992 24639 20995
rect 24670 20992 24676 21004
rect 24627 20964 24676 20992
rect 24627 20961 24639 20964
rect 24581 20955 24639 20961
rect 24670 20952 24676 20964
rect 24728 20952 24734 21004
rect 11330 20924 11336 20936
rect 11291 20896 11336 20924
rect 11330 20884 11336 20896
rect 11388 20884 11394 20936
rect 11790 20924 11796 20936
rect 11751 20896 11796 20924
rect 11790 20884 11796 20896
rect 11848 20884 11854 20936
rect 13173 20927 13231 20933
rect 13173 20893 13185 20927
rect 13219 20893 13231 20927
rect 13173 20887 13231 20893
rect 12526 20816 12532 20868
rect 12584 20856 12590 20868
rect 12986 20856 12992 20868
rect 12584 20828 12992 20856
rect 12584 20816 12590 20828
rect 12986 20816 12992 20828
rect 13044 20856 13050 20868
rect 13188 20856 13216 20887
rect 13044 20828 13216 20856
rect 13044 20816 13050 20828
rect 12710 20788 12716 20800
rect 12671 20760 12716 20788
rect 12710 20748 12716 20760
rect 12768 20748 12774 20800
rect 15654 20748 15660 20800
rect 15712 20788 15718 20800
rect 24719 20791 24777 20797
rect 24719 20788 24731 20791
rect 15712 20760 24731 20788
rect 15712 20748 15718 20760
rect 24719 20757 24731 20760
rect 24765 20757 24777 20791
rect 24719 20751 24777 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 11241 20587 11299 20593
rect 11241 20553 11253 20587
rect 11287 20584 11299 20587
rect 11330 20584 11336 20596
rect 11287 20556 11336 20584
rect 11287 20553 11299 20556
rect 11241 20547 11299 20553
rect 11330 20544 11336 20556
rect 11388 20544 11394 20596
rect 11514 20544 11520 20596
rect 11572 20584 11578 20596
rect 11793 20587 11851 20593
rect 11793 20584 11805 20587
rect 11572 20556 11805 20584
rect 11572 20544 11578 20556
rect 11793 20553 11805 20556
rect 11839 20553 11851 20587
rect 24670 20584 24676 20596
rect 24631 20556 24676 20584
rect 11793 20547 11851 20553
rect 24670 20544 24676 20556
rect 24728 20544 24734 20596
rect 11348 20457 11376 20544
rect 11333 20451 11391 20457
rect 11333 20417 11345 20451
rect 11379 20417 11391 20451
rect 12710 20448 12716 20460
rect 12671 20420 12716 20448
rect 11333 20411 11391 20417
rect 12710 20408 12716 20420
rect 12768 20408 12774 20460
rect 12986 20448 12992 20460
rect 12947 20420 12992 20448
rect 12986 20408 12992 20420
rect 13044 20408 13050 20460
rect 12805 20315 12863 20321
rect 12805 20312 12817 20315
rect 12176 20284 12817 20312
rect 12176 20256 12204 20284
rect 12805 20281 12817 20284
rect 12851 20281 12863 20315
rect 12805 20275 12863 20281
rect 12158 20244 12164 20256
rect 12119 20216 12164 20244
rect 12158 20204 12164 20216
rect 12216 20204 12222 20256
rect 13078 20204 13084 20256
rect 13136 20244 13142 20256
rect 13633 20247 13691 20253
rect 13633 20244 13645 20247
rect 13136 20216 13645 20244
rect 13136 20204 13142 20216
rect 13633 20213 13645 20216
rect 13679 20213 13691 20247
rect 13633 20207 13691 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 12894 20000 12900 20052
rect 12952 20040 12958 20052
rect 13357 20043 13415 20049
rect 13357 20040 13369 20043
rect 12952 20012 13369 20040
rect 12952 20000 12958 20012
rect 13357 20009 13369 20012
rect 13403 20009 13415 20043
rect 13357 20003 13415 20009
rect 13078 19972 13084 19984
rect 13039 19944 13084 19972
rect 13078 19932 13084 19944
rect 13136 19932 13142 19984
rect 12158 19864 12164 19916
rect 12216 19904 12222 19916
rect 12437 19907 12495 19913
rect 12437 19904 12449 19907
rect 12216 19876 12449 19904
rect 12216 19864 12222 19876
rect 12437 19873 12449 19876
rect 12483 19873 12495 19907
rect 12437 19867 12495 19873
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 12158 19116 12164 19168
rect 12216 19156 12222 19168
rect 12621 19159 12679 19165
rect 12621 19156 12633 19159
rect 12216 19128 12633 19156
rect 12216 19116 12222 19128
rect 12621 19125 12633 19128
rect 12667 19125 12679 19159
rect 12621 19119 12679 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 11514 17864 11520 17876
rect 11475 17836 11520 17864
rect 11514 17824 11520 17836
rect 11572 17824 11578 17876
rect 24762 17864 24768 17876
rect 24723 17836 24768 17864
rect 24762 17824 24768 17836
rect 24820 17824 24826 17876
rect 11333 17731 11391 17737
rect 11333 17697 11345 17731
rect 11379 17728 11391 17731
rect 11606 17728 11612 17740
rect 11379 17700 11612 17728
rect 11379 17697 11391 17700
rect 11333 17691 11391 17697
rect 11606 17688 11612 17700
rect 11664 17688 11670 17740
rect 24210 17688 24216 17740
rect 24268 17728 24274 17740
rect 24581 17731 24639 17737
rect 24581 17728 24593 17731
rect 24268 17700 24593 17728
rect 24268 17688 24274 17700
rect 24581 17697 24593 17700
rect 24627 17697 24639 17731
rect 24581 17691 24639 17697
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 11425 16983 11483 16989
rect 11425 16949 11437 16983
rect 11471 16980 11483 16983
rect 11606 16980 11612 16992
rect 11471 16952 11612 16980
rect 11471 16949 11483 16952
rect 11425 16943 11483 16949
rect 11606 16940 11612 16952
rect 11664 16940 11670 16992
rect 24210 16940 24216 16992
rect 24268 16980 24274 16992
rect 24581 16983 24639 16989
rect 24581 16980 24593 16983
rect 24268 16952 24593 16980
rect 24268 16940 24274 16952
rect 24581 16949 24593 16952
rect 24627 16949 24639 16983
rect 24581 16943 24639 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 198 16600 204 16652
rect 256 16640 262 16652
rect 6362 16640 6368 16652
rect 6420 16649 6426 16652
rect 6420 16643 6458 16649
rect 256 16612 6368 16640
rect 256 16600 262 16612
rect 6362 16600 6368 16612
rect 6446 16609 6458 16643
rect 8202 16640 8208 16652
rect 8163 16612 8208 16640
rect 6420 16603 6458 16609
rect 6420 16600 6426 16603
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 7558 16572 7564 16584
rect 7519 16544 7564 16572
rect 7558 16532 7564 16544
rect 7616 16532 7622 16584
rect 6503 16439 6561 16445
rect 6503 16405 6515 16439
rect 6549 16436 6561 16439
rect 7466 16436 7472 16448
rect 6549 16408 7472 16436
rect 6549 16405 6561 16408
rect 6503 16399 6561 16405
rect 7466 16396 7472 16408
rect 7524 16396 7530 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 6362 16232 6368 16244
rect 6323 16204 6368 16232
rect 6362 16192 6368 16204
rect 6420 16192 6426 16244
rect 25133 16235 25191 16241
rect 25133 16201 25145 16235
rect 25179 16232 25191 16235
rect 26418 16232 26424 16244
rect 25179 16204 26424 16232
rect 25179 16201 25191 16204
rect 25133 16195 25191 16201
rect 7926 16124 7932 16176
rect 7984 16164 7990 16176
rect 8757 16167 8815 16173
rect 8757 16164 8769 16167
rect 7984 16136 8769 16164
rect 7984 16124 7990 16136
rect 8757 16133 8769 16136
rect 8803 16133 8815 16167
rect 8757 16127 8815 16133
rect 8205 16099 8263 16105
rect 8205 16065 8217 16099
rect 8251 16096 8263 16099
rect 8478 16096 8484 16108
rect 8251 16068 8484 16096
rect 8251 16065 8263 16068
rect 8205 16059 8263 16065
rect 8478 16056 8484 16068
rect 8536 16056 8542 16108
rect 7098 16028 7104 16040
rect 7059 16000 7104 16028
rect 7098 15988 7104 16000
rect 7156 15988 7162 16040
rect 24648 16031 24706 16037
rect 24648 15997 24660 16031
rect 24694 16028 24706 16031
rect 25148 16028 25176 16195
rect 26418 16192 26424 16204
rect 26476 16192 26482 16244
rect 24694 16000 25176 16028
rect 24694 15997 24706 16000
rect 24648 15991 24706 15997
rect 7239 15963 7297 15969
rect 7239 15960 7251 15963
rect 4126 15932 7251 15960
rect 2406 15852 2412 15904
rect 2464 15892 2470 15904
rect 4126 15892 4154 15932
rect 7239 15929 7251 15932
rect 7285 15929 7297 15963
rect 7239 15923 7297 15929
rect 7653 15963 7711 15969
rect 7653 15929 7665 15963
rect 7699 15960 7711 15963
rect 8021 15963 8079 15969
rect 8021 15960 8033 15963
rect 7699 15932 8033 15960
rect 7699 15929 7711 15932
rect 7653 15923 7711 15929
rect 8021 15929 8033 15932
rect 8067 15960 8079 15963
rect 8202 15960 8208 15972
rect 8067 15932 8208 15960
rect 8067 15929 8079 15932
rect 8021 15923 8079 15929
rect 8202 15920 8208 15932
rect 8260 15960 8266 15972
rect 8297 15963 8355 15969
rect 8297 15960 8309 15963
rect 8260 15932 8309 15960
rect 8260 15920 8266 15932
rect 8297 15929 8309 15932
rect 8343 15929 8355 15963
rect 8297 15923 8355 15929
rect 2464 15864 4154 15892
rect 2464 15852 2470 15864
rect 15654 15852 15660 15904
rect 15712 15892 15718 15904
rect 24719 15895 24777 15901
rect 24719 15892 24731 15895
rect 15712 15864 24731 15892
rect 15712 15852 15718 15864
rect 24719 15861 24731 15864
rect 24765 15861 24777 15895
rect 24719 15855 24777 15861
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 18414 15648 18420 15700
rect 18472 15688 18478 15700
rect 19426 15688 19432 15700
rect 18472 15660 19432 15688
rect 18472 15648 18478 15660
rect 19426 15648 19432 15660
rect 19484 15648 19490 15700
rect 7558 15620 7564 15632
rect 7519 15592 7564 15620
rect 7558 15580 7564 15592
rect 7616 15580 7622 15632
rect 6086 15552 6092 15564
rect 6047 15524 6092 15552
rect 6086 15512 6092 15524
rect 6144 15512 6150 15564
rect 6549 15487 6607 15493
rect 6549 15453 6561 15487
rect 6595 15484 6607 15487
rect 6730 15484 6736 15496
rect 6595 15456 6736 15484
rect 6595 15453 6607 15456
rect 6549 15447 6607 15453
rect 6730 15444 6736 15456
rect 6788 15444 6794 15496
rect 7466 15484 7472 15496
rect 7427 15456 7472 15484
rect 7466 15444 7472 15456
rect 7524 15444 7530 15496
rect 7926 15484 7932 15496
rect 7887 15456 7932 15484
rect 7926 15444 7932 15456
rect 7984 15444 7990 15496
rect 7098 15308 7104 15360
rect 7156 15348 7162 15360
rect 7193 15351 7251 15357
rect 7193 15348 7205 15351
rect 7156 15320 7205 15348
rect 7156 15308 7162 15320
rect 7193 15317 7205 15320
rect 7239 15348 7251 15351
rect 8294 15348 8300 15360
rect 7239 15320 8300 15348
rect 7239 15317 7251 15320
rect 7193 15311 7251 15317
rect 8294 15308 8300 15320
rect 8352 15308 8358 15360
rect 8478 15348 8484 15360
rect 8439 15320 8484 15348
rect 8478 15308 8484 15320
rect 8536 15308 8542 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 6086 15144 6092 15156
rect 6047 15116 6092 15144
rect 6086 15104 6092 15116
rect 6144 15104 6150 15156
rect 7469 15147 7527 15153
rect 7469 15113 7481 15147
rect 7515 15144 7527 15147
rect 7558 15144 7564 15156
rect 7515 15116 7564 15144
rect 7515 15113 7527 15116
rect 7469 15107 7527 15113
rect 7558 15104 7564 15116
rect 7616 15104 7622 15156
rect 14182 15144 14188 15156
rect 14143 15116 14188 15144
rect 14182 15104 14188 15116
rect 14240 15104 14246 15156
rect 24762 15144 24768 15156
rect 24723 15116 24768 15144
rect 24762 15104 24768 15116
rect 24820 15104 24826 15156
rect 8294 15076 8300 15088
rect 8255 15048 8300 15076
rect 8294 15036 8300 15048
rect 8352 15036 8358 15088
rect 7466 14968 7472 15020
rect 7524 15008 7530 15020
rect 8665 15011 8723 15017
rect 8665 15008 8677 15011
rect 7524 14980 8677 15008
rect 7524 14968 7530 14980
rect 8665 14977 8677 14980
rect 8711 14977 8723 15011
rect 24486 15008 24492 15020
rect 24447 14980 24492 15008
rect 8665 14971 8723 14977
rect 24486 14968 24492 14980
rect 24544 15008 24550 15020
rect 25133 15011 25191 15017
rect 25133 15008 25145 15011
rect 24544 14980 25145 15008
rect 24544 14968 24550 14980
rect 25133 14977 25145 14980
rect 25179 14977 25191 15011
rect 25133 14971 25191 14977
rect 5696 14943 5754 14949
rect 5696 14909 5708 14943
rect 5742 14940 5754 14943
rect 9122 14940 9128 14952
rect 5742 14912 6316 14940
rect 9035 14912 9128 14940
rect 5742 14909 5754 14912
rect 5696 14903 5754 14909
rect 6288 14816 6316 14912
rect 9122 14900 9128 14912
rect 9180 14940 9186 14952
rect 9309 14943 9367 14949
rect 9309 14940 9321 14943
rect 9180 14912 9321 14940
rect 9180 14900 9186 14912
rect 9309 14909 9321 14912
rect 9355 14909 9367 14943
rect 9309 14903 9367 14909
rect 14001 14943 14059 14949
rect 14001 14909 14013 14943
rect 14047 14940 14059 14943
rect 14047 14912 14688 14940
rect 14047 14909 14059 14912
rect 14001 14903 14059 14909
rect 7745 14875 7803 14881
rect 7745 14872 7757 14875
rect 7024 14844 7757 14872
rect 7024 14816 7052 14844
rect 7745 14841 7757 14844
rect 7791 14841 7803 14875
rect 7745 14835 7803 14841
rect 7846 14875 7904 14881
rect 7846 14841 7858 14875
rect 7892 14872 7904 14875
rect 8018 14872 8024 14884
rect 7892 14844 8024 14872
rect 7892 14841 7904 14844
rect 7846 14835 7904 14841
rect 8018 14832 8024 14844
rect 8076 14872 8082 14884
rect 9217 14875 9275 14881
rect 9217 14872 9229 14875
rect 8076 14844 9229 14872
rect 8076 14832 8082 14844
rect 9217 14841 9229 14844
rect 9263 14841 9275 14875
rect 9217 14835 9275 14841
rect 5767 14807 5825 14813
rect 5767 14773 5779 14807
rect 5813 14804 5825 14807
rect 6178 14804 6184 14816
rect 5813 14776 6184 14804
rect 5813 14773 5825 14776
rect 5767 14767 5825 14773
rect 6178 14764 6184 14776
rect 6236 14764 6242 14816
rect 6270 14764 6276 14816
rect 6328 14804 6334 14816
rect 6457 14807 6515 14813
rect 6457 14804 6469 14807
rect 6328 14776 6469 14804
rect 6328 14764 6334 14776
rect 6457 14773 6469 14776
rect 6503 14773 6515 14807
rect 7006 14804 7012 14816
rect 6967 14776 7012 14804
rect 6457 14767 6515 14773
rect 7006 14764 7012 14776
rect 7064 14764 7070 14816
rect 14660 14813 14688 14912
rect 14645 14807 14703 14813
rect 14645 14773 14657 14807
rect 14691 14804 14703 14807
rect 15838 14804 15844 14816
rect 14691 14776 15844 14804
rect 14691 14773 14703 14776
rect 14645 14767 14703 14773
rect 15838 14764 15844 14776
rect 15896 14764 15902 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 6178 14560 6184 14612
rect 6236 14600 6242 14612
rect 6457 14603 6515 14609
rect 6457 14600 6469 14603
rect 6236 14572 6469 14600
rect 6236 14560 6242 14572
rect 6457 14569 6469 14572
rect 6503 14569 6515 14603
rect 6457 14563 6515 14569
rect 8570 14560 8576 14612
rect 8628 14600 8634 14612
rect 9769 14603 9827 14609
rect 9769 14600 9781 14603
rect 8628 14572 9781 14600
rect 8628 14560 8634 14572
rect 9769 14569 9781 14572
rect 9815 14569 9827 14603
rect 9769 14563 9827 14569
rect 5077 14535 5135 14541
rect 5077 14501 5089 14535
rect 5123 14532 5135 14535
rect 7006 14532 7012 14544
rect 5123 14504 7012 14532
rect 5123 14501 5135 14504
rect 5077 14495 5135 14501
rect 7006 14492 7012 14504
rect 7064 14492 7070 14544
rect 8021 14535 8079 14541
rect 8021 14501 8033 14535
rect 8067 14532 8079 14535
rect 8386 14532 8392 14544
rect 8067 14504 8392 14532
rect 8067 14501 8079 14504
rect 8021 14495 8079 14501
rect 8386 14492 8392 14504
rect 8444 14532 8450 14544
rect 9122 14532 9128 14544
rect 8444 14504 9128 14532
rect 8444 14492 8450 14504
rect 9122 14492 9128 14504
rect 9180 14492 9186 14544
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14464 1455 14467
rect 2406 14464 2412 14476
rect 1443 14436 2412 14464
rect 1443 14433 1455 14436
rect 1397 14427 1455 14433
rect 2406 14424 2412 14436
rect 2464 14424 2470 14476
rect 9674 14464 9680 14476
rect 9635 14436 9680 14464
rect 9674 14424 9680 14436
rect 9732 14424 9738 14476
rect 10134 14464 10140 14476
rect 10095 14436 10140 14464
rect 10134 14424 10140 14436
rect 10192 14424 10198 14476
rect 24581 14467 24639 14473
rect 24581 14433 24593 14467
rect 24627 14464 24639 14467
rect 24670 14464 24676 14476
rect 24627 14436 24676 14464
rect 24627 14433 24639 14436
rect 24581 14427 24639 14433
rect 24670 14424 24676 14436
rect 24728 14424 24734 14476
rect 6089 14399 6147 14405
rect 6089 14365 6101 14399
rect 6135 14396 6147 14399
rect 6546 14396 6552 14408
rect 6135 14368 6552 14396
rect 6135 14365 6147 14368
rect 6089 14359 6147 14365
rect 6546 14356 6552 14368
rect 6604 14356 6610 14408
rect 7466 14356 7472 14408
rect 7524 14396 7530 14408
rect 7926 14396 7932 14408
rect 7524 14368 7932 14396
rect 7524 14356 7530 14368
rect 7926 14356 7932 14368
rect 7984 14356 7990 14408
rect 8294 14396 8300 14408
rect 8255 14368 8300 14396
rect 8294 14356 8300 14368
rect 8352 14356 8358 14408
rect 1578 14328 1584 14340
rect 1539 14300 1584 14328
rect 1578 14288 1584 14300
rect 1636 14288 1642 14340
rect 7009 14331 7067 14337
rect 7009 14297 7021 14331
rect 7055 14328 7067 14331
rect 7374 14328 7380 14340
rect 7055 14300 7380 14328
rect 7055 14297 7067 14300
rect 7009 14291 7067 14297
rect 7374 14288 7380 14300
rect 7432 14288 7438 14340
rect 7745 14331 7803 14337
rect 7745 14297 7757 14331
rect 7791 14328 7803 14331
rect 8018 14328 8024 14340
rect 7791 14300 8024 14328
rect 7791 14297 7803 14300
rect 7745 14291 7803 14297
rect 8018 14288 8024 14300
rect 8076 14288 8082 14340
rect 22002 14220 22008 14272
rect 22060 14260 22066 14272
rect 24719 14263 24777 14269
rect 24719 14260 24731 14263
rect 22060 14232 24731 14260
rect 22060 14220 22066 14232
rect 24719 14229 24731 14232
rect 24765 14229 24777 14263
rect 24719 14223 24777 14229
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 2406 14056 2412 14068
rect 2367 14028 2412 14056
rect 2406 14016 2412 14028
rect 2464 14016 2470 14068
rect 7101 14059 7159 14065
rect 7101 14025 7113 14059
rect 7147 14056 7159 14059
rect 8386 14056 8392 14068
rect 7147 14028 8392 14056
rect 7147 14025 7159 14028
rect 7101 14019 7159 14025
rect 8386 14016 8392 14028
rect 8444 14056 8450 14068
rect 8481 14059 8539 14065
rect 8481 14056 8493 14059
rect 8444 14028 8493 14056
rect 8444 14016 8450 14028
rect 8481 14025 8493 14028
rect 8527 14025 8539 14059
rect 11422 14056 11428 14068
rect 11383 14028 11428 14056
rect 8481 14019 8539 14025
rect 11422 14016 11428 14028
rect 11480 14016 11486 14068
rect 24670 14056 24676 14068
rect 24631 14028 24676 14056
rect 24670 14016 24676 14028
rect 24728 14016 24734 14068
rect 14 13880 20 13932
rect 72 13920 78 13932
rect 4246 13920 4252 13932
rect 72 13892 4252 13920
rect 72 13880 78 13892
rect 4246 13880 4252 13892
rect 4304 13880 4310 13932
rect 7561 13923 7619 13929
rect 7561 13889 7573 13923
rect 7607 13920 7619 13923
rect 8754 13920 8760 13932
rect 7607 13892 8760 13920
rect 7607 13889 7619 13892
rect 7561 13883 7619 13889
rect 8754 13880 8760 13892
rect 8812 13880 8818 13932
rect 10962 13880 10968 13932
rect 11020 13920 11026 13932
rect 11020 13892 12515 13920
rect 11020 13880 11026 13892
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13852 1455 13855
rect 1670 13852 1676 13864
rect 1443 13824 1676 13852
rect 1443 13821 1455 13824
rect 1397 13815 1455 13821
rect 1670 13812 1676 13824
rect 1728 13852 1734 13864
rect 1949 13855 2007 13861
rect 1949 13852 1961 13855
rect 1728 13824 1961 13852
rect 1728 13812 1734 13824
rect 1949 13821 1961 13824
rect 1995 13821 2007 13855
rect 1949 13815 2007 13821
rect 3053 13855 3111 13861
rect 3053 13821 3065 13855
rect 3099 13821 3111 13855
rect 3053 13815 3111 13821
rect 5077 13855 5135 13861
rect 5077 13821 5089 13855
rect 5123 13852 5135 13855
rect 5350 13852 5356 13864
rect 5123 13824 5356 13852
rect 5123 13821 5135 13824
rect 5077 13815 5135 13821
rect 2958 13784 2964 13796
rect 2919 13756 2964 13784
rect 2958 13744 2964 13756
rect 3016 13744 3022 13796
rect 1578 13716 1584 13728
rect 1539 13688 1584 13716
rect 1578 13676 1584 13688
rect 1636 13676 1642 13728
rect 2682 13676 2688 13728
rect 2740 13716 2746 13728
rect 2777 13719 2835 13725
rect 2777 13716 2789 13719
rect 2740 13688 2789 13716
rect 2740 13676 2746 13688
rect 2777 13685 2789 13688
rect 2823 13716 2835 13719
rect 3068 13716 3096 13815
rect 5350 13812 5356 13824
rect 5408 13812 5414 13864
rect 5718 13852 5724 13864
rect 5679 13824 5724 13852
rect 5718 13812 5724 13824
rect 5776 13812 5782 13864
rect 9214 13812 9220 13864
rect 9272 13852 9278 13864
rect 9344 13855 9402 13861
rect 9344 13852 9356 13855
rect 9272 13824 9356 13852
rect 9272 13812 9278 13824
rect 9344 13821 9356 13824
rect 9390 13821 9402 13855
rect 9344 13815 9402 13821
rect 10505 13855 10563 13861
rect 10505 13821 10517 13855
rect 10551 13852 10563 13855
rect 10686 13852 10692 13864
rect 10551 13824 10692 13852
rect 10551 13821 10563 13824
rect 10505 13815 10563 13821
rect 10686 13812 10692 13824
rect 10744 13812 10750 13864
rect 12487 13861 12515 13892
rect 13722 13880 13728 13932
rect 13780 13920 13786 13932
rect 14734 13920 14740 13932
rect 13780 13892 14740 13920
rect 13780 13880 13786 13892
rect 14734 13880 14740 13892
rect 14792 13880 14798 13932
rect 12472 13855 12530 13861
rect 12472 13821 12484 13855
rect 12518 13852 12530 13855
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 12518 13824 12909 13852
rect 12518 13821 12530 13824
rect 12472 13815 12530 13821
rect 12897 13821 12909 13824
rect 12943 13821 12955 13855
rect 12897 13815 12955 13821
rect 7926 13793 7932 13796
rect 7377 13787 7435 13793
rect 7377 13784 7389 13787
rect 6196 13756 7389 13784
rect 6196 13728 6224 13756
rect 7377 13753 7389 13756
rect 7423 13784 7435 13787
rect 7882 13787 7932 13793
rect 7882 13784 7894 13787
rect 7423 13756 7894 13784
rect 7423 13753 7435 13756
rect 7377 13747 7435 13753
rect 7882 13753 7894 13756
rect 7928 13753 7932 13787
rect 7882 13747 7932 13753
rect 7926 13744 7932 13747
rect 7984 13784 7990 13796
rect 7984 13756 9628 13784
rect 7984 13744 7990 13756
rect 5258 13716 5264 13728
rect 2823 13688 3096 13716
rect 5219 13688 5264 13716
rect 2823 13685 2835 13688
rect 2777 13679 2835 13685
rect 5258 13676 5264 13688
rect 5316 13676 5322 13728
rect 6178 13716 6184 13728
rect 6139 13688 6184 13716
rect 6178 13676 6184 13688
rect 6236 13676 6242 13728
rect 6546 13716 6552 13728
rect 6507 13688 6552 13716
rect 6546 13676 6552 13688
rect 6604 13676 6610 13728
rect 9030 13676 9036 13728
rect 9088 13716 9094 13728
rect 9125 13719 9183 13725
rect 9125 13716 9137 13719
rect 9088 13688 9137 13716
rect 9088 13676 9094 13688
rect 9125 13685 9137 13688
rect 9171 13685 9183 13719
rect 9125 13679 9183 13685
rect 9306 13676 9312 13728
rect 9364 13716 9370 13728
rect 9447 13719 9505 13725
rect 9447 13716 9459 13719
rect 9364 13688 9459 13716
rect 9364 13676 9370 13688
rect 9447 13685 9459 13688
rect 9493 13685 9505 13719
rect 9600 13716 9628 13756
rect 9674 13744 9680 13796
rect 9732 13784 9738 13796
rect 9769 13787 9827 13793
rect 9769 13784 9781 13787
rect 9732 13756 9781 13784
rect 9732 13744 9738 13756
rect 9769 13753 9781 13756
rect 9815 13753 9827 13787
rect 10826 13787 10884 13793
rect 10826 13784 10838 13787
rect 9769 13747 9827 13753
rect 10336 13756 10838 13784
rect 10336 13725 10364 13756
rect 10826 13753 10838 13756
rect 10872 13753 10884 13787
rect 10826 13747 10884 13753
rect 14829 13787 14887 13793
rect 14829 13753 14841 13787
rect 14875 13753 14887 13787
rect 14829 13747 14887 13753
rect 15381 13787 15439 13793
rect 15381 13753 15393 13787
rect 15427 13784 15439 13787
rect 15930 13784 15936 13796
rect 15427 13756 15936 13784
rect 15427 13753 15439 13756
rect 15381 13747 15439 13753
rect 10321 13719 10379 13725
rect 10321 13716 10333 13719
rect 9600 13688 10333 13716
rect 9447 13679 9505 13685
rect 10321 13685 10333 13688
rect 10367 13685 10379 13719
rect 10321 13679 10379 13685
rect 12575 13719 12633 13725
rect 12575 13685 12587 13719
rect 12621 13716 12633 13719
rect 14182 13716 14188 13728
rect 12621 13688 14188 13716
rect 12621 13685 12633 13688
rect 12575 13679 12633 13685
rect 14182 13676 14188 13688
rect 14240 13676 14246 13728
rect 14458 13716 14464 13728
rect 14419 13688 14464 13716
rect 14458 13676 14464 13688
rect 14516 13716 14522 13728
rect 14844 13716 14872 13747
rect 15930 13744 15936 13756
rect 15988 13744 15994 13796
rect 14516 13688 14872 13716
rect 14516 13676 14522 13688
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1535 13515 1593 13521
rect 1535 13481 1547 13515
rect 1581 13512 1593 13515
rect 1670 13512 1676 13524
rect 1581 13484 1676 13512
rect 1581 13481 1593 13484
rect 1535 13475 1593 13481
rect 1670 13472 1676 13484
rect 1728 13472 1734 13524
rect 5074 13472 5080 13524
rect 5132 13512 5138 13524
rect 6457 13515 6515 13521
rect 6457 13512 6469 13515
rect 5132 13484 6469 13512
rect 5132 13472 5138 13484
rect 6457 13481 6469 13484
rect 6503 13481 6515 13515
rect 7466 13512 7472 13524
rect 7427 13484 7472 13512
rect 6457 13475 6515 13481
rect 7466 13472 7472 13484
rect 7524 13472 7530 13524
rect 7926 13512 7932 13524
rect 7887 13484 7932 13512
rect 7926 13472 7932 13484
rect 7984 13472 7990 13524
rect 8202 13472 8208 13524
rect 8260 13512 8266 13524
rect 8481 13515 8539 13521
rect 8481 13512 8493 13515
rect 8260 13484 8493 13512
rect 8260 13472 8266 13484
rect 8481 13481 8493 13484
rect 8527 13481 8539 13515
rect 8481 13475 8539 13481
rect 8754 13472 8760 13524
rect 8812 13512 8818 13524
rect 9769 13515 9827 13521
rect 9769 13512 9781 13515
rect 8812 13484 9781 13512
rect 8812 13472 8818 13484
rect 9769 13481 9781 13484
rect 9815 13481 9827 13515
rect 9769 13475 9827 13481
rect 11609 13515 11667 13521
rect 11609 13481 11621 13515
rect 11655 13512 11667 13515
rect 11698 13512 11704 13524
rect 11655 13484 11704 13512
rect 11655 13481 11667 13484
rect 11609 13475 11667 13481
rect 11698 13472 11704 13484
rect 11756 13472 11762 13524
rect 12158 13512 12164 13524
rect 12119 13484 12164 13512
rect 12158 13472 12164 13484
rect 12216 13472 12222 13524
rect 14734 13512 14740 13524
rect 14695 13484 14740 13512
rect 14734 13472 14740 13484
rect 14792 13472 14798 13524
rect 2590 13444 2596 13456
rect 2551 13416 2596 13444
rect 2590 13404 2596 13416
rect 2648 13404 2654 13456
rect 5899 13447 5957 13453
rect 5899 13413 5911 13447
rect 5945 13444 5957 13447
rect 6178 13444 6184 13456
rect 5945 13416 6184 13444
rect 5945 13413 5957 13416
rect 5899 13407 5957 13413
rect 6178 13404 6184 13416
rect 6236 13404 6242 13456
rect 14369 13447 14427 13453
rect 14369 13413 14381 13447
rect 14415 13444 14427 13447
rect 14458 13444 14464 13456
rect 14415 13416 14464 13444
rect 14415 13413 14427 13416
rect 14369 13407 14427 13413
rect 14458 13404 14464 13416
rect 14516 13404 14522 13456
rect 15470 13444 15476 13456
rect 15431 13416 15476 13444
rect 15470 13404 15476 13416
rect 15528 13404 15534 13456
rect 1464 13379 1522 13385
rect 1464 13345 1476 13379
rect 1510 13376 1522 13379
rect 9674 13376 9680 13388
rect 1510 13348 1992 13376
rect 9635 13348 9680 13376
rect 1510 13345 1522 13348
rect 1464 13339 1522 13345
rect 1964 13181 1992 13348
rect 9674 13336 9680 13348
rect 9732 13336 9738 13388
rect 10134 13376 10140 13388
rect 10047 13348 10140 13376
rect 10134 13336 10140 13348
rect 10192 13336 10198 13388
rect 13722 13376 13728 13388
rect 13683 13348 13728 13376
rect 13722 13336 13728 13348
rect 13780 13336 13786 13388
rect 2314 13268 2320 13320
rect 2372 13308 2378 13320
rect 2498 13308 2504 13320
rect 2372 13280 2504 13308
rect 2372 13268 2378 13280
rect 2498 13268 2504 13280
rect 2556 13268 2562 13320
rect 2866 13308 2872 13320
rect 2827 13280 2872 13308
rect 2866 13268 2872 13280
rect 2924 13268 2930 13320
rect 4062 13308 4068 13320
rect 4023 13280 4068 13308
rect 4062 13268 4068 13280
rect 4120 13268 4126 13320
rect 5534 13308 5540 13320
rect 5495 13280 5540 13308
rect 5534 13268 5540 13280
rect 5592 13268 5598 13320
rect 7561 13311 7619 13317
rect 7561 13277 7573 13311
rect 7607 13308 7619 13311
rect 8570 13308 8576 13320
rect 7607 13280 8576 13308
rect 7607 13277 7619 13280
rect 7561 13271 7619 13277
rect 8570 13268 8576 13280
rect 8628 13268 8634 13320
rect 9030 13268 9036 13320
rect 9088 13308 9094 13320
rect 10152 13308 10180 13336
rect 11238 13308 11244 13320
rect 9088 13280 10180 13308
rect 11199 13280 11244 13308
rect 9088 13268 9094 13280
rect 11238 13268 11244 13280
rect 11296 13268 11302 13320
rect 15381 13311 15439 13317
rect 15381 13277 15393 13311
rect 15427 13308 15439 13311
rect 15746 13308 15752 13320
rect 15427 13280 15752 13308
rect 15427 13277 15439 13280
rect 15381 13271 15439 13277
rect 15746 13268 15752 13280
rect 15804 13308 15810 13320
rect 22002 13308 22008 13320
rect 15804 13280 22008 13308
rect 15804 13268 15810 13280
rect 22002 13268 22008 13280
rect 22060 13268 22066 13320
rect 2225 13243 2283 13249
rect 2225 13209 2237 13243
rect 2271 13240 2283 13243
rect 2884 13240 2912 13268
rect 2271 13212 2912 13240
rect 2271 13209 2283 13212
rect 2225 13203 2283 13209
rect 5718 13200 5724 13252
rect 5776 13200 5782 13252
rect 15930 13240 15936 13252
rect 15891 13212 15936 13240
rect 15930 13200 15936 13212
rect 15988 13200 15994 13252
rect 1949 13175 2007 13181
rect 1949 13141 1961 13175
rect 1995 13172 2007 13175
rect 3142 13172 3148 13184
rect 1995 13144 3148 13172
rect 1995 13141 2007 13144
rect 1949 13135 2007 13141
rect 3142 13132 3148 13144
rect 3200 13132 3206 13184
rect 5261 13175 5319 13181
rect 5261 13141 5273 13175
rect 5307 13172 5319 13175
rect 5736 13172 5764 13200
rect 7282 13172 7288 13184
rect 5307 13144 7288 13172
rect 5307 13141 5319 13144
rect 5261 13135 5319 13141
rect 7282 13132 7288 13144
rect 7340 13132 7346 13184
rect 7742 13132 7748 13184
rect 7800 13172 7806 13184
rect 9214 13172 9220 13184
rect 7800 13144 9220 13172
rect 7800 13132 7806 13144
rect 9214 13132 9220 13144
rect 9272 13172 9278 13184
rect 9309 13175 9367 13181
rect 9309 13172 9321 13175
rect 9272 13144 9321 13172
rect 9272 13132 9278 13144
rect 9309 13141 9321 13144
rect 9355 13141 9367 13175
rect 9309 13135 9367 13141
rect 10502 13132 10508 13184
rect 10560 13172 10566 13184
rect 10686 13172 10692 13184
rect 10560 13144 10692 13172
rect 10560 13132 10566 13144
rect 10686 13132 10692 13144
rect 10744 13132 10750 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 5350 12928 5356 12980
rect 5408 12968 5414 12980
rect 5408 12940 5625 12968
rect 5408 12928 5414 12940
rect 2682 12860 2688 12912
rect 2740 12900 2746 12912
rect 4249 12903 4307 12909
rect 4249 12900 4261 12903
rect 2740 12872 4261 12900
rect 2740 12860 2746 12872
rect 4249 12869 4261 12872
rect 4295 12869 4307 12903
rect 4249 12863 4307 12869
rect 4709 12903 4767 12909
rect 4709 12869 4721 12903
rect 4755 12900 4767 12903
rect 5597 12900 5625 12940
rect 6178 12928 6184 12980
rect 6236 12968 6242 12980
rect 7837 12971 7895 12977
rect 7837 12968 7849 12971
rect 6236 12940 7849 12968
rect 6236 12928 6242 12940
rect 7837 12937 7849 12940
rect 7883 12937 7895 12971
rect 7837 12931 7895 12937
rect 8297 12971 8355 12977
rect 8297 12937 8309 12971
rect 8343 12968 8355 12971
rect 8570 12968 8576 12980
rect 8343 12940 8576 12968
rect 8343 12937 8355 12940
rect 8297 12931 8355 12937
rect 8570 12928 8576 12940
rect 8628 12928 8634 12980
rect 11606 12928 11612 12980
rect 11664 12968 11670 12980
rect 12575 12971 12633 12977
rect 12575 12968 12587 12971
rect 11664 12940 12587 12968
rect 11664 12928 11670 12940
rect 12575 12937 12587 12940
rect 12621 12937 12633 12971
rect 12575 12931 12633 12937
rect 13633 12971 13691 12977
rect 13633 12937 13645 12971
rect 13679 12968 13691 12971
rect 13722 12968 13728 12980
rect 13679 12940 13728 12968
rect 13679 12937 13691 12940
rect 13633 12931 13691 12937
rect 13722 12928 13728 12940
rect 13780 12968 13786 12980
rect 15013 12971 15071 12977
rect 15013 12968 15025 12971
rect 13780 12940 15025 12968
rect 13780 12928 13786 12940
rect 15013 12937 15025 12940
rect 15059 12968 15071 12971
rect 15289 12971 15347 12977
rect 15289 12968 15301 12971
rect 15059 12940 15301 12968
rect 15059 12937 15071 12940
rect 15013 12931 15071 12937
rect 15289 12937 15301 12940
rect 15335 12968 15347 12971
rect 15470 12968 15476 12980
rect 15335 12940 15476 12968
rect 15335 12937 15347 12940
rect 15289 12931 15347 12937
rect 15470 12928 15476 12940
rect 15528 12928 15534 12980
rect 15746 12968 15752 12980
rect 15707 12940 15752 12968
rect 15746 12928 15752 12940
rect 15804 12928 15810 12980
rect 15838 12928 15844 12980
rect 15896 12968 15902 12980
rect 15979 12971 16037 12977
rect 15979 12968 15991 12971
rect 15896 12940 15991 12968
rect 15896 12928 15902 12940
rect 15979 12937 15991 12940
rect 16025 12937 16037 12971
rect 15979 12931 16037 12937
rect 8941 12903 8999 12909
rect 8941 12900 8953 12903
rect 4755 12872 5488 12900
rect 5597 12872 8953 12900
rect 4755 12869 4767 12872
rect 4709 12863 4767 12869
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12832 2559 12835
rect 2590 12832 2596 12844
rect 2547 12804 2596 12832
rect 2547 12801 2559 12804
rect 2501 12795 2559 12801
rect 2590 12792 2596 12804
rect 2648 12832 2654 12844
rect 2777 12835 2835 12841
rect 2777 12832 2789 12835
rect 2648 12804 2789 12832
rect 2648 12792 2654 12804
rect 2777 12801 2789 12804
rect 2823 12801 2835 12835
rect 4982 12832 4988 12844
rect 2777 12795 2835 12801
rect 2884 12804 4988 12832
rect 1673 12767 1731 12773
rect 1673 12733 1685 12767
rect 1719 12764 1731 12767
rect 2409 12767 2467 12773
rect 2409 12764 2421 12767
rect 1719 12736 2421 12764
rect 1719 12733 1731 12736
rect 1673 12727 1731 12733
rect 2409 12733 2421 12736
rect 2455 12764 2467 12767
rect 2884 12764 2912 12804
rect 4982 12792 4988 12804
rect 5040 12792 5046 12844
rect 3326 12764 3332 12776
rect 2455 12736 2912 12764
rect 3287 12736 3332 12764
rect 2455 12733 2467 12736
rect 2409 12727 2467 12733
rect 3326 12724 3332 12736
rect 3384 12724 3390 12776
rect 5353 12767 5411 12773
rect 5353 12733 5365 12767
rect 5399 12733 5411 12767
rect 5460 12764 5488 12872
rect 8941 12869 8953 12872
rect 8987 12900 8999 12903
rect 9490 12900 9496 12912
rect 8987 12872 9496 12900
rect 8987 12869 8999 12872
rect 8941 12863 8999 12869
rect 9490 12860 9496 12872
rect 9548 12860 9554 12912
rect 11698 12860 11704 12912
rect 11756 12900 11762 12912
rect 11793 12903 11851 12909
rect 11793 12900 11805 12903
rect 11756 12872 11805 12900
rect 11756 12860 11762 12872
rect 11793 12869 11805 12872
rect 11839 12900 11851 12903
rect 13909 12903 13967 12909
rect 13909 12900 13921 12903
rect 11839 12872 13921 12900
rect 11839 12869 11851 12872
rect 11793 12863 11851 12869
rect 13909 12869 13921 12872
rect 13955 12869 13967 12903
rect 13909 12863 13967 12869
rect 5534 12792 5540 12844
rect 5592 12832 5598 12844
rect 5721 12835 5779 12841
rect 5721 12832 5733 12835
rect 5592 12804 5733 12832
rect 5592 12792 5598 12804
rect 5721 12801 5733 12804
rect 5767 12801 5779 12835
rect 5721 12795 5779 12801
rect 6641 12835 6699 12841
rect 6641 12801 6653 12835
rect 6687 12832 6699 12835
rect 7650 12832 7656 12844
rect 6687 12804 7656 12832
rect 6687 12801 6699 12804
rect 6641 12795 6699 12801
rect 5629 12767 5687 12773
rect 5629 12764 5641 12767
rect 5460 12736 5641 12764
rect 5353 12727 5411 12733
rect 5629 12733 5641 12736
rect 5675 12764 5687 12767
rect 6362 12764 6368 12776
rect 5675 12736 6368 12764
rect 5675 12733 5687 12736
rect 5629 12727 5687 12733
rect 3237 12699 3295 12705
rect 3237 12665 3249 12699
rect 3283 12696 3295 12699
rect 3650 12699 3708 12705
rect 3650 12696 3662 12699
rect 3283 12668 3662 12696
rect 3283 12665 3295 12668
rect 3237 12659 3295 12665
rect 3650 12665 3662 12668
rect 3696 12696 3708 12699
rect 4430 12696 4436 12708
rect 3696 12668 4436 12696
rect 3696 12665 3708 12668
rect 3650 12659 3708 12665
rect 4430 12656 4436 12668
rect 4488 12656 4494 12708
rect 5368 12696 5396 12727
rect 6362 12724 6368 12736
rect 6420 12724 6426 12776
rect 7116 12773 7144 12804
rect 7650 12792 7656 12804
rect 7708 12832 7714 12844
rect 9585 12835 9643 12841
rect 9585 12832 9597 12835
rect 7708 12804 9597 12832
rect 7708 12792 7714 12804
rect 9585 12801 9597 12804
rect 9631 12832 9643 12835
rect 9674 12832 9680 12844
rect 9631 12804 9680 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 9674 12792 9680 12804
rect 9732 12832 9738 12844
rect 10502 12832 10508 12844
rect 9732 12804 9812 12832
rect 10463 12804 10508 12832
rect 9732 12792 9738 12804
rect 7101 12767 7159 12773
rect 7101 12764 7113 12767
rect 7079 12736 7113 12764
rect 7101 12733 7113 12736
rect 7147 12733 7159 12767
rect 7282 12764 7288 12776
rect 7243 12736 7288 12764
rect 7101 12727 7159 12733
rect 7282 12724 7288 12736
rect 7340 12724 7346 12776
rect 8754 12764 8760 12776
rect 8715 12736 8760 12764
rect 8754 12724 8760 12736
rect 8812 12764 8818 12776
rect 9217 12767 9275 12773
rect 9217 12764 9229 12767
rect 8812 12736 9229 12764
rect 8812 12724 8818 12736
rect 9217 12733 9229 12736
rect 9263 12764 9275 12767
rect 9398 12764 9404 12776
rect 9263 12736 9404 12764
rect 9263 12733 9275 12736
rect 9217 12727 9275 12733
rect 9398 12724 9404 12736
rect 9456 12724 9462 12776
rect 9784 12773 9812 12804
rect 10502 12792 10508 12804
rect 10560 12792 10566 12844
rect 13924 12832 13952 12863
rect 13924 12804 14457 12832
rect 9769 12767 9827 12773
rect 9769 12733 9781 12767
rect 9815 12733 9827 12767
rect 9769 12727 9827 12733
rect 8018 12696 8024 12708
rect 5368 12668 8024 12696
rect 4154 12588 4160 12640
rect 4212 12628 4218 12640
rect 5077 12631 5135 12637
rect 5077 12628 5089 12631
rect 4212 12600 5089 12628
rect 4212 12588 4218 12600
rect 5077 12597 5089 12600
rect 5123 12628 5135 12631
rect 5368 12628 5396 12668
rect 8018 12656 8024 12668
rect 8076 12656 8082 12708
rect 9784 12696 9812 12727
rect 10134 12724 10140 12776
rect 10192 12764 10198 12776
rect 10229 12767 10287 12773
rect 10229 12764 10241 12767
rect 10192 12736 10241 12764
rect 10192 12724 10198 12736
rect 10229 12733 10241 12736
rect 10275 12764 10287 12767
rect 11149 12767 11207 12773
rect 11149 12764 11161 12767
rect 10275 12736 11161 12764
rect 10275 12733 10287 12736
rect 10229 12727 10287 12733
rect 11149 12733 11161 12736
rect 11195 12733 11207 12767
rect 12472 12767 12530 12773
rect 12472 12764 12484 12767
rect 11149 12727 11207 12733
rect 12452 12733 12484 12764
rect 12518 12733 12530 12767
rect 12452 12727 12530 12733
rect 13265 12767 13323 12773
rect 13265 12733 13277 12767
rect 13311 12764 13323 12767
rect 14090 12764 14096 12776
rect 13311 12736 14096 12764
rect 13311 12733 13323 12736
rect 13265 12727 13323 12733
rect 10781 12699 10839 12705
rect 10781 12696 10793 12699
rect 9784 12668 10793 12696
rect 10781 12665 10793 12668
rect 10827 12665 10839 12699
rect 10781 12659 10839 12665
rect 11054 12656 11060 12708
rect 11112 12696 11118 12708
rect 11333 12699 11391 12705
rect 11333 12696 11345 12699
rect 11112 12668 11345 12696
rect 11112 12656 11118 12668
rect 11333 12665 11345 12668
rect 11379 12665 11391 12699
rect 11333 12659 11391 12665
rect 6178 12628 6184 12640
rect 5123 12600 5396 12628
rect 6139 12600 6184 12628
rect 5123 12597 5135 12600
rect 5077 12591 5135 12597
rect 6178 12588 6184 12600
rect 6236 12588 6242 12640
rect 6914 12628 6920 12640
rect 6875 12600 6920 12628
rect 6914 12588 6920 12600
rect 6972 12588 6978 12640
rect 12253 12631 12311 12637
rect 12253 12597 12265 12631
rect 12299 12628 12311 12631
rect 12452 12628 12480 12727
rect 14090 12724 14096 12736
rect 14148 12724 14154 12776
rect 14429 12708 14457 12804
rect 15908 12767 15966 12773
rect 15908 12733 15920 12767
rect 15954 12764 15966 12767
rect 16022 12764 16028 12776
rect 15954 12736 16028 12764
rect 15954 12733 15966 12736
rect 15908 12727 15966 12733
rect 16022 12724 16028 12736
rect 16080 12764 16086 12776
rect 16301 12767 16359 12773
rect 16301 12764 16313 12767
rect 16080 12736 16313 12764
rect 16080 12724 16086 12736
rect 16301 12733 16313 12736
rect 16347 12733 16359 12767
rect 16301 12727 16359 12733
rect 14366 12696 14372 12708
rect 14324 12668 14372 12696
rect 14366 12656 14372 12668
rect 14424 12705 14457 12708
rect 14424 12699 14472 12705
rect 14424 12665 14426 12699
rect 14460 12665 14472 12699
rect 14424 12659 14472 12665
rect 14424 12656 14430 12659
rect 13354 12628 13360 12640
rect 12299 12600 13360 12628
rect 12299 12597 12311 12600
rect 12253 12591 12311 12597
rect 13354 12588 13360 12600
rect 13412 12588 13418 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 2314 12424 2320 12436
rect 2275 12396 2320 12424
rect 2314 12384 2320 12396
rect 2372 12384 2378 12436
rect 4430 12424 4436 12436
rect 4391 12396 4436 12424
rect 4430 12384 4436 12396
rect 4488 12384 4494 12436
rect 4982 12424 4988 12436
rect 4943 12396 4988 12424
rect 4982 12384 4988 12396
rect 5040 12384 5046 12436
rect 5534 12424 5540 12436
rect 5495 12396 5540 12424
rect 5534 12384 5540 12396
rect 5592 12384 5598 12436
rect 8110 12384 8116 12436
rect 8168 12424 8174 12436
rect 9033 12427 9091 12433
rect 9033 12424 9045 12427
rect 8168 12396 9045 12424
rect 8168 12384 8174 12396
rect 9033 12393 9045 12396
rect 9079 12424 9091 12427
rect 9122 12424 9128 12436
rect 9079 12396 9128 12424
rect 9079 12393 9091 12396
rect 9033 12387 9091 12393
rect 9122 12384 9128 12396
rect 9180 12384 9186 12436
rect 11054 12424 11060 12436
rect 11015 12396 11060 12424
rect 11054 12384 11060 12396
rect 11112 12384 11118 12436
rect 24762 12424 24768 12436
rect 24723 12396 24768 12424
rect 24762 12384 24768 12396
rect 24820 12384 24826 12436
rect 2590 12356 2596 12368
rect 2551 12328 2596 12356
rect 2590 12316 2596 12328
rect 2648 12316 2654 12368
rect 3326 12316 3332 12368
rect 3384 12356 3390 12368
rect 3513 12359 3571 12365
rect 3513 12356 3525 12359
rect 3384 12328 3525 12356
rect 3384 12316 3390 12328
rect 3513 12325 3525 12328
rect 3559 12356 3571 12359
rect 4448 12356 4476 12384
rect 6178 12356 6184 12368
rect 3559 12328 3832 12356
rect 4448 12328 6184 12356
rect 3559 12325 3571 12328
rect 3513 12319 3571 12325
rect 3142 12248 3148 12300
rect 3200 12288 3206 12300
rect 3694 12288 3700 12300
rect 3200 12260 3700 12288
rect 3200 12248 3206 12260
rect 3694 12248 3700 12260
rect 3752 12248 3758 12300
rect 3804 12288 3832 12328
rect 6178 12316 6184 12328
rect 6236 12316 6242 12368
rect 6546 12356 6552 12368
rect 6507 12328 6552 12356
rect 6546 12316 6552 12328
rect 6604 12316 6610 12368
rect 10689 12359 10747 12365
rect 10689 12325 10701 12359
rect 10735 12356 10747 12359
rect 11238 12356 11244 12368
rect 10735 12328 11244 12356
rect 10735 12325 10747 12328
rect 10689 12319 10747 12325
rect 11238 12316 11244 12328
rect 11296 12356 11302 12368
rect 11333 12359 11391 12365
rect 11333 12356 11345 12359
rect 11296 12328 11345 12356
rect 11296 12316 11302 12328
rect 11333 12325 11345 12328
rect 11379 12325 11391 12359
rect 11333 12319 11391 12325
rect 5994 12288 6000 12300
rect 3804 12260 5902 12288
rect 5955 12260 6000 12288
rect 2501 12223 2559 12229
rect 2501 12189 2513 12223
rect 2547 12220 2559 12223
rect 2866 12220 2872 12232
rect 2547 12192 2872 12220
rect 2547 12189 2559 12192
rect 2501 12183 2559 12189
rect 2866 12180 2872 12192
rect 2924 12220 2930 12232
rect 2924 12192 3188 12220
rect 2924 12180 2930 12192
rect 3160 12152 3188 12192
rect 3878 12180 3884 12232
rect 3936 12220 3942 12232
rect 4065 12223 4123 12229
rect 4065 12220 4077 12223
rect 3936 12192 4077 12220
rect 3936 12180 3942 12192
rect 4065 12189 4077 12192
rect 4111 12220 4123 12223
rect 5258 12220 5264 12232
rect 4111 12192 5264 12220
rect 4111 12189 4123 12192
rect 4065 12183 4123 12189
rect 5258 12180 5264 12192
rect 5316 12180 5322 12232
rect 5874 12220 5902 12260
rect 5994 12248 6000 12260
rect 6052 12248 6058 12300
rect 6362 12288 6368 12300
rect 6323 12260 6368 12288
rect 6362 12248 6368 12260
rect 6420 12248 6426 12300
rect 8110 12288 8116 12300
rect 8071 12260 8116 12288
rect 8110 12248 8116 12260
rect 8168 12248 8174 12300
rect 8294 12288 8300 12300
rect 8255 12260 8300 12288
rect 8294 12248 8300 12260
rect 8352 12248 8358 12300
rect 9490 12248 9496 12300
rect 9548 12288 9554 12300
rect 9953 12291 10011 12297
rect 9953 12288 9965 12291
rect 9548 12260 9965 12288
rect 9548 12248 9554 12260
rect 9953 12257 9965 12260
rect 9999 12257 10011 12291
rect 9953 12251 10011 12257
rect 10134 12248 10140 12300
rect 10192 12288 10198 12300
rect 10413 12291 10471 12297
rect 10413 12288 10425 12291
rect 10192 12260 10425 12288
rect 10192 12248 10198 12260
rect 10413 12257 10425 12260
rect 10459 12257 10471 12291
rect 11606 12288 11612 12300
rect 11567 12260 11612 12288
rect 10413 12251 10471 12257
rect 11606 12248 11612 12260
rect 11664 12248 11670 12300
rect 14160 12291 14218 12297
rect 14160 12257 14172 12291
rect 14206 12288 14218 12291
rect 14274 12288 14280 12300
rect 14206 12260 14280 12288
rect 14206 12257 14218 12260
rect 14160 12251 14218 12257
rect 14274 12248 14280 12260
rect 14332 12248 14338 12300
rect 15378 12288 15384 12300
rect 15339 12260 15384 12288
rect 15378 12248 15384 12260
rect 15436 12248 15442 12300
rect 24026 12248 24032 12300
rect 24084 12288 24090 12300
rect 24581 12291 24639 12297
rect 24581 12288 24593 12291
rect 24084 12260 24593 12288
rect 24084 12248 24090 12260
rect 24581 12257 24593 12260
rect 24627 12257 24639 12291
rect 24581 12251 24639 12257
rect 6914 12220 6920 12232
rect 5874 12192 6920 12220
rect 6914 12180 6920 12192
rect 6972 12180 6978 12232
rect 8386 12220 8392 12232
rect 8347 12192 8392 12220
rect 8386 12180 8392 12192
rect 8444 12180 8450 12232
rect 8846 12180 8852 12232
rect 8904 12220 8910 12232
rect 11517 12223 11575 12229
rect 11517 12220 11529 12223
rect 8904 12192 11529 12220
rect 8904 12180 8910 12192
rect 11517 12189 11529 12192
rect 11563 12189 11575 12223
rect 13078 12220 13084 12232
rect 13039 12192 13084 12220
rect 11517 12183 11575 12189
rect 13078 12180 13084 12192
rect 13136 12180 13142 12232
rect 4890 12152 4896 12164
rect 3160 12124 4896 12152
rect 4890 12112 4896 12124
rect 4948 12112 4954 12164
rect 7098 12112 7104 12164
rect 7156 12152 7162 12164
rect 9030 12152 9036 12164
rect 7156 12124 9036 12152
rect 7156 12112 7162 12124
rect 9030 12112 9036 12124
rect 9088 12152 9094 12164
rect 9401 12155 9459 12161
rect 9401 12152 9413 12155
rect 9088 12124 9413 12152
rect 9088 12112 9094 12124
rect 9401 12121 9413 12124
rect 9447 12121 9459 12155
rect 9401 12115 9459 12121
rect 1670 12084 1676 12096
rect 1631 12056 1676 12084
rect 1670 12044 1676 12056
rect 1728 12044 1734 12096
rect 3881 12087 3939 12093
rect 3881 12053 3893 12087
rect 3927 12084 3939 12087
rect 4614 12084 4620 12096
rect 3927 12056 4620 12084
rect 3927 12053 3939 12056
rect 3881 12047 3939 12053
rect 4614 12044 4620 12056
rect 4672 12044 4678 12096
rect 6917 12087 6975 12093
rect 6917 12053 6929 12087
rect 6963 12084 6975 12087
rect 7282 12084 7288 12096
rect 6963 12056 7288 12084
rect 6963 12053 6975 12056
rect 6917 12047 6975 12053
rect 7282 12044 7288 12056
rect 7340 12084 7346 12096
rect 7926 12084 7932 12096
rect 7340 12056 7932 12084
rect 7340 12044 7346 12056
rect 7926 12044 7932 12056
rect 7984 12044 7990 12096
rect 14231 12087 14289 12093
rect 14231 12053 14243 12087
rect 14277 12084 14289 12087
rect 15286 12084 15292 12096
rect 14277 12056 15292 12084
rect 14277 12053 14289 12056
rect 14231 12047 14289 12053
rect 15286 12044 15292 12056
rect 15344 12044 15350 12096
rect 15562 12084 15568 12096
rect 15523 12056 15568 12084
rect 15562 12044 15568 12056
rect 15620 12044 15626 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2869 11883 2927 11889
rect 2869 11849 2881 11883
rect 2915 11880 2927 11883
rect 2958 11880 2964 11892
rect 2915 11852 2964 11880
rect 2915 11849 2927 11852
rect 2869 11843 2927 11849
rect 2958 11840 2964 11852
rect 3016 11840 3022 11892
rect 8110 11840 8116 11892
rect 8168 11880 8174 11892
rect 8665 11883 8723 11889
rect 8665 11880 8677 11883
rect 8168 11852 8677 11880
rect 8168 11840 8174 11852
rect 8665 11849 8677 11852
rect 8711 11849 8723 11883
rect 8665 11843 8723 11849
rect 9214 11840 9220 11892
rect 9272 11880 9278 11892
rect 11606 11880 11612 11892
rect 9272 11852 11612 11880
rect 9272 11840 9278 11852
rect 11606 11840 11612 11852
rect 11664 11840 11670 11892
rect 14185 11883 14243 11889
rect 14185 11849 14197 11883
rect 14231 11880 14243 11883
rect 14274 11880 14280 11892
rect 14231 11852 14280 11880
rect 14231 11849 14243 11852
rect 14185 11843 14243 11849
rect 14274 11840 14280 11852
rect 14332 11840 14338 11892
rect 15378 11880 15384 11892
rect 15339 11852 15384 11880
rect 15378 11840 15384 11852
rect 15436 11840 15442 11892
rect 1670 11772 1676 11824
rect 1728 11812 1734 11824
rect 4154 11812 4160 11824
rect 1728 11784 4160 11812
rect 1728 11772 1734 11784
rect 1673 11679 1731 11685
rect 1673 11645 1685 11679
rect 1719 11676 1731 11679
rect 1780 11676 1808 11784
rect 4154 11772 4160 11784
rect 4212 11772 4218 11824
rect 10962 11772 10968 11824
rect 11020 11812 11026 11824
rect 11241 11815 11299 11821
rect 11241 11812 11253 11815
rect 11020 11784 11253 11812
rect 11020 11772 11026 11784
rect 11241 11781 11253 11784
rect 11287 11781 11299 11815
rect 16485 11815 16543 11821
rect 16485 11812 16497 11815
rect 11241 11775 11299 11781
rect 15717 11784 16497 11812
rect 2501 11747 2559 11753
rect 2501 11713 2513 11747
rect 2547 11744 2559 11747
rect 3053 11747 3111 11753
rect 3053 11744 3065 11747
rect 2547 11716 3065 11744
rect 2547 11713 2559 11716
rect 2501 11707 2559 11713
rect 3053 11713 3065 11716
rect 3099 11744 3111 11747
rect 4062 11744 4068 11756
rect 3099 11716 4068 11744
rect 3099 11713 3111 11716
rect 3053 11707 3111 11713
rect 4062 11704 4068 11716
rect 4120 11704 4126 11756
rect 4890 11744 4896 11756
rect 4851 11716 4896 11744
rect 4890 11704 4896 11716
rect 4948 11704 4954 11756
rect 5534 11704 5540 11756
rect 5592 11744 5598 11756
rect 5905 11747 5963 11753
rect 5905 11744 5917 11747
rect 5592 11716 5917 11744
rect 5592 11704 5598 11716
rect 5905 11713 5917 11716
rect 5951 11744 5963 11747
rect 5994 11744 6000 11756
rect 5951 11716 6000 11744
rect 5951 11713 5963 11716
rect 5905 11707 5963 11713
rect 5994 11704 6000 11716
rect 6052 11744 6058 11756
rect 7466 11744 7472 11756
rect 6052 11716 7472 11744
rect 6052 11704 6058 11716
rect 7466 11704 7472 11716
rect 7524 11704 7530 11756
rect 7742 11744 7748 11756
rect 7703 11716 7748 11744
rect 7742 11704 7748 11716
rect 7800 11704 7806 11756
rect 9122 11744 9128 11756
rect 9083 11716 9128 11744
rect 9122 11704 9128 11716
rect 9180 11704 9186 11756
rect 10505 11747 10563 11753
rect 10505 11713 10517 11747
rect 10551 11744 10563 11747
rect 10778 11744 10784 11756
rect 10551 11716 10784 11744
rect 10551 11713 10563 11716
rect 10505 11707 10563 11713
rect 10778 11704 10784 11716
rect 10836 11744 10842 11756
rect 12437 11747 12495 11753
rect 12437 11744 12449 11747
rect 10836 11716 12449 11744
rect 10836 11704 10842 11716
rect 12437 11713 12449 11716
rect 12483 11713 12495 11747
rect 12437 11707 12495 11713
rect 15565 11747 15623 11753
rect 15565 11713 15577 11747
rect 15611 11744 15623 11747
rect 15717 11744 15745 11784
rect 16485 11781 16497 11784
rect 16531 11812 16543 11815
rect 17218 11812 17224 11824
rect 16531 11784 17224 11812
rect 16531 11781 16543 11784
rect 16485 11775 16543 11781
rect 17218 11772 17224 11784
rect 17276 11772 17282 11824
rect 16022 11744 16028 11756
rect 15611 11716 15745 11744
rect 15983 11716 16028 11744
rect 15611 11713 15623 11716
rect 15565 11707 15623 11713
rect 16022 11704 16028 11716
rect 16080 11704 16086 11756
rect 1946 11676 1952 11688
rect 1719 11648 1808 11676
rect 1907 11648 1952 11676
rect 1719 11645 1731 11648
rect 1673 11639 1731 11645
rect 1946 11636 1952 11648
rect 2004 11636 2010 11688
rect 3694 11636 3700 11688
rect 3752 11676 3758 11688
rect 3752 11648 3797 11676
rect 3752 11636 3758 11648
rect 11330 11636 11336 11688
rect 11388 11676 11394 11688
rect 12253 11679 12311 11685
rect 12253 11676 12265 11679
rect 11388 11648 12265 11676
rect 11388 11636 11394 11648
rect 12253 11645 12265 11648
rect 12299 11676 12311 11679
rect 12529 11679 12587 11685
rect 12529 11676 12541 11679
rect 12299 11648 12541 11676
rect 12299 11645 12311 11648
rect 12253 11639 12311 11645
rect 12529 11645 12541 11648
rect 12575 11645 12587 11679
rect 12529 11639 12587 11645
rect 23728 11679 23786 11685
rect 23728 11645 23740 11679
rect 23774 11676 23786 11679
rect 23774 11648 23980 11676
rect 23774 11645 23786 11648
rect 23728 11639 23786 11645
rect 2130 11608 2136 11620
rect 2091 11580 2136 11608
rect 2130 11568 2136 11580
rect 2188 11568 2194 11620
rect 3145 11611 3203 11617
rect 3145 11577 3157 11611
rect 3191 11577 3203 11611
rect 4614 11608 4620 11620
rect 4575 11580 4620 11608
rect 3145 11571 3203 11577
rect 2958 11500 2964 11552
rect 3016 11540 3022 11552
rect 3160 11540 3188 11571
rect 4614 11568 4620 11580
rect 4672 11568 4678 11620
rect 4709 11611 4767 11617
rect 4709 11577 4721 11611
rect 4755 11608 4767 11611
rect 4982 11608 4988 11620
rect 4755 11580 4988 11608
rect 4755 11577 4767 11580
rect 4709 11571 4767 11577
rect 4982 11568 4988 11580
rect 5040 11568 5046 11620
rect 7374 11608 7380 11620
rect 7335 11580 7380 11608
rect 7374 11568 7380 11580
rect 7432 11568 7438 11620
rect 7469 11611 7527 11617
rect 7469 11577 7481 11611
rect 7515 11608 7527 11611
rect 8018 11608 8024 11620
rect 7515 11580 8024 11608
rect 7515 11577 7527 11580
rect 7469 11571 7527 11577
rect 3016 11512 3188 11540
rect 4157 11543 4215 11549
rect 3016 11500 3022 11512
rect 4157 11509 4169 11543
rect 4203 11540 4215 11543
rect 4430 11540 4436 11552
rect 4203 11512 4436 11540
rect 4203 11509 4215 11512
rect 4157 11503 4215 11509
rect 4430 11500 4436 11512
rect 4488 11500 4494 11552
rect 6273 11543 6331 11549
rect 6273 11509 6285 11543
rect 6319 11540 6331 11543
rect 6362 11540 6368 11552
rect 6319 11512 6368 11540
rect 6319 11509 6331 11512
rect 6273 11503 6331 11509
rect 6362 11500 6368 11512
rect 6420 11500 6426 11552
rect 7193 11543 7251 11549
rect 7193 11509 7205 11543
rect 7239 11540 7251 11543
rect 7484 11540 7512 11571
rect 8018 11568 8024 11580
rect 8076 11568 8082 11620
rect 9214 11608 9220 11620
rect 9175 11580 9220 11608
rect 9214 11568 9220 11580
rect 9272 11568 9278 11620
rect 9766 11608 9772 11620
rect 9727 11580 9772 11608
rect 9766 11568 9772 11580
rect 9824 11568 9830 11620
rect 10689 11611 10747 11617
rect 10689 11577 10701 11611
rect 10735 11577 10747 11611
rect 10689 11571 10747 11577
rect 8294 11540 8300 11552
rect 7239 11512 7512 11540
rect 8255 11512 8300 11540
rect 7239 11509 7251 11512
rect 7193 11503 7251 11509
rect 8294 11500 8300 11512
rect 8352 11500 8358 11552
rect 10134 11540 10140 11552
rect 10095 11512 10140 11540
rect 10134 11500 10140 11512
rect 10192 11500 10198 11552
rect 10704 11540 10732 11571
rect 10778 11568 10784 11620
rect 10836 11608 10842 11620
rect 15657 11611 15715 11617
rect 10836 11580 10881 11608
rect 10836 11568 10842 11580
rect 15657 11577 15669 11611
rect 15703 11577 15715 11611
rect 15657 11571 15715 11577
rect 11054 11540 11060 11552
rect 10704 11512 11060 11540
rect 11054 11500 11060 11512
rect 11112 11500 11118 11552
rect 13170 11500 13176 11552
rect 13228 11540 13234 11552
rect 14274 11540 14280 11552
rect 13228 11512 14280 11540
rect 13228 11500 13234 11512
rect 14274 11500 14280 11512
rect 14332 11500 14338 11552
rect 14458 11540 14464 11552
rect 14419 11512 14464 11540
rect 14458 11500 14464 11512
rect 14516 11500 14522 11552
rect 15013 11543 15071 11549
rect 15013 11509 15025 11543
rect 15059 11540 15071 11543
rect 15378 11540 15384 11552
rect 15059 11512 15384 11540
rect 15059 11509 15071 11512
rect 15013 11503 15071 11509
rect 15378 11500 15384 11512
rect 15436 11540 15442 11552
rect 15672 11540 15700 11571
rect 15436 11512 15700 11540
rect 15436 11500 15442 11512
rect 18598 11500 18604 11552
rect 18656 11540 18662 11552
rect 23799 11543 23857 11549
rect 23799 11540 23811 11543
rect 18656 11512 23811 11540
rect 18656 11500 18662 11512
rect 23799 11509 23811 11512
rect 23845 11509 23857 11543
rect 23952 11540 23980 11648
rect 24026 11568 24032 11620
rect 24084 11608 24090 11620
rect 24581 11611 24639 11617
rect 24581 11608 24593 11611
rect 24084 11580 24593 11608
rect 24084 11568 24090 11580
rect 24581 11577 24593 11580
rect 24627 11577 24639 11611
rect 24581 11571 24639 11577
rect 24213 11543 24271 11549
rect 24213 11540 24225 11543
rect 23952 11512 24225 11540
rect 23799 11503 23857 11509
rect 24213 11509 24225 11512
rect 24259 11540 24271 11543
rect 24762 11540 24768 11552
rect 24259 11512 24768 11540
rect 24259 11509 24271 11512
rect 24213 11503 24271 11509
rect 24762 11500 24768 11512
rect 24820 11500 24826 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 2317 11339 2375 11345
rect 2317 11305 2329 11339
rect 2363 11336 2375 11339
rect 2590 11336 2596 11348
rect 2363 11308 2596 11336
rect 2363 11305 2375 11308
rect 2317 11299 2375 11305
rect 2590 11296 2596 11308
rect 2648 11296 2654 11348
rect 3878 11336 3884 11348
rect 3839 11308 3884 11336
rect 3878 11296 3884 11308
rect 3936 11296 3942 11348
rect 4982 11296 4988 11348
rect 5040 11336 5046 11348
rect 5353 11339 5411 11345
rect 5353 11336 5365 11339
rect 5040 11308 5365 11336
rect 5040 11296 5046 11308
rect 5353 11305 5365 11308
rect 5399 11305 5411 11339
rect 7374 11336 7380 11348
rect 7335 11308 7380 11336
rect 5353 11299 5411 11305
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 9125 11339 9183 11345
rect 9125 11305 9137 11339
rect 9171 11336 9183 11339
rect 9214 11336 9220 11348
rect 9171 11308 9220 11336
rect 9171 11305 9183 11308
rect 9125 11299 9183 11305
rect 9214 11296 9220 11308
rect 9272 11296 9278 11348
rect 9490 11296 9496 11348
rect 9548 11336 9554 11348
rect 9953 11339 10011 11345
rect 9953 11336 9965 11339
rect 9548 11308 9965 11336
rect 9548 11296 9554 11308
rect 9953 11305 9965 11308
rect 9999 11305 10011 11339
rect 11330 11336 11336 11348
rect 9953 11299 10011 11305
rect 10428 11308 11336 11336
rect 5077 11271 5135 11277
rect 5077 11237 5089 11271
rect 5123 11268 5135 11271
rect 5994 11268 6000 11280
rect 5123 11240 6000 11268
rect 5123 11237 5135 11240
rect 5077 11231 5135 11237
rect 5994 11228 6000 11240
rect 6052 11268 6058 11280
rect 6089 11271 6147 11277
rect 6089 11268 6101 11271
rect 6052 11240 6101 11268
rect 6052 11228 6058 11240
rect 6089 11237 6101 11240
rect 6135 11237 6147 11271
rect 6089 11231 6147 11237
rect 7834 11228 7840 11280
rect 7892 11268 7898 11280
rect 8205 11271 8263 11277
rect 8205 11268 8217 11271
rect 7892 11240 8217 11268
rect 7892 11228 7898 11240
rect 8205 11237 8217 11240
rect 8251 11268 8263 11271
rect 8846 11268 8852 11280
rect 8251 11240 8852 11268
rect 8251 11237 8263 11240
rect 8205 11231 8263 11237
rect 8846 11228 8852 11240
rect 8904 11228 8910 11280
rect 10428 11277 10456 11308
rect 11330 11296 11336 11308
rect 11388 11296 11394 11348
rect 22738 11336 22744 11348
rect 16960 11308 22744 11336
rect 16960 11280 16988 11308
rect 22738 11296 22744 11308
rect 22796 11296 22802 11348
rect 10413 11271 10471 11277
rect 10413 11237 10425 11271
rect 10459 11237 10471 11271
rect 10962 11268 10968 11280
rect 10923 11240 10968 11268
rect 10413 11231 10471 11237
rect 10962 11228 10968 11240
rect 11020 11228 11026 11280
rect 14458 11228 14464 11280
rect 14516 11268 14522 11280
rect 15381 11271 15439 11277
rect 15381 11268 15393 11271
rect 14516 11240 15393 11268
rect 14516 11228 14522 11240
rect 15381 11237 15393 11240
rect 15427 11237 15439 11271
rect 15381 11231 15439 11237
rect 15473 11271 15531 11277
rect 15473 11237 15485 11271
rect 15519 11268 15531 11271
rect 15562 11268 15568 11280
rect 15519 11240 15568 11268
rect 15519 11237 15531 11240
rect 15473 11231 15531 11237
rect 15562 11228 15568 11240
rect 15620 11228 15626 11280
rect 16022 11268 16028 11280
rect 15983 11240 16028 11268
rect 16022 11228 16028 11240
rect 16080 11228 16086 11280
rect 16942 11268 16948 11280
rect 16855 11240 16948 11268
rect 16942 11228 16948 11240
rect 17000 11228 17006 11280
rect 17037 11271 17095 11277
rect 17037 11237 17049 11271
rect 17083 11268 17095 11271
rect 17402 11268 17408 11280
rect 17083 11240 17408 11268
rect 17083 11237 17095 11240
rect 17037 11231 17095 11237
rect 17402 11228 17408 11240
rect 17460 11228 17466 11280
rect 1464 11203 1522 11209
rect 1464 11169 1476 11203
rect 1510 11200 1522 11203
rect 1762 11200 1768 11212
rect 1510 11172 1768 11200
rect 1510 11169 1522 11172
rect 1464 11163 1522 11169
rect 1762 11160 1768 11172
rect 1820 11160 1826 11212
rect 2682 11200 2688 11212
rect 2643 11172 2688 11200
rect 2682 11160 2688 11172
rect 2740 11160 2746 11212
rect 2866 11200 2872 11212
rect 2827 11172 2872 11200
rect 2866 11160 2872 11172
rect 2924 11160 2930 11212
rect 4522 11200 4528 11212
rect 4483 11172 4528 11200
rect 4522 11160 4528 11172
rect 4580 11160 4586 11212
rect 11882 11200 11888 11212
rect 11843 11172 11888 11200
rect 11882 11160 11888 11172
rect 11940 11160 11946 11212
rect 13630 11200 13636 11212
rect 13591 11172 13636 11200
rect 13630 11160 13636 11172
rect 13688 11160 13694 11212
rect 1946 11132 1952 11144
rect 1859 11104 1952 11132
rect 1946 11092 1952 11104
rect 2004 11132 2010 11144
rect 2884 11132 2912 11160
rect 2004 11104 2912 11132
rect 3145 11135 3203 11141
rect 2004 11092 2010 11104
rect 3145 11101 3157 11135
rect 3191 11132 3203 11135
rect 3602 11132 3608 11144
rect 3191 11104 3608 11132
rect 3191 11101 3203 11104
rect 3145 11095 3203 11101
rect 3602 11092 3608 11104
rect 3660 11092 3666 11144
rect 5997 11135 6055 11141
rect 5997 11101 6009 11135
rect 6043 11132 6055 11135
rect 6086 11132 6092 11144
rect 6043 11104 6092 11132
rect 6043 11101 6055 11104
rect 5997 11095 6055 11101
rect 6086 11092 6092 11104
rect 6144 11092 6150 11144
rect 6270 11132 6276 11144
rect 6231 11104 6276 11132
rect 6270 11092 6276 11104
rect 6328 11092 6334 11144
rect 8113 11135 8171 11141
rect 8113 11132 8125 11135
rect 7852 11104 8125 11132
rect 1535 11067 1593 11073
rect 1535 11033 1547 11067
rect 1581 11064 1593 11067
rect 3234 11064 3240 11076
rect 1581 11036 3240 11064
rect 1581 11033 1593 11036
rect 1535 11027 1593 11033
rect 3234 11024 3240 11036
rect 3292 11024 3298 11076
rect 2406 10956 2412 11008
rect 2464 10996 2470 11008
rect 3421 10999 3479 11005
rect 3421 10996 3433 10999
rect 2464 10968 3433 10996
rect 2464 10956 2470 10968
rect 3421 10965 3433 10968
rect 3467 10965 3479 10999
rect 3421 10959 3479 10965
rect 5166 10956 5172 11008
rect 5224 10996 5230 11008
rect 7852 11005 7880 11104
rect 8113 11101 8125 11104
rect 8159 11101 8171 11135
rect 8113 11095 8171 11101
rect 8757 11135 8815 11141
rect 8757 11101 8769 11135
rect 8803 11132 8815 11135
rect 9766 11132 9772 11144
rect 8803 11104 9772 11132
rect 8803 11101 8815 11104
rect 8757 11095 8815 11101
rect 9766 11092 9772 11104
rect 9824 11132 9830 11144
rect 10318 11132 10324 11144
rect 9824 11104 10324 11132
rect 9824 11092 9830 11104
rect 10318 11092 10324 11104
rect 10376 11092 10382 11144
rect 12529 11135 12587 11141
rect 12529 11101 12541 11135
rect 12575 11132 12587 11135
rect 12618 11132 12624 11144
rect 12575 11104 12624 11132
rect 12575 11101 12587 11104
rect 12529 11095 12587 11101
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 12802 11092 12808 11144
rect 12860 11132 12866 11144
rect 13357 11135 13415 11141
rect 13357 11132 13369 11135
rect 12860 11104 13369 11132
rect 12860 11092 12866 11104
rect 13357 11101 13369 11104
rect 13403 11101 13415 11135
rect 17218 11132 17224 11144
rect 17179 11104 17224 11132
rect 13357 11095 13415 11101
rect 17218 11092 17224 11104
rect 17276 11092 17282 11144
rect 7837 10999 7895 11005
rect 7837 10996 7849 10999
rect 5224 10968 7849 10996
rect 5224 10956 5230 10968
rect 7837 10965 7849 10968
rect 7883 10965 7895 10999
rect 16482 10996 16488 11008
rect 16443 10968 16488 10996
rect 7837 10959 7895 10965
rect 16482 10956 16488 10968
rect 16540 10956 16546 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 2682 10792 2688 10804
rect 2643 10764 2688 10792
rect 2682 10752 2688 10764
rect 2740 10792 2746 10804
rect 3694 10792 3700 10804
rect 2740 10764 3700 10792
rect 2740 10752 2746 10764
rect 3694 10752 3700 10764
rect 3752 10792 3758 10804
rect 4522 10792 4528 10804
rect 3752 10764 4154 10792
rect 4483 10764 4528 10792
rect 3752 10752 3758 10764
rect 4126 10724 4154 10764
rect 4522 10752 4528 10764
rect 4580 10752 4586 10804
rect 5994 10792 6000 10804
rect 5955 10764 6000 10792
rect 5994 10752 6000 10764
rect 6052 10752 6058 10804
rect 7834 10792 7840 10804
rect 7795 10764 7840 10792
rect 7834 10752 7840 10764
rect 7892 10752 7898 10804
rect 9214 10792 9220 10804
rect 9175 10764 9220 10792
rect 9214 10752 9220 10764
rect 9272 10752 9278 10804
rect 10318 10752 10324 10804
rect 10376 10792 10382 10804
rect 11241 10795 11299 10801
rect 11241 10792 11253 10795
rect 10376 10764 11253 10792
rect 10376 10752 10382 10764
rect 11241 10761 11253 10764
rect 11287 10761 11299 10795
rect 11882 10792 11888 10804
rect 11843 10764 11888 10792
rect 11241 10755 11299 10761
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 13630 10792 13636 10804
rect 13591 10764 13636 10792
rect 13630 10752 13636 10764
rect 13688 10752 13694 10804
rect 14366 10792 14372 10804
rect 14327 10764 14372 10792
rect 14366 10752 14372 10764
rect 14424 10752 14430 10804
rect 15378 10792 15384 10804
rect 15339 10764 15384 10792
rect 15378 10752 15384 10764
rect 15436 10752 15442 10804
rect 15562 10752 15568 10804
rect 15620 10792 15626 10804
rect 15657 10795 15715 10801
rect 15657 10792 15669 10795
rect 15620 10764 15669 10792
rect 15620 10752 15626 10764
rect 15657 10761 15669 10764
rect 15703 10761 15715 10795
rect 15657 10755 15715 10761
rect 24765 10795 24823 10801
rect 24765 10761 24777 10795
rect 24811 10792 24823 10795
rect 25222 10792 25228 10804
rect 24811 10764 25228 10792
rect 24811 10761 24823 10764
rect 24765 10755 24823 10761
rect 25222 10752 25228 10764
rect 25280 10752 25286 10804
rect 5534 10724 5540 10736
rect 4126 10696 5540 10724
rect 5534 10684 5540 10696
rect 5592 10684 5598 10736
rect 9585 10727 9643 10733
rect 9585 10693 9597 10727
rect 9631 10724 9643 10727
rect 10965 10727 11023 10733
rect 10965 10724 10977 10727
rect 9631 10696 10977 10724
rect 9631 10693 9643 10696
rect 9585 10687 9643 10693
rect 10965 10693 10977 10696
rect 11011 10724 11023 10727
rect 11330 10724 11336 10736
rect 11011 10696 11336 10724
rect 11011 10693 11023 10696
rect 10965 10687 11023 10693
rect 11330 10684 11336 10696
rect 11388 10684 11394 10736
rect 1670 10656 1676 10668
rect 1583 10628 1676 10656
rect 1670 10616 1676 10628
rect 1728 10656 1734 10668
rect 3329 10659 3387 10665
rect 3329 10656 3341 10659
rect 1728 10628 3341 10656
rect 1728 10616 1734 10628
rect 3329 10625 3341 10628
rect 3375 10625 3387 10659
rect 3329 10619 3387 10625
rect 3605 10659 3663 10665
rect 3605 10625 3617 10659
rect 3651 10656 3663 10659
rect 6086 10656 6092 10668
rect 3651 10628 6092 10656
rect 3651 10625 3663 10628
rect 3605 10619 3663 10625
rect 6086 10616 6092 10628
rect 6144 10656 6150 10668
rect 6273 10659 6331 10665
rect 6273 10656 6285 10659
rect 6144 10628 6285 10656
rect 6144 10616 6150 10628
rect 6273 10625 6285 10628
rect 6319 10625 6331 10659
rect 6273 10619 6331 10625
rect 7101 10659 7159 10665
rect 7101 10625 7113 10659
rect 7147 10656 7159 10659
rect 7374 10656 7380 10668
rect 7147 10628 7380 10656
rect 7147 10625 7159 10628
rect 7101 10619 7159 10625
rect 7374 10616 7380 10628
rect 7432 10616 7438 10668
rect 8297 10659 8355 10665
rect 8297 10625 8309 10659
rect 8343 10656 8355 10659
rect 8386 10656 8392 10668
rect 8343 10628 8392 10656
rect 8343 10625 8355 10628
rect 8297 10619 8355 10625
rect 8386 10616 8392 10628
rect 8444 10616 8450 10668
rect 12710 10656 12716 10668
rect 12623 10628 12716 10656
rect 12710 10616 12716 10628
rect 12768 10656 12774 10668
rect 13078 10656 13084 10668
rect 12768 10628 13084 10656
rect 12768 10616 12774 10628
rect 13078 10616 13084 10628
rect 13136 10616 13142 10668
rect 14461 10659 14519 10665
rect 14461 10625 14473 10659
rect 14507 10656 14519 10659
rect 14734 10656 14740 10668
rect 14507 10628 14740 10656
rect 14507 10625 14519 10628
rect 14461 10619 14519 10625
rect 14734 10616 14740 10628
rect 14792 10616 14798 10668
rect 16482 10656 16488 10668
rect 16443 10628 16488 10656
rect 16482 10616 16488 10628
rect 16540 10616 16546 10668
rect 17129 10659 17187 10665
rect 17129 10625 17141 10659
rect 17175 10656 17187 10659
rect 17218 10656 17224 10668
rect 17175 10628 17224 10656
rect 17175 10625 17187 10628
rect 17129 10619 17187 10625
rect 17218 10616 17224 10628
rect 17276 10616 17282 10668
rect 10042 10588 10048 10600
rect 10003 10560 10048 10588
rect 10042 10548 10048 10560
rect 10100 10548 10106 10600
rect 18141 10591 18199 10597
rect 18141 10557 18153 10591
rect 18187 10557 18199 10591
rect 18141 10551 18199 10557
rect 1765 10523 1823 10529
rect 1765 10489 1777 10523
rect 1811 10489 1823 10523
rect 1765 10483 1823 10489
rect 2317 10523 2375 10529
rect 2317 10489 2329 10523
rect 2363 10520 2375 10523
rect 2406 10520 2412 10532
rect 2363 10492 2412 10520
rect 2363 10489 2375 10492
rect 2317 10483 2375 10489
rect 1780 10452 1808 10483
rect 2406 10480 2412 10492
rect 2464 10480 2470 10532
rect 4706 10520 4712 10532
rect 4667 10492 4712 10520
rect 4706 10480 4712 10492
rect 4764 10480 4770 10532
rect 4801 10523 4859 10529
rect 4801 10489 4813 10523
rect 4847 10489 4859 10523
rect 4801 10483 4859 10489
rect 5353 10523 5411 10529
rect 5353 10489 5365 10523
rect 5399 10520 5411 10523
rect 6270 10520 6276 10532
rect 5399 10492 6276 10520
rect 5399 10489 5411 10492
rect 5353 10483 5411 10489
rect 2222 10452 2228 10464
rect 1780 10424 2228 10452
rect 2222 10412 2228 10424
rect 2280 10412 2286 10464
rect 2866 10412 2872 10464
rect 2924 10452 2930 10464
rect 2961 10455 3019 10461
rect 2961 10452 2973 10455
rect 2924 10424 2973 10452
rect 2924 10412 2930 10424
rect 2961 10421 2973 10424
rect 3007 10421 3019 10455
rect 2961 10415 3019 10421
rect 4157 10455 4215 10461
rect 4157 10421 4169 10455
rect 4203 10452 4215 10455
rect 4522 10452 4528 10464
rect 4203 10424 4528 10452
rect 4203 10421 4215 10424
rect 4157 10415 4215 10421
rect 4522 10412 4528 10424
rect 4580 10452 4586 10464
rect 4816 10452 4844 10483
rect 6270 10480 6276 10492
rect 6328 10480 6334 10532
rect 8202 10520 8208 10532
rect 8115 10492 8208 10520
rect 8202 10480 8208 10492
rect 8260 10520 8266 10532
rect 8659 10523 8717 10529
rect 8659 10520 8671 10523
rect 8260 10492 8671 10520
rect 8260 10480 8266 10492
rect 8659 10489 8671 10492
rect 8705 10520 8717 10523
rect 10366 10523 10424 10529
rect 10366 10520 10378 10523
rect 8705 10492 10378 10520
rect 8705 10489 8717 10492
rect 8659 10483 8717 10489
rect 4580 10424 4844 10452
rect 4580 10412 4586 10424
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 9876 10461 9904 10492
rect 10366 10489 10378 10492
rect 10412 10489 10424 10523
rect 10366 10483 10424 10489
rect 12802 10480 12808 10532
rect 12860 10520 12866 10532
rect 13354 10520 13360 10532
rect 12860 10492 12905 10520
rect 13315 10492 13360 10520
rect 12860 10480 12866 10492
rect 13354 10480 13360 10492
rect 13412 10480 13418 10532
rect 14366 10480 14372 10532
rect 14424 10520 14430 10532
rect 14782 10523 14840 10529
rect 14782 10520 14794 10523
rect 14424 10492 14794 10520
rect 14424 10480 14430 10492
rect 14782 10489 14794 10492
rect 14828 10520 14840 10523
rect 15654 10520 15660 10532
rect 14828 10492 15660 10520
rect 14828 10489 14840 10492
rect 14782 10483 14840 10489
rect 15654 10480 15660 10492
rect 15712 10480 15718 10532
rect 16577 10523 16635 10529
rect 16577 10489 16589 10523
rect 16623 10489 16635 10523
rect 18049 10523 18107 10529
rect 18049 10520 18061 10523
rect 16577 10483 16635 10489
rect 17236 10492 18061 10520
rect 9861 10455 9919 10461
rect 9861 10452 9873 10455
rect 9824 10424 9873 10452
rect 9824 10412 9830 10424
rect 9861 10421 9873 10424
rect 9907 10421 9919 10455
rect 9861 10415 9919 10421
rect 12253 10455 12311 10461
rect 12253 10421 12265 10455
rect 12299 10452 12311 10455
rect 12820 10452 12848 10480
rect 12299 10424 12848 10452
rect 16301 10455 16359 10461
rect 12299 10421 12311 10424
rect 12253 10415 12311 10421
rect 16301 10421 16313 10455
rect 16347 10452 16359 10455
rect 16592 10452 16620 10483
rect 17236 10452 17264 10492
rect 18049 10489 18061 10492
rect 18095 10489 18107 10523
rect 18049 10483 18107 10489
rect 17402 10452 17408 10464
rect 16347 10424 17264 10452
rect 17363 10424 17408 10452
rect 16347 10421 16359 10424
rect 16301 10415 16359 10421
rect 17402 10412 17408 10424
rect 17460 10452 17466 10464
rect 17773 10455 17831 10461
rect 17773 10452 17785 10455
rect 17460 10424 17785 10452
rect 17460 10412 17466 10424
rect 17773 10421 17785 10424
rect 17819 10452 17831 10455
rect 18156 10452 18184 10551
rect 24118 10548 24124 10600
rect 24176 10588 24182 10600
rect 24581 10591 24639 10597
rect 24581 10588 24593 10591
rect 24176 10560 24593 10588
rect 24176 10548 24182 10560
rect 24581 10557 24593 10560
rect 24627 10588 24639 10591
rect 25133 10591 25191 10597
rect 25133 10588 25145 10591
rect 24627 10560 25145 10588
rect 24627 10557 24639 10560
rect 24581 10551 24639 10557
rect 25133 10557 25145 10560
rect 25179 10557 25191 10591
rect 25133 10551 25191 10557
rect 17819 10424 18184 10452
rect 17819 10421 17831 10424
rect 17773 10415 17831 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 4706 10208 4712 10260
rect 4764 10248 4770 10260
rect 5261 10251 5319 10257
rect 5261 10248 5273 10251
rect 4764 10220 5273 10248
rect 4764 10208 4770 10220
rect 5261 10217 5273 10220
rect 5307 10217 5319 10251
rect 8386 10248 8392 10260
rect 8347 10220 8392 10248
rect 5261 10211 5319 10217
rect 8386 10208 8392 10220
rect 8444 10208 8450 10260
rect 9953 10251 10011 10257
rect 9953 10217 9965 10251
rect 9999 10248 10011 10251
rect 10042 10248 10048 10260
rect 9999 10220 10048 10248
rect 9999 10217 10011 10220
rect 9953 10211 10011 10217
rect 10042 10208 10048 10220
rect 10100 10248 10106 10260
rect 10689 10251 10747 10257
rect 10689 10248 10701 10251
rect 10100 10220 10701 10248
rect 10100 10208 10106 10220
rect 10689 10217 10701 10220
rect 10735 10217 10747 10251
rect 12710 10248 12716 10260
rect 12671 10220 12716 10248
rect 10689 10211 10747 10217
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 13630 10248 13636 10260
rect 13188 10220 13636 10248
rect 2593 10183 2651 10189
rect 2593 10149 2605 10183
rect 2639 10180 2651 10183
rect 2774 10180 2780 10192
rect 2639 10152 2780 10180
rect 2639 10149 2651 10152
rect 2593 10143 2651 10149
rect 2774 10140 2780 10152
rect 2832 10180 2838 10192
rect 4430 10189 4436 10192
rect 3421 10183 3479 10189
rect 3421 10180 3433 10183
rect 2832 10152 3433 10180
rect 2832 10140 2838 10152
rect 3421 10149 3433 10152
rect 3467 10149 3479 10183
rect 4427 10180 4436 10189
rect 4343 10152 4436 10180
rect 3421 10143 3479 10149
rect 4427 10143 4436 10152
rect 4488 10180 4494 10192
rect 5534 10180 5540 10192
rect 4488 10152 5540 10180
rect 4430 10140 4436 10143
rect 4488 10140 4494 10152
rect 5534 10140 5540 10152
rect 5592 10140 5598 10192
rect 7190 10180 7196 10192
rect 7151 10152 7196 10180
rect 7190 10140 7196 10152
rect 7248 10140 7254 10192
rect 7742 10180 7748 10192
rect 7703 10152 7748 10180
rect 7742 10140 7748 10152
rect 7800 10140 7806 10192
rect 8018 10140 8024 10192
rect 8076 10180 8082 10192
rect 13188 10189 13216 10220
rect 13630 10208 13636 10220
rect 13688 10208 13694 10260
rect 14458 10208 14464 10260
rect 14516 10248 14522 10260
rect 15013 10251 15071 10257
rect 15013 10248 15025 10251
rect 14516 10220 15025 10248
rect 14516 10208 14522 10220
rect 15013 10217 15025 10220
rect 15059 10217 15071 10251
rect 15654 10248 15660 10260
rect 15615 10220 15660 10248
rect 15013 10211 15071 10217
rect 15654 10208 15660 10220
rect 15712 10208 15718 10260
rect 16482 10208 16488 10260
rect 16540 10248 16546 10260
rect 17451 10251 17509 10257
rect 17451 10248 17463 10251
rect 16540 10220 17463 10248
rect 16540 10208 16546 10220
rect 17451 10217 17463 10220
rect 17497 10217 17509 10251
rect 17451 10211 17509 10217
rect 23707 10251 23765 10257
rect 23707 10217 23719 10251
rect 23753 10248 23765 10251
rect 24210 10248 24216 10260
rect 23753 10220 24216 10248
rect 23753 10217 23765 10220
rect 23707 10211 23765 10217
rect 24210 10208 24216 10220
rect 24268 10208 24274 10260
rect 11241 10183 11299 10189
rect 11241 10180 11253 10183
rect 8076 10152 11253 10180
rect 8076 10140 8082 10152
rect 11241 10149 11253 10152
rect 11287 10149 11299 10183
rect 11241 10143 11299 10149
rect 13173 10183 13231 10189
rect 13173 10149 13185 10183
rect 13219 10149 13231 10183
rect 13173 10143 13231 10149
rect 13354 10140 13360 10192
rect 13412 10180 13418 10192
rect 13725 10183 13783 10189
rect 13725 10180 13737 10183
rect 13412 10152 13737 10180
rect 13412 10140 13418 10152
rect 13725 10149 13737 10152
rect 13771 10149 13783 10183
rect 16942 10180 16948 10192
rect 16903 10152 16948 10180
rect 13725 10143 13783 10149
rect 16942 10140 16948 10152
rect 17000 10140 17006 10192
rect 18414 10180 18420 10192
rect 18375 10152 18420 10180
rect 18414 10140 18420 10152
rect 18472 10140 18478 10192
rect 18509 10183 18567 10189
rect 18509 10149 18521 10183
rect 18555 10180 18567 10183
rect 18598 10180 18604 10192
rect 18555 10152 18604 10180
rect 18555 10149 18567 10152
rect 18509 10143 18567 10149
rect 18598 10140 18604 10152
rect 18656 10140 18662 10192
rect 4522 10072 4528 10124
rect 4580 10112 4586 10124
rect 4985 10115 5043 10121
rect 4985 10112 4997 10115
rect 4580 10084 4997 10112
rect 4580 10072 4586 10084
rect 4985 10081 4997 10084
rect 5031 10081 5043 10115
rect 8570 10112 8576 10124
rect 8531 10084 8576 10112
rect 4985 10075 5043 10081
rect 8570 10072 8576 10084
rect 8628 10072 8634 10124
rect 9861 10115 9919 10121
rect 9861 10081 9873 10115
rect 9907 10081 9919 10115
rect 9861 10075 9919 10081
rect 1397 10047 1455 10053
rect 1397 10013 1409 10047
rect 1443 10044 1455 10047
rect 2222 10044 2228 10056
rect 1443 10016 2228 10044
rect 1443 10013 1455 10016
rect 1397 10007 1455 10013
rect 2222 10004 2228 10016
rect 2280 10004 2286 10056
rect 2501 10047 2559 10053
rect 2501 10013 2513 10047
rect 2547 10013 2559 10047
rect 3142 10044 3148 10056
rect 3103 10016 3148 10044
rect 2501 10007 2559 10013
rect 2406 9936 2412 9988
rect 2464 9976 2470 9988
rect 2516 9976 2544 10007
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 3970 10004 3976 10056
rect 4028 10044 4034 10056
rect 4065 10047 4123 10053
rect 4065 10044 4077 10047
rect 4028 10016 4077 10044
rect 4028 10004 4034 10016
rect 4065 10013 4077 10016
rect 4111 10013 4123 10047
rect 4065 10007 4123 10013
rect 7101 10047 7159 10053
rect 7101 10013 7113 10047
rect 7147 10013 7159 10047
rect 9876 10044 9904 10075
rect 9950 10072 9956 10124
rect 10008 10112 10014 10124
rect 10137 10115 10195 10121
rect 10137 10112 10149 10115
rect 10008 10084 10149 10112
rect 10008 10072 10014 10084
rect 10137 10081 10149 10084
rect 10183 10081 10195 10115
rect 11606 10112 11612 10124
rect 11567 10084 11612 10112
rect 10137 10075 10195 10081
rect 11606 10072 11612 10084
rect 11664 10072 11670 10124
rect 17310 10112 17316 10124
rect 17271 10084 17316 10112
rect 17310 10072 17316 10084
rect 17368 10072 17374 10124
rect 23636 10115 23694 10121
rect 23636 10081 23648 10115
rect 23682 10112 23694 10115
rect 23842 10112 23848 10124
rect 23682 10084 23848 10112
rect 23682 10081 23694 10084
rect 23636 10075 23694 10081
rect 23842 10072 23848 10084
rect 23900 10072 23906 10124
rect 10870 10044 10876 10056
rect 9876 10016 10876 10044
rect 7101 10007 7159 10013
rect 2464 9948 2544 9976
rect 2464 9936 2470 9948
rect 3326 9936 3332 9988
rect 3384 9976 3390 9988
rect 4706 9976 4712 9988
rect 3384 9948 4712 9976
rect 3384 9936 3390 9948
rect 4706 9936 4712 9948
rect 4764 9936 4770 9988
rect 1762 9868 1768 9920
rect 1820 9908 1826 9920
rect 1857 9911 1915 9917
rect 1857 9908 1869 9911
rect 1820 9880 1869 9908
rect 1820 9868 1826 9880
rect 1857 9877 1869 9880
rect 1903 9877 1915 9911
rect 2314 9908 2320 9920
rect 2275 9880 2320 9908
rect 1857 9871 1915 9877
rect 2314 9868 2320 9880
rect 2372 9868 2378 9920
rect 2590 9868 2596 9920
rect 2648 9908 2654 9920
rect 3789 9911 3847 9917
rect 3789 9908 3801 9911
rect 2648 9880 3801 9908
rect 2648 9868 2654 9880
rect 3789 9877 3801 9880
rect 3835 9877 3847 9911
rect 3789 9871 3847 9877
rect 6917 9911 6975 9917
rect 6917 9877 6929 9911
rect 6963 9908 6975 9911
rect 7116 9908 7144 10007
rect 10870 10004 10876 10016
rect 10928 10004 10934 10056
rect 13081 10047 13139 10053
rect 13081 10013 13093 10047
rect 13127 10044 13139 10047
rect 15289 10047 15347 10053
rect 13127 10016 13814 10044
rect 13127 10013 13139 10016
rect 13081 10007 13139 10013
rect 13786 9988 13814 10016
rect 15289 10013 15301 10047
rect 15335 10044 15347 10047
rect 15838 10044 15844 10056
rect 15335 10016 15844 10044
rect 15335 10013 15347 10016
rect 15289 10007 15347 10013
rect 15838 10004 15844 10016
rect 15896 10004 15902 10056
rect 19058 10044 19064 10056
rect 19019 10016 19064 10044
rect 19058 10004 19064 10016
rect 19116 10004 19122 10056
rect 13722 9936 13728 9988
rect 13780 9948 13814 9988
rect 16209 9979 16267 9985
rect 13780 9936 13786 9948
rect 16209 9945 16221 9979
rect 16255 9976 16267 9979
rect 17402 9976 17408 9988
rect 16255 9948 17408 9976
rect 16255 9945 16267 9948
rect 16209 9939 16267 9945
rect 17402 9936 17408 9948
rect 17460 9936 17466 9988
rect 7374 9908 7380 9920
rect 6963 9880 7380 9908
rect 6963 9877 6975 9880
rect 6917 9871 6975 9877
rect 7374 9868 7380 9880
rect 7432 9868 7438 9920
rect 7650 9868 7656 9920
rect 7708 9908 7714 9920
rect 8757 9911 8815 9917
rect 8757 9908 8769 9911
rect 7708 9880 8769 9908
rect 7708 9868 7714 9880
rect 8757 9877 8769 9880
rect 8803 9877 8815 9911
rect 8757 9871 8815 9877
rect 14553 9911 14611 9917
rect 14553 9877 14565 9911
rect 14599 9908 14611 9911
rect 14734 9908 14740 9920
rect 14599 9880 14740 9908
rect 14599 9877 14611 9880
rect 14553 9871 14611 9877
rect 14734 9868 14740 9880
rect 14792 9868 14798 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 1535 9707 1593 9713
rect 1535 9673 1547 9707
rect 1581 9704 1593 9707
rect 1670 9704 1676 9716
rect 1581 9676 1676 9704
rect 1581 9673 1593 9676
rect 1535 9667 1593 9673
rect 1670 9664 1676 9676
rect 1728 9664 1734 9716
rect 3142 9664 3148 9716
rect 3200 9704 3206 9716
rect 3200 9676 4154 9704
rect 3200 9664 3206 9676
rect 4126 9636 4154 9676
rect 7190 9664 7196 9716
rect 7248 9704 7254 9716
rect 7745 9707 7803 9713
rect 7745 9704 7757 9707
rect 7248 9676 7757 9704
rect 7248 9664 7254 9676
rect 7745 9673 7757 9676
rect 7791 9704 7803 9707
rect 8113 9707 8171 9713
rect 8113 9704 8125 9707
rect 7791 9676 8125 9704
rect 7791 9673 7803 9676
rect 7745 9667 7803 9673
rect 8113 9673 8125 9676
rect 8159 9704 8171 9707
rect 11606 9704 11612 9716
rect 8159 9676 11612 9704
rect 8159 9673 8171 9676
rect 8113 9667 8171 9673
rect 11606 9664 11612 9676
rect 11664 9664 11670 9716
rect 13357 9707 13415 9713
rect 13357 9673 13369 9707
rect 13403 9704 13415 9707
rect 13630 9704 13636 9716
rect 13403 9676 13636 9704
rect 13403 9673 13415 9676
rect 13357 9667 13415 9673
rect 13630 9664 13636 9676
rect 13688 9664 13694 9716
rect 15381 9707 15439 9713
rect 15381 9673 15393 9707
rect 15427 9704 15439 9707
rect 15654 9704 15660 9716
rect 15427 9676 15660 9704
rect 15427 9673 15439 9676
rect 15381 9667 15439 9673
rect 15654 9664 15660 9676
rect 15712 9664 15718 9716
rect 17865 9707 17923 9713
rect 17865 9673 17877 9707
rect 17911 9704 17923 9707
rect 18414 9704 18420 9716
rect 17911 9676 18420 9704
rect 17911 9673 17923 9676
rect 17865 9667 17923 9673
rect 18414 9664 18420 9676
rect 18472 9664 18478 9716
rect 23842 9704 23848 9716
rect 23803 9676 23848 9704
rect 23842 9664 23848 9676
rect 23900 9664 23906 9716
rect 4614 9636 4620 9648
rect 4126 9608 4620 9636
rect 4614 9596 4620 9608
rect 4672 9596 4678 9648
rect 5626 9596 5632 9648
rect 5684 9636 5690 9648
rect 6641 9639 6699 9645
rect 6641 9636 6653 9639
rect 5684 9608 6653 9636
rect 5684 9596 5690 9608
rect 6641 9605 6653 9608
rect 6687 9636 6699 9639
rect 8481 9639 8539 9645
rect 6687 9608 7328 9636
rect 6687 9605 6699 9608
rect 6641 9599 6699 9605
rect 2222 9528 2228 9580
rect 2280 9568 2286 9580
rect 4065 9571 4123 9577
rect 4065 9568 4077 9571
rect 2280 9540 4077 9568
rect 2280 9528 2286 9540
rect 4065 9537 4077 9540
rect 4111 9568 4123 9571
rect 4985 9571 5043 9577
rect 4985 9568 4997 9571
rect 4111 9540 4997 9568
rect 4111 9537 4123 9540
rect 4065 9531 4123 9537
rect 4985 9537 4997 9540
rect 5031 9537 5043 9571
rect 4985 9531 5043 9537
rect 6730 9528 6736 9580
rect 6788 9568 6794 9580
rect 7190 9568 7196 9580
rect 6788 9540 7196 9568
rect 6788 9528 6794 9540
rect 7190 9528 7196 9540
rect 7248 9528 7254 9580
rect 1464 9503 1522 9509
rect 1464 9469 1476 9503
rect 1510 9500 1522 9503
rect 1854 9500 1860 9512
rect 1510 9472 1860 9500
rect 1510 9469 1522 9472
rect 1464 9463 1522 9469
rect 1854 9460 1860 9472
rect 1912 9460 1918 9512
rect 2317 9503 2375 9509
rect 2317 9469 2329 9503
rect 2363 9500 2375 9503
rect 2774 9500 2780 9512
rect 2363 9472 2780 9500
rect 2363 9469 2375 9472
rect 2317 9463 2375 9469
rect 2774 9460 2780 9472
rect 2832 9460 2838 9512
rect 5788 9503 5846 9509
rect 5788 9469 5800 9503
rect 5834 9500 5846 9503
rect 6822 9500 6828 9512
rect 5834 9472 6316 9500
rect 6783 9472 6828 9500
rect 5834 9469 5846 9472
rect 5788 9463 5846 9469
rect 6288 9441 6316 9472
rect 6822 9460 6828 9472
rect 6880 9460 6886 9512
rect 3145 9435 3203 9441
rect 3145 9401 3157 9435
rect 3191 9432 3203 9435
rect 3421 9435 3479 9441
rect 3421 9432 3433 9435
rect 3191 9404 3433 9432
rect 3191 9401 3203 9404
rect 3145 9395 3203 9401
rect 3421 9401 3433 9404
rect 3467 9432 3479 9435
rect 4157 9435 4215 9441
rect 3467 9404 3924 9432
rect 3467 9401 3479 9404
rect 3421 9395 3479 9401
rect 2682 9324 2688 9376
rect 2740 9364 2746 9376
rect 3789 9367 3847 9373
rect 3789 9364 3801 9367
rect 2740 9336 3801 9364
rect 2740 9324 2746 9336
rect 3789 9333 3801 9336
rect 3835 9333 3847 9367
rect 3896 9364 3924 9404
rect 4157 9401 4169 9435
rect 4203 9401 4215 9435
rect 4157 9395 4215 9401
rect 6273 9435 6331 9441
rect 6273 9401 6285 9435
rect 6319 9432 6331 9435
rect 7187 9435 7245 9441
rect 6319 9404 6868 9432
rect 6319 9401 6331 9404
rect 6273 9395 6331 9401
rect 4172 9364 4200 9395
rect 3896 9336 4200 9364
rect 3789 9327 3847 9333
rect 4706 9324 4712 9376
rect 4764 9364 4770 9376
rect 5353 9367 5411 9373
rect 5353 9364 5365 9367
rect 4764 9336 5365 9364
rect 4764 9324 4770 9336
rect 5353 9333 5365 9336
rect 5399 9333 5411 9367
rect 5353 9327 5411 9333
rect 5859 9367 5917 9373
rect 5859 9333 5871 9367
rect 5905 9364 5917 9367
rect 6086 9364 6092 9376
rect 5905 9336 6092 9364
rect 5905 9333 5917 9336
rect 5859 9327 5917 9333
rect 6086 9324 6092 9336
rect 6144 9324 6150 9376
rect 6840 9364 6868 9404
rect 7187 9401 7199 9435
rect 7233 9432 7245 9435
rect 7300 9432 7328 9608
rect 8481 9605 8493 9639
rect 8527 9636 8539 9639
rect 8570 9636 8576 9648
rect 8527 9608 8576 9636
rect 8527 9605 8539 9608
rect 8481 9599 8539 9605
rect 8496 9500 8524 9599
rect 8570 9596 8576 9608
rect 8628 9636 8634 9648
rect 9398 9636 9404 9648
rect 8628 9608 9168 9636
rect 9359 9608 9404 9636
rect 8628 9596 8634 9608
rect 8565 9503 8623 9509
rect 8565 9500 8577 9503
rect 8496 9472 8577 9500
rect 8565 9469 8577 9472
rect 8611 9469 8623 9503
rect 8565 9463 8623 9469
rect 8202 9432 8208 9444
rect 7233 9404 8208 9432
rect 7233 9401 7245 9404
rect 7187 9395 7245 9401
rect 8202 9392 8208 9404
rect 8260 9392 8266 9444
rect 9140 9441 9168 9608
rect 9398 9596 9404 9608
rect 9456 9596 9462 9648
rect 9766 9596 9772 9648
rect 9824 9636 9830 9648
rect 12161 9639 12219 9645
rect 12161 9636 12173 9639
rect 9824 9608 12173 9636
rect 9824 9596 9830 9608
rect 12161 9605 12173 9608
rect 12207 9605 12219 9639
rect 12161 9599 12219 9605
rect 9416 9500 9444 9596
rect 12176 9568 12204 9599
rect 13722 9596 13728 9648
rect 13780 9636 13786 9648
rect 19058 9636 19064 9648
rect 13780 9608 19064 9636
rect 13780 9596 13786 9608
rect 19058 9596 19064 9608
rect 19116 9636 19122 9648
rect 19153 9639 19211 9645
rect 19153 9636 19165 9639
rect 19116 9608 19165 9636
rect 19116 9596 19122 9608
rect 19153 9605 19165 9608
rect 19199 9605 19211 9639
rect 19153 9599 19211 9605
rect 14734 9568 14740 9580
rect 12176 9540 12801 9568
rect 14695 9540 14740 9568
rect 9677 9503 9735 9509
rect 9677 9500 9689 9503
rect 9416 9472 9689 9500
rect 9677 9469 9689 9472
rect 9723 9500 9735 9503
rect 9858 9500 9864 9512
rect 9723 9472 9864 9500
rect 9723 9469 9735 9472
rect 9677 9463 9735 9469
rect 9858 9460 9864 9472
rect 9916 9460 9922 9512
rect 12158 9460 12164 9512
rect 12216 9500 12222 9512
rect 12437 9503 12495 9509
rect 12437 9500 12449 9503
rect 12216 9472 12449 9500
rect 12216 9460 12222 9472
rect 12437 9469 12449 9472
rect 12483 9469 12495 9503
rect 12437 9463 12495 9469
rect 12773 9444 12801 9540
rect 14734 9528 14740 9540
rect 14792 9528 14798 9580
rect 18601 9571 18659 9577
rect 15672 9540 16252 9568
rect 13906 9460 13912 9512
rect 13964 9500 13970 9512
rect 14185 9503 14243 9509
rect 14185 9500 14197 9503
rect 13964 9472 14197 9500
rect 13964 9460 13970 9472
rect 14185 9469 14197 9472
rect 14231 9469 14243 9503
rect 14185 9463 14243 9469
rect 14642 9460 14648 9512
rect 14700 9500 14706 9512
rect 15672 9500 15700 9540
rect 16224 9509 16252 9540
rect 18601 9537 18613 9571
rect 18647 9568 18659 9571
rect 19518 9568 19524 9580
rect 18647 9540 19524 9568
rect 18647 9537 18659 9540
rect 18601 9531 18659 9537
rect 19518 9528 19524 9540
rect 19576 9528 19582 9580
rect 14700 9472 15700 9500
rect 16025 9503 16083 9509
rect 14700 9460 14706 9472
rect 16025 9469 16037 9503
rect 16071 9469 16083 9503
rect 16025 9463 16083 9469
rect 16209 9503 16267 9509
rect 16209 9469 16221 9503
rect 16255 9500 16267 9503
rect 16482 9500 16488 9512
rect 16255 9472 16488 9500
rect 16255 9469 16267 9472
rect 16209 9463 16267 9469
rect 9125 9435 9183 9441
rect 9125 9401 9137 9435
rect 9171 9432 9183 9435
rect 9585 9435 9643 9441
rect 9585 9432 9597 9435
rect 9171 9404 9597 9432
rect 9171 9401 9183 9404
rect 9125 9395 9183 9401
rect 9585 9401 9597 9404
rect 9631 9401 9643 9435
rect 12710 9432 12716 9444
rect 12668 9404 12716 9432
rect 9585 9395 9643 9401
rect 12710 9392 12716 9404
rect 12768 9441 12801 9444
rect 12768 9435 12816 9441
rect 12768 9401 12770 9435
rect 12804 9401 12816 9435
rect 12768 9395 12816 9401
rect 12768 9392 12774 9395
rect 13630 9392 13636 9444
rect 13688 9432 13694 9444
rect 16040 9432 16068 9463
rect 16482 9460 16488 9472
rect 16540 9460 16546 9512
rect 16761 9435 16819 9441
rect 16761 9432 16773 9435
rect 13688 9404 16773 9432
rect 13688 9392 13694 9404
rect 16761 9401 16773 9404
rect 16807 9401 16819 9435
rect 16761 9395 16819 9401
rect 18690 9392 18696 9444
rect 18748 9432 18754 9444
rect 18748 9404 18793 9432
rect 18748 9392 18754 9404
rect 7282 9364 7288 9376
rect 6840 9336 7288 9364
rect 7282 9324 7288 9336
rect 7340 9324 7346 9376
rect 7466 9324 7472 9376
rect 7524 9364 7530 9376
rect 8757 9367 8815 9373
rect 8757 9364 8769 9367
rect 7524 9336 8769 9364
rect 7524 9324 7530 9336
rect 8757 9333 8769 9336
rect 8803 9364 8815 9367
rect 10689 9367 10747 9373
rect 10689 9364 10701 9367
rect 8803 9336 10701 9364
rect 8803 9333 8815 9336
rect 8757 9327 8815 9333
rect 10689 9333 10701 9336
rect 10735 9364 10747 9367
rect 10870 9364 10876 9376
rect 10735 9336 10876 9364
rect 10735 9333 10747 9336
rect 10689 9327 10747 9333
rect 10870 9324 10876 9336
rect 10928 9324 10934 9376
rect 11146 9364 11152 9376
rect 11107 9336 11152 9364
rect 11146 9324 11152 9336
rect 11204 9324 11210 9376
rect 13906 9324 13912 9376
rect 13964 9364 13970 9376
rect 14001 9367 14059 9373
rect 14001 9364 14013 9367
rect 13964 9336 14013 9364
rect 13964 9324 13970 9336
rect 14001 9333 14013 9336
rect 14047 9333 14059 9367
rect 15838 9364 15844 9376
rect 15799 9336 15844 9364
rect 14001 9327 14059 9333
rect 15838 9324 15844 9336
rect 15896 9324 15902 9376
rect 17310 9364 17316 9376
rect 17271 9336 17316 9364
rect 17310 9324 17316 9336
rect 17368 9324 17374 9376
rect 18417 9367 18475 9373
rect 18417 9333 18429 9367
rect 18463 9364 18475 9367
rect 18708 9364 18736 9392
rect 18463 9336 18736 9364
rect 18463 9333 18475 9336
rect 18417 9327 18475 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 2593 9163 2651 9169
rect 2593 9129 2605 9163
rect 2639 9160 2651 9163
rect 2682 9160 2688 9172
rect 2639 9132 2688 9160
rect 2639 9129 2651 9132
rect 2593 9123 2651 9129
rect 2682 9120 2688 9132
rect 2740 9120 2746 9172
rect 2774 9120 2780 9172
rect 2832 9160 2838 9172
rect 3145 9163 3203 9169
rect 3145 9160 3157 9163
rect 2832 9132 3157 9160
rect 2832 9120 2838 9132
rect 3145 9129 3157 9132
rect 3191 9129 3203 9163
rect 3145 9123 3203 9129
rect 3234 9120 3240 9172
rect 3292 9160 3298 9172
rect 5077 9163 5135 9169
rect 5077 9160 5089 9163
rect 3292 9132 5089 9160
rect 3292 9120 3298 9132
rect 5077 9129 5089 9132
rect 5123 9160 5135 9163
rect 5258 9160 5264 9172
rect 5123 9132 5264 9160
rect 5123 9129 5135 9132
rect 5077 9123 5135 9129
rect 5258 9120 5264 9132
rect 5316 9120 5322 9172
rect 5626 9160 5632 9172
rect 5587 9132 5632 9160
rect 5626 9120 5632 9132
rect 5684 9120 5690 9172
rect 6086 9120 6092 9172
rect 6144 9160 6150 9172
rect 6457 9163 6515 9169
rect 6457 9160 6469 9163
rect 6144 9132 6469 9160
rect 6144 9120 6150 9132
rect 6457 9129 6469 9132
rect 6503 9160 6515 9163
rect 11882 9160 11888 9172
rect 6503 9132 7144 9160
rect 6503 9129 6515 9132
rect 6457 9123 6515 9129
rect 6822 9092 6828 9104
rect 6783 9064 6828 9092
rect 6822 9052 6828 9064
rect 6880 9052 6886 9104
rect 7116 9101 7144 9132
rect 11072 9132 11888 9160
rect 11072 9104 11100 9132
rect 11882 9120 11888 9132
rect 11940 9120 11946 9172
rect 13541 9163 13599 9169
rect 13541 9129 13553 9163
rect 13587 9160 13599 9163
rect 13722 9160 13728 9172
rect 13587 9132 13728 9160
rect 13587 9129 13599 9132
rect 13541 9123 13599 9129
rect 13722 9120 13728 9132
rect 13780 9120 13786 9172
rect 15105 9163 15163 9169
rect 15105 9129 15117 9163
rect 15151 9160 15163 9163
rect 15838 9160 15844 9172
rect 15151 9132 15844 9160
rect 15151 9129 15163 9132
rect 15105 9123 15163 9129
rect 15838 9120 15844 9132
rect 15896 9120 15902 9172
rect 16482 9160 16488 9172
rect 16443 9132 16488 9160
rect 16482 9120 16488 9132
rect 16540 9120 16546 9172
rect 18690 9120 18696 9172
rect 18748 9160 18754 9172
rect 18877 9163 18935 9169
rect 18877 9160 18889 9163
rect 18748 9132 18889 9160
rect 18748 9120 18754 9132
rect 18877 9129 18889 9132
rect 18923 9129 18935 9163
rect 18877 9123 18935 9129
rect 7101 9095 7159 9101
rect 7101 9061 7113 9095
rect 7147 9061 7159 9095
rect 7101 9055 7159 9061
rect 7190 9052 7196 9104
rect 7248 9092 7254 9104
rect 11054 9092 11060 9104
rect 7248 9064 7293 9092
rect 10967 9064 11060 9092
rect 7248 9052 7254 9064
rect 11054 9052 11060 9064
rect 11112 9052 11118 9104
rect 11146 9052 11152 9104
rect 11204 9092 11210 9104
rect 12250 9092 12256 9104
rect 11204 9064 12256 9092
rect 11204 9052 11210 9064
rect 12250 9052 12256 9064
rect 12308 9092 12314 9104
rect 12529 9095 12587 9101
rect 12529 9092 12541 9095
rect 12308 9064 12541 9092
rect 12308 9052 12314 9064
rect 12529 9061 12541 9064
rect 12575 9061 12587 9095
rect 12529 9055 12587 9061
rect 12618 9052 12624 9104
rect 12676 9092 12682 9104
rect 13170 9092 13176 9104
rect 12676 9064 12721 9092
rect 13131 9064 13176 9092
rect 12676 9052 12682 9064
rect 13170 9052 13176 9064
rect 13228 9052 13234 9104
rect 15470 9052 15476 9104
rect 15528 9092 15534 9104
rect 15654 9101 15660 9104
rect 15610 9095 15660 9101
rect 15610 9092 15622 9095
rect 15528 9064 15622 9092
rect 15528 9052 15534 9064
rect 15610 9061 15622 9064
rect 15656 9061 15660 9095
rect 15610 9055 15660 9061
rect 15654 9052 15660 9055
rect 15712 9052 15718 9104
rect 3602 8984 3608 9036
rect 3660 9024 3666 9036
rect 4065 9027 4123 9033
rect 3660 8996 3924 9024
rect 3660 8984 3666 8996
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8956 2283 8959
rect 2271 8928 3832 8956
rect 2271 8925 2283 8928
rect 2225 8919 2283 8925
rect 3804 8832 3832 8928
rect 1394 8780 1400 8832
rect 1452 8820 1458 8832
rect 1581 8823 1639 8829
rect 1581 8820 1593 8823
rect 1452 8792 1593 8820
rect 1452 8780 1458 8792
rect 1581 8789 1593 8792
rect 1627 8789 1639 8823
rect 2038 8820 2044 8832
rect 1999 8792 2044 8820
rect 1581 8783 1639 8789
rect 2038 8780 2044 8792
rect 2096 8780 2102 8832
rect 3510 8820 3516 8832
rect 3471 8792 3516 8820
rect 3510 8780 3516 8792
rect 3568 8780 3574 8832
rect 3786 8820 3792 8832
rect 3747 8792 3792 8820
rect 3786 8780 3792 8792
rect 3844 8780 3850 8832
rect 3896 8820 3924 8996
rect 4065 8993 4077 9027
rect 4111 9024 4123 9027
rect 4246 9024 4252 9036
rect 4111 8996 4252 9024
rect 4111 8993 4123 8996
rect 4065 8987 4123 8993
rect 3970 8916 3976 8968
rect 4028 8956 4034 8968
rect 4172 8956 4200 8996
rect 4246 8984 4252 8996
rect 4304 8984 4310 9036
rect 5074 8984 5080 9036
rect 5132 9024 5138 9036
rect 5261 9027 5319 9033
rect 5261 9024 5273 9027
rect 5132 8996 5273 9024
rect 5132 8984 5138 8996
rect 5261 8993 5273 8996
rect 5307 9024 5319 9027
rect 5994 9024 6000 9036
rect 5307 8996 6000 9024
rect 5307 8993 5319 8996
rect 5261 8987 5319 8993
rect 5994 8984 6000 8996
rect 6052 8984 6058 9036
rect 8570 9024 8576 9036
rect 8531 8996 8576 9024
rect 8570 8984 8576 8996
rect 8628 8984 8634 9036
rect 9858 9024 9864 9036
rect 9819 8996 9864 9024
rect 9858 8984 9864 8996
rect 9916 8984 9922 9036
rect 7374 8956 7380 8968
rect 4028 8928 4200 8956
rect 7335 8928 7380 8956
rect 4028 8916 4034 8928
rect 7374 8916 7380 8928
rect 7432 8916 7438 8968
rect 7742 8916 7748 8968
rect 7800 8956 7806 8968
rect 8113 8959 8171 8965
rect 8113 8956 8125 8959
rect 7800 8928 8125 8956
rect 7800 8916 7806 8928
rect 8113 8925 8125 8928
rect 8159 8956 8171 8959
rect 9122 8956 9128 8968
rect 8159 8928 9128 8956
rect 8159 8925 8171 8928
rect 8113 8919 8171 8925
rect 9122 8916 9128 8928
rect 9180 8916 9186 8968
rect 10962 8956 10968 8968
rect 10923 8928 10968 8956
rect 10962 8916 10968 8928
rect 11020 8916 11026 8968
rect 11609 8959 11667 8965
rect 11609 8925 11621 8959
rect 11655 8956 11667 8959
rect 13188 8956 13216 9052
rect 17126 9024 17132 9036
rect 17087 8996 17132 9024
rect 17126 8984 17132 8996
rect 17184 8984 17190 9036
rect 18598 9024 18604 9036
rect 18340 8996 18604 9024
rect 11655 8928 13216 8956
rect 11655 8925 11667 8928
rect 11609 8919 11667 8925
rect 14642 8916 14648 8968
rect 14700 8956 14706 8968
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 14700 8928 15301 8956
rect 14700 8916 14706 8928
rect 15289 8925 15301 8928
rect 15335 8925 15347 8959
rect 15289 8919 15347 8925
rect 16206 8916 16212 8968
rect 16264 8956 16270 8968
rect 17037 8959 17095 8965
rect 17037 8956 17049 8959
rect 16264 8928 17049 8956
rect 16264 8916 16270 8928
rect 17037 8925 17049 8928
rect 17083 8925 17095 8959
rect 17037 8919 17095 8925
rect 8294 8848 8300 8900
rect 8352 8888 8358 8900
rect 9950 8888 9956 8900
rect 8352 8860 9956 8888
rect 8352 8848 8358 8860
rect 9950 8848 9956 8860
rect 10008 8888 10014 8900
rect 10321 8891 10379 8897
rect 10321 8888 10333 8891
rect 10008 8860 10333 8888
rect 10008 8848 10014 8860
rect 10321 8857 10333 8860
rect 10367 8857 10379 8891
rect 13630 8888 13636 8900
rect 10321 8851 10379 8857
rect 10520 8860 13636 8888
rect 4249 8823 4307 8829
rect 4249 8820 4261 8823
rect 3896 8792 4261 8820
rect 4249 8789 4261 8792
rect 4295 8789 4307 8823
rect 4249 8783 4307 8789
rect 4338 8780 4344 8832
rect 4396 8820 4402 8832
rect 4525 8823 4583 8829
rect 4525 8820 4537 8823
rect 4396 8792 4537 8820
rect 4396 8780 4402 8792
rect 4525 8789 4537 8792
rect 4571 8789 4583 8823
rect 4525 8783 4583 8789
rect 6086 8780 6092 8832
rect 6144 8820 6150 8832
rect 6181 8823 6239 8829
rect 6181 8820 6193 8823
rect 6144 8792 6193 8820
rect 6144 8780 6150 8792
rect 6181 8789 6193 8792
rect 6227 8789 6239 8823
rect 8386 8820 8392 8832
rect 8347 8792 8392 8820
rect 6181 8783 6239 8789
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 8754 8820 8760 8832
rect 8715 8792 8760 8820
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 10045 8823 10103 8829
rect 10045 8789 10057 8823
rect 10091 8820 10103 8823
rect 10520 8820 10548 8860
rect 13630 8848 13636 8860
rect 13688 8848 13694 8900
rect 10686 8820 10692 8832
rect 10091 8792 10548 8820
rect 10647 8792 10692 8820
rect 10091 8789 10103 8792
rect 10045 8783 10103 8789
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 12158 8780 12164 8832
rect 12216 8820 12222 8832
rect 12253 8823 12311 8829
rect 12253 8820 12265 8823
rect 12216 8792 12265 8820
rect 12216 8780 12222 8792
rect 12253 8789 12265 8792
rect 12299 8789 12311 8823
rect 14182 8820 14188 8832
rect 14143 8792 14188 8820
rect 12253 8783 12311 8789
rect 14182 8780 14188 8792
rect 14240 8820 14246 8832
rect 14550 8820 14556 8832
rect 14240 8792 14556 8820
rect 14240 8780 14246 8792
rect 14550 8780 14556 8792
rect 14608 8780 14614 8832
rect 18340 8829 18368 8996
rect 18598 8984 18604 8996
rect 18656 9024 18662 9036
rect 18693 9027 18751 9033
rect 18693 9024 18705 9027
rect 18656 8996 18705 9024
rect 18656 8984 18662 8996
rect 18693 8993 18705 8996
rect 18739 8993 18751 9027
rect 18693 8987 18751 8993
rect 16209 8823 16267 8829
rect 16209 8789 16221 8823
rect 16255 8820 16267 8823
rect 18325 8823 18383 8829
rect 18325 8820 18337 8823
rect 16255 8792 18337 8820
rect 16255 8789 16267 8792
rect 16209 8783 16267 8789
rect 18325 8789 18337 8792
rect 18371 8789 18383 8823
rect 18325 8783 18383 8789
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 3970 8576 3976 8628
rect 4028 8616 4034 8628
rect 4249 8619 4307 8625
rect 4249 8616 4261 8619
rect 4028 8588 4261 8616
rect 4028 8576 4034 8588
rect 4249 8585 4261 8588
rect 4295 8585 4307 8619
rect 4249 8579 4307 8585
rect 5077 8619 5135 8625
rect 5077 8585 5089 8619
rect 5123 8616 5135 8619
rect 5534 8616 5540 8628
rect 5123 8588 5540 8616
rect 5123 8585 5135 8588
rect 5077 8579 5135 8585
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 5994 8576 6000 8628
rect 6052 8616 6058 8628
rect 6181 8619 6239 8625
rect 6181 8616 6193 8619
rect 6052 8588 6193 8616
rect 6052 8576 6058 8588
rect 6181 8585 6193 8588
rect 6227 8585 6239 8619
rect 6181 8579 6239 8585
rect 7101 8619 7159 8625
rect 7101 8585 7113 8619
rect 7147 8616 7159 8619
rect 7190 8616 7196 8628
rect 7147 8588 7196 8616
rect 7147 8585 7159 8588
rect 7101 8579 7159 8585
rect 7190 8576 7196 8588
rect 7248 8576 7254 8628
rect 8570 8616 8576 8628
rect 8531 8588 8576 8616
rect 8570 8576 8576 8588
rect 8628 8576 8634 8628
rect 9769 8619 9827 8625
rect 9769 8585 9781 8619
rect 9815 8616 9827 8619
rect 9858 8616 9864 8628
rect 9815 8588 9864 8616
rect 9815 8585 9827 8588
rect 9769 8579 9827 8585
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 10781 8619 10839 8625
rect 10781 8585 10793 8619
rect 10827 8616 10839 8619
rect 11054 8616 11060 8628
rect 10827 8588 11060 8616
rect 10827 8585 10839 8588
rect 10781 8579 10839 8585
rect 11054 8576 11060 8588
rect 11112 8576 11118 8628
rect 12250 8616 12256 8628
rect 12211 8588 12256 8616
rect 12250 8576 12256 8588
rect 12308 8576 12314 8628
rect 12618 8616 12624 8628
rect 12579 8588 12624 8616
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 14642 8616 14648 8628
rect 14603 8588 14648 8616
rect 14642 8576 14648 8588
rect 14700 8576 14706 8628
rect 17126 8616 17132 8628
rect 17087 8588 17132 8616
rect 17126 8576 17132 8588
rect 17184 8576 17190 8628
rect 18598 8616 18604 8628
rect 18559 8588 18604 8616
rect 18598 8576 18604 8588
rect 18656 8576 18662 8628
rect 19518 8576 19524 8628
rect 19576 8616 19582 8628
rect 19613 8619 19671 8625
rect 19613 8616 19625 8619
rect 19576 8588 19625 8616
rect 19576 8576 19582 8588
rect 19613 8585 19625 8588
rect 19659 8585 19671 8619
rect 19613 8579 19671 8585
rect 3786 8548 3792 8560
rect 3747 8520 3792 8548
rect 3786 8508 3792 8520
rect 3844 8508 3850 8560
rect 6641 8551 6699 8557
rect 6641 8517 6653 8551
rect 6687 8548 6699 8551
rect 7742 8548 7748 8560
rect 6687 8520 7512 8548
rect 7703 8520 7748 8548
rect 6687 8517 6699 8520
rect 6641 8511 6699 8517
rect 7484 8492 7512 8520
rect 7742 8508 7748 8520
rect 7800 8508 7806 8560
rect 7926 8548 7932 8560
rect 7887 8520 7932 8548
rect 7926 8508 7932 8520
rect 7984 8508 7990 8560
rect 15930 8548 15936 8560
rect 15764 8520 15936 8548
rect 1946 8440 1952 8492
rect 2004 8480 2010 8492
rect 2682 8480 2688 8492
rect 2004 8452 2688 8480
rect 2004 8440 2010 8452
rect 2682 8440 2688 8452
rect 2740 8440 2746 8492
rect 4614 8480 4620 8492
rect 3528 8452 4620 8480
rect 3528 8424 3556 8452
rect 4614 8440 4620 8452
rect 4672 8440 4678 8492
rect 5258 8480 5264 8492
rect 5219 8452 5264 8480
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8480 5963 8483
rect 7374 8480 7380 8492
rect 5951 8452 7380 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 7374 8440 7380 8452
rect 7432 8440 7438 8492
rect 7466 8440 7472 8492
rect 7524 8480 7530 8492
rect 7837 8483 7895 8489
rect 7837 8480 7849 8483
rect 7524 8452 7849 8480
rect 7524 8440 7530 8452
rect 7837 8449 7849 8452
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 8846 8440 8852 8492
rect 8904 8480 8910 8492
rect 13173 8483 13231 8489
rect 13173 8480 13185 8483
rect 8904 8452 13185 8480
rect 8904 8440 8910 8452
rect 13173 8449 13185 8452
rect 13219 8480 13231 8483
rect 14090 8480 14096 8492
rect 13219 8452 13814 8480
rect 14051 8452 14096 8480
rect 13219 8449 13231 8452
rect 13173 8443 13231 8449
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8412 1731 8415
rect 3145 8415 3203 8421
rect 1719 8384 2452 8412
rect 1719 8381 1731 8384
rect 1673 8375 1731 8381
rect 1394 8304 1400 8356
rect 1452 8344 1458 8356
rect 1489 8347 1547 8353
rect 1489 8344 1501 8347
rect 1452 8316 1501 8344
rect 1452 8304 1458 8316
rect 1489 8313 1501 8316
rect 1535 8313 1547 8347
rect 1489 8307 1547 8313
rect 1762 8276 1768 8288
rect 1723 8248 1768 8276
rect 1762 8236 1768 8248
rect 1820 8236 1826 8288
rect 2424 8285 2452 8384
rect 3145 8381 3157 8415
rect 3191 8381 3203 8415
rect 3510 8412 3516 8424
rect 3471 8384 3516 8412
rect 3145 8375 3203 8381
rect 2958 8304 2964 8356
rect 3016 8344 3022 8356
rect 3160 8344 3188 8375
rect 3510 8372 3516 8384
rect 3568 8372 3574 8424
rect 3694 8412 3700 8424
rect 3655 8384 3700 8412
rect 3694 8372 3700 8384
rect 3752 8372 3758 8424
rect 7616 8415 7674 8421
rect 7616 8381 7628 8415
rect 7662 8412 7674 8415
rect 8941 8415 8999 8421
rect 8941 8412 8953 8415
rect 7662 8384 8953 8412
rect 7662 8381 7674 8384
rect 7616 8375 7674 8381
rect 8941 8381 8953 8384
rect 8987 8412 8999 8415
rect 9674 8412 9680 8424
rect 8987 8384 9680 8412
rect 8987 8381 8999 8384
rect 8941 8375 8999 8381
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 9861 8415 9919 8421
rect 9861 8381 9873 8415
rect 9907 8412 9919 8415
rect 10686 8412 10692 8424
rect 9907 8384 10692 8412
rect 9907 8381 9919 8384
rect 9861 8375 9919 8381
rect 10686 8372 10692 8384
rect 10744 8372 10750 8424
rect 13630 8412 13636 8424
rect 13591 8384 13636 8412
rect 13630 8372 13636 8384
rect 13688 8372 13694 8424
rect 13786 8412 13814 8452
rect 14090 8440 14096 8452
rect 14148 8440 14154 8492
rect 15764 8489 15792 8520
rect 15930 8508 15936 8520
rect 15988 8548 15994 8560
rect 16669 8551 16727 8557
rect 16669 8548 16681 8551
rect 15988 8520 16681 8548
rect 15988 8508 15994 8520
rect 16669 8517 16681 8520
rect 16715 8517 16727 8551
rect 16669 8511 16727 8517
rect 15749 8483 15807 8489
rect 15749 8449 15761 8483
rect 15795 8449 15807 8483
rect 15749 8443 15807 8449
rect 16114 8440 16120 8492
rect 16172 8480 16178 8492
rect 18049 8483 18107 8489
rect 18049 8480 18061 8483
rect 16172 8452 18061 8480
rect 16172 8440 16178 8452
rect 18049 8449 18061 8452
rect 18095 8449 18107 8483
rect 18049 8443 18107 8449
rect 13909 8415 13967 8421
rect 13909 8412 13921 8415
rect 13786 8384 13921 8412
rect 13909 8381 13921 8384
rect 13955 8412 13967 8415
rect 15378 8412 15384 8424
rect 13955 8384 15384 8412
rect 13955 8381 13967 8384
rect 13909 8375 13967 8381
rect 15378 8372 15384 8384
rect 15436 8372 15442 8424
rect 19404 8415 19462 8421
rect 19404 8381 19416 8415
rect 19450 8412 19462 8415
rect 19450 8384 19932 8412
rect 19450 8381 19462 8384
rect 19404 8375 19462 8381
rect 5353 8347 5411 8353
rect 3016 8316 4752 8344
rect 3016 8304 3022 8316
rect 2409 8279 2467 8285
rect 2409 8245 2421 8279
rect 2455 8276 2467 8279
rect 2498 8276 2504 8288
rect 2455 8248 2504 8276
rect 2455 8245 2467 8248
rect 2409 8239 2467 8245
rect 2498 8236 2504 8248
rect 2556 8236 2562 8288
rect 4614 8276 4620 8288
rect 4575 8248 4620 8276
rect 4614 8236 4620 8248
rect 4672 8236 4678 8288
rect 4724 8276 4752 8316
rect 5353 8313 5365 8347
rect 5399 8344 5411 8347
rect 5534 8344 5540 8356
rect 5399 8316 5540 8344
rect 5399 8313 5411 8316
rect 5353 8307 5411 8313
rect 5534 8304 5540 8316
rect 5592 8344 5598 8356
rect 6086 8344 6092 8356
rect 5592 8316 6092 8344
rect 5592 8304 5598 8316
rect 6086 8304 6092 8316
rect 6144 8304 6150 8356
rect 7466 8344 7472 8356
rect 7427 8316 7472 8344
rect 7466 8304 7472 8316
rect 7524 8304 7530 8356
rect 9401 8347 9459 8353
rect 9401 8313 9413 8347
rect 9447 8344 9459 8347
rect 9766 8344 9772 8356
rect 9447 8316 9772 8344
rect 9447 8313 9459 8316
rect 9401 8307 9459 8313
rect 9766 8304 9772 8316
rect 9824 8344 9830 8356
rect 10182 8347 10240 8353
rect 10182 8344 10194 8347
rect 9824 8316 10194 8344
rect 9824 8304 9830 8316
rect 10182 8313 10194 8316
rect 10228 8313 10240 8347
rect 10182 8307 10240 8313
rect 15013 8347 15071 8353
rect 15013 8313 15025 8347
rect 15059 8344 15071 8347
rect 15059 8316 15700 8344
rect 15059 8313 15071 8316
rect 15013 8307 15071 8313
rect 7484 8276 7512 8304
rect 4724 8248 7512 8276
rect 10962 8236 10968 8288
rect 11020 8276 11026 8288
rect 11425 8279 11483 8285
rect 11425 8276 11437 8279
rect 11020 8248 11437 8276
rect 11020 8236 11026 8248
rect 11425 8245 11437 8248
rect 11471 8245 11483 8279
rect 11425 8239 11483 8245
rect 12710 8236 12716 8288
rect 12768 8276 12774 8288
rect 15289 8279 15347 8285
rect 15289 8276 15301 8279
rect 12768 8248 15301 8276
rect 12768 8236 12774 8248
rect 15289 8245 15301 8248
rect 15335 8276 15347 8279
rect 15470 8276 15476 8288
rect 15335 8248 15476 8276
rect 15335 8245 15347 8248
rect 15289 8239 15347 8245
rect 15470 8236 15476 8248
rect 15528 8236 15534 8288
rect 15672 8276 15700 8316
rect 15838 8304 15844 8356
rect 15896 8344 15902 8356
rect 16390 8344 16396 8356
rect 15896 8316 15941 8344
rect 16351 8316 16396 8344
rect 15896 8304 15902 8316
rect 16390 8304 16396 8316
rect 16448 8304 16454 8356
rect 15856 8276 15884 8304
rect 19904 8285 19932 8384
rect 15672 8248 15884 8276
rect 19889 8279 19947 8285
rect 19889 8245 19901 8279
rect 19935 8276 19947 8279
rect 21174 8276 21180 8288
rect 19935 8248 21180 8276
rect 19935 8245 19947 8248
rect 19889 8239 19947 8245
rect 21174 8236 21180 8248
rect 21232 8236 21238 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 3329 8075 3387 8081
rect 3329 8041 3341 8075
rect 3375 8072 3387 8075
rect 3694 8072 3700 8084
rect 3375 8044 3700 8072
rect 3375 8041 3387 8044
rect 3329 8035 3387 8041
rect 3694 8032 3700 8044
rect 3752 8032 3758 8084
rect 4338 8072 4344 8084
rect 4299 8044 4344 8072
rect 4338 8032 4344 8044
rect 4396 8032 4402 8084
rect 5534 8072 5540 8084
rect 5495 8044 5540 8072
rect 5534 8032 5540 8044
rect 5592 8032 5598 8084
rect 10781 8075 10839 8081
rect 10781 8072 10793 8075
rect 9968 8044 10793 8072
rect 1851 8007 1909 8013
rect 1851 7973 1863 8007
rect 1897 8004 1909 8007
rect 1946 8004 1952 8016
rect 1897 7976 1952 8004
rect 1897 7973 1909 7976
rect 1851 7967 1909 7973
rect 1946 7964 1952 7976
rect 2004 7964 2010 8016
rect 3712 8004 3740 8032
rect 4430 8004 4436 8016
rect 3712 7976 4436 8004
rect 4430 7964 4436 7976
rect 4488 8004 4494 8016
rect 8294 8004 8300 8016
rect 4488 7976 4936 8004
rect 8255 7976 8300 8004
rect 4488 7964 4494 7976
rect 4154 7896 4160 7948
rect 4212 7936 4218 7948
rect 4614 7936 4620 7948
rect 4212 7908 4257 7936
rect 4575 7908 4620 7936
rect 4212 7896 4218 7908
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 4908 7945 4936 7976
rect 8294 7964 8300 7976
rect 8352 7964 8358 8016
rect 4893 7939 4951 7945
rect 4893 7905 4905 7939
rect 4939 7905 4951 7939
rect 6178 7936 6184 7948
rect 6139 7908 6184 7936
rect 4893 7899 4951 7905
rect 6178 7896 6184 7908
rect 6236 7896 6242 7948
rect 7561 7939 7619 7945
rect 7561 7905 7573 7939
rect 7607 7936 7619 7939
rect 7742 7936 7748 7948
rect 7607 7908 7748 7936
rect 7607 7905 7619 7908
rect 7561 7899 7619 7905
rect 7742 7896 7748 7908
rect 7800 7896 7806 7948
rect 9968 7945 9996 8044
rect 10781 8041 10793 8044
rect 10827 8072 10839 8075
rect 10870 8072 10876 8084
rect 10827 8044 10876 8072
rect 10827 8041 10839 8044
rect 10781 8035 10839 8041
rect 10870 8032 10876 8044
rect 10928 8032 10934 8084
rect 12158 8072 12164 8084
rect 12119 8044 12164 8072
rect 12158 8032 12164 8044
rect 12216 8032 12222 8084
rect 17129 8075 17187 8081
rect 17129 8072 17141 8075
rect 15304 8044 17141 8072
rect 10413 8007 10471 8013
rect 10413 7973 10425 8007
rect 10459 8004 10471 8007
rect 10686 8004 10692 8016
rect 10459 7976 10692 8004
rect 10459 7973 10471 7976
rect 10413 7967 10471 7973
rect 10686 7964 10692 7976
rect 10744 7964 10750 8016
rect 14277 8007 14335 8013
rect 14277 7973 14289 8007
rect 14323 8004 14335 8007
rect 14642 8004 14648 8016
rect 14323 7976 14648 8004
rect 14323 7973 14335 7976
rect 14277 7967 14335 7973
rect 14642 7964 14648 7976
rect 14700 7964 14706 8016
rect 15304 7948 15332 8044
rect 17129 8041 17141 8044
rect 17175 8041 17187 8075
rect 17129 8035 17187 8041
rect 15470 7964 15476 8016
rect 15528 8004 15534 8016
rect 15610 8007 15668 8013
rect 15610 8004 15622 8007
rect 15528 7976 15622 8004
rect 15528 7964 15534 7976
rect 15610 7973 15622 7976
rect 15656 7973 15668 8007
rect 15610 7967 15668 7973
rect 15717 7976 17540 8004
rect 9953 7939 10011 7945
rect 9953 7905 9965 7939
rect 9999 7905 10011 7939
rect 9953 7899 10011 7905
rect 10042 7896 10048 7948
rect 10100 7936 10106 7948
rect 10137 7939 10195 7945
rect 10137 7936 10149 7939
rect 10100 7908 10149 7936
rect 10100 7896 10106 7908
rect 10137 7905 10149 7908
rect 10183 7936 10195 7939
rect 11057 7939 11115 7945
rect 11057 7936 11069 7939
rect 10183 7908 11069 7936
rect 10183 7905 10195 7908
rect 10137 7899 10195 7905
rect 11057 7905 11069 7908
rect 11103 7905 11115 7939
rect 11057 7899 11115 7905
rect 11977 7939 12035 7945
rect 11977 7905 11989 7939
rect 12023 7905 12035 7939
rect 12342 7936 12348 7948
rect 12303 7908 12348 7936
rect 11977 7899 12035 7905
rect 1489 7871 1547 7877
rect 1489 7837 1501 7871
rect 1535 7868 1547 7871
rect 2038 7868 2044 7880
rect 1535 7840 2044 7868
rect 1535 7837 1547 7840
rect 1489 7831 1547 7837
rect 2038 7828 2044 7840
rect 2096 7868 2102 7880
rect 2774 7868 2780 7880
rect 2096 7840 2780 7868
rect 2096 7828 2102 7840
rect 2774 7828 2780 7840
rect 2832 7828 2838 7880
rect 3694 7868 3700 7880
rect 3607 7840 3700 7868
rect 3694 7828 3700 7840
rect 3752 7868 3758 7880
rect 4632 7868 4660 7896
rect 3752 7840 4660 7868
rect 3752 7828 3758 7840
rect 7006 7828 7012 7880
rect 7064 7868 7070 7880
rect 7929 7871 7987 7877
rect 7929 7868 7941 7871
rect 7064 7840 7941 7868
rect 7064 7828 7070 7840
rect 7929 7837 7941 7840
rect 7975 7868 7987 7871
rect 7975 7840 8248 7868
rect 7975 7837 7987 7840
rect 7929 7831 7987 7837
rect 7726 7803 7784 7809
rect 7726 7769 7738 7803
rect 7772 7800 7784 7803
rect 8110 7800 8116 7812
rect 7772 7772 8116 7800
rect 7772 7769 7784 7772
rect 7726 7763 7784 7769
rect 8110 7760 8116 7772
rect 8168 7760 8174 7812
rect 8220 7800 8248 7840
rect 8754 7828 8760 7880
rect 8812 7868 8818 7880
rect 8812 7840 9674 7868
rect 8812 7828 8818 7840
rect 8386 7800 8392 7812
rect 8220 7772 8392 7800
rect 8386 7760 8392 7772
rect 8444 7800 8450 7812
rect 9646 7800 9674 7840
rect 11992 7812 12020 7899
rect 12342 7896 12348 7908
rect 12400 7896 12406 7948
rect 13449 7939 13507 7945
rect 13449 7905 13461 7939
rect 13495 7936 13507 7939
rect 13630 7936 13636 7948
rect 13495 7908 13636 7936
rect 13495 7905 13507 7908
rect 13449 7899 13507 7905
rect 13630 7896 13636 7908
rect 13688 7896 13694 7948
rect 14001 7939 14059 7945
rect 14001 7936 14013 7939
rect 13786 7908 14013 7936
rect 12360 7868 12388 7896
rect 13786 7868 13814 7908
rect 14001 7905 14013 7908
rect 14047 7905 14059 7939
rect 15286 7936 15292 7948
rect 15199 7908 15292 7936
rect 14001 7899 14059 7905
rect 15286 7896 15292 7908
rect 15344 7896 15350 7948
rect 15378 7896 15384 7948
rect 15436 7936 15442 7948
rect 15717 7936 15745 7976
rect 17512 7948 17540 7976
rect 15436 7908 15745 7936
rect 15436 7896 15442 7908
rect 17034 7896 17040 7948
rect 17092 7936 17098 7948
rect 17129 7939 17187 7945
rect 17129 7936 17141 7939
rect 17092 7908 17141 7936
rect 17092 7896 17098 7908
rect 17129 7905 17141 7908
rect 17175 7905 17187 7939
rect 17494 7936 17500 7948
rect 17455 7908 17500 7936
rect 17129 7899 17187 7905
rect 17494 7896 17500 7908
rect 17552 7896 17558 7948
rect 12360 7840 13814 7868
rect 11974 7800 11980 7812
rect 8444 7772 9076 7800
rect 9646 7772 11980 7800
rect 8444 7760 8450 7772
rect 9048 7744 9076 7772
rect 11974 7760 11980 7772
rect 12032 7760 12038 7812
rect 15838 7760 15844 7812
rect 15896 7800 15902 7812
rect 16209 7803 16267 7809
rect 16209 7800 16221 7803
rect 15896 7772 16221 7800
rect 15896 7760 15902 7772
rect 16209 7769 16221 7772
rect 16255 7800 16267 7803
rect 17126 7800 17132 7812
rect 16255 7772 17132 7800
rect 16255 7769 16267 7772
rect 16209 7763 16267 7769
rect 17126 7760 17132 7772
rect 17184 7760 17190 7812
rect 2222 7692 2228 7744
rect 2280 7732 2286 7744
rect 2409 7735 2467 7741
rect 2409 7732 2421 7735
rect 2280 7704 2421 7732
rect 2280 7692 2286 7704
rect 2409 7701 2421 7704
rect 2455 7701 2467 7735
rect 2958 7732 2964 7744
rect 2919 7704 2964 7732
rect 2409 7695 2467 7701
rect 2958 7692 2964 7704
rect 3016 7692 3022 7744
rect 5905 7735 5963 7741
rect 5905 7701 5917 7735
rect 5951 7732 5963 7735
rect 5994 7732 6000 7744
rect 5951 7704 6000 7732
rect 5951 7701 5963 7704
rect 5905 7695 5963 7701
rect 5994 7692 6000 7704
rect 6052 7692 6058 7744
rect 6270 7732 6276 7744
rect 6231 7704 6276 7732
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 7101 7735 7159 7741
rect 7101 7701 7113 7735
rect 7147 7732 7159 7735
rect 7466 7732 7472 7744
rect 7147 7704 7472 7732
rect 7147 7701 7159 7704
rect 7101 7695 7159 7701
rect 7466 7692 7472 7704
rect 7524 7692 7530 7744
rect 7834 7732 7840 7744
rect 7795 7704 7840 7732
rect 7834 7692 7840 7704
rect 7892 7692 7898 7744
rect 8570 7732 8576 7744
rect 8531 7704 8576 7732
rect 8570 7692 8576 7704
rect 8628 7692 8634 7744
rect 8938 7732 8944 7744
rect 8899 7704 8944 7732
rect 8938 7692 8944 7704
rect 8996 7692 9002 7744
rect 9030 7692 9036 7744
rect 9088 7732 9094 7744
rect 9401 7735 9459 7741
rect 9401 7732 9413 7735
rect 9088 7704 9413 7732
rect 9088 7692 9094 7704
rect 9401 7701 9413 7704
rect 9447 7732 9459 7735
rect 9858 7732 9864 7744
rect 9447 7704 9864 7732
rect 9447 7701 9459 7704
rect 9401 7695 9459 7701
rect 9858 7692 9864 7704
rect 9916 7692 9922 7744
rect 13906 7692 13912 7744
rect 13964 7732 13970 7744
rect 17034 7732 17040 7744
rect 13964 7704 17040 7732
rect 13964 7692 13970 7704
rect 17034 7692 17040 7704
rect 17092 7692 17098 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 4430 7528 4436 7540
rect 4391 7500 4436 7528
rect 4430 7488 4436 7500
rect 4488 7488 4494 7540
rect 6730 7488 6736 7540
rect 6788 7528 6794 7540
rect 7653 7531 7711 7537
rect 7653 7528 7665 7531
rect 6788 7500 7665 7528
rect 6788 7488 6794 7500
rect 7653 7497 7665 7500
rect 7699 7528 7711 7531
rect 7834 7528 7840 7540
rect 7699 7500 7840 7528
rect 7699 7497 7711 7500
rect 7653 7491 7711 7497
rect 7834 7488 7840 7500
rect 7892 7488 7898 7540
rect 8662 7528 8668 7540
rect 8623 7500 8668 7528
rect 8662 7488 8668 7500
rect 8720 7488 8726 7540
rect 9122 7488 9128 7540
rect 9180 7528 9186 7540
rect 9766 7537 9772 7540
rect 9750 7531 9772 7537
rect 9750 7528 9762 7531
rect 9180 7500 9628 7528
rect 9679 7500 9762 7528
rect 9180 7488 9186 7500
rect 1857 7463 1915 7469
rect 1857 7429 1869 7463
rect 1903 7460 1915 7463
rect 2958 7460 2964 7472
rect 1903 7432 2964 7460
rect 1903 7429 1915 7432
rect 1857 7423 1915 7429
rect 2958 7420 2964 7432
rect 3016 7420 3022 7472
rect 8297 7463 8355 7469
rect 8297 7429 8309 7463
rect 8343 7460 8355 7463
rect 8938 7460 8944 7472
rect 8343 7432 8944 7460
rect 8343 7429 8355 7432
rect 8297 7423 8355 7429
rect 8938 7420 8944 7432
rect 8996 7460 9002 7472
rect 9306 7460 9312 7472
rect 8996 7432 9312 7460
rect 8996 7420 9002 7432
rect 9306 7420 9312 7432
rect 9364 7420 9370 7472
rect 9600 7460 9628 7500
rect 9750 7497 9762 7500
rect 9824 7528 9830 7540
rect 9824 7500 10088 7528
rect 9750 7491 9772 7497
rect 9766 7488 9772 7491
rect 9824 7488 9830 7500
rect 9861 7463 9919 7469
rect 9861 7460 9873 7463
rect 9600 7432 9873 7460
rect 9861 7429 9873 7432
rect 9907 7429 9919 7463
rect 9861 7423 9919 7429
rect 8389 7395 8447 7401
rect 8389 7361 8401 7395
rect 8435 7392 8447 7395
rect 9030 7392 9036 7404
rect 8435 7364 9036 7392
rect 8435 7361 8447 7364
rect 8389 7355 8447 7361
rect 9030 7352 9036 7364
rect 9088 7352 9094 7404
rect 9398 7352 9404 7404
rect 9456 7392 9462 7404
rect 9953 7395 10011 7401
rect 9953 7392 9965 7395
rect 9456 7364 9965 7392
rect 9456 7352 9462 7364
rect 9953 7361 9965 7364
rect 9999 7361 10011 7395
rect 10060 7392 10088 7500
rect 10134 7488 10140 7540
rect 10192 7528 10198 7540
rect 10229 7531 10287 7537
rect 10229 7528 10241 7531
rect 10192 7500 10241 7528
rect 10192 7488 10198 7500
rect 10229 7497 10241 7500
rect 10275 7497 10287 7531
rect 11974 7528 11980 7540
rect 11935 7500 11980 7528
rect 10229 7491 10287 7497
rect 11974 7488 11980 7500
rect 12032 7488 12038 7540
rect 13630 7488 13636 7540
rect 13688 7528 13694 7540
rect 13814 7528 13820 7540
rect 13688 7500 13820 7528
rect 13688 7488 13694 7500
rect 13814 7488 13820 7500
rect 13872 7528 13878 7540
rect 14277 7531 14335 7537
rect 14277 7528 14289 7531
rect 13872 7500 14289 7528
rect 13872 7488 13878 7500
rect 14277 7497 14289 7500
rect 14323 7497 14335 7531
rect 14277 7491 14335 7497
rect 14921 7531 14979 7537
rect 14921 7497 14933 7531
rect 14967 7528 14979 7531
rect 15286 7528 15292 7540
rect 14967 7500 15292 7528
rect 14967 7497 14979 7500
rect 14921 7491 14979 7497
rect 15286 7488 15292 7500
rect 15344 7488 15350 7540
rect 15470 7528 15476 7540
rect 15431 7500 15476 7528
rect 15470 7488 15476 7500
rect 15528 7488 15534 7540
rect 17034 7528 17040 7540
rect 16995 7500 17040 7528
rect 17034 7488 17040 7500
rect 17092 7488 17098 7540
rect 17494 7528 17500 7540
rect 17455 7500 17500 7528
rect 17494 7488 17500 7500
rect 17552 7488 17558 7540
rect 25130 7528 25136 7540
rect 25091 7500 25136 7528
rect 25130 7488 25136 7500
rect 25188 7488 25194 7540
rect 13446 7420 13452 7472
rect 13504 7460 13510 7472
rect 17773 7463 17831 7469
rect 17773 7460 17785 7463
rect 13504 7432 17785 7460
rect 13504 7420 13510 7432
rect 17773 7429 17785 7432
rect 17819 7429 17831 7463
rect 17773 7423 17831 7429
rect 10597 7395 10655 7401
rect 10597 7392 10609 7395
rect 10060 7364 10609 7392
rect 9953 7355 10011 7361
rect 10597 7361 10609 7364
rect 10643 7392 10655 7395
rect 10686 7392 10692 7404
rect 10643 7364 10692 7392
rect 10643 7361 10655 7364
rect 10597 7355 10655 7361
rect 10686 7352 10692 7364
rect 10744 7352 10750 7404
rect 13998 7392 14004 7404
rect 13959 7364 14004 7392
rect 13998 7352 14004 7364
rect 14056 7352 14062 7404
rect 16390 7392 16396 7404
rect 15095 7364 16396 7392
rect 15095 7336 15123 7364
rect 16390 7352 16396 7364
rect 16448 7352 16454 7404
rect 1673 7327 1731 7333
rect 1673 7293 1685 7327
rect 1719 7324 1731 7327
rect 1854 7324 1860 7336
rect 1719 7296 1860 7324
rect 1719 7293 1731 7296
rect 1673 7287 1731 7293
rect 1854 7284 1860 7296
rect 1912 7324 1918 7336
rect 2501 7327 2559 7333
rect 2501 7324 2513 7327
rect 1912 7296 2513 7324
rect 1912 7284 1918 7296
rect 2501 7293 2513 7296
rect 2547 7293 2559 7327
rect 2958 7324 2964 7336
rect 2919 7296 2964 7324
rect 2501 7287 2559 7293
rect 2958 7284 2964 7296
rect 3016 7284 3022 7336
rect 3510 7324 3516 7336
rect 3471 7296 3516 7324
rect 3510 7284 3516 7296
rect 3568 7284 3574 7336
rect 3694 7324 3700 7336
rect 3655 7296 3700 7324
rect 3694 7284 3700 7296
rect 3752 7284 3758 7336
rect 3878 7284 3884 7336
rect 3936 7324 3942 7336
rect 5077 7327 5135 7333
rect 5077 7324 5089 7327
rect 3936 7296 5089 7324
rect 3936 7284 3942 7296
rect 5077 7293 5089 7296
rect 5123 7324 5135 7327
rect 5813 7327 5871 7333
rect 5813 7324 5825 7327
rect 5123 7296 5825 7324
rect 5123 7293 5135 7296
rect 5077 7287 5135 7293
rect 5813 7293 5825 7296
rect 5859 7324 5871 7327
rect 6730 7324 6736 7336
rect 5859 7296 6736 7324
rect 5859 7293 5871 7296
rect 5813 7287 5871 7293
rect 6730 7284 6736 7296
rect 6788 7284 6794 7336
rect 6825 7327 6883 7333
rect 6825 7293 6837 7327
rect 6871 7293 6883 7327
rect 6825 7287 6883 7293
rect 8168 7327 8226 7333
rect 8168 7293 8180 7327
rect 8214 7324 8226 7327
rect 8570 7324 8576 7336
rect 8214 7296 8576 7324
rect 8214 7293 8226 7296
rect 8168 7287 8226 7293
rect 4154 7216 4160 7268
rect 4212 7256 4218 7268
rect 4212 7228 4257 7256
rect 4212 7216 4218 7228
rect 5350 7216 5356 7268
rect 5408 7256 5414 7268
rect 6270 7256 6276 7268
rect 5408 7228 6276 7256
rect 5408 7216 5414 7228
rect 6270 7216 6276 7228
rect 6328 7256 6334 7268
rect 6549 7259 6607 7265
rect 6549 7256 6561 7259
rect 6328 7228 6561 7256
rect 6328 7216 6334 7228
rect 6549 7225 6561 7228
rect 6595 7256 6607 7259
rect 6840 7256 6868 7287
rect 8570 7284 8576 7296
rect 8628 7284 8634 7336
rect 8754 7284 8760 7336
rect 8812 7324 8818 7336
rect 12342 7324 12348 7336
rect 8812 7296 12348 7324
rect 8812 7284 8818 7296
rect 12342 7284 12348 7296
rect 12400 7324 12406 7336
rect 15095 7333 15108 7336
rect 12621 7327 12679 7333
rect 12621 7324 12633 7327
rect 12400 7296 12633 7324
rect 12400 7284 12406 7296
rect 12621 7293 12633 7296
rect 12667 7324 12679 7327
rect 13081 7327 13139 7333
rect 13081 7324 13093 7327
rect 12667 7296 13093 7324
rect 12667 7293 12679 7296
rect 12621 7287 12679 7293
rect 13081 7293 13093 7296
rect 13127 7293 13139 7327
rect 15080 7327 15108 7333
rect 15080 7324 15092 7327
rect 15015 7296 15092 7324
rect 13081 7287 13139 7293
rect 15080 7293 15092 7296
rect 15080 7287 15108 7293
rect 15102 7284 15108 7287
rect 15160 7284 15166 7336
rect 17788 7324 17816 7423
rect 18141 7327 18199 7333
rect 18141 7324 18153 7327
rect 17788 7296 18153 7324
rect 18141 7293 18153 7296
rect 18187 7293 18199 7327
rect 18141 7287 18199 7293
rect 24648 7327 24706 7333
rect 24648 7293 24660 7327
rect 24694 7324 24706 7327
rect 25130 7324 25136 7336
rect 24694 7296 25136 7324
rect 24694 7293 24706 7296
rect 24648 7287 24706 7293
rect 25130 7284 25136 7296
rect 25188 7284 25194 7336
rect 6595 7228 6868 7256
rect 6595 7225 6607 7228
rect 6549 7219 6607 7225
rect 7466 7216 7472 7268
rect 7524 7256 7530 7268
rect 8021 7259 8079 7265
rect 8021 7256 8033 7259
rect 7524 7228 8033 7256
rect 7524 7216 7530 7228
rect 8021 7225 8033 7228
rect 8067 7256 8079 7259
rect 8478 7256 8484 7268
rect 8067 7228 8484 7256
rect 8067 7225 8079 7228
rect 8021 7219 8079 7225
rect 8478 7216 8484 7228
rect 8536 7216 8542 7268
rect 8588 7256 8616 7284
rect 9214 7256 9220 7268
rect 8588 7228 9220 7256
rect 9214 7216 9220 7228
rect 9272 7216 9278 7268
rect 9582 7256 9588 7268
rect 9543 7228 9588 7256
rect 9582 7216 9588 7228
rect 9640 7256 9646 7268
rect 10965 7259 11023 7265
rect 10965 7256 10977 7259
rect 9640 7228 10977 7256
rect 9640 7216 9646 7228
rect 10965 7225 10977 7228
rect 11011 7225 11023 7259
rect 13354 7256 13360 7268
rect 13315 7228 13360 7256
rect 10965 7219 11023 7225
rect 13354 7216 13360 7228
rect 13412 7216 13418 7268
rect 13446 7216 13452 7268
rect 13504 7256 13510 7268
rect 16114 7256 16120 7268
rect 13504 7228 13549 7256
rect 16075 7228 16120 7256
rect 13504 7216 13510 7228
rect 16114 7216 16120 7228
rect 16172 7216 16178 7268
rect 16206 7216 16212 7268
rect 16264 7256 16270 7268
rect 18046 7256 18052 7268
rect 16264 7228 16309 7256
rect 18007 7228 18052 7256
rect 16264 7216 16270 7228
rect 18046 7216 18052 7228
rect 18104 7216 18110 7268
rect 2038 7148 2044 7200
rect 2096 7188 2102 7200
rect 2133 7191 2191 7197
rect 2133 7188 2145 7191
rect 2096 7160 2145 7188
rect 2096 7148 2102 7160
rect 2133 7157 2145 7160
rect 2179 7157 2191 7191
rect 2774 7188 2780 7200
rect 2735 7160 2780 7188
rect 2133 7151 2191 7157
rect 2774 7148 2780 7160
rect 2832 7148 2838 7200
rect 5442 7188 5448 7200
rect 5403 7160 5448 7188
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 6178 7188 6184 7200
rect 6139 7160 6184 7188
rect 6178 7148 6184 7160
rect 6236 7148 6242 7200
rect 7006 7188 7012 7200
rect 6967 7160 7012 7188
rect 7006 7148 7012 7160
rect 7064 7148 7070 7200
rect 9122 7188 9128 7200
rect 9083 7160 9128 7188
rect 9122 7148 9128 7160
rect 9180 7148 9186 7200
rect 9398 7188 9404 7200
rect 9359 7160 9404 7188
rect 9398 7148 9404 7160
rect 9456 7148 9462 7200
rect 11330 7188 11336 7200
rect 11291 7160 11336 7188
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 15151 7191 15209 7197
rect 15151 7157 15163 7191
rect 15197 7188 15209 7191
rect 15286 7188 15292 7200
rect 15197 7160 15292 7188
rect 15197 7157 15209 7160
rect 15151 7151 15209 7157
rect 15286 7148 15292 7160
rect 15344 7148 15350 7200
rect 15933 7191 15991 7197
rect 15933 7157 15945 7191
rect 15979 7188 15991 7191
rect 16224 7188 16252 7216
rect 15979 7160 16252 7188
rect 24719 7191 24777 7197
rect 15979 7157 15991 7160
rect 15933 7151 15991 7157
rect 24719 7157 24731 7191
rect 24765 7188 24777 7191
rect 25130 7188 25136 7200
rect 24765 7160 25136 7188
rect 24765 7157 24777 7160
rect 24719 7151 24777 7157
rect 25130 7148 25136 7160
rect 25188 7148 25194 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 2777 6987 2835 6993
rect 2777 6953 2789 6987
rect 2823 6984 2835 6987
rect 2958 6984 2964 6996
rect 2823 6956 2964 6984
rect 2823 6953 2835 6956
rect 2777 6947 2835 6953
rect 2958 6944 2964 6956
rect 3016 6944 3022 6996
rect 3145 6987 3203 6993
rect 3145 6953 3157 6987
rect 3191 6984 3203 6987
rect 3694 6984 3700 6996
rect 3191 6956 3700 6984
rect 3191 6953 3203 6956
rect 3145 6947 3203 6953
rect 3694 6944 3700 6956
rect 3752 6984 3758 6996
rect 3789 6987 3847 6993
rect 3789 6984 3801 6987
rect 3752 6956 3801 6984
rect 3752 6944 3758 6956
rect 3789 6953 3801 6956
rect 3835 6953 3847 6987
rect 3789 6947 3847 6953
rect 4246 6944 4252 6996
rect 4304 6984 4310 6996
rect 8846 6984 8852 6996
rect 4304 6956 8852 6984
rect 4304 6944 4310 6956
rect 8846 6944 8852 6956
rect 8904 6944 8910 6996
rect 8938 6944 8944 6996
rect 8996 6984 9002 6996
rect 9769 6987 9827 6993
rect 9769 6984 9781 6987
rect 8996 6956 9781 6984
rect 8996 6944 9002 6956
rect 9769 6953 9781 6956
rect 9815 6953 9827 6987
rect 9769 6947 9827 6953
rect 13173 6987 13231 6993
rect 13173 6953 13185 6987
rect 13219 6984 13231 6987
rect 13446 6984 13452 6996
rect 13219 6956 13452 6984
rect 13219 6953 13231 6956
rect 13173 6947 13231 6953
rect 13446 6944 13452 6956
rect 13504 6944 13510 6996
rect 15102 6984 15108 6996
rect 15063 6956 15108 6984
rect 15102 6944 15108 6956
rect 15160 6944 15166 6996
rect 16114 6944 16120 6996
rect 16172 6984 16178 6996
rect 16301 6987 16359 6993
rect 16301 6984 16313 6987
rect 16172 6956 16313 6984
rect 16172 6944 16178 6956
rect 16301 6953 16313 6956
rect 16347 6953 16359 6987
rect 16301 6947 16359 6953
rect 16482 6944 16488 6996
rect 16540 6984 16546 6996
rect 18509 6987 18567 6993
rect 18509 6984 18521 6987
rect 16540 6956 18521 6984
rect 16540 6944 16546 6956
rect 18509 6953 18521 6956
rect 18555 6953 18567 6987
rect 18509 6947 18567 6953
rect 3510 6916 3516 6928
rect 3471 6888 3516 6916
rect 3510 6876 3516 6888
rect 3568 6876 3574 6928
rect 5074 6916 5080 6928
rect 4356 6888 5080 6916
rect 2041 6851 2099 6857
rect 2041 6817 2053 6851
rect 2087 6848 2099 6851
rect 2222 6848 2228 6860
rect 2087 6820 2228 6848
rect 2087 6817 2099 6820
rect 2041 6811 2099 6817
rect 2222 6808 2228 6820
rect 2280 6808 2286 6860
rect 2961 6851 3019 6857
rect 2961 6817 2973 6851
rect 3007 6848 3019 6851
rect 3142 6848 3148 6860
rect 3007 6820 3148 6848
rect 3007 6817 3019 6820
rect 2961 6811 3019 6817
rect 3142 6808 3148 6820
rect 3200 6808 3206 6860
rect 3878 6808 3884 6860
rect 3936 6848 3942 6860
rect 4065 6851 4123 6857
rect 4065 6848 4077 6851
rect 3936 6820 4077 6848
rect 3936 6808 3942 6820
rect 4065 6817 4077 6820
rect 4111 6817 4123 6851
rect 4065 6811 4123 6817
rect 1854 6740 1860 6792
rect 1912 6780 1918 6792
rect 4356 6780 4384 6888
rect 5074 6876 5080 6888
rect 5132 6916 5138 6928
rect 6454 6916 6460 6928
rect 5132 6888 6460 6916
rect 5132 6876 5138 6888
rect 6454 6876 6460 6888
rect 6512 6876 6518 6928
rect 8754 6916 8760 6928
rect 8715 6888 8760 6916
rect 8754 6876 8760 6888
rect 8812 6876 8818 6928
rect 11057 6919 11115 6925
rect 11057 6916 11069 6919
rect 9692 6888 11069 6916
rect 9692 6860 9720 6888
rect 11057 6885 11069 6888
rect 11103 6885 11115 6919
rect 11057 6879 11115 6885
rect 12615 6919 12673 6925
rect 12615 6885 12627 6919
rect 12661 6916 12673 6919
rect 12710 6916 12716 6928
rect 12661 6888 12716 6916
rect 12661 6885 12673 6888
rect 12615 6879 12673 6885
rect 12710 6876 12716 6888
rect 12768 6876 12774 6928
rect 14550 6876 14556 6928
rect 14608 6916 14614 6928
rect 15473 6919 15531 6925
rect 15473 6916 15485 6919
rect 14608 6888 15485 6916
rect 14608 6876 14614 6888
rect 15473 6885 15485 6888
rect 15519 6916 15531 6919
rect 18046 6916 18052 6928
rect 15519 6888 18052 6916
rect 15519 6885 15531 6888
rect 15473 6879 15531 6885
rect 18046 6876 18052 6888
rect 18104 6876 18110 6928
rect 4614 6848 4620 6860
rect 4575 6820 4620 6848
rect 4614 6808 4620 6820
rect 4672 6808 4678 6860
rect 4982 6808 4988 6860
rect 5040 6848 5046 6860
rect 5040 6820 6408 6848
rect 5040 6808 5046 6820
rect 6380 6789 6408 6820
rect 7742 6808 7748 6860
rect 7800 6848 7806 6860
rect 8021 6851 8079 6857
rect 8021 6848 8033 6851
rect 7800 6820 8033 6848
rect 7800 6808 7806 6820
rect 8021 6817 8033 6820
rect 8067 6817 8079 6851
rect 8021 6811 8079 6817
rect 8110 6808 8116 6860
rect 8168 6857 8174 6860
rect 8168 6851 8226 6857
rect 8168 6817 8180 6851
rect 8214 6848 8226 6851
rect 9490 6848 9496 6860
rect 8214 6820 9496 6848
rect 8214 6817 8226 6820
rect 8168 6811 8226 6817
rect 8168 6808 8174 6811
rect 9490 6808 9496 6820
rect 9548 6808 9554 6860
rect 9674 6848 9680 6860
rect 9635 6820 9680 6848
rect 9674 6808 9680 6820
rect 9732 6808 9738 6860
rect 10137 6851 10195 6857
rect 10137 6817 10149 6851
rect 10183 6817 10195 6851
rect 11238 6848 11244 6860
rect 11199 6820 11244 6848
rect 10137 6811 10195 6817
rect 1912 6752 4384 6780
rect 4433 6783 4491 6789
rect 1912 6740 1918 6752
rect 4433 6749 4445 6783
rect 4479 6780 4491 6783
rect 6365 6783 6423 6789
rect 4479 6752 5580 6780
rect 4479 6749 4491 6752
rect 4433 6743 4491 6749
rect 5552 6656 5580 6752
rect 6365 6749 6377 6783
rect 6411 6780 6423 6783
rect 6825 6783 6883 6789
rect 6825 6780 6837 6783
rect 6411 6752 6837 6780
rect 6411 6749 6423 6752
rect 6365 6743 6423 6749
rect 6825 6749 6837 6752
rect 6871 6780 6883 6783
rect 7006 6780 7012 6792
rect 6871 6752 7012 6780
rect 6871 6749 6883 6752
rect 6825 6743 6883 6749
rect 7006 6740 7012 6752
rect 7064 6740 7070 6792
rect 7558 6740 7564 6792
rect 7616 6780 7622 6792
rect 8389 6783 8447 6789
rect 8389 6780 8401 6783
rect 7616 6752 8401 6780
rect 7616 6740 7622 6752
rect 8389 6749 8401 6752
rect 8435 6749 8447 6783
rect 10042 6780 10048 6792
rect 8389 6743 8447 6749
rect 9600 6752 10048 6780
rect 5994 6712 6000 6724
rect 5907 6684 6000 6712
rect 5994 6672 6000 6684
rect 6052 6712 6058 6724
rect 6730 6712 6736 6724
rect 6052 6684 6647 6712
rect 6691 6684 6736 6712
rect 6052 6672 6058 6684
rect 1670 6644 1676 6656
rect 1631 6616 1676 6644
rect 1670 6604 1676 6616
rect 1728 6604 1734 6656
rect 5261 6647 5319 6653
rect 5261 6613 5273 6647
rect 5307 6644 5319 6647
rect 5442 6644 5448 6656
rect 5307 6616 5448 6644
rect 5307 6613 5319 6616
rect 5261 6607 5319 6613
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 5534 6604 5540 6656
rect 5592 6644 5598 6656
rect 6619 6653 6647 6684
rect 6730 6672 6736 6684
rect 6788 6672 6794 6724
rect 7101 6715 7159 6721
rect 7101 6681 7113 6715
rect 7147 6712 7159 6715
rect 9600 6712 9628 6752
rect 10042 6740 10048 6752
rect 10100 6780 10106 6792
rect 10152 6780 10180 6811
rect 11238 6808 11244 6820
rect 11296 6808 11302 6860
rect 11330 6808 11336 6860
rect 11388 6848 11394 6860
rect 11388 6820 15056 6848
rect 11388 6808 11394 6820
rect 11701 6783 11759 6789
rect 11701 6780 11713 6783
rect 10100 6752 11713 6780
rect 10100 6740 10106 6752
rect 11701 6749 11713 6752
rect 11747 6749 11759 6783
rect 12250 6780 12256 6792
rect 12211 6752 12256 6780
rect 11701 6743 11759 6749
rect 12250 6740 12256 6752
rect 12308 6740 12314 6792
rect 14185 6783 14243 6789
rect 14185 6749 14197 6783
rect 14231 6780 14243 6783
rect 14642 6780 14648 6792
rect 14231 6752 14648 6780
rect 14231 6749 14243 6752
rect 14185 6743 14243 6749
rect 14642 6740 14648 6752
rect 14700 6740 14706 6792
rect 15028 6780 15056 6820
rect 16206 6808 16212 6860
rect 16264 6848 16270 6860
rect 16853 6851 16911 6857
rect 16853 6848 16865 6851
rect 16264 6820 16865 6848
rect 16264 6808 16270 6820
rect 16853 6817 16865 6820
rect 16899 6817 16911 6851
rect 18414 6848 18420 6860
rect 18375 6820 18420 6848
rect 16853 6811 16911 6817
rect 18414 6808 18420 6820
rect 18472 6808 18478 6860
rect 18874 6848 18880 6860
rect 18835 6820 18880 6848
rect 18874 6808 18880 6820
rect 18932 6808 18938 6860
rect 23198 6808 23204 6860
rect 23256 6848 23262 6860
rect 23753 6851 23811 6857
rect 23753 6848 23765 6851
rect 23256 6820 23765 6848
rect 23256 6808 23262 6820
rect 23753 6817 23765 6820
rect 23799 6817 23811 6851
rect 23753 6811 23811 6817
rect 15378 6780 15384 6792
rect 15028 6752 15384 6780
rect 15378 6740 15384 6752
rect 15436 6740 15442 6792
rect 15657 6783 15715 6789
rect 15657 6749 15669 6783
rect 15703 6749 15715 6783
rect 15657 6743 15715 6749
rect 17221 6783 17279 6789
rect 17221 6749 17233 6783
rect 17267 6780 17279 6783
rect 17494 6780 17500 6792
rect 17267 6752 17500 6780
rect 17267 6749 17279 6752
rect 17221 6743 17279 6749
rect 7147 6684 9628 6712
rect 7147 6681 7159 6684
rect 7101 6675 7159 6681
rect 13446 6672 13452 6724
rect 13504 6712 13510 6724
rect 13817 6715 13875 6721
rect 13817 6712 13829 6715
rect 13504 6684 13829 6712
rect 13504 6672 13510 6684
rect 13817 6681 13829 6684
rect 13863 6681 13875 6715
rect 13817 6675 13875 6681
rect 13998 6672 14004 6724
rect 14056 6712 14062 6724
rect 15672 6712 15700 6743
rect 17494 6740 17500 6752
rect 17552 6740 17558 6792
rect 17589 6783 17647 6789
rect 17589 6749 17601 6783
rect 17635 6780 17647 6783
rect 18141 6783 18199 6789
rect 18141 6780 18153 6783
rect 17635 6752 18153 6780
rect 17635 6749 17647 6752
rect 17589 6743 17647 6749
rect 18141 6749 18153 6752
rect 18187 6780 18199 6783
rect 18892 6780 18920 6808
rect 18187 6752 18920 6780
rect 18187 6749 18199 6752
rect 18141 6743 18199 6749
rect 14056 6684 15700 6712
rect 15764 6684 16896 6712
rect 14056 6672 14062 6684
rect 6619 6647 6680 6653
rect 5592 6616 5637 6644
rect 6619 6616 6634 6647
rect 5592 6604 5598 6616
rect 6622 6613 6634 6616
rect 6668 6644 6680 6647
rect 7006 6644 7012 6656
rect 6668 6616 7012 6644
rect 6668 6613 6680 6616
rect 6622 6607 6680 6613
rect 7006 6604 7012 6616
rect 7064 6604 7070 6656
rect 7653 6647 7711 6653
rect 7653 6613 7665 6647
rect 7699 6644 7711 6647
rect 7742 6644 7748 6656
rect 7699 6616 7748 6644
rect 7699 6613 7711 6616
rect 7653 6607 7711 6613
rect 7742 6604 7748 6616
rect 7800 6604 7806 6656
rect 8294 6644 8300 6656
rect 8255 6616 8300 6644
rect 8294 6604 8300 6616
rect 8352 6604 8358 6656
rect 8570 6604 8576 6656
rect 8628 6644 8634 6656
rect 9033 6647 9091 6653
rect 9033 6644 9045 6647
rect 8628 6616 9045 6644
rect 8628 6604 8634 6616
rect 9033 6613 9045 6616
rect 9079 6613 9091 6647
rect 9033 6607 9091 6613
rect 9306 6604 9312 6656
rect 9364 6644 9370 6656
rect 9401 6647 9459 6653
rect 9401 6644 9413 6647
rect 9364 6616 9413 6644
rect 9364 6604 9370 6616
rect 9401 6613 9413 6616
rect 9447 6613 9459 6647
rect 9401 6607 9459 6613
rect 9490 6604 9496 6656
rect 9548 6644 9554 6656
rect 10689 6647 10747 6653
rect 10689 6644 10701 6647
rect 9548 6616 10701 6644
rect 9548 6604 9554 6616
rect 10689 6613 10701 6616
rect 10735 6613 10747 6647
rect 10689 6607 10747 6613
rect 10778 6604 10784 6656
rect 10836 6644 10842 6656
rect 11425 6647 11483 6653
rect 11425 6644 11437 6647
rect 10836 6616 11437 6644
rect 10836 6604 10842 6616
rect 11425 6613 11437 6616
rect 11471 6644 11483 6647
rect 15764 6644 15792 6684
rect 16868 6656 16896 6684
rect 16758 6644 16764 6656
rect 11471 6616 15792 6644
rect 16719 6616 16764 6644
rect 11471 6613 11483 6616
rect 11425 6607 11483 6613
rect 16758 6604 16764 6616
rect 16816 6604 16822 6656
rect 16850 6604 16856 6656
rect 16908 6644 16914 6656
rect 16991 6647 17049 6653
rect 16991 6644 17003 6647
rect 16908 6616 17003 6644
rect 16908 6604 16914 6616
rect 16991 6613 17003 6616
rect 17037 6613 17049 6647
rect 16991 6607 17049 6613
rect 17129 6647 17187 6653
rect 17129 6613 17141 6647
rect 17175 6644 17187 6647
rect 17218 6644 17224 6656
rect 17175 6616 17224 6644
rect 17175 6613 17187 6616
rect 17129 6607 17187 6613
rect 17218 6604 17224 6616
rect 17276 6604 17282 6656
rect 23934 6644 23940 6656
rect 23895 6616 23940 6644
rect 23934 6604 23940 6616
rect 23992 6604 23998 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 5334 6443 5392 6449
rect 5334 6409 5346 6443
rect 5380 6440 5392 6443
rect 5534 6440 5540 6452
rect 5380 6412 5540 6440
rect 5380 6409 5392 6412
rect 5334 6403 5392 6409
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 5813 6443 5871 6449
rect 5813 6409 5825 6443
rect 5859 6440 5871 6443
rect 6362 6440 6368 6452
rect 5859 6412 6368 6440
rect 5859 6409 5871 6412
rect 5813 6403 5871 6409
rect 6362 6400 6368 6412
rect 6420 6400 6426 6452
rect 6549 6443 6607 6449
rect 6549 6409 6561 6443
rect 6595 6440 6607 6443
rect 6730 6440 6736 6452
rect 6595 6412 6736 6440
rect 6595 6409 6607 6412
rect 6549 6403 6607 6409
rect 6730 6400 6736 6412
rect 6788 6400 6794 6452
rect 7558 6440 7564 6452
rect 7519 6412 7564 6440
rect 7558 6400 7564 6412
rect 7616 6440 7622 6452
rect 7837 6443 7895 6449
rect 7837 6440 7849 6443
rect 7616 6412 7849 6440
rect 7616 6400 7622 6412
rect 7837 6409 7849 6412
rect 7883 6409 7895 6443
rect 8294 6440 8300 6452
rect 8207 6412 8300 6440
rect 7837 6403 7895 6409
rect 5442 6332 5448 6384
rect 5500 6372 5506 6384
rect 6914 6372 6920 6384
rect 5500 6344 6920 6372
rect 5500 6332 5506 6344
rect 6914 6332 6920 6344
rect 6972 6332 6978 6384
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6304 2283 6307
rect 2406 6304 2412 6316
rect 2271 6276 2412 6304
rect 2271 6273 2283 6276
rect 2225 6267 2283 6273
rect 2406 6264 2412 6276
rect 2464 6264 2470 6316
rect 4706 6304 4712 6316
rect 3436 6276 4712 6304
rect 2961 6239 3019 6245
rect 2961 6205 2973 6239
rect 3007 6236 3019 6239
rect 3234 6236 3240 6248
rect 3007 6208 3240 6236
rect 3007 6205 3019 6208
rect 2961 6199 3019 6205
rect 3234 6196 3240 6208
rect 3292 6196 3298 6248
rect 1578 6168 1584 6180
rect 1539 6140 1584 6168
rect 1578 6128 1584 6140
rect 1636 6128 1642 6180
rect 1670 6128 1676 6180
rect 1728 6168 1734 6180
rect 3436 6168 3464 6276
rect 4706 6264 4712 6276
rect 4764 6264 4770 6316
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6273 5595 6307
rect 7852 6304 7880 6403
rect 8294 6400 8300 6412
rect 8352 6440 8358 6452
rect 9122 6440 9128 6452
rect 8352 6412 9128 6440
rect 8352 6400 8358 6412
rect 9122 6400 9128 6412
rect 9180 6400 9186 6452
rect 9306 6400 9312 6452
rect 9364 6440 9370 6452
rect 9861 6443 9919 6449
rect 9861 6440 9873 6443
rect 9364 6412 9873 6440
rect 9364 6400 9370 6412
rect 9861 6409 9873 6412
rect 9907 6440 9919 6443
rect 9950 6440 9956 6452
rect 9907 6412 9956 6440
rect 9907 6409 9919 6412
rect 9861 6403 9919 6409
rect 9950 6400 9956 6412
rect 10008 6400 10014 6452
rect 10686 6440 10692 6452
rect 10647 6412 10692 6440
rect 10686 6400 10692 6412
rect 10744 6400 10750 6452
rect 12253 6443 12311 6449
rect 12253 6409 12265 6443
rect 12299 6440 12311 6443
rect 12710 6440 12716 6452
rect 12299 6412 12716 6440
rect 12299 6409 12311 6412
rect 12253 6403 12311 6409
rect 12710 6400 12716 6412
rect 12768 6400 12774 6452
rect 14550 6440 14556 6452
rect 14511 6412 14556 6440
rect 14550 6400 14556 6412
rect 14608 6400 14614 6452
rect 16669 6443 16727 6449
rect 16669 6409 16681 6443
rect 16715 6440 16727 6443
rect 16850 6440 16856 6452
rect 16715 6412 16856 6440
rect 16715 6409 16727 6412
rect 16669 6403 16727 6409
rect 16850 6400 16856 6412
rect 16908 6400 16914 6452
rect 17218 6440 17224 6452
rect 17179 6412 17224 6440
rect 17218 6400 17224 6412
rect 17276 6400 17282 6452
rect 18414 6400 18420 6452
rect 18472 6440 18478 6452
rect 19061 6443 19119 6449
rect 19061 6440 19073 6443
rect 18472 6412 19073 6440
rect 18472 6400 18478 6412
rect 19061 6409 19073 6412
rect 19107 6409 19119 6443
rect 23934 6440 23940 6452
rect 23895 6412 23940 6440
rect 19061 6403 19119 6409
rect 23934 6400 23940 6412
rect 23992 6400 23998 6452
rect 25130 6440 25136 6452
rect 25091 6412 25136 6440
rect 25130 6400 25136 6412
rect 25188 6400 25194 6452
rect 8110 6332 8116 6384
rect 8168 6381 8174 6384
rect 8168 6375 8217 6381
rect 8168 6341 8171 6375
rect 8205 6341 8217 6375
rect 8168 6335 8217 6341
rect 8168 6332 8174 6335
rect 8478 6332 8484 6384
rect 8536 6372 8542 6384
rect 9674 6372 9680 6384
rect 8536 6344 9680 6372
rect 8536 6332 8542 6344
rect 9674 6332 9680 6344
rect 9732 6332 9738 6384
rect 11333 6375 11391 6381
rect 11333 6372 11345 6375
rect 10060 6344 11345 6372
rect 10060 6316 10088 6344
rect 11333 6341 11345 6344
rect 11379 6341 11391 6375
rect 11333 6335 11391 6341
rect 8389 6307 8447 6313
rect 8389 6304 8401 6307
rect 7852 6276 8401 6304
rect 5537 6267 5595 6273
rect 8389 6273 8401 6276
rect 8435 6304 8447 6307
rect 9398 6304 9404 6316
rect 8435 6276 9404 6304
rect 8435 6273 8447 6276
rect 8389 6267 8447 6273
rect 3694 6236 3700 6248
rect 3655 6208 3700 6236
rect 3694 6196 3700 6208
rect 3752 6196 3758 6248
rect 3881 6239 3939 6245
rect 3881 6205 3893 6239
rect 3927 6236 3939 6239
rect 3970 6236 3976 6248
rect 3927 6208 3976 6236
rect 3927 6205 3939 6208
rect 3881 6199 3939 6205
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 5350 6196 5356 6248
rect 5408 6236 5414 6248
rect 5552 6236 5580 6267
rect 9398 6264 9404 6276
rect 9456 6304 9462 6316
rect 9953 6307 10011 6313
rect 9953 6304 9965 6307
rect 9456 6276 9965 6304
rect 9456 6264 9462 6276
rect 9953 6273 9965 6276
rect 9999 6304 10011 6307
rect 10042 6304 10048 6316
rect 9999 6276 10048 6304
rect 9999 6273 10011 6276
rect 9953 6267 10011 6273
rect 10042 6264 10048 6276
rect 10100 6264 10106 6316
rect 15013 6307 15071 6313
rect 15013 6273 15025 6307
rect 15059 6304 15071 6307
rect 15102 6304 15108 6316
rect 15059 6276 15108 6304
rect 15059 6273 15071 6276
rect 15013 6267 15071 6273
rect 15102 6264 15108 6276
rect 15160 6304 15166 6316
rect 18509 6307 18567 6313
rect 18509 6304 18521 6307
rect 15160 6276 18521 6304
rect 15160 6264 15166 6276
rect 18509 6273 18521 6276
rect 18555 6273 18567 6307
rect 18509 6267 18567 6273
rect 24213 6307 24271 6313
rect 24213 6273 24225 6307
rect 24259 6304 24271 6307
rect 25148 6304 25176 6400
rect 24259 6276 25176 6304
rect 24259 6273 24271 6276
rect 24213 6267 24271 6273
rect 5408 6208 5580 6236
rect 5408 6196 5414 6208
rect 5626 6196 5632 6248
rect 5684 6236 5690 6248
rect 6825 6239 6883 6245
rect 6825 6236 6837 6239
rect 5684 6208 6837 6236
rect 5684 6196 5690 6208
rect 6825 6205 6837 6208
rect 6871 6205 6883 6239
rect 9582 6236 9588 6248
rect 9543 6208 9588 6236
rect 6825 6199 6883 6205
rect 9582 6196 9588 6208
rect 9640 6196 9646 6248
rect 9766 6245 9772 6248
rect 9732 6239 9772 6245
rect 9732 6205 9744 6239
rect 9824 6236 9830 6248
rect 10686 6236 10692 6248
rect 9824 6208 10692 6236
rect 9732 6199 9772 6205
rect 9766 6196 9772 6199
rect 9824 6196 9830 6208
rect 10686 6196 10692 6208
rect 10744 6196 10750 6248
rect 11146 6236 11152 6248
rect 11107 6208 11152 6236
rect 11146 6196 11152 6208
rect 11204 6236 11210 6248
rect 11609 6239 11667 6245
rect 11609 6236 11621 6239
rect 11204 6208 11621 6236
rect 11204 6196 11210 6208
rect 11609 6205 11621 6208
rect 11655 6205 11667 6239
rect 11609 6199 11667 6205
rect 12437 6239 12495 6245
rect 12437 6205 12449 6239
rect 12483 6236 12495 6239
rect 13633 6239 13691 6245
rect 13633 6236 13645 6239
rect 12483 6208 13645 6236
rect 12483 6205 12495 6208
rect 12437 6199 12495 6205
rect 13633 6205 13645 6208
rect 13679 6236 13691 6239
rect 16482 6236 16488 6248
rect 13679 6208 16488 6236
rect 13679 6205 13691 6208
rect 13633 6199 13691 6205
rect 16482 6196 16488 6208
rect 16540 6196 16546 6248
rect 16758 6236 16764 6248
rect 16722 6208 16764 6236
rect 16758 6196 16764 6208
rect 16816 6245 16822 6248
rect 16816 6239 16870 6245
rect 16816 6205 16824 6239
rect 16858 6236 16870 6239
rect 17126 6236 17132 6248
rect 16858 6208 17132 6236
rect 16858 6205 16870 6208
rect 16816 6199 16870 6205
rect 16816 6196 16822 6199
rect 17126 6196 17132 6208
rect 17184 6196 17190 6248
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 17788 6208 18061 6236
rect 1728 6140 1773 6168
rect 2424 6140 3464 6168
rect 1728 6128 1734 6140
rect 1596 6100 1624 6128
rect 2424 6100 2452 6140
rect 3510 6128 3516 6180
rect 3568 6168 3574 6180
rect 5077 6171 5135 6177
rect 5077 6168 5089 6171
rect 3568 6140 5089 6168
rect 3568 6128 3574 6140
rect 5077 6137 5089 6140
rect 5123 6168 5135 6171
rect 5169 6171 5227 6177
rect 5169 6168 5181 6171
rect 5123 6140 5181 6168
rect 5123 6137 5135 6140
rect 5077 6131 5135 6137
rect 5169 6137 5181 6140
rect 5215 6168 5227 6171
rect 7742 6168 7748 6180
rect 5215 6140 7748 6168
rect 5215 6137 5227 6140
rect 5169 6131 5227 6137
rect 7742 6128 7748 6140
rect 7800 6128 7806 6180
rect 8018 6168 8024 6180
rect 7979 6140 8024 6168
rect 8018 6128 8024 6140
rect 8076 6168 8082 6180
rect 8570 6168 8576 6180
rect 8076 6140 8576 6168
rect 8076 6128 8082 6140
rect 8570 6128 8576 6140
rect 8628 6128 8634 6180
rect 8754 6168 8760 6180
rect 8715 6140 8760 6168
rect 8754 6128 8760 6140
rect 8812 6128 8818 6180
rect 9306 6128 9312 6180
rect 9364 6168 9370 6180
rect 10965 6171 11023 6177
rect 10965 6168 10977 6171
rect 9364 6140 10977 6168
rect 9364 6128 9370 6140
rect 10965 6137 10977 6140
rect 11011 6168 11023 6171
rect 11238 6168 11244 6180
rect 11011 6140 11244 6168
rect 11011 6137 11023 6140
rect 10965 6131 11023 6137
rect 11238 6128 11244 6140
rect 11296 6128 11302 6180
rect 14734 6168 14740 6180
rect 12820 6140 14740 6168
rect 1596 6072 2452 6100
rect 2593 6103 2651 6109
rect 2593 6069 2605 6103
rect 2639 6100 2651 6103
rect 3970 6100 3976 6112
rect 2639 6072 3976 6100
rect 2639 6069 2651 6072
rect 2593 6063 2651 6069
rect 3970 6060 3976 6072
rect 4028 6060 4034 6112
rect 4062 6060 4068 6112
rect 4120 6100 4126 6112
rect 4157 6103 4215 6109
rect 4157 6100 4169 6103
rect 4120 6072 4169 6100
rect 4120 6060 4126 6072
rect 4157 6069 4169 6072
rect 4203 6069 4215 6103
rect 4157 6063 4215 6069
rect 4525 6103 4583 6109
rect 4525 6069 4537 6103
rect 4571 6100 4583 6103
rect 4614 6100 4620 6112
rect 4571 6072 4620 6100
rect 4571 6069 4583 6072
rect 4525 6063 4583 6069
rect 4614 6060 4620 6072
rect 4672 6100 4678 6112
rect 4890 6100 4896 6112
rect 4672 6072 4896 6100
rect 4672 6060 4678 6072
rect 4890 6060 4896 6072
rect 4948 6100 4954 6112
rect 6178 6100 6184 6112
rect 4948 6072 6184 6100
rect 4948 6060 4954 6072
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 7006 6100 7012 6112
rect 6919 6072 7012 6100
rect 7006 6060 7012 6072
rect 7064 6100 7070 6112
rect 8110 6100 8116 6112
rect 7064 6072 8116 6100
rect 7064 6060 7070 6072
rect 8110 6060 8116 6072
rect 8168 6060 8174 6112
rect 8202 6060 8208 6112
rect 8260 6100 8266 6112
rect 10229 6103 10287 6109
rect 10229 6100 10241 6103
rect 8260 6072 10241 6100
rect 8260 6060 8266 6072
rect 10229 6069 10241 6072
rect 10275 6069 10287 6103
rect 10229 6063 10287 6069
rect 12710 6060 12716 6112
rect 12768 6100 12774 6112
rect 12820 6109 12848 6140
rect 14734 6128 14740 6140
rect 14792 6168 14798 6180
rect 14829 6171 14887 6177
rect 14829 6168 14841 6171
rect 14792 6140 14841 6168
rect 14792 6128 14798 6140
rect 14829 6137 14841 6140
rect 14875 6168 14887 6171
rect 15334 6171 15392 6177
rect 15334 6168 15346 6171
rect 14875 6140 15346 6168
rect 14875 6137 14887 6140
rect 14829 6131 14887 6137
rect 15334 6137 15346 6140
rect 15380 6137 15392 6171
rect 15334 6131 15392 6137
rect 15470 6128 15476 6180
rect 15528 6168 15534 6180
rect 16899 6171 16957 6177
rect 16899 6168 16911 6171
rect 15528 6140 16911 6168
rect 15528 6128 15534 6140
rect 16899 6137 16911 6140
rect 16945 6137 16957 6171
rect 16899 6131 16957 6137
rect 12805 6103 12863 6109
rect 12805 6100 12817 6103
rect 12768 6072 12817 6100
rect 12768 6060 12774 6072
rect 12805 6069 12817 6072
rect 12851 6069 12863 6103
rect 13354 6100 13360 6112
rect 13315 6072 13360 6100
rect 12805 6063 12863 6069
rect 13354 6060 13360 6072
rect 13412 6060 13418 6112
rect 13998 6100 14004 6112
rect 13959 6072 14004 6100
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 15930 6100 15936 6112
rect 15891 6072 15936 6100
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 16206 6100 16212 6112
rect 16167 6072 16212 6100
rect 16206 6060 16212 6072
rect 16264 6060 16270 6112
rect 17034 6060 17040 6112
rect 17092 6100 17098 6112
rect 17788 6109 17816 6208
rect 18049 6205 18061 6208
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 18601 6239 18659 6245
rect 18601 6205 18613 6239
rect 18647 6236 18659 6239
rect 18874 6236 18880 6248
rect 18647 6208 18880 6236
rect 18647 6205 18659 6208
rect 18601 6199 18659 6205
rect 18874 6196 18880 6208
rect 18932 6236 18938 6248
rect 19429 6239 19487 6245
rect 19429 6236 19441 6239
rect 18932 6208 19441 6236
rect 18932 6196 18938 6208
rect 19429 6205 19441 6208
rect 19475 6205 19487 6239
rect 19429 6199 19487 6205
rect 24305 6171 24363 6177
rect 24305 6137 24317 6171
rect 24351 6137 24363 6171
rect 24854 6168 24860 6180
rect 24815 6140 24860 6168
rect 24305 6131 24363 6137
rect 17773 6103 17831 6109
rect 17773 6100 17785 6103
rect 17092 6072 17785 6100
rect 17092 6060 17098 6072
rect 17773 6069 17785 6072
rect 17819 6069 17831 6103
rect 17773 6063 17831 6069
rect 23198 6060 23204 6112
rect 23256 6100 23262 6112
rect 23385 6103 23443 6109
rect 23385 6100 23397 6103
rect 23256 6072 23397 6100
rect 23256 6060 23262 6072
rect 23385 6069 23397 6072
rect 23431 6069 23443 6103
rect 23385 6063 23443 6069
rect 23934 6060 23940 6112
rect 23992 6100 23998 6112
rect 24320 6100 24348 6131
rect 24854 6128 24860 6140
rect 24912 6128 24918 6180
rect 23992 6072 24348 6100
rect 23992 6060 23998 6072
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1670 5856 1676 5908
rect 1728 5896 1734 5908
rect 1857 5899 1915 5905
rect 1857 5896 1869 5899
rect 1728 5868 1869 5896
rect 1728 5856 1734 5868
rect 1857 5865 1869 5868
rect 1903 5865 1915 5899
rect 2222 5896 2228 5908
rect 2183 5868 2228 5896
rect 1857 5859 1915 5865
rect 2222 5856 2228 5868
rect 2280 5856 2286 5908
rect 3510 5896 3516 5908
rect 2516 5868 3516 5896
rect 2516 5828 2544 5868
rect 3510 5856 3516 5868
rect 3568 5856 3574 5908
rect 3878 5896 3884 5908
rect 3839 5868 3884 5896
rect 3878 5856 3884 5868
rect 3936 5856 3942 5908
rect 5813 5899 5871 5905
rect 5813 5865 5825 5899
rect 5859 5896 5871 5899
rect 5994 5896 6000 5908
rect 5859 5868 6000 5896
rect 5859 5865 5871 5868
rect 5813 5859 5871 5865
rect 5994 5856 6000 5868
rect 6052 5856 6058 5908
rect 6454 5856 6460 5908
rect 6512 5896 6518 5908
rect 7285 5899 7343 5905
rect 7285 5896 7297 5899
rect 6512 5868 7297 5896
rect 6512 5856 6518 5868
rect 7285 5865 7297 5868
rect 7331 5896 7343 5899
rect 8018 5896 8024 5908
rect 7331 5868 8024 5896
rect 7331 5865 7343 5868
rect 7285 5859 7343 5865
rect 8018 5856 8024 5868
rect 8076 5856 8082 5908
rect 8754 5856 8760 5908
rect 8812 5896 8818 5908
rect 11149 5899 11207 5905
rect 11149 5896 11161 5899
rect 8812 5868 11161 5896
rect 8812 5856 8818 5868
rect 11149 5865 11161 5868
rect 11195 5896 11207 5899
rect 11238 5896 11244 5908
rect 11195 5868 11244 5896
rect 11195 5865 11207 5868
rect 11149 5859 11207 5865
rect 11238 5856 11244 5868
rect 11296 5856 11302 5908
rect 11606 5856 11612 5908
rect 11664 5896 11670 5908
rect 12529 5899 12587 5905
rect 12529 5896 12541 5899
rect 11664 5868 12541 5896
rect 11664 5856 11670 5868
rect 12529 5865 12541 5868
rect 12575 5896 12587 5899
rect 12710 5896 12716 5908
rect 12575 5868 12716 5896
rect 12575 5865 12587 5868
rect 12529 5859 12587 5865
rect 12710 5856 12716 5868
rect 12768 5856 12774 5908
rect 15102 5896 15108 5908
rect 15063 5868 15108 5896
rect 15102 5856 15108 5868
rect 15160 5856 15166 5908
rect 15378 5856 15384 5908
rect 15436 5896 15442 5908
rect 15933 5899 15991 5905
rect 15933 5896 15945 5899
rect 15436 5868 15945 5896
rect 15436 5856 15442 5868
rect 15933 5865 15945 5868
rect 15979 5865 15991 5899
rect 15933 5859 15991 5865
rect 1780 5800 2544 5828
rect 2593 5831 2651 5837
rect 1780 5772 1808 5800
rect 2593 5797 2605 5831
rect 2639 5828 2651 5831
rect 2866 5828 2872 5840
rect 2639 5800 2872 5828
rect 2639 5797 2651 5800
rect 2593 5791 2651 5797
rect 2866 5788 2872 5800
rect 2924 5828 2930 5840
rect 2924 5800 3188 5828
rect 2924 5788 2930 5800
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5760 1455 5763
rect 1762 5760 1768 5772
rect 1443 5732 1768 5760
rect 1443 5729 1455 5732
rect 1397 5723 1455 5729
rect 1762 5720 1768 5732
rect 1820 5720 1826 5772
rect 3160 5760 3188 5800
rect 3418 5788 3424 5840
rect 3476 5828 3482 5840
rect 4338 5828 4344 5840
rect 3476 5800 4344 5828
rect 3476 5788 3482 5800
rect 4338 5788 4344 5800
rect 4396 5837 4402 5840
rect 4396 5831 4444 5837
rect 4396 5797 4398 5831
rect 4432 5797 4444 5831
rect 8202 5828 8208 5840
rect 4396 5791 4444 5797
rect 6748 5800 8208 5828
rect 4396 5788 4402 5791
rect 4522 5760 4528 5772
rect 3160 5732 4528 5760
rect 4522 5720 4528 5732
rect 4580 5760 4586 5772
rect 4985 5763 5043 5769
rect 4985 5760 4997 5763
rect 4580 5732 4997 5760
rect 4580 5720 4586 5732
rect 4985 5729 4997 5732
rect 5031 5729 5043 5763
rect 6362 5760 6368 5772
rect 6323 5732 6368 5760
rect 4985 5723 5043 5729
rect 6362 5720 6368 5732
rect 6420 5720 6426 5772
rect 6454 5720 6460 5772
rect 6512 5760 6518 5772
rect 6748 5769 6776 5800
rect 8202 5788 8208 5800
rect 8260 5788 8266 5840
rect 9490 5828 9496 5840
rect 9451 5800 9496 5828
rect 9490 5788 9496 5800
rect 9548 5788 9554 5840
rect 11256 5828 11284 5856
rect 12161 5831 12219 5837
rect 11256 5800 11928 5828
rect 6733 5763 6791 5769
rect 6733 5760 6745 5763
rect 6512 5732 6745 5760
rect 6512 5720 6518 5732
rect 6733 5729 6745 5732
rect 6779 5729 6791 5763
rect 6733 5723 6791 5729
rect 7742 5720 7748 5772
rect 7800 5760 7806 5772
rect 7837 5763 7895 5769
rect 7837 5760 7849 5763
rect 7800 5732 7849 5760
rect 7800 5720 7806 5732
rect 7837 5729 7849 5732
rect 7883 5729 7895 5763
rect 7837 5723 7895 5729
rect 7926 5720 7932 5772
rect 7984 5769 7990 5772
rect 7984 5763 8042 5769
rect 7984 5729 7996 5763
rect 8030 5760 8042 5763
rect 8110 5760 8116 5772
rect 8030 5732 8116 5760
rect 8030 5729 8042 5732
rect 7984 5723 8042 5729
rect 7984 5720 7990 5723
rect 8110 5720 8116 5732
rect 8168 5720 8174 5772
rect 9674 5760 9680 5772
rect 9587 5732 9680 5760
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 9766 5720 9772 5772
rect 9824 5769 9830 5772
rect 11900 5769 11928 5800
rect 12161 5797 12173 5831
rect 12207 5828 12219 5831
rect 12250 5828 12256 5840
rect 12207 5800 12256 5828
rect 12207 5797 12219 5800
rect 12161 5791 12219 5797
rect 12250 5788 12256 5800
rect 12308 5828 12314 5840
rect 12805 5831 12863 5837
rect 12805 5828 12817 5831
rect 12308 5800 12817 5828
rect 12308 5788 12314 5800
rect 12805 5797 12817 5800
rect 12851 5797 12863 5831
rect 16666 5828 16672 5840
rect 16627 5800 16672 5828
rect 12805 5791 12863 5797
rect 16666 5788 16672 5800
rect 16724 5788 16730 5840
rect 17770 5788 17776 5840
rect 17828 5828 17834 5840
rect 18233 5831 18291 5837
rect 18233 5828 18245 5831
rect 17828 5800 18245 5828
rect 17828 5788 17834 5800
rect 18233 5797 18245 5800
rect 18279 5797 18291 5831
rect 18233 5791 18291 5797
rect 23198 5788 23204 5840
rect 23256 5828 23262 5840
rect 24213 5831 24271 5837
rect 24213 5828 24225 5831
rect 23256 5800 24225 5828
rect 23256 5788 23262 5800
rect 24213 5797 24225 5800
rect 24259 5797 24271 5831
rect 24213 5791 24271 5797
rect 9824 5763 9882 5769
rect 9824 5729 9836 5763
rect 9870 5729 9882 5763
rect 9824 5723 9882 5729
rect 11701 5763 11759 5769
rect 11701 5729 11713 5763
rect 11747 5729 11759 5763
rect 11701 5723 11759 5729
rect 11885 5763 11943 5769
rect 11885 5729 11897 5763
rect 11931 5729 11943 5763
rect 13906 5760 13912 5772
rect 13867 5732 13912 5760
rect 11885 5723 11943 5729
rect 9824 5720 9830 5723
rect 2501 5695 2559 5701
rect 2501 5661 2513 5695
rect 2547 5692 2559 5695
rect 2590 5692 2596 5704
rect 2547 5664 2596 5692
rect 2547 5661 2559 5664
rect 2501 5655 2559 5661
rect 2590 5652 2596 5664
rect 2648 5652 2654 5704
rect 3145 5695 3203 5701
rect 3145 5661 3157 5695
rect 3191 5692 3203 5695
rect 3326 5692 3332 5704
rect 3191 5664 3332 5692
rect 3191 5661 3203 5664
rect 3145 5655 3203 5661
rect 3326 5652 3332 5664
rect 3384 5652 3390 5704
rect 4062 5692 4068 5704
rect 4023 5664 4068 5692
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 6822 5692 6828 5704
rect 6783 5664 6828 5692
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 8202 5692 8208 5704
rect 8163 5664 8208 5692
rect 8202 5652 8208 5664
rect 8260 5652 8266 5704
rect 8941 5695 8999 5701
rect 8941 5661 8953 5695
rect 8987 5692 8999 5695
rect 9122 5692 9128 5704
rect 8987 5664 9128 5692
rect 8987 5661 8999 5664
rect 8941 5655 8999 5661
rect 9122 5652 9128 5664
rect 9180 5652 9186 5704
rect 9692 5692 9720 5720
rect 10042 5692 10048 5704
rect 9692 5664 9904 5692
rect 10003 5664 10048 5692
rect 1581 5627 1639 5633
rect 1581 5593 1593 5627
rect 1627 5624 1639 5627
rect 3234 5624 3240 5636
rect 1627 5596 3240 5624
rect 1627 5593 1639 5596
rect 1581 5587 1639 5593
rect 3234 5584 3240 5596
rect 3292 5584 3298 5636
rect 5534 5584 5540 5636
rect 5592 5624 5598 5636
rect 6089 5627 6147 5633
rect 6089 5624 6101 5627
rect 5592 5596 6101 5624
rect 5592 5584 5598 5596
rect 6089 5593 6101 5596
rect 6135 5593 6147 5627
rect 6089 5587 6147 5593
rect 6178 5584 6184 5636
rect 6236 5624 6242 5636
rect 9674 5624 9680 5636
rect 6236 5596 9680 5624
rect 6236 5584 6242 5596
rect 9674 5584 9680 5596
rect 9732 5584 9738 5636
rect 9876 5624 9904 5664
rect 10042 5652 10048 5664
rect 10100 5652 10106 5704
rect 11716 5692 11744 5723
rect 13906 5720 13912 5732
rect 13964 5720 13970 5772
rect 14093 5763 14151 5769
rect 14093 5729 14105 5763
rect 14139 5729 14151 5763
rect 14093 5723 14151 5729
rect 14737 5763 14795 5769
rect 14737 5729 14749 5763
rect 14783 5760 14795 5763
rect 15381 5763 15439 5769
rect 15381 5760 15393 5763
rect 14783 5732 15393 5760
rect 14783 5729 14795 5732
rect 14737 5723 14795 5729
rect 15381 5729 15393 5732
rect 15427 5760 15439 5763
rect 15470 5760 15476 5772
rect 15427 5732 15476 5760
rect 15427 5729 15439 5732
rect 15381 5723 15439 5729
rect 11974 5692 11980 5704
rect 11716 5664 11980 5692
rect 11974 5652 11980 5664
rect 12032 5652 12038 5704
rect 13630 5652 13636 5704
rect 13688 5692 13694 5704
rect 14108 5692 14136 5723
rect 15470 5720 15476 5732
rect 15528 5720 15534 5772
rect 17494 5760 17500 5772
rect 17455 5732 17500 5760
rect 17494 5720 17500 5732
rect 17552 5720 17558 5772
rect 23017 5763 23075 5769
rect 23017 5729 23029 5763
rect 23063 5760 23075 5763
rect 23106 5760 23112 5772
rect 23063 5732 23112 5760
rect 23063 5729 23075 5732
rect 23017 5723 23075 5729
rect 23106 5720 23112 5732
rect 23164 5720 23170 5772
rect 14366 5692 14372 5704
rect 13688 5664 14136 5692
rect 14327 5664 14372 5692
rect 13688 5652 13694 5664
rect 14366 5652 14372 5664
rect 14424 5652 14430 5704
rect 14642 5652 14648 5704
rect 14700 5692 14706 5704
rect 16577 5695 16635 5701
rect 16577 5692 16589 5695
rect 14700 5664 16589 5692
rect 14700 5652 14706 5664
rect 16577 5661 16589 5664
rect 16623 5692 16635 5695
rect 16942 5692 16948 5704
rect 16623 5664 16948 5692
rect 16623 5661 16635 5664
rect 16577 5655 16635 5661
rect 16942 5652 16948 5664
rect 17000 5652 17006 5704
rect 18138 5692 18144 5704
rect 18099 5664 18144 5692
rect 18138 5652 18144 5664
rect 18196 5652 18202 5704
rect 18417 5695 18475 5701
rect 18417 5692 18429 5695
rect 18248 5664 18429 5692
rect 10686 5624 10692 5636
rect 9876 5596 10692 5624
rect 10686 5584 10692 5596
rect 10744 5584 10750 5636
rect 10870 5624 10876 5636
rect 10783 5596 10876 5624
rect 10870 5584 10876 5596
rect 10928 5624 10934 5636
rect 13814 5624 13820 5636
rect 10928 5596 13820 5624
rect 10928 5584 10934 5596
rect 13814 5584 13820 5596
rect 13872 5584 13878 5636
rect 15565 5627 15623 5633
rect 15565 5593 15577 5627
rect 15611 5624 15623 5627
rect 16758 5624 16764 5636
rect 15611 5596 16764 5624
rect 15611 5593 15623 5596
rect 15565 5587 15623 5593
rect 16758 5584 16764 5596
rect 16816 5584 16822 5636
rect 17126 5624 17132 5636
rect 17039 5596 17132 5624
rect 17126 5584 17132 5596
rect 17184 5624 17190 5636
rect 18248 5624 18276 5664
rect 18417 5661 18429 5664
rect 18463 5661 18475 5695
rect 18417 5655 18475 5661
rect 24121 5695 24179 5701
rect 24121 5661 24133 5695
rect 24167 5692 24179 5695
rect 25038 5692 25044 5704
rect 24167 5664 25044 5692
rect 24167 5661 24179 5664
rect 24121 5655 24179 5661
rect 25038 5652 25044 5664
rect 25096 5652 25102 5704
rect 17184 5596 18276 5624
rect 17184 5584 17190 5596
rect 24026 5584 24032 5636
rect 24084 5624 24090 5636
rect 24673 5627 24731 5633
rect 24673 5624 24685 5627
rect 24084 5596 24685 5624
rect 24084 5584 24090 5596
rect 24673 5593 24685 5596
rect 24719 5624 24731 5627
rect 24854 5624 24860 5636
rect 24719 5596 24860 5624
rect 24719 5593 24731 5596
rect 24673 5587 24731 5593
rect 24854 5584 24860 5596
rect 24912 5584 24918 5636
rect 3142 5516 3148 5568
rect 3200 5556 3206 5568
rect 3421 5559 3479 5565
rect 3421 5556 3433 5559
rect 3200 5528 3433 5556
rect 3200 5516 3206 5528
rect 3421 5525 3433 5528
rect 3467 5525 3479 5559
rect 5350 5556 5356 5568
rect 5311 5528 5356 5556
rect 3421 5519 3479 5525
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 5994 5516 6000 5568
rect 6052 5556 6058 5568
rect 7098 5556 7104 5568
rect 6052 5528 7104 5556
rect 6052 5516 6058 5528
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 7742 5556 7748 5568
rect 7703 5528 7748 5556
rect 7742 5516 7748 5528
rect 7800 5516 7806 5568
rect 8110 5556 8116 5568
rect 8071 5528 8116 5556
rect 8110 5516 8116 5528
rect 8168 5516 8174 5568
rect 8478 5556 8484 5568
rect 8439 5528 8484 5556
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 9950 5556 9956 5568
rect 9911 5528 9956 5556
rect 9950 5516 9956 5528
rect 10008 5516 10014 5568
rect 10134 5556 10140 5568
rect 10095 5528 10140 5556
rect 10134 5516 10140 5528
rect 10192 5516 10198 5568
rect 13541 5559 13599 5565
rect 13541 5525 13553 5559
rect 13587 5556 13599 5559
rect 13722 5556 13728 5568
rect 13587 5528 13728 5556
rect 13587 5525 13599 5528
rect 13541 5519 13599 5525
rect 13722 5516 13728 5528
rect 13780 5516 13786 5568
rect 23155 5559 23213 5565
rect 23155 5525 23167 5559
rect 23201 5556 23213 5559
rect 23842 5556 23848 5568
rect 23201 5528 23848 5556
rect 23201 5525 23213 5528
rect 23155 5519 23213 5525
rect 23842 5516 23848 5528
rect 23900 5516 23906 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1673 5355 1731 5361
rect 1673 5321 1685 5355
rect 1719 5352 1731 5355
rect 1762 5352 1768 5364
rect 1719 5324 1768 5352
rect 1719 5321 1731 5324
rect 1673 5315 1731 5321
rect 1762 5312 1768 5324
rect 1820 5312 1826 5364
rect 9217 5355 9275 5361
rect 9217 5352 9229 5355
rect 2424 5324 9229 5352
rect 2424 5157 2452 5324
rect 9217 5321 9229 5324
rect 9263 5321 9275 5355
rect 9217 5315 9275 5321
rect 4338 5244 4344 5296
rect 4396 5284 4402 5296
rect 4985 5287 5043 5293
rect 4985 5284 4997 5287
rect 4396 5256 4997 5284
rect 4396 5244 4402 5256
rect 4985 5253 4997 5256
rect 5031 5284 5043 5287
rect 5810 5284 5816 5296
rect 5031 5256 5816 5284
rect 5031 5253 5043 5256
rect 4985 5247 5043 5253
rect 5810 5244 5816 5256
rect 5868 5244 5874 5296
rect 5905 5287 5963 5293
rect 5905 5253 5917 5287
rect 5951 5284 5963 5287
rect 6086 5284 6092 5296
rect 5951 5256 6092 5284
rect 5951 5253 5963 5256
rect 5905 5247 5963 5253
rect 6086 5244 6092 5256
rect 6144 5244 6150 5296
rect 6273 5287 6331 5293
rect 6273 5253 6285 5287
rect 6319 5284 6331 5287
rect 6730 5284 6736 5296
rect 6319 5256 6736 5284
rect 6319 5253 6331 5256
rect 6273 5247 6331 5253
rect 3053 5219 3111 5225
rect 3053 5185 3065 5219
rect 3099 5216 3111 5219
rect 3878 5216 3884 5228
rect 3099 5188 3884 5216
rect 3099 5185 3111 5188
rect 3053 5179 3111 5185
rect 2409 5151 2467 5157
rect 2409 5148 2421 5151
rect 2148 5120 2421 5148
rect 106 4972 112 5024
rect 164 5012 170 5024
rect 2148 5021 2176 5120
rect 2409 5117 2421 5120
rect 2455 5117 2467 5151
rect 2409 5111 2467 5117
rect 2590 5108 2596 5160
rect 2648 5148 2654 5160
rect 3068 5148 3096 5179
rect 3878 5176 3884 5188
rect 3936 5176 3942 5228
rect 4126 5188 5764 5216
rect 2648 5120 3096 5148
rect 2648 5108 2654 5120
rect 3050 5040 3056 5092
rect 3108 5080 3114 5092
rect 4126 5080 4154 5188
rect 4522 5148 4528 5160
rect 4483 5120 4528 5148
rect 4522 5108 4528 5120
rect 4580 5108 4586 5160
rect 5736 5157 5764 5188
rect 5721 5151 5779 5157
rect 5721 5117 5733 5151
rect 5767 5148 5779 5151
rect 6288 5148 6316 5247
rect 6730 5244 6736 5256
rect 6788 5244 6794 5296
rect 7926 5244 7932 5296
rect 7984 5293 7990 5296
rect 7984 5287 8033 5293
rect 7984 5253 7987 5287
rect 8021 5253 8033 5287
rect 7984 5247 8033 5253
rect 7984 5244 7990 5247
rect 8110 5244 8116 5296
rect 8168 5284 8174 5296
rect 8168 5256 8261 5284
rect 8168 5244 8174 5256
rect 7006 5176 7012 5228
rect 7064 5216 7070 5228
rect 8128 5216 8156 5244
rect 7064 5188 8156 5216
rect 7064 5176 7070 5188
rect 8202 5176 8208 5228
rect 8260 5216 8266 5228
rect 8260 5188 8353 5216
rect 8260 5176 8266 5188
rect 5767 5120 6316 5148
rect 6825 5151 6883 5157
rect 5767 5117 5779 5120
rect 5721 5111 5779 5117
rect 6825 5117 6837 5151
rect 6871 5148 6883 5151
rect 6914 5148 6920 5160
rect 6871 5120 6920 5148
rect 6871 5117 6883 5120
rect 6825 5111 6883 5117
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 7374 5108 7380 5160
rect 7432 5148 7438 5160
rect 7837 5151 7895 5157
rect 7837 5148 7849 5151
rect 7432 5120 7849 5148
rect 7432 5108 7438 5120
rect 7837 5117 7849 5120
rect 7883 5148 7895 5151
rect 8018 5148 8024 5160
rect 7883 5120 8024 5148
rect 7883 5117 7895 5120
rect 7837 5111 7895 5117
rect 8018 5108 8024 5120
rect 8076 5108 8082 5160
rect 4614 5080 4620 5092
rect 3108 5052 4154 5080
rect 4575 5052 4620 5080
rect 3108 5040 3114 5052
rect 4614 5040 4620 5052
rect 4672 5040 4678 5092
rect 5629 5083 5687 5089
rect 5629 5049 5641 5083
rect 5675 5080 5687 5083
rect 6454 5080 6460 5092
rect 5675 5052 6460 5080
rect 5675 5049 5687 5052
rect 5629 5043 5687 5049
rect 6454 5040 6460 5052
rect 6512 5040 6518 5092
rect 7190 5040 7196 5092
rect 7248 5080 7254 5092
rect 7285 5083 7343 5089
rect 7285 5080 7297 5083
rect 7248 5052 7297 5080
rect 7248 5040 7254 5052
rect 7285 5049 7297 5052
rect 7331 5080 7343 5083
rect 7653 5083 7711 5089
rect 7653 5080 7665 5083
rect 7331 5052 7665 5080
rect 7331 5049 7343 5052
rect 7285 5043 7343 5049
rect 7653 5049 7665 5052
rect 7699 5080 7711 5083
rect 8220 5080 8248 5176
rect 9232 5148 9260 5315
rect 9306 5312 9312 5364
rect 9364 5352 9370 5364
rect 9677 5355 9735 5361
rect 9677 5352 9689 5355
rect 9364 5324 9689 5352
rect 9364 5312 9370 5324
rect 9677 5321 9689 5324
rect 9723 5321 9735 5355
rect 9677 5315 9735 5321
rect 11790 5312 11796 5364
rect 11848 5352 11854 5364
rect 12526 5352 12532 5364
rect 11848 5324 12532 5352
rect 11848 5312 11854 5324
rect 12526 5312 12532 5324
rect 12584 5352 12590 5364
rect 12621 5355 12679 5361
rect 12621 5352 12633 5355
rect 12584 5324 12633 5352
rect 12584 5312 12590 5324
rect 12621 5321 12633 5324
rect 12667 5321 12679 5355
rect 12621 5315 12679 5321
rect 13081 5355 13139 5361
rect 13081 5321 13093 5355
rect 13127 5352 13139 5355
rect 16206 5352 16212 5364
rect 13127 5324 16212 5352
rect 13127 5321 13139 5324
rect 13081 5315 13139 5321
rect 16206 5312 16212 5324
rect 16264 5312 16270 5364
rect 16942 5352 16948 5364
rect 16903 5324 16948 5352
rect 16942 5312 16948 5324
rect 17000 5312 17006 5364
rect 17497 5355 17555 5361
rect 17497 5321 17509 5355
rect 17543 5352 17555 5355
rect 18138 5352 18144 5364
rect 17543 5324 18144 5352
rect 17543 5321 17555 5324
rect 17497 5315 17555 5321
rect 18138 5312 18144 5324
rect 18196 5312 18202 5364
rect 23106 5352 23112 5364
rect 23067 5324 23112 5352
rect 23106 5312 23112 5324
rect 23164 5312 23170 5364
rect 23198 5312 23204 5364
rect 23256 5352 23262 5364
rect 24673 5355 24731 5361
rect 24673 5352 24685 5355
rect 23256 5324 24685 5352
rect 23256 5312 23262 5324
rect 24673 5321 24685 5324
rect 24719 5321 24731 5355
rect 25038 5352 25044 5364
rect 24999 5324 25044 5352
rect 24673 5315 24731 5321
rect 25038 5312 25044 5324
rect 25096 5352 25102 5364
rect 25363 5355 25421 5361
rect 25363 5352 25375 5355
rect 25096 5324 25375 5352
rect 25096 5312 25102 5324
rect 25363 5321 25375 5324
rect 25409 5321 25421 5355
rect 25363 5315 25421 5321
rect 11885 5287 11943 5293
rect 11885 5253 11897 5287
rect 11931 5284 11943 5287
rect 11974 5284 11980 5296
rect 11931 5256 11980 5284
rect 11931 5253 11943 5256
rect 11885 5247 11943 5253
rect 11974 5244 11980 5256
rect 12032 5244 12038 5296
rect 12943 5287 13001 5293
rect 12943 5253 12955 5287
rect 12989 5284 13001 5287
rect 16022 5284 16028 5296
rect 12989 5256 16028 5284
rect 12989 5253 13001 5256
rect 12943 5247 13001 5253
rect 16022 5244 16028 5256
rect 16080 5244 16086 5296
rect 16301 5287 16359 5293
rect 16301 5253 16313 5287
rect 16347 5284 16359 5287
rect 16347 5256 19334 5284
rect 16347 5253 16359 5256
rect 16301 5247 16359 5253
rect 11054 5176 11060 5228
rect 11112 5216 11118 5228
rect 17034 5216 17040 5228
rect 11112 5188 17040 5216
rect 11112 5176 11118 5188
rect 17034 5176 17040 5188
rect 17092 5176 17098 5228
rect 19306 5216 19334 5256
rect 23385 5219 23443 5225
rect 23385 5216 23397 5219
rect 19306 5188 23397 5216
rect 23385 5185 23397 5188
rect 23431 5216 23443 5219
rect 23431 5188 23796 5216
rect 23431 5185 23443 5188
rect 23385 5179 23443 5185
rect 9401 5151 9459 5157
rect 9401 5148 9413 5151
rect 9232 5120 9413 5148
rect 9401 5117 9413 5120
rect 9447 5117 9459 5151
rect 9401 5111 9459 5117
rect 9585 5151 9643 5157
rect 9585 5117 9597 5151
rect 9631 5148 9643 5151
rect 9674 5148 9680 5160
rect 9631 5120 9680 5148
rect 9631 5117 9643 5120
rect 9585 5111 9643 5117
rect 9674 5108 9680 5120
rect 9732 5148 9738 5160
rect 10229 5151 10287 5157
rect 10229 5148 10241 5151
rect 9732 5120 10241 5148
rect 9732 5108 9738 5120
rect 10229 5117 10241 5120
rect 10275 5117 10287 5151
rect 10870 5148 10876 5160
rect 10831 5120 10876 5148
rect 10229 5111 10287 5117
rect 10870 5108 10876 5120
rect 10928 5108 10934 5160
rect 11238 5148 11244 5160
rect 11199 5120 11244 5148
rect 11238 5108 11244 5120
rect 11296 5148 11302 5160
rect 12161 5151 12219 5157
rect 12161 5148 12173 5151
rect 11296 5120 12173 5148
rect 11296 5108 11302 5120
rect 12161 5117 12173 5120
rect 12207 5117 12219 5151
rect 12161 5111 12219 5117
rect 12434 5108 12440 5160
rect 12492 5148 12498 5160
rect 12840 5151 12898 5157
rect 12840 5148 12852 5151
rect 12492 5120 12852 5148
rect 12492 5108 12498 5120
rect 12840 5117 12852 5120
rect 12886 5148 12898 5151
rect 13265 5151 13323 5157
rect 13265 5148 13277 5151
rect 12886 5120 13277 5148
rect 12886 5117 12898 5120
rect 12840 5111 12898 5117
rect 13265 5117 13277 5120
rect 13311 5117 13323 5151
rect 13817 5151 13875 5157
rect 13817 5148 13829 5151
rect 13265 5111 13323 5117
rect 13648 5120 13829 5148
rect 7699 5052 8248 5080
rect 8573 5083 8631 5089
rect 7699 5049 7711 5052
rect 7653 5043 7711 5049
rect 8573 5049 8585 5083
rect 8619 5080 8631 5083
rect 11330 5080 11336 5092
rect 8619 5052 11336 5080
rect 8619 5049 8631 5052
rect 8573 5043 8631 5049
rect 11330 5040 11336 5052
rect 11388 5040 11394 5092
rect 11514 5080 11520 5092
rect 11475 5052 11520 5080
rect 11514 5040 11520 5052
rect 11572 5040 11578 5092
rect 11974 5040 11980 5092
rect 12032 5080 12038 5092
rect 13648 5089 13676 5120
rect 13817 5117 13829 5120
rect 13863 5148 13875 5151
rect 13906 5148 13912 5160
rect 13863 5120 13912 5148
rect 13863 5117 13875 5120
rect 13817 5111 13875 5117
rect 13906 5108 13912 5120
rect 13964 5108 13970 5160
rect 14274 5148 14280 5160
rect 14235 5120 14280 5148
rect 14274 5108 14280 5120
rect 14332 5108 14338 5160
rect 14550 5148 14556 5160
rect 14511 5120 14556 5148
rect 14550 5108 14556 5120
rect 14608 5108 14614 5160
rect 14734 5108 14740 5160
rect 14792 5148 14798 5160
rect 15194 5148 15200 5160
rect 14792 5120 15200 5148
rect 14792 5108 14798 5120
rect 15194 5108 15200 5120
rect 15252 5108 15258 5160
rect 15378 5148 15384 5160
rect 15339 5120 15384 5148
rect 15378 5108 15384 5120
rect 15436 5108 15442 5160
rect 16850 5108 16856 5160
rect 16908 5148 16914 5160
rect 18049 5151 18107 5157
rect 18049 5148 18061 5151
rect 16908 5120 18061 5148
rect 16908 5108 16914 5120
rect 18049 5117 18061 5120
rect 18095 5117 18107 5151
rect 18690 5148 18696 5160
rect 18651 5120 18696 5148
rect 18049 5111 18107 5117
rect 18690 5108 18696 5120
rect 18748 5108 18754 5160
rect 23768 5157 23796 5188
rect 23753 5151 23811 5157
rect 23753 5117 23765 5151
rect 23799 5148 23811 5151
rect 24118 5148 24124 5160
rect 23799 5120 24124 5148
rect 23799 5117 23811 5120
rect 23753 5111 23811 5117
rect 24118 5108 24124 5120
rect 24176 5108 24182 5160
rect 25292 5151 25350 5157
rect 25292 5117 25304 5151
rect 25338 5148 25350 5151
rect 25338 5120 25820 5148
rect 25338 5117 25350 5120
rect 25292 5111 25350 5117
rect 13633 5083 13691 5089
rect 13633 5080 13645 5083
rect 12032 5052 13645 5080
rect 12032 5040 12038 5052
rect 13633 5049 13645 5052
rect 13679 5049 13691 5083
rect 13924 5080 13952 5108
rect 14829 5083 14887 5089
rect 14829 5080 14841 5083
rect 13924 5052 14841 5080
rect 13633 5043 13691 5049
rect 14829 5049 14841 5052
rect 14875 5049 14887 5083
rect 15212 5080 15240 5108
rect 15702 5083 15760 5089
rect 15702 5080 15714 5083
rect 15212 5052 15714 5080
rect 14829 5043 14887 5049
rect 15702 5049 15714 5052
rect 15748 5049 15760 5083
rect 15702 5043 15760 5049
rect 17954 5040 17960 5092
rect 18012 5080 18018 5092
rect 19613 5083 19671 5089
rect 19613 5080 19625 5083
rect 18012 5052 19625 5080
rect 18012 5040 18018 5052
rect 19613 5049 19625 5052
rect 19659 5049 19671 5083
rect 19613 5043 19671 5049
rect 2133 5015 2191 5021
rect 2133 5012 2145 5015
rect 164 4984 2145 5012
rect 164 4972 170 4984
rect 2133 4981 2145 4984
rect 2179 4981 2191 5015
rect 2133 4975 2191 4981
rect 3697 5015 3755 5021
rect 3697 4981 3709 5015
rect 3743 5012 3755 5015
rect 3970 5012 3976 5024
rect 3743 4984 3976 5012
rect 3743 4981 3755 4984
rect 3697 4975 3755 4981
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 5258 4972 5264 5024
rect 5316 5012 5322 5024
rect 6362 5012 6368 5024
rect 5316 4984 6368 5012
rect 5316 4972 5322 4984
rect 6362 4972 6368 4984
rect 6420 5012 6426 5024
rect 6549 5015 6607 5021
rect 6549 5012 6561 5015
rect 6420 4984 6561 5012
rect 6420 4972 6426 4984
rect 6549 4981 6561 4984
rect 6595 4981 6607 5015
rect 7006 5012 7012 5024
rect 6967 4984 7012 5012
rect 6549 4975 6607 4981
rect 7006 4972 7012 4984
rect 7064 4972 7070 5024
rect 8754 4972 8760 5024
rect 8812 5012 8818 5024
rect 8941 5015 8999 5021
rect 8941 5012 8953 5015
rect 8812 4984 8953 5012
rect 8812 4972 8818 4984
rect 8941 4981 8953 4984
rect 8987 5012 8999 5015
rect 9766 5012 9772 5024
rect 8987 4984 9772 5012
rect 8987 4981 8999 4984
rect 8941 4975 8999 4981
rect 9766 4972 9772 4984
rect 9824 4972 9830 5024
rect 10686 5012 10692 5024
rect 10599 4984 10692 5012
rect 10686 4972 10692 4984
rect 10744 5012 10750 5024
rect 13081 5015 13139 5021
rect 13081 5012 13093 5015
rect 10744 4984 13093 5012
rect 10744 4972 10750 4984
rect 13081 4981 13093 4984
rect 13127 4981 13139 5015
rect 16666 5012 16672 5024
rect 16627 4984 16672 5012
rect 13081 4975 13139 4981
rect 16666 4972 16672 4984
rect 16724 4972 16730 5024
rect 17770 5012 17776 5024
rect 17731 4984 17776 5012
rect 17770 4972 17776 4984
rect 17828 4972 17834 5024
rect 22278 5012 22284 5024
rect 22239 4984 22284 5012
rect 22278 4972 22284 4984
rect 22336 4972 22342 5024
rect 23934 5012 23940 5024
rect 23895 4984 23940 5012
rect 23934 4972 23940 4984
rect 23992 4972 23998 5024
rect 25792 5021 25820 5120
rect 25777 5015 25835 5021
rect 25777 4981 25789 5015
rect 25823 5012 25835 5015
rect 27062 5012 27068 5024
rect 25823 4984 27068 5012
rect 25823 4981 25835 4984
rect 25777 4975 25835 4981
rect 27062 4972 27068 4984
rect 27120 4972 27126 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 2501 4811 2559 4817
rect 2501 4777 2513 4811
rect 2547 4808 2559 4811
rect 2866 4808 2872 4820
rect 2547 4780 2872 4808
rect 2547 4777 2559 4780
rect 2501 4771 2559 4777
rect 2866 4768 2872 4780
rect 2924 4768 2930 4820
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 5721 4811 5779 4817
rect 5721 4808 5733 4811
rect 4120 4780 5733 4808
rect 4120 4768 4126 4780
rect 5721 4777 5733 4780
rect 5767 4777 5779 4811
rect 5721 4771 5779 4777
rect 5810 4768 5816 4820
rect 5868 4808 5874 4820
rect 6730 4808 6736 4820
rect 5868 4780 6736 4808
rect 5868 4768 5874 4780
rect 6730 4768 6736 4780
rect 6788 4768 6794 4820
rect 7374 4808 7380 4820
rect 7335 4780 7380 4808
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 7558 4808 7564 4820
rect 7484 4780 7564 4808
rect 1394 4740 1400 4752
rect 1355 4712 1400 4740
rect 1394 4700 1400 4712
rect 1452 4700 1458 4752
rect 2682 4700 2688 4752
rect 2740 4740 2746 4752
rect 3099 4743 3157 4749
rect 3099 4740 3111 4743
rect 2740 4712 3111 4740
rect 2740 4700 2746 4712
rect 3099 4709 3111 4712
rect 3145 4709 3157 4743
rect 3099 4703 3157 4709
rect 4525 4743 4583 4749
rect 4525 4709 4537 4743
rect 4571 4740 4583 4743
rect 4614 4740 4620 4752
rect 4571 4712 4620 4740
rect 4571 4709 4583 4712
rect 4525 4703 4583 4709
rect 4614 4700 4620 4712
rect 4672 4700 4678 4752
rect 7484 4740 7512 4780
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 7742 4768 7748 4820
rect 7800 4808 7806 4820
rect 8481 4811 8539 4817
rect 8481 4808 8493 4811
rect 7800 4780 8493 4808
rect 7800 4768 7806 4780
rect 8481 4777 8493 4780
rect 8527 4777 8539 4811
rect 8481 4771 8539 4777
rect 9953 4811 10011 4817
rect 9953 4777 9965 4811
rect 9999 4808 10011 4811
rect 10042 4808 10048 4820
rect 9999 4780 10048 4808
rect 9999 4777 10011 4780
rect 9953 4771 10011 4777
rect 10042 4768 10048 4780
rect 10100 4768 10106 4820
rect 11422 4768 11428 4820
rect 11480 4808 11486 4820
rect 13081 4811 13139 4817
rect 13081 4808 13093 4811
rect 11480 4780 13093 4808
rect 11480 4768 11486 4780
rect 13081 4777 13093 4780
rect 13127 4777 13139 4811
rect 13081 4771 13139 4777
rect 13357 4811 13415 4817
rect 13357 4777 13369 4811
rect 13403 4808 13415 4811
rect 13630 4808 13636 4820
rect 13403 4780 13636 4808
rect 13403 4777 13415 4780
rect 13357 4771 13415 4777
rect 13630 4768 13636 4780
rect 13688 4808 13694 4820
rect 14734 4808 14740 4820
rect 13688 4780 14740 4808
rect 13688 4768 13694 4780
rect 14734 4768 14740 4780
rect 14792 4768 14798 4820
rect 14826 4768 14832 4820
rect 14884 4808 14890 4820
rect 15105 4811 15163 4817
rect 15105 4808 15117 4811
rect 14884 4780 15117 4808
rect 14884 4768 14890 4780
rect 15105 4777 15117 4780
rect 15151 4808 15163 4811
rect 15378 4808 15384 4820
rect 15151 4780 15384 4808
rect 15151 4777 15163 4780
rect 15105 4771 15163 4777
rect 15378 4768 15384 4780
rect 15436 4768 15442 4820
rect 15930 4768 15936 4820
rect 15988 4808 15994 4820
rect 16945 4811 17003 4817
rect 16945 4808 16957 4811
rect 15988 4780 16957 4808
rect 15988 4768 15994 4780
rect 16945 4777 16957 4780
rect 16991 4808 17003 4811
rect 17770 4808 17776 4820
rect 16991 4780 17776 4808
rect 16991 4777 17003 4780
rect 16945 4771 17003 4777
rect 7650 4740 7656 4752
rect 6196 4712 7512 4740
rect 7611 4712 7656 4740
rect 6196 4684 6224 4712
rect 7650 4700 7656 4712
rect 7708 4700 7714 4752
rect 7926 4700 7932 4752
rect 7984 4740 7990 4752
rect 9217 4743 9275 4749
rect 9217 4740 9229 4743
rect 7984 4712 9229 4740
rect 7984 4700 7990 4712
rect 9217 4709 9229 4712
rect 9263 4709 9275 4743
rect 9217 4703 9275 4709
rect 10410 4700 10416 4752
rect 10468 4740 10474 4752
rect 10867 4743 10925 4749
rect 10867 4740 10879 4743
rect 10468 4712 10879 4740
rect 10468 4700 10474 4712
rect 10867 4709 10879 4712
rect 10913 4740 10925 4743
rect 11606 4740 11612 4752
rect 10913 4712 11612 4740
rect 10913 4709 10925 4712
rect 10867 4703 10925 4709
rect 11606 4700 11612 4712
rect 11664 4700 11670 4752
rect 11793 4743 11851 4749
rect 11793 4709 11805 4743
rect 11839 4740 11851 4743
rect 12894 4740 12900 4752
rect 11839 4712 12900 4740
rect 11839 4709 11851 4712
rect 11793 4703 11851 4709
rect 12894 4700 12900 4712
rect 12952 4700 12958 4752
rect 15194 4700 15200 4752
rect 15252 4740 15258 4752
rect 15702 4743 15760 4749
rect 15702 4740 15714 4743
rect 15252 4712 15714 4740
rect 15252 4700 15258 4712
rect 15702 4709 15714 4712
rect 15748 4709 15760 4743
rect 15702 4703 15760 4709
rect 16666 4700 16672 4752
rect 16724 4740 16730 4752
rect 17129 4743 17187 4749
rect 17129 4740 17141 4743
rect 16724 4712 17141 4740
rect 16724 4700 16730 4712
rect 17129 4709 17141 4712
rect 17175 4709 17187 4743
rect 17129 4703 17187 4709
rect 1762 4672 1768 4684
rect 1723 4644 1768 4672
rect 1762 4632 1768 4644
rect 1820 4632 1826 4684
rect 2958 4672 2964 4684
rect 2919 4644 2964 4672
rect 2958 4632 2964 4644
rect 3016 4632 3022 4684
rect 6178 4672 6184 4684
rect 6139 4644 6184 4672
rect 6178 4632 6184 4644
rect 6236 4632 6242 4684
rect 6454 4672 6460 4684
rect 6415 4644 6460 4672
rect 6454 4632 6460 4644
rect 6512 4632 6518 4684
rect 8205 4675 8263 4681
rect 8205 4641 8217 4675
rect 8251 4672 8263 4675
rect 8294 4672 8300 4684
rect 8251 4644 8300 4672
rect 8251 4641 8263 4644
rect 8205 4635 8263 4641
rect 8294 4632 8300 4644
rect 8352 4672 8358 4684
rect 11425 4675 11483 4681
rect 8352 4644 11284 4672
rect 8352 4632 8358 4644
rect 4430 4604 4436 4616
rect 4391 4576 4436 4604
rect 4430 4564 4436 4576
rect 4488 4564 4494 4616
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4573 4767 4607
rect 6638 4604 6644 4616
rect 6599 4576 6644 4604
rect 4709 4567 4767 4573
rect 3326 4496 3332 4548
rect 3384 4536 3390 4548
rect 4724 4536 4752 4567
rect 6638 4564 6644 4576
rect 6696 4564 6702 4616
rect 7558 4604 7564 4616
rect 7519 4576 7564 4604
rect 7558 4564 7564 4576
rect 7616 4564 7622 4616
rect 10502 4604 10508 4616
rect 10463 4576 10508 4604
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 11256 4604 11284 4644
rect 11425 4641 11437 4675
rect 11471 4672 11483 4675
rect 12342 4672 12348 4684
rect 11471 4644 12348 4672
rect 11471 4641 11483 4644
rect 11425 4635 11483 4641
rect 12342 4632 12348 4644
rect 12400 4632 12406 4684
rect 12672 4675 12730 4681
rect 12672 4641 12684 4675
rect 12718 4672 12730 4675
rect 13262 4672 13268 4684
rect 12718 4644 13268 4672
rect 12718 4641 12730 4644
rect 12672 4635 12730 4641
rect 13262 4632 13268 4644
rect 13320 4632 13326 4684
rect 13814 4672 13820 4684
rect 13775 4644 13820 4672
rect 13814 4632 13820 4644
rect 13872 4632 13878 4684
rect 14093 4675 14151 4681
rect 14093 4641 14105 4675
rect 14139 4672 14151 4675
rect 14274 4672 14280 4684
rect 14139 4644 14280 4672
rect 14139 4641 14151 4644
rect 14093 4635 14151 4641
rect 14274 4632 14280 4644
rect 14332 4672 14338 4684
rect 17236 4681 17264 4780
rect 17770 4768 17776 4780
rect 17828 4768 17834 4820
rect 22554 4740 22560 4752
rect 22515 4712 22560 4740
rect 22554 4700 22560 4712
rect 22612 4700 22618 4752
rect 24118 4740 24124 4752
rect 24079 4712 24124 4740
rect 24118 4700 24124 4712
rect 24176 4700 24182 4752
rect 14645 4675 14703 4681
rect 14645 4672 14657 4675
rect 14332 4644 14657 4672
rect 14332 4632 14338 4644
rect 14645 4641 14657 4644
rect 14691 4641 14703 4675
rect 14645 4635 14703 4641
rect 17221 4675 17279 4681
rect 17221 4641 17233 4675
rect 17267 4641 17279 4675
rect 18782 4672 18788 4684
rect 18743 4644 18788 4672
rect 17221 4635 17279 4641
rect 18782 4632 18788 4644
rect 18840 4632 18846 4684
rect 12069 4607 12127 4613
rect 12069 4604 12081 4607
rect 11256 4576 12081 4604
rect 12069 4573 12081 4576
rect 12115 4573 12127 4607
rect 12069 4567 12127 4573
rect 12759 4607 12817 4613
rect 12759 4573 12771 4607
rect 12805 4604 12817 4607
rect 13906 4604 13912 4616
rect 12805 4576 13912 4604
rect 12805 4573 12817 4576
rect 12759 4567 12817 4573
rect 13906 4564 13912 4576
rect 13964 4564 13970 4616
rect 14182 4604 14188 4616
rect 14143 4576 14188 4604
rect 14182 4564 14188 4576
rect 14240 4564 14246 4616
rect 14366 4564 14372 4616
rect 14424 4604 14430 4616
rect 15381 4607 15439 4613
rect 15381 4604 15393 4607
rect 14424 4576 15393 4604
rect 14424 4564 14430 4576
rect 15381 4573 15393 4576
rect 15427 4604 15439 4607
rect 16666 4604 16672 4616
rect 15427 4576 16672 4604
rect 15427 4573 15439 4576
rect 15381 4567 15439 4573
rect 16666 4564 16672 4576
rect 16724 4564 16730 4616
rect 18693 4607 18751 4613
rect 18693 4604 18705 4607
rect 16868 4576 18705 4604
rect 7006 4536 7012 4548
rect 3384 4508 4752 4536
rect 5276 4508 7012 4536
rect 3384 4496 3390 4508
rect 3697 4471 3755 4477
rect 3697 4437 3709 4471
rect 3743 4468 3755 4471
rect 3878 4468 3884 4480
rect 3743 4440 3884 4468
rect 3743 4437 3755 4440
rect 3697 4431 3755 4437
rect 3878 4428 3884 4440
rect 3936 4468 3942 4480
rect 5276 4468 5304 4508
rect 7006 4496 7012 4508
rect 7064 4536 7070 4548
rect 8662 4536 8668 4548
rect 7064 4508 8668 4536
rect 7064 4496 7070 4508
rect 8662 4496 8668 4508
rect 8720 4536 8726 4548
rect 8849 4539 8907 4545
rect 8849 4536 8861 4539
rect 8720 4508 8861 4536
rect 8720 4496 8726 4508
rect 8849 4505 8861 4508
rect 8895 4536 8907 4539
rect 9950 4536 9956 4548
rect 8895 4508 9956 4536
rect 8895 4505 8907 4508
rect 8849 4499 8907 4505
rect 9950 4496 9956 4508
rect 10008 4536 10014 4548
rect 10229 4539 10287 4545
rect 10229 4536 10241 4539
rect 10008 4508 10241 4536
rect 10008 4496 10014 4508
rect 10229 4505 10241 4508
rect 10275 4505 10287 4539
rect 10229 4499 10287 4505
rect 11882 4496 11888 4548
rect 11940 4536 11946 4548
rect 12437 4539 12495 4545
rect 12437 4536 12449 4539
rect 11940 4508 12449 4536
rect 11940 4496 11946 4508
rect 12437 4505 12449 4508
rect 12483 4505 12495 4539
rect 12437 4499 12495 4505
rect 12618 4496 12624 4548
rect 12676 4536 12682 4548
rect 16868 4536 16896 4576
rect 18693 4573 18705 4576
rect 18739 4573 18751 4607
rect 22462 4604 22468 4616
rect 22423 4576 22468 4604
rect 18693 4567 18751 4573
rect 22462 4564 22468 4576
rect 22520 4564 22526 4616
rect 22738 4604 22744 4616
rect 22699 4576 22744 4604
rect 22738 4564 22744 4576
rect 22796 4564 22802 4616
rect 23842 4564 23848 4616
rect 23900 4604 23906 4616
rect 24026 4604 24032 4616
rect 23900 4576 24032 4604
rect 23900 4564 23906 4576
rect 24026 4564 24032 4576
rect 24084 4564 24090 4616
rect 24210 4564 24216 4616
rect 24268 4604 24274 4616
rect 24305 4607 24363 4613
rect 24305 4604 24317 4607
rect 24268 4576 24317 4604
rect 24268 4564 24274 4576
rect 24305 4573 24317 4576
rect 24351 4573 24363 4607
rect 24305 4567 24363 4573
rect 12676 4508 16896 4536
rect 22480 4536 22508 4564
rect 24228 4536 24256 4564
rect 22480 4508 24256 4536
rect 12676 4496 12682 4508
rect 5442 4468 5448 4480
rect 3936 4440 5304 4468
rect 5403 4440 5448 4468
rect 3936 4428 3942 4440
rect 5442 4428 5448 4440
rect 5500 4428 5506 4480
rect 6914 4468 6920 4480
rect 6875 4440 6920 4468
rect 6914 4428 6920 4440
rect 6972 4428 6978 4480
rect 11330 4428 11336 4480
rect 11388 4468 11394 4480
rect 13357 4471 13415 4477
rect 13357 4468 13369 4471
rect 11388 4440 13369 4468
rect 11388 4428 11394 4440
rect 13357 4437 13369 4440
rect 13403 4468 13415 4471
rect 13449 4471 13507 4477
rect 13449 4468 13461 4471
rect 13403 4440 13461 4468
rect 13403 4437 13415 4440
rect 13357 4431 13415 4437
rect 13449 4437 13461 4440
rect 13495 4437 13507 4471
rect 16298 4468 16304 4480
rect 16259 4440 16304 4468
rect 13449 4431 13507 4437
rect 16298 4428 16304 4440
rect 16356 4428 16362 4480
rect 18233 4471 18291 4477
rect 18233 4437 18245 4471
rect 18279 4468 18291 4471
rect 18690 4468 18696 4480
rect 18279 4440 18696 4468
rect 18279 4437 18291 4440
rect 18233 4431 18291 4437
rect 18690 4428 18696 4440
rect 18748 4428 18754 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1854 4264 1860 4276
rect 1815 4236 1860 4264
rect 1854 4224 1860 4236
rect 1912 4224 1918 4276
rect 2958 4264 2964 4276
rect 2919 4236 2964 4264
rect 2958 4224 2964 4236
rect 3016 4224 3022 4276
rect 3513 4267 3571 4273
rect 3513 4233 3525 4267
rect 3559 4264 3571 4267
rect 3694 4264 3700 4276
rect 3559 4236 3700 4264
rect 3559 4233 3571 4236
rect 3513 4227 3571 4233
rect 3694 4224 3700 4236
rect 3752 4273 3758 4276
rect 3752 4267 3801 4273
rect 3752 4233 3755 4267
rect 3789 4233 3801 4267
rect 3878 4264 3884 4276
rect 3839 4236 3884 4264
rect 3752 4227 3801 4233
rect 3752 4224 3758 4227
rect 3878 4224 3884 4236
rect 3936 4224 3942 4276
rect 4246 4264 4252 4276
rect 4207 4236 4252 4264
rect 4246 4224 4252 4236
rect 4304 4224 4310 4276
rect 4614 4264 4620 4276
rect 4575 4236 4620 4264
rect 4614 4224 4620 4236
rect 4672 4224 4678 4276
rect 5166 4224 5172 4276
rect 5224 4224 5230 4276
rect 8110 4264 8116 4276
rect 6472 4236 8116 4264
rect 4522 4156 4528 4208
rect 4580 4196 4586 4208
rect 5184 4196 5212 4224
rect 6178 4196 6184 4208
rect 4580 4168 5212 4196
rect 6139 4168 6184 4196
rect 4580 4156 4586 4168
rect 6178 4156 6184 4168
rect 6236 4156 6242 4208
rect 3970 4128 3976 4140
rect 3931 4100 3976 4128
rect 3970 4088 3976 4100
rect 4028 4088 4034 4140
rect 4798 4088 4804 4140
rect 4856 4128 4862 4140
rect 5718 4128 5724 4140
rect 4856 4100 5724 4128
rect 4856 4088 4862 4100
rect 5718 4088 5724 4100
rect 5776 4088 5782 4140
rect 1762 4060 1768 4072
rect 1723 4032 1768 4060
rect 1762 4020 1768 4032
rect 1820 4020 1826 4072
rect 2498 4060 2504 4072
rect 2459 4032 2504 4060
rect 2498 4020 2504 4032
rect 2556 4020 2562 4072
rect 3234 4020 3240 4072
rect 3292 4060 3298 4072
rect 3602 4060 3608 4072
rect 3292 4032 3608 4060
rect 3292 4020 3298 4032
rect 3602 4020 3608 4032
rect 3660 4020 3666 4072
rect 5077 4063 5135 4069
rect 5077 4029 5089 4063
rect 5123 4060 5135 4063
rect 5258 4060 5264 4072
rect 5123 4032 5264 4060
rect 5123 4029 5135 4032
rect 5077 4023 5135 4029
rect 5258 4020 5264 4032
rect 5316 4020 5322 4072
rect 5442 4020 5448 4072
rect 5500 4060 5506 4072
rect 5629 4063 5687 4069
rect 5629 4060 5641 4063
rect 5500 4032 5641 4060
rect 5500 4020 5506 4032
rect 5629 4029 5641 4032
rect 5675 4060 5687 4063
rect 6472 4060 6500 4236
rect 8110 4224 8116 4236
rect 8168 4224 8174 4276
rect 8202 4224 8208 4276
rect 8260 4264 8266 4276
rect 10502 4264 10508 4276
rect 8260 4236 10508 4264
rect 8260 4224 8266 4236
rect 10502 4224 10508 4236
rect 10560 4264 10566 4276
rect 10870 4264 10876 4276
rect 10560 4236 10876 4264
rect 10560 4224 10566 4236
rect 10870 4224 10876 4236
rect 10928 4224 10934 4276
rect 13262 4224 13268 4276
rect 13320 4264 13326 4276
rect 13998 4264 14004 4276
rect 13320 4236 14004 4264
rect 13320 4224 13326 4236
rect 13998 4224 14004 4236
rect 14056 4264 14062 4276
rect 16577 4267 16635 4273
rect 16577 4264 16589 4267
rect 14056 4236 16589 4264
rect 14056 4224 14062 4236
rect 16577 4233 16589 4236
rect 16623 4233 16635 4267
rect 16850 4264 16856 4276
rect 16811 4236 16856 4264
rect 16577 4227 16635 4233
rect 16850 4224 16856 4236
rect 16908 4224 16914 4276
rect 21545 4267 21603 4273
rect 21545 4233 21557 4267
rect 21591 4264 21603 4267
rect 22462 4264 22468 4276
rect 21591 4236 22468 4264
rect 21591 4233 21603 4236
rect 21545 4227 21603 4233
rect 22462 4224 22468 4236
rect 22520 4224 22526 4276
rect 23934 4264 23940 4276
rect 23895 4236 23940 4264
rect 23934 4224 23940 4236
rect 23992 4224 23998 4276
rect 6730 4156 6736 4208
rect 6788 4196 6794 4208
rect 7374 4196 7380 4208
rect 6788 4168 7380 4196
rect 6788 4156 6794 4168
rect 7374 4156 7380 4168
rect 7432 4156 7438 4208
rect 8662 4196 8668 4208
rect 8623 4168 8668 4196
rect 8662 4156 8668 4168
rect 8720 4156 8726 4208
rect 9723 4199 9781 4205
rect 9723 4165 9735 4199
rect 9769 4196 9781 4199
rect 11422 4196 11428 4208
rect 9769 4168 11428 4196
rect 9769 4165 9781 4168
rect 9723 4159 9781 4165
rect 11422 4156 11428 4168
rect 11480 4156 11486 4208
rect 13538 4156 13544 4208
rect 13596 4196 13602 4208
rect 17034 4196 17040 4208
rect 13596 4168 17040 4196
rect 13596 4156 13602 4168
rect 17034 4156 17040 4168
rect 17092 4156 17098 4208
rect 17218 4156 17224 4208
rect 17276 4196 17282 4208
rect 18782 4196 18788 4208
rect 17276 4168 18788 4196
rect 17276 4156 17282 4168
rect 18782 4156 18788 4168
rect 18840 4196 18846 4208
rect 19061 4199 19119 4205
rect 19061 4196 19073 4199
rect 18840 4168 19073 4196
rect 18840 4156 18846 4168
rect 19061 4165 19073 4168
rect 19107 4165 19119 4199
rect 19061 4159 19119 4165
rect 23477 4199 23535 4205
rect 23477 4165 23489 4199
rect 23523 4196 23535 4199
rect 24118 4196 24124 4208
rect 23523 4168 24124 4196
rect 23523 4165 23535 4168
rect 23477 4159 23535 4165
rect 24118 4156 24124 4168
rect 24176 4156 24182 4208
rect 8202 4128 8208 4140
rect 5675 4032 6500 4060
rect 6564 4100 8208 4128
rect 5675 4029 5687 4032
rect 5629 4023 5687 4029
rect 1673 3995 1731 4001
rect 1673 3961 1685 3995
rect 1719 3992 1731 3995
rect 2516 3992 2544 4020
rect 1719 3964 2544 3992
rect 1719 3961 1731 3964
rect 1673 3955 1731 3961
rect 4798 3952 4804 4004
rect 4856 3992 4862 4004
rect 5905 3995 5963 4001
rect 4856 3964 5764 3992
rect 4856 3952 4862 3964
rect 5736 3924 5764 3964
rect 5905 3961 5917 3995
rect 5951 3992 5963 3995
rect 6564 3992 6592 4100
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 11882 4128 11888 4140
rect 10244 4100 11888 4128
rect 6638 4020 6644 4072
rect 6696 4060 6702 4072
rect 9674 4069 9680 4072
rect 7469 4063 7527 4069
rect 7469 4060 7481 4063
rect 6696 4032 7481 4060
rect 6696 4020 6702 4032
rect 7469 4029 7481 4032
rect 7515 4060 7527 4063
rect 9493 4063 9551 4069
rect 9493 4060 9505 4063
rect 7515 4032 9505 4060
rect 7515 4029 7527 4032
rect 7469 4023 7527 4029
rect 9493 4029 9505 4032
rect 9539 4029 9551 4063
rect 9652 4063 9680 4069
rect 9652 4060 9664 4063
rect 9587 4032 9664 4060
rect 9493 4023 9551 4029
rect 9652 4029 9664 4032
rect 9732 4060 9738 4072
rect 10244 4060 10272 4100
rect 11882 4088 11888 4100
rect 11940 4088 11946 4140
rect 12526 4128 12532 4140
rect 12487 4100 12532 4128
rect 12526 4088 12532 4100
rect 12584 4088 12590 4140
rect 13814 4088 13820 4140
rect 13872 4128 13878 4140
rect 13909 4131 13967 4137
rect 13909 4128 13921 4131
rect 13872 4100 13921 4128
rect 13872 4088 13878 4100
rect 13909 4097 13921 4100
rect 13955 4128 13967 4131
rect 14001 4131 14059 4137
rect 14001 4128 14013 4131
rect 13955 4100 14013 4128
rect 13955 4097 13967 4100
rect 13909 4091 13967 4097
rect 14001 4097 14013 4100
rect 14047 4097 14059 4131
rect 14826 4128 14832 4140
rect 14787 4100 14832 4128
rect 14001 4091 14059 4097
rect 10410 4060 10416 4072
rect 9732 4032 10272 4060
rect 10371 4032 10416 4060
rect 9652 4023 9680 4029
rect 9674 4020 9680 4023
rect 9732 4020 9738 4032
rect 10410 4020 10416 4032
rect 10468 4020 10474 4072
rect 10597 4063 10655 4069
rect 10597 4029 10609 4063
rect 10643 4060 10655 4063
rect 10686 4060 10692 4072
rect 10643 4032 10692 4060
rect 10643 4029 10655 4032
rect 10597 4023 10655 4029
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 11517 4063 11575 4069
rect 11517 4029 11529 4063
rect 11563 4060 11575 4063
rect 11974 4060 11980 4072
rect 11563 4032 11980 4060
rect 11563 4029 11575 4032
rect 11517 4023 11575 4029
rect 11974 4020 11980 4032
rect 12032 4020 12038 4072
rect 14016 4060 14044 4091
rect 14826 4088 14832 4100
rect 14884 4088 14890 4140
rect 15286 4088 15292 4140
rect 15344 4128 15350 4140
rect 15381 4131 15439 4137
rect 15381 4128 15393 4131
rect 15344 4100 15393 4128
rect 15344 4088 15350 4100
rect 15381 4097 15393 4100
rect 15427 4097 15439 4131
rect 15381 4091 15439 4097
rect 16485 4131 16543 4137
rect 16485 4097 16497 4131
rect 16531 4128 16543 4131
rect 16577 4131 16635 4137
rect 16577 4128 16589 4131
rect 16531 4100 16589 4128
rect 16531 4097 16543 4100
rect 16485 4091 16543 4097
rect 16577 4097 16589 4100
rect 16623 4128 16635 4131
rect 18966 4128 18972 4140
rect 16623 4100 18972 4128
rect 16623 4097 16635 4100
rect 16577 4091 16635 4097
rect 18966 4088 18972 4100
rect 19024 4088 19030 4140
rect 22097 4131 22155 4137
rect 22097 4097 22109 4131
rect 22143 4128 22155 4131
rect 22278 4128 22284 4140
rect 22143 4100 22284 4128
rect 22143 4097 22155 4100
rect 22097 4091 22155 4097
rect 22278 4088 22284 4100
rect 22336 4088 22342 4140
rect 22738 4128 22744 4140
rect 22699 4100 22744 4128
rect 22738 4088 22744 4100
rect 22796 4088 22802 4140
rect 24210 4088 24216 4140
rect 24268 4128 24274 4140
rect 24489 4131 24547 4137
rect 24489 4128 24501 4131
rect 24268 4100 24501 4128
rect 24268 4088 24274 4100
rect 24489 4097 24501 4100
rect 24535 4097 24547 4131
rect 24489 4091 24547 4097
rect 14185 4063 14243 4069
rect 14185 4060 14197 4063
rect 14016 4032 14197 4060
rect 14185 4029 14197 4032
rect 14231 4029 14243 4063
rect 14734 4060 14740 4072
rect 14695 4032 14740 4060
rect 14185 4023 14243 4029
rect 14734 4020 14740 4032
rect 14792 4020 14798 4072
rect 16666 4020 16672 4072
rect 16724 4060 16730 4072
rect 17129 4063 17187 4069
rect 17129 4060 17141 4063
rect 16724 4032 17141 4060
rect 16724 4020 16730 4032
rect 17129 4029 17141 4032
rect 17175 4029 17187 4063
rect 17129 4023 17187 4029
rect 17218 4020 17224 4072
rect 17276 4060 17282 4072
rect 17865 4063 17923 4069
rect 17865 4060 17877 4063
rect 17276 4032 17877 4060
rect 17276 4020 17282 4032
rect 17865 4029 17877 4032
rect 17911 4060 17923 4063
rect 18141 4063 18199 4069
rect 18141 4060 18153 4063
rect 17911 4032 18153 4060
rect 17911 4029 17923 4032
rect 17865 4023 17923 4029
rect 18141 4029 18153 4032
rect 18187 4029 18199 4063
rect 18141 4023 18199 4029
rect 20692 4063 20750 4069
rect 20692 4029 20704 4063
rect 20738 4060 20750 4063
rect 21082 4060 21088 4072
rect 20738 4032 21088 4060
rect 20738 4029 20750 4032
rect 20692 4023 20750 4029
rect 21082 4020 21088 4032
rect 21140 4020 21146 4072
rect 7650 3992 7656 4004
rect 5951 3964 6592 3992
rect 7300 3964 7656 3992
rect 5951 3961 5963 3964
rect 5905 3955 5963 3961
rect 6549 3927 6607 3933
rect 6549 3924 6561 3927
rect 5736 3896 6561 3924
rect 6549 3893 6561 3896
rect 6595 3924 6607 3927
rect 7300 3924 7328 3964
rect 7650 3952 7656 3964
rect 7708 3952 7714 4004
rect 7810 3995 7868 4001
rect 7810 3961 7822 3995
rect 7856 3992 7868 3995
rect 9122 3992 9128 4004
rect 7856 3964 9128 3992
rect 7856 3961 7868 3964
rect 7810 3955 7868 3961
rect 9122 3952 9128 3964
rect 9180 3992 9186 4004
rect 10137 3995 10195 4001
rect 10137 3992 10149 3995
rect 9180 3964 10149 3992
rect 9180 3952 9186 3964
rect 10137 3961 10149 3964
rect 10183 3992 10195 3995
rect 10428 3992 10456 4020
rect 10918 3995 10976 4001
rect 10918 3992 10930 3995
rect 10183 3964 10930 3992
rect 10183 3961 10195 3964
rect 10137 3955 10195 3961
rect 10918 3961 10930 3964
rect 10964 3961 10976 3995
rect 10918 3955 10976 3961
rect 12253 3995 12311 4001
rect 12253 3961 12265 3995
rect 12299 3992 12311 3995
rect 12618 3992 12624 4004
rect 12299 3964 12624 3992
rect 12299 3961 12311 3964
rect 12253 3955 12311 3961
rect 12618 3952 12624 3964
rect 12676 3952 12682 4004
rect 13173 3995 13231 4001
rect 13173 3961 13185 3995
rect 13219 3992 13231 3995
rect 13814 3992 13820 4004
rect 13219 3964 13820 3992
rect 13219 3961 13231 3964
rect 13173 3955 13231 3961
rect 13814 3952 13820 3964
rect 13872 3992 13878 4004
rect 15838 3992 15844 4004
rect 13872 3964 15745 3992
rect 15799 3964 15844 3992
rect 13872 3952 13878 3964
rect 6595 3896 7328 3924
rect 6595 3893 6607 3896
rect 6549 3887 6607 3893
rect 7374 3884 7380 3936
rect 7432 3924 7438 3936
rect 8389 3927 8447 3933
rect 8389 3924 8401 3927
rect 7432 3896 8401 3924
rect 7432 3884 7438 3896
rect 8389 3893 8401 3896
rect 8435 3924 8447 3927
rect 9033 3927 9091 3933
rect 9033 3924 9045 3927
rect 8435 3896 9045 3924
rect 8435 3893 8447 3896
rect 8389 3887 8447 3893
rect 9033 3893 9045 3896
rect 9079 3924 9091 3927
rect 9306 3924 9312 3936
rect 9079 3896 9312 3924
rect 9079 3893 9091 3896
rect 9033 3887 9091 3893
rect 9306 3884 9312 3896
rect 9364 3884 9370 3936
rect 9398 3884 9404 3936
rect 9456 3924 9462 3936
rect 11793 3927 11851 3933
rect 11793 3924 11805 3927
rect 9456 3896 11805 3924
rect 9456 3884 9462 3896
rect 11793 3893 11805 3896
rect 11839 3893 11851 3927
rect 11793 3887 11851 3893
rect 12342 3884 12348 3936
rect 12400 3924 12406 3936
rect 13538 3924 13544 3936
rect 12400 3896 13544 3924
rect 12400 3884 12406 3896
rect 13538 3884 13544 3896
rect 13596 3884 13602 3936
rect 13725 3927 13783 3933
rect 13725 3893 13737 3927
rect 13771 3924 13783 3927
rect 13909 3927 13967 3933
rect 13909 3924 13921 3927
rect 13771 3896 13921 3924
rect 13771 3893 13783 3896
rect 13725 3887 13783 3893
rect 13909 3893 13921 3896
rect 13955 3893 13967 3927
rect 15717 3924 15745 3964
rect 15838 3952 15844 3964
rect 15896 3952 15902 4004
rect 15933 3995 15991 4001
rect 15933 3961 15945 3995
rect 15979 3992 15991 3995
rect 16850 3992 16856 4004
rect 15979 3964 16856 3992
rect 15979 3961 15991 3964
rect 15933 3955 15991 3961
rect 16850 3952 16856 3964
rect 16908 3952 16914 4004
rect 17770 3992 17776 4004
rect 17052 3964 17776 3992
rect 17052 3924 17080 3964
rect 17770 3952 17776 3964
rect 17828 3952 17834 4004
rect 18046 3992 18052 4004
rect 18007 3964 18052 3992
rect 18046 3952 18052 3964
rect 18104 3952 18110 4004
rect 21913 3995 21971 4001
rect 21913 3961 21925 3995
rect 21959 3992 21971 3995
rect 22186 3992 22192 4004
rect 21959 3964 22192 3992
rect 21959 3961 21971 3964
rect 21913 3955 21971 3961
rect 22186 3952 22192 3964
rect 22244 3952 22250 4004
rect 24210 3992 24216 4004
rect 24171 3964 24216 3992
rect 24210 3952 24216 3964
rect 24268 3952 24274 4004
rect 24305 3995 24363 4001
rect 24305 3961 24317 3995
rect 24351 3961 24363 3995
rect 24305 3955 24363 3961
rect 15717 3896 17080 3924
rect 13909 3887 13967 3893
rect 18138 3884 18144 3936
rect 18196 3924 18202 3936
rect 19613 3927 19671 3933
rect 19613 3924 19625 3927
rect 18196 3896 19625 3924
rect 18196 3884 18202 3896
rect 19613 3893 19625 3896
rect 19659 3893 19671 3927
rect 19613 3887 19671 3893
rect 19978 3884 19984 3936
rect 20036 3924 20042 3936
rect 20763 3927 20821 3933
rect 20763 3924 20775 3927
rect 20036 3896 20775 3924
rect 20036 3884 20042 3896
rect 20763 3893 20775 3896
rect 20809 3893 20821 3927
rect 20763 3887 20821 3893
rect 22554 3884 22560 3936
rect 22612 3924 22618 3936
rect 23017 3927 23075 3933
rect 23017 3924 23029 3927
rect 22612 3896 23029 3924
rect 22612 3884 22618 3896
rect 23017 3893 23029 3896
rect 23063 3893 23075 3927
rect 23017 3887 23075 3893
rect 23934 3884 23940 3936
rect 23992 3924 23998 3936
rect 24320 3924 24348 3955
rect 23992 3896 24348 3924
rect 23992 3884 23998 3896
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1578 3680 1584 3732
rect 1636 3720 1642 3732
rect 1673 3723 1731 3729
rect 1673 3720 1685 3723
rect 1636 3692 1685 3720
rect 1636 3680 1642 3692
rect 1673 3689 1685 3692
rect 1719 3689 1731 3723
rect 3602 3720 3608 3732
rect 3563 3692 3608 3720
rect 1673 3683 1731 3689
rect 3602 3680 3608 3692
rect 3660 3680 3666 3732
rect 3970 3680 3976 3732
rect 4028 3720 4034 3732
rect 4982 3720 4988 3732
rect 4028 3692 4988 3720
rect 4028 3680 4034 3692
rect 4982 3680 4988 3692
rect 5040 3680 5046 3732
rect 6273 3723 6331 3729
rect 6273 3689 6285 3723
rect 6319 3720 6331 3723
rect 6454 3720 6460 3732
rect 6319 3692 6460 3720
rect 6319 3689 6331 3692
rect 6273 3683 6331 3689
rect 6454 3680 6460 3692
rect 6512 3680 6518 3732
rect 6638 3680 6644 3732
rect 6696 3720 6702 3732
rect 7926 3720 7932 3732
rect 6696 3692 7211 3720
rect 7887 3692 7932 3720
rect 6696 3680 6702 3692
rect 2409 3655 2467 3661
rect 2409 3621 2421 3655
rect 2455 3652 2467 3655
rect 2590 3652 2596 3664
rect 2455 3624 2596 3652
rect 2455 3621 2467 3624
rect 2409 3615 2467 3621
rect 2590 3612 2596 3624
rect 2648 3612 2654 3664
rect 3142 3652 3148 3664
rect 3103 3624 3148 3652
rect 3142 3612 3148 3624
rect 3200 3612 3206 3664
rect 3234 3612 3240 3664
rect 3292 3652 3298 3664
rect 5353 3655 5411 3661
rect 5353 3652 5365 3655
rect 3292 3624 5365 3652
rect 3292 3612 3298 3624
rect 5353 3621 5365 3624
rect 5399 3652 5411 3655
rect 6549 3655 6607 3661
rect 6549 3652 6561 3655
rect 5399 3624 6561 3652
rect 5399 3621 5411 3624
rect 5353 3615 5411 3621
rect 6549 3621 6561 3624
rect 6595 3621 6607 3655
rect 6549 3615 6607 3621
rect 1302 3544 1308 3596
rect 1360 3584 1366 3596
rect 1464 3587 1522 3593
rect 1464 3584 1476 3587
rect 1360 3556 1476 3584
rect 1360 3544 1366 3556
rect 1464 3553 1476 3556
rect 1510 3584 1522 3587
rect 1854 3584 1860 3596
rect 1510 3556 1860 3584
rect 1510 3553 1522 3556
rect 1464 3547 1522 3553
rect 1854 3544 1860 3556
rect 1912 3544 1918 3596
rect 4224 3587 4282 3593
rect 4224 3553 4236 3587
rect 4270 3584 4282 3587
rect 4706 3584 4712 3596
rect 4270 3556 4712 3584
rect 4270 3553 4282 3556
rect 4224 3547 4282 3553
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 6564 3584 6592 3615
rect 6730 3612 6736 3664
rect 6788 3652 6794 3664
rect 7054 3655 7112 3661
rect 7054 3652 7066 3655
rect 6788 3624 7066 3652
rect 6788 3612 6794 3624
rect 7054 3621 7066 3624
rect 7100 3621 7112 3655
rect 7183 3652 7211 3692
rect 7926 3680 7932 3692
rect 7984 3680 7990 3732
rect 9306 3720 9312 3732
rect 9267 3692 9312 3720
rect 9306 3680 9312 3692
rect 9364 3680 9370 3732
rect 10870 3720 10876 3732
rect 10831 3692 10876 3720
rect 10870 3680 10876 3692
rect 10928 3680 10934 3732
rect 14274 3680 14280 3732
rect 14332 3720 14338 3732
rect 14461 3723 14519 3729
rect 14461 3720 14473 3723
rect 14332 3692 14473 3720
rect 14332 3680 14338 3692
rect 14461 3689 14473 3692
rect 14507 3689 14519 3723
rect 14461 3683 14519 3689
rect 14734 3680 14740 3732
rect 14792 3720 14798 3732
rect 14829 3723 14887 3729
rect 14829 3720 14841 3723
rect 14792 3692 14841 3720
rect 14792 3680 14798 3692
rect 14829 3689 14841 3692
rect 14875 3689 14887 3723
rect 14829 3683 14887 3689
rect 15838 3680 15844 3732
rect 15896 3720 15902 3732
rect 16577 3723 16635 3729
rect 16577 3720 16589 3723
rect 15896 3692 16589 3720
rect 15896 3680 15902 3692
rect 16577 3689 16589 3692
rect 16623 3720 16635 3723
rect 17954 3720 17960 3732
rect 16623 3692 17960 3720
rect 16623 3689 16635 3692
rect 16577 3683 16635 3689
rect 17954 3680 17960 3692
rect 18012 3680 18018 3732
rect 22097 3723 22155 3729
rect 22097 3689 22109 3723
rect 22143 3720 22155 3723
rect 22278 3720 22284 3732
rect 22143 3692 22284 3720
rect 22143 3689 22155 3692
rect 22097 3683 22155 3689
rect 22278 3680 22284 3692
rect 22336 3680 22342 3732
rect 24026 3680 24032 3732
rect 24084 3720 24090 3732
rect 24213 3723 24271 3729
rect 24213 3720 24225 3723
rect 24084 3692 24225 3720
rect 24084 3680 24090 3692
rect 24213 3689 24225 3692
rect 24259 3689 24271 3723
rect 24903 3723 24961 3729
rect 24903 3720 24915 3723
rect 24213 3683 24271 3689
rect 24596 3692 24915 3720
rect 10597 3655 10655 3661
rect 7183 3624 10456 3652
rect 7054 3615 7112 3621
rect 7653 3587 7711 3593
rect 7653 3584 7665 3587
rect 6564 3556 7665 3584
rect 7653 3553 7665 3556
rect 7699 3584 7711 3587
rect 8297 3587 8355 3593
rect 8297 3584 8309 3587
rect 7699 3556 8309 3584
rect 7699 3553 7711 3556
rect 7653 3547 7711 3553
rect 8297 3553 8309 3556
rect 8343 3553 8355 3587
rect 9858 3584 9864 3596
rect 9819 3556 9864 3584
rect 8297 3547 8355 3553
rect 9858 3544 9864 3556
rect 9916 3544 9922 3596
rect 10318 3584 10324 3596
rect 10279 3556 10324 3584
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 10428 3584 10456 3624
rect 10597 3621 10609 3655
rect 10643 3652 10655 3655
rect 10686 3652 10692 3664
rect 10643 3624 10692 3652
rect 10643 3621 10655 3624
rect 10597 3615 10655 3621
rect 10686 3612 10692 3624
rect 10744 3652 10750 3664
rect 11241 3655 11299 3661
rect 11241 3652 11253 3655
rect 10744 3624 11253 3652
rect 10744 3612 10750 3624
rect 11241 3621 11253 3624
rect 11287 3621 11299 3655
rect 11241 3615 11299 3621
rect 11606 3612 11612 3664
rect 11664 3652 11670 3664
rect 12022 3655 12080 3661
rect 12022 3652 12034 3655
rect 11664 3624 12034 3652
rect 11664 3612 11670 3624
rect 12022 3621 12034 3624
rect 12068 3621 12080 3655
rect 12022 3615 12080 3621
rect 13538 3612 13544 3664
rect 13596 3652 13602 3664
rect 13633 3655 13691 3661
rect 13633 3652 13645 3655
rect 13596 3624 13645 3652
rect 13596 3612 13602 3624
rect 13633 3621 13645 3624
rect 13679 3621 13691 3655
rect 13633 3615 13691 3621
rect 15286 3612 15292 3664
rect 15344 3652 15350 3664
rect 15610 3655 15668 3661
rect 15610 3652 15622 3655
rect 15344 3624 15622 3652
rect 15344 3612 15350 3624
rect 15610 3621 15622 3624
rect 15656 3621 15668 3655
rect 17218 3652 17224 3664
rect 15610 3615 15668 3621
rect 16224 3624 17224 3652
rect 16224 3593 16252 3624
rect 17218 3612 17224 3624
rect 17276 3612 17282 3664
rect 17770 3612 17776 3664
rect 17828 3652 17834 3664
rect 18417 3655 18475 3661
rect 18417 3652 18429 3655
rect 17828 3624 18429 3652
rect 17828 3612 17834 3624
rect 18417 3621 18429 3624
rect 18463 3621 18475 3655
rect 18417 3615 18475 3621
rect 13265 3587 13323 3593
rect 13265 3584 13277 3587
rect 10428 3556 13277 3584
rect 13265 3553 13277 3556
rect 13311 3553 13323 3587
rect 13265 3547 13323 3553
rect 16209 3587 16267 3593
rect 16209 3553 16221 3587
rect 16255 3553 16267 3587
rect 18432 3584 18460 3615
rect 18690 3612 18696 3664
rect 18748 3652 18754 3664
rect 18785 3655 18843 3661
rect 18785 3652 18797 3655
rect 18748 3624 18797 3652
rect 18748 3612 18754 3624
rect 18785 3621 18797 3624
rect 18831 3652 18843 3655
rect 19058 3652 19064 3664
rect 18831 3624 19064 3652
rect 18831 3621 18843 3624
rect 18785 3615 18843 3621
rect 19058 3612 19064 3624
rect 19116 3612 19122 3664
rect 22186 3652 22192 3664
rect 22147 3624 22192 3652
rect 22186 3612 22192 3624
rect 22244 3612 22250 3664
rect 20809 3587 20867 3593
rect 18432 3556 18552 3584
rect 16209 3547 16267 3553
rect 1946 3476 1952 3528
rect 2004 3516 2010 3528
rect 2777 3519 2835 3525
rect 2777 3516 2789 3519
rect 2004 3488 2789 3516
rect 2004 3476 2010 3488
rect 2777 3485 2789 3488
rect 2823 3516 2835 3519
rect 3786 3516 3792 3528
rect 2823 3488 3792 3516
rect 2823 3485 2835 3488
rect 2777 3479 2835 3485
rect 3786 3476 3792 3488
rect 3844 3476 3850 3528
rect 4525 3519 4583 3525
rect 4525 3516 4537 3519
rect 4356 3488 4537 3516
rect 2685 3451 2743 3457
rect 2685 3417 2697 3451
rect 2731 3448 2743 3451
rect 3050 3448 3056 3460
rect 2731 3420 3056 3448
rect 2731 3417 2743 3420
rect 2685 3411 2743 3417
rect 3050 3408 3056 3420
rect 3108 3408 3114 3460
rect 4246 3408 4252 3460
rect 4304 3448 4310 3460
rect 4356 3448 4384 3488
rect 4525 3485 4537 3488
rect 4571 3485 4583 3519
rect 4525 3479 4583 3485
rect 5261 3519 5319 3525
rect 5261 3485 5273 3519
rect 5307 3516 5319 3519
rect 5905 3519 5963 3525
rect 5307 3488 5672 3516
rect 5307 3485 5319 3488
rect 5261 3479 5319 3485
rect 4304 3420 4384 3448
rect 4304 3408 4310 3420
rect 4430 3408 4436 3460
rect 4488 3448 4494 3460
rect 5534 3448 5540 3460
rect 4488 3420 5540 3448
rect 4488 3408 4494 3420
rect 5534 3408 5540 3420
rect 5592 3408 5598 3460
rect 5644 3448 5672 3488
rect 5905 3485 5917 3519
rect 5951 3516 5963 3519
rect 6086 3516 6092 3528
rect 5951 3488 6092 3516
rect 5951 3485 5963 3488
rect 5905 3479 5963 3485
rect 6086 3476 6092 3488
rect 6144 3476 6150 3528
rect 6733 3519 6791 3525
rect 6733 3485 6745 3519
rect 6779 3485 6791 3519
rect 6733 3479 6791 3485
rect 5718 3448 5724 3460
rect 5631 3420 5724 3448
rect 5718 3408 5724 3420
rect 5776 3448 5782 3460
rect 6638 3448 6644 3460
rect 5776 3420 6644 3448
rect 5776 3408 5782 3420
rect 6638 3408 6644 3420
rect 6696 3408 6702 3460
rect 6748 3448 6776 3479
rect 8202 3476 8208 3528
rect 8260 3516 8266 3528
rect 8481 3519 8539 3525
rect 8481 3516 8493 3519
rect 8260 3488 8493 3516
rect 8260 3476 8266 3488
rect 8481 3485 8493 3488
rect 8527 3485 8539 3519
rect 8481 3479 8539 3485
rect 11514 3476 11520 3528
rect 11572 3516 11578 3528
rect 11701 3519 11759 3525
rect 11701 3516 11713 3519
rect 11572 3488 11713 3516
rect 11572 3476 11578 3488
rect 11701 3485 11713 3488
rect 11747 3516 11759 3519
rect 11974 3516 11980 3528
rect 11747 3488 11980 3516
rect 11747 3485 11759 3488
rect 11701 3479 11759 3485
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3516 13599 3519
rect 13630 3516 13636 3528
rect 13587 3488 13636 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 13630 3476 13636 3488
rect 13688 3476 13694 3528
rect 13814 3516 13820 3528
rect 13775 3488 13820 3516
rect 13814 3476 13820 3488
rect 13872 3476 13878 3528
rect 14550 3476 14556 3528
rect 14608 3516 14614 3528
rect 15289 3519 15347 3525
rect 15289 3516 15301 3519
rect 14608 3488 15301 3516
rect 14608 3476 14614 3488
rect 15289 3485 15301 3488
rect 15335 3485 15347 3519
rect 17129 3519 17187 3525
rect 17129 3516 17141 3519
rect 15289 3479 15347 3485
rect 16868 3488 17141 3516
rect 6822 3448 6828 3460
rect 6735 3420 6828 3448
rect 6822 3408 6828 3420
rect 6880 3448 6886 3460
rect 8941 3451 8999 3457
rect 8941 3448 8953 3451
rect 6880 3420 8953 3448
rect 6880 3408 6886 3420
rect 8941 3417 8953 3420
rect 8987 3417 8999 3451
rect 8941 3411 8999 3417
rect 12526 3408 12532 3460
rect 12584 3448 12590 3460
rect 12897 3451 12955 3457
rect 12897 3448 12909 3451
rect 12584 3420 12909 3448
rect 12584 3408 12590 3420
rect 12897 3417 12909 3420
rect 12943 3417 12955 3451
rect 12897 3411 12955 3417
rect 842 3340 848 3392
rect 900 3380 906 3392
rect 1762 3380 1768 3392
rect 900 3352 1768 3380
rect 900 3340 906 3352
rect 1762 3340 1768 3352
rect 1820 3380 1826 3392
rect 1857 3383 1915 3389
rect 1857 3380 1869 3383
rect 1820 3352 1869 3380
rect 1820 3340 1826 3352
rect 1857 3349 1869 3352
rect 1903 3380 1915 3383
rect 2225 3383 2283 3389
rect 2225 3380 2237 3383
rect 1903 3352 2237 3380
rect 1903 3349 1915 3352
rect 1857 3343 1915 3349
rect 2225 3349 2237 3352
rect 2271 3349 2283 3383
rect 2225 3343 2283 3349
rect 2574 3383 2632 3389
rect 2574 3349 2586 3383
rect 2620 3380 2632 3383
rect 3418 3380 3424 3392
rect 2620 3352 3424 3380
rect 2620 3349 2632 3352
rect 2574 3343 2632 3349
rect 3418 3340 3424 3352
rect 3476 3340 3482 3392
rect 4614 3380 4620 3392
rect 4575 3352 4620 3380
rect 4614 3340 4620 3352
rect 4672 3340 4678 3392
rect 4982 3380 4988 3392
rect 4943 3352 4988 3380
rect 4982 3340 4988 3352
rect 5040 3340 5046 3392
rect 6270 3340 6276 3392
rect 6328 3380 6334 3392
rect 8754 3380 8760 3392
rect 6328 3352 8760 3380
rect 6328 3340 6334 3352
rect 8754 3340 8760 3352
rect 8812 3340 8818 3392
rect 12621 3383 12679 3389
rect 12621 3349 12633 3383
rect 12667 3380 12679 3383
rect 12802 3380 12808 3392
rect 12667 3352 12808 3380
rect 12667 3349 12679 3352
rect 12621 3343 12679 3349
rect 12802 3340 12808 3352
rect 12860 3340 12866 3392
rect 16666 3340 16672 3392
rect 16724 3380 16730 3392
rect 16868 3389 16896 3488
rect 17129 3485 17141 3488
rect 17175 3485 17187 3519
rect 17129 3479 17187 3485
rect 17773 3519 17831 3525
rect 17773 3485 17785 3519
rect 17819 3516 17831 3519
rect 18414 3516 18420 3528
rect 17819 3488 18420 3516
rect 17819 3485 17831 3488
rect 17773 3479 17831 3485
rect 18414 3476 18420 3488
rect 18472 3476 18478 3528
rect 18524 3516 18552 3556
rect 20809 3553 20821 3587
rect 20855 3584 20867 3587
rect 20898 3584 20904 3596
rect 20855 3556 20904 3584
rect 20855 3553 20867 3556
rect 20809 3547 20867 3553
rect 20898 3544 20904 3556
rect 20956 3544 20962 3596
rect 22554 3584 22560 3596
rect 22515 3556 22560 3584
rect 22554 3544 22560 3556
rect 22612 3544 22618 3596
rect 22738 3544 22744 3596
rect 22796 3584 22802 3596
rect 23474 3584 23480 3596
rect 22796 3556 23480 3584
rect 22796 3544 22802 3556
rect 23474 3544 23480 3556
rect 23532 3584 23538 3596
rect 23788 3587 23846 3593
rect 23788 3584 23800 3587
rect 23532 3556 23800 3584
rect 23532 3544 23538 3556
rect 23788 3553 23800 3556
rect 23834 3553 23846 3587
rect 23788 3547 23846 3553
rect 24210 3544 24216 3596
rect 24268 3584 24274 3596
rect 24596 3593 24624 3692
rect 24903 3689 24915 3692
rect 24949 3689 24961 3723
rect 24903 3683 24961 3689
rect 24581 3587 24639 3593
rect 24581 3584 24593 3587
rect 24268 3556 24593 3584
rect 24268 3544 24274 3556
rect 24581 3553 24593 3556
rect 24627 3553 24639 3587
rect 24581 3547 24639 3553
rect 24832 3587 24890 3593
rect 24832 3553 24844 3587
rect 24878 3584 24890 3587
rect 24946 3584 24952 3596
rect 24878 3556 24952 3584
rect 24878 3553 24890 3556
rect 24832 3547 24890 3553
rect 24946 3544 24952 3556
rect 25004 3544 25010 3596
rect 18693 3519 18751 3525
rect 18693 3516 18705 3519
rect 18524 3488 18705 3516
rect 18693 3485 18705 3488
rect 18739 3485 18751 3519
rect 18966 3516 18972 3528
rect 18927 3488 18972 3516
rect 18693 3479 18751 3485
rect 18966 3476 18972 3488
rect 19024 3476 19030 3528
rect 16853 3383 16911 3389
rect 16853 3380 16865 3383
rect 16724 3352 16865 3380
rect 16724 3340 16730 3352
rect 16853 3349 16865 3352
rect 16899 3349 16911 3383
rect 16853 3343 16911 3349
rect 17402 3340 17408 3392
rect 17460 3380 17466 3392
rect 21039 3383 21097 3389
rect 21039 3380 21051 3383
rect 17460 3352 21051 3380
rect 17460 3340 17466 3352
rect 21039 3349 21051 3352
rect 21085 3349 21097 3383
rect 21039 3343 21097 3349
rect 23382 3340 23388 3392
rect 23440 3380 23446 3392
rect 23891 3383 23949 3389
rect 23891 3380 23903 3383
rect 23440 3352 23903 3380
rect 23440 3340 23446 3352
rect 23891 3349 23903 3352
rect 23937 3349 23949 3383
rect 23891 3343 23949 3349
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1946 3176 1952 3188
rect 1907 3148 1952 3176
rect 1946 3136 1952 3148
rect 2004 3136 2010 3188
rect 3050 3176 3056 3188
rect 3011 3148 3056 3176
rect 3050 3136 3056 3148
rect 3108 3136 3114 3188
rect 3418 3176 3424 3188
rect 3379 3148 3424 3176
rect 3418 3136 3424 3148
rect 3476 3136 3482 3188
rect 5077 3179 5135 3185
rect 5077 3145 5089 3179
rect 5123 3176 5135 3179
rect 5166 3176 5172 3188
rect 5123 3148 5172 3176
rect 5123 3145 5135 3148
rect 5077 3139 5135 3145
rect 5166 3136 5172 3148
rect 5224 3176 5230 3188
rect 5445 3179 5503 3185
rect 5445 3176 5457 3179
rect 5224 3148 5457 3176
rect 5224 3136 5230 3148
rect 5445 3145 5457 3148
rect 5491 3145 5503 3179
rect 5445 3139 5503 3145
rect 5813 3179 5871 3185
rect 5813 3145 5825 3179
rect 5859 3176 5871 3179
rect 5994 3176 6000 3188
rect 5859 3148 6000 3176
rect 5859 3145 5871 3148
rect 5813 3139 5871 3145
rect 5994 3136 6000 3148
rect 6052 3136 6058 3188
rect 6270 3176 6276 3188
rect 6231 3148 6276 3176
rect 6270 3136 6276 3148
rect 6328 3136 6334 3188
rect 6730 3136 6736 3188
rect 6788 3176 6794 3188
rect 7101 3179 7159 3185
rect 7101 3176 7113 3179
rect 6788 3148 7113 3176
rect 6788 3136 6794 3148
rect 7101 3145 7113 3148
rect 7147 3145 7159 3179
rect 8294 3176 8300 3188
rect 7101 3139 7159 3145
rect 7484 3148 8300 3176
rect 3602 3068 3608 3120
rect 3660 3108 3666 3120
rect 5334 3111 5392 3117
rect 3660 3080 4936 3108
rect 3660 3068 3666 3080
rect 4614 3040 4620 3052
rect 4172 3012 4620 3040
rect 2682 2972 2688 2984
rect 2643 2944 2688 2972
rect 2682 2932 2688 2944
rect 2740 2932 2746 2984
rect 4172 2981 4200 3012
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 4157 2975 4215 2981
rect 4157 2941 4169 2975
rect 4203 2941 4215 2975
rect 4908 2972 4936 3080
rect 5334 3077 5346 3111
rect 5380 3108 5392 3111
rect 6288 3108 6316 3136
rect 5380 3080 6316 3108
rect 5380 3077 5392 3080
rect 5334 3071 5392 3077
rect 4982 3000 4988 3052
rect 5040 3040 5046 3052
rect 5537 3043 5595 3049
rect 5537 3040 5549 3043
rect 5040 3012 5549 3040
rect 5040 3000 5046 3012
rect 5537 3009 5549 3012
rect 5583 3009 5595 3043
rect 5537 3003 5595 3009
rect 6086 3000 6092 3052
rect 6144 3040 6150 3052
rect 7285 3043 7343 3049
rect 7285 3040 7297 3043
rect 6144 3012 7297 3040
rect 6144 3000 6150 3012
rect 7285 3009 7297 3012
rect 7331 3040 7343 3043
rect 7484 3040 7512 3148
rect 8294 3136 8300 3148
rect 8352 3136 8358 3188
rect 9582 3136 9588 3188
rect 9640 3176 9646 3188
rect 9677 3179 9735 3185
rect 9677 3176 9689 3179
rect 9640 3148 9689 3176
rect 9640 3136 9646 3148
rect 9677 3145 9689 3148
rect 9723 3145 9735 3179
rect 9677 3139 9735 3145
rect 9692 3108 9720 3139
rect 9858 3136 9864 3188
rect 9916 3176 9922 3188
rect 9953 3179 10011 3185
rect 9953 3176 9965 3179
rect 9916 3148 9965 3176
rect 9916 3136 9922 3148
rect 9953 3145 9965 3148
rect 9999 3145 10011 3179
rect 10318 3176 10324 3188
rect 10279 3148 10324 3176
rect 9953 3139 10011 3145
rect 10318 3136 10324 3148
rect 10376 3136 10382 3188
rect 11606 3136 11612 3188
rect 11664 3176 11670 3188
rect 11701 3179 11759 3185
rect 11701 3176 11713 3179
rect 11664 3148 11713 3176
rect 11664 3136 11670 3148
rect 11701 3145 11713 3148
rect 11747 3145 11759 3179
rect 13538 3176 13544 3188
rect 13499 3148 13544 3176
rect 11701 3139 11759 3145
rect 10686 3108 10692 3120
rect 9692 3080 10692 3108
rect 10686 3068 10692 3080
rect 10744 3068 10750 3120
rect 11716 3108 11744 3139
rect 13538 3136 13544 3148
rect 13596 3136 13602 3188
rect 14093 3179 14151 3185
rect 14093 3145 14105 3179
rect 14139 3176 14151 3179
rect 14182 3176 14188 3188
rect 14139 3148 14188 3176
rect 14139 3145 14151 3148
rect 14093 3139 14151 3145
rect 14182 3136 14188 3148
rect 14240 3176 14246 3188
rect 14240 3148 14596 3176
rect 14240 3136 14246 3148
rect 14369 3111 14427 3117
rect 14369 3108 14381 3111
rect 11716 3080 14381 3108
rect 14369 3077 14381 3080
rect 14415 3077 14427 3111
rect 14369 3071 14427 3077
rect 7331 3012 7512 3040
rect 8297 3043 8355 3049
rect 7331 3009 7343 3012
rect 7285 3003 7343 3009
rect 8297 3009 8309 3043
rect 8343 3040 8355 3043
rect 8757 3043 8815 3049
rect 8757 3040 8769 3043
rect 8343 3012 8769 3040
rect 8343 3009 8355 3012
rect 8297 3003 8355 3009
rect 8757 3009 8769 3012
rect 8803 3040 8815 3043
rect 8938 3040 8944 3052
rect 8803 3012 8944 3040
rect 8803 3009 8815 3012
rect 8757 3003 8815 3009
rect 8938 3000 8944 3012
rect 8996 3000 9002 3052
rect 10870 3040 10876 3052
rect 10831 3012 10876 3040
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3040 13231 3043
rect 13354 3040 13360 3052
rect 13219 3012 13360 3040
rect 13219 3009 13231 3012
rect 13173 3003 13231 3009
rect 13354 3000 13360 3012
rect 13412 3000 13418 3052
rect 5169 2975 5227 2981
rect 5169 2972 5181 2975
rect 4908 2944 5181 2972
rect 4157 2935 4215 2941
rect 5169 2941 5181 2944
rect 5215 2972 5227 2975
rect 6549 2975 6607 2981
rect 6549 2972 6561 2975
rect 5215 2944 6561 2972
rect 5215 2941 5227 2944
rect 5169 2935 5227 2941
rect 6549 2941 6561 2944
rect 6595 2941 6607 2975
rect 6549 2935 6607 2941
rect 8110 2932 8116 2984
rect 8168 2972 8174 2984
rect 8168 2944 9674 2972
rect 8168 2932 8174 2944
rect 2774 2904 2780 2916
rect 2735 2876 2780 2904
rect 2774 2864 2780 2876
rect 2832 2864 2838 2916
rect 3418 2864 3424 2916
rect 3476 2904 3482 2916
rect 4338 2904 4344 2916
rect 3476 2876 4154 2904
rect 4299 2876 4344 2904
rect 3476 2864 3482 2876
rect 4126 2836 4154 2876
rect 4338 2864 4344 2876
rect 4396 2864 4402 2916
rect 4890 2904 4896 2916
rect 4448 2876 4896 2904
rect 4448 2836 4476 2876
rect 4890 2864 4896 2876
rect 4948 2864 4954 2916
rect 7374 2904 7380 2916
rect 5828 2876 7144 2904
rect 7335 2876 7380 2904
rect 4706 2836 4712 2848
rect 4126 2808 4476 2836
rect 4619 2808 4712 2836
rect 4706 2796 4712 2808
rect 4764 2836 4770 2848
rect 5828 2836 5856 2876
rect 4764 2808 5856 2836
rect 7116 2836 7144 2876
rect 7374 2864 7380 2876
rect 7432 2864 7438 2916
rect 7929 2907 7987 2913
rect 7929 2873 7941 2907
rect 7975 2904 7987 2907
rect 8846 2904 8852 2916
rect 7975 2876 8852 2904
rect 7975 2873 7987 2876
rect 7929 2867 7987 2873
rect 8846 2864 8852 2876
rect 8904 2864 8910 2916
rect 9646 2904 9674 2944
rect 10597 2907 10655 2913
rect 10597 2904 10609 2907
rect 9646 2876 10609 2904
rect 10597 2873 10609 2876
rect 10643 2873 10655 2907
rect 10597 2867 10655 2873
rect 8386 2836 8392 2848
rect 7116 2808 8392 2836
rect 4764 2796 4770 2808
rect 8386 2796 8392 2808
rect 8444 2796 8450 2848
rect 8665 2839 8723 2845
rect 8665 2805 8677 2839
rect 8711 2836 8723 2839
rect 9122 2836 9128 2848
rect 8711 2808 9128 2836
rect 8711 2805 8723 2808
rect 8665 2799 8723 2805
rect 9122 2796 9128 2808
rect 9180 2796 9186 2848
rect 10612 2836 10640 2867
rect 10686 2864 10692 2916
rect 10744 2904 10750 2916
rect 12526 2904 12532 2916
rect 10744 2876 10789 2904
rect 12487 2876 12532 2904
rect 10744 2864 10750 2876
rect 12526 2864 12532 2876
rect 12584 2864 12590 2916
rect 12621 2907 12679 2913
rect 12621 2873 12633 2907
rect 12667 2904 12679 2907
rect 14384 2904 14412 3071
rect 14568 3049 14596 3148
rect 15378 3136 15384 3188
rect 15436 3176 15442 3188
rect 17034 3176 17040 3188
rect 15436 3148 17040 3176
rect 15436 3136 15442 3148
rect 17034 3136 17040 3148
rect 17092 3136 17098 3188
rect 17218 3136 17224 3188
rect 17276 3176 17282 3188
rect 17313 3179 17371 3185
rect 17313 3176 17325 3179
rect 17276 3148 17325 3176
rect 17276 3136 17282 3148
rect 17313 3145 17325 3148
rect 17359 3145 17371 3179
rect 17313 3139 17371 3145
rect 17865 3179 17923 3185
rect 17865 3145 17877 3179
rect 17911 3176 17923 3179
rect 18046 3176 18052 3188
rect 17911 3148 18052 3176
rect 17911 3145 17923 3148
rect 17865 3139 17923 3145
rect 18046 3136 18052 3148
rect 18104 3136 18110 3188
rect 19058 3176 19064 3188
rect 19019 3148 19064 3176
rect 19058 3136 19064 3148
rect 19116 3136 19122 3188
rect 22554 3136 22560 3188
rect 22612 3176 22618 3188
rect 23017 3179 23075 3185
rect 23017 3176 23029 3179
rect 22612 3148 23029 3176
rect 22612 3136 22618 3148
rect 23017 3145 23029 3148
rect 23063 3145 23075 3179
rect 23017 3139 23075 3145
rect 23474 3136 23480 3188
rect 23532 3176 23538 3188
rect 24857 3179 24915 3185
rect 23532 3148 23577 3176
rect 23532 3136 23538 3148
rect 24857 3145 24869 3179
rect 24903 3176 24915 3179
rect 24946 3176 24952 3188
rect 24903 3148 24952 3176
rect 24903 3145 24915 3148
rect 24857 3139 24915 3145
rect 24946 3136 24952 3148
rect 25004 3176 25010 3188
rect 26970 3176 26976 3188
rect 25004 3148 26976 3176
rect 25004 3136 25010 3148
rect 26970 3136 26976 3148
rect 27028 3136 27034 3188
rect 15286 3068 15292 3120
rect 15344 3108 15350 3120
rect 19889 3111 19947 3117
rect 19889 3108 19901 3111
rect 15344 3080 19901 3108
rect 15344 3068 15350 3080
rect 19889 3077 19901 3080
rect 19935 3077 19947 3111
rect 19889 3071 19947 3077
rect 14553 3043 14611 3049
rect 14553 3009 14565 3043
rect 14599 3009 14611 3043
rect 16666 3040 16672 3052
rect 16627 3012 16672 3040
rect 14553 3003 14611 3009
rect 16666 3000 16672 3012
rect 16724 3000 16730 3052
rect 18138 3040 18144 3052
rect 18099 3012 18144 3040
rect 18138 3000 18144 3012
rect 18196 3000 18202 3052
rect 18414 3040 18420 3052
rect 18375 3012 18420 3040
rect 18414 3000 18420 3012
rect 18472 3040 18478 3052
rect 21637 3043 21695 3049
rect 21637 3040 21649 3043
rect 18472 3012 21649 3040
rect 18472 3000 18478 3012
rect 21227 2981 21255 3012
rect 21637 3009 21649 3012
rect 21683 3009 21695 3043
rect 22646 3040 22652 3052
rect 22607 3012 22652 3040
rect 21637 3003 21695 3009
rect 22646 3000 22652 3012
rect 22704 3000 22710 3052
rect 19705 2975 19763 2981
rect 19705 2972 19717 2975
rect 19444 2944 19717 2972
rect 14874 2907 14932 2913
rect 14874 2904 14886 2907
rect 12667 2876 13814 2904
rect 14384 2876 14886 2904
rect 12667 2873 12679 2876
rect 12621 2867 12679 2873
rect 11146 2836 11152 2848
rect 10612 2808 11152 2836
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 12253 2839 12311 2845
rect 12253 2805 12265 2839
rect 12299 2836 12311 2839
rect 12636 2836 12664 2867
rect 12299 2808 12664 2836
rect 13786 2836 13814 2876
rect 14874 2873 14886 2876
rect 14920 2904 14932 2907
rect 15749 2907 15807 2913
rect 15749 2904 15761 2907
rect 14920 2876 15761 2904
rect 14920 2873 14932 2876
rect 14874 2867 14932 2873
rect 15749 2873 15761 2876
rect 15795 2873 15807 2907
rect 16390 2904 16396 2916
rect 16351 2876 16396 2904
rect 15749 2867 15807 2873
rect 16390 2864 16396 2876
rect 16448 2864 16454 2916
rect 16485 2907 16543 2913
rect 16485 2873 16497 2907
rect 16531 2904 16543 2907
rect 17862 2904 17868 2916
rect 16531 2876 17868 2904
rect 16531 2873 16543 2876
rect 16485 2867 16543 2873
rect 15286 2836 15292 2848
rect 13786 2808 15292 2836
rect 12299 2805 12311 2808
rect 12253 2799 12311 2805
rect 15286 2796 15292 2808
rect 15344 2796 15350 2848
rect 15378 2796 15384 2848
rect 15436 2836 15442 2848
rect 15473 2839 15531 2845
rect 15473 2836 15485 2839
rect 15436 2808 15485 2836
rect 15436 2796 15442 2808
rect 15473 2805 15485 2808
rect 15519 2805 15531 2839
rect 15473 2799 15531 2805
rect 16209 2839 16267 2845
rect 16209 2805 16221 2839
rect 16255 2836 16267 2839
rect 16500 2836 16528 2867
rect 17862 2864 17868 2876
rect 17920 2864 17926 2916
rect 18233 2907 18291 2913
rect 18233 2873 18245 2907
rect 18279 2873 18291 2907
rect 18233 2867 18291 2873
rect 16255 2808 16528 2836
rect 16255 2805 16267 2808
rect 16209 2799 16267 2805
rect 18046 2796 18052 2848
rect 18104 2836 18110 2848
rect 18248 2836 18276 2867
rect 19444 2848 19472 2944
rect 19705 2941 19717 2944
rect 19751 2941 19763 2975
rect 19705 2935 19763 2941
rect 21212 2975 21270 2981
rect 21212 2941 21224 2975
rect 21258 2941 21270 2975
rect 21212 2935 21270 2941
rect 22256 2975 22314 2981
rect 22256 2941 22268 2975
rect 22302 2972 22314 2975
rect 22664 2972 22692 3000
rect 22302 2944 22692 2972
rect 24121 2975 24179 2981
rect 22302 2941 22314 2944
rect 22256 2935 22314 2941
rect 24121 2941 24133 2975
rect 24167 2972 24179 2975
rect 24264 2975 24322 2981
rect 24264 2972 24276 2975
rect 24167 2944 24276 2972
rect 24167 2941 24179 2944
rect 24121 2935 24179 2941
rect 24264 2941 24276 2944
rect 24310 2972 24322 2975
rect 25774 2972 25780 2984
rect 24310 2944 25780 2972
rect 24310 2941 24322 2944
rect 24264 2935 24322 2941
rect 25774 2932 25780 2944
rect 25832 2932 25838 2984
rect 24351 2907 24409 2913
rect 24351 2904 24363 2907
rect 23446 2876 24363 2904
rect 19426 2836 19432 2848
rect 18104 2808 18276 2836
rect 19387 2808 19432 2836
rect 18104 2796 18110 2808
rect 19426 2796 19432 2808
rect 19484 2796 19490 2848
rect 20898 2836 20904 2848
rect 20859 2808 20904 2836
rect 20898 2796 20904 2808
rect 20956 2796 20962 2848
rect 20990 2796 20996 2848
rect 21048 2836 21054 2848
rect 21315 2839 21373 2845
rect 21315 2836 21327 2839
rect 21048 2808 21327 2836
rect 21048 2796 21054 2808
rect 21315 2805 21327 2808
rect 21361 2805 21373 2839
rect 21315 2799 21373 2805
rect 21450 2796 21456 2848
rect 21508 2836 21514 2848
rect 22327 2839 22385 2845
rect 22327 2836 22339 2839
rect 21508 2808 22339 2836
rect 21508 2796 21514 2808
rect 22327 2805 22339 2808
rect 22373 2805 22385 2839
rect 22327 2799 22385 2805
rect 23106 2796 23112 2848
rect 23164 2836 23170 2848
rect 23446 2836 23474 2876
rect 24351 2873 24363 2876
rect 24397 2873 24409 2907
rect 24351 2867 24409 2873
rect 23164 2808 23474 2836
rect 23164 2796 23170 2808
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1854 2632 1860 2644
rect 1815 2604 1860 2632
rect 1854 2592 1860 2604
rect 1912 2592 1918 2644
rect 2774 2592 2780 2644
rect 2832 2632 2838 2644
rect 4387 2635 4445 2641
rect 2832 2604 4154 2632
rect 2832 2592 2838 2604
rect 2222 2564 2228 2576
rect 2183 2536 2228 2564
rect 2222 2524 2228 2536
rect 2280 2524 2286 2576
rect 3234 2564 3240 2576
rect 3068 2536 3240 2564
rect 1464 2499 1522 2505
rect 1464 2465 1476 2499
rect 1510 2496 1522 2499
rect 2240 2496 2268 2524
rect 3068 2505 3096 2536
rect 3234 2524 3240 2536
rect 3292 2524 3298 2576
rect 4126 2564 4154 2604
rect 4387 2601 4399 2635
rect 4433 2632 4445 2635
rect 4522 2632 4528 2644
rect 4433 2604 4528 2632
rect 4433 2601 4445 2604
rect 4387 2595 4445 2601
rect 4522 2592 4528 2604
rect 4580 2592 4586 2644
rect 5074 2632 5080 2644
rect 5035 2604 5080 2632
rect 5074 2592 5080 2604
rect 5132 2632 5138 2644
rect 5902 2632 5908 2644
rect 5132 2604 5304 2632
rect 5863 2604 5908 2632
rect 5132 2592 5138 2604
rect 5166 2564 5172 2576
rect 4126 2536 5172 2564
rect 5166 2524 5172 2536
rect 5224 2524 5230 2576
rect 5276 2573 5304 2604
rect 5902 2592 5908 2604
rect 5960 2592 5966 2644
rect 6089 2635 6147 2641
rect 6089 2601 6101 2635
rect 6135 2632 6147 2635
rect 6365 2635 6423 2641
rect 6365 2632 6377 2635
rect 6135 2604 6377 2632
rect 6135 2601 6147 2604
rect 6089 2595 6147 2601
rect 6365 2601 6377 2604
rect 6411 2632 6423 2635
rect 6914 2632 6920 2644
rect 6411 2604 6920 2632
rect 6411 2601 6423 2604
rect 6365 2595 6423 2601
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 7239 2635 7297 2641
rect 7239 2601 7251 2635
rect 7285 2632 7297 2635
rect 8110 2632 8116 2644
rect 7285 2604 8116 2632
rect 7285 2601 7297 2604
rect 7239 2595 7297 2601
rect 8110 2592 8116 2604
rect 8168 2592 8174 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 8220 2604 9137 2632
rect 8220 2576 8248 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 9125 2595 9183 2601
rect 10686 2592 10692 2644
rect 10744 2632 10750 2644
rect 10781 2635 10839 2641
rect 10781 2632 10793 2635
rect 10744 2604 10793 2632
rect 10744 2592 10750 2604
rect 10781 2601 10793 2604
rect 10827 2601 10839 2635
rect 11146 2632 11152 2644
rect 11107 2604 11152 2632
rect 10781 2595 10839 2601
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 11609 2635 11667 2641
rect 11609 2601 11621 2635
rect 11655 2601 11667 2635
rect 11974 2632 11980 2644
rect 11935 2604 11980 2632
rect 11609 2595 11667 2601
rect 5261 2567 5319 2573
rect 5261 2533 5273 2567
rect 5307 2533 5319 2567
rect 5261 2527 5319 2533
rect 5350 2524 5356 2576
rect 5408 2564 5414 2576
rect 7929 2567 7987 2573
rect 7929 2564 7941 2567
rect 5408 2536 7941 2564
rect 5408 2524 5414 2536
rect 7929 2533 7941 2536
rect 7975 2533 7987 2567
rect 8202 2564 8208 2576
rect 8163 2536 8208 2564
rect 7929 2527 7987 2533
rect 1510 2468 2268 2496
rect 3053 2499 3111 2505
rect 1510 2465 1522 2468
rect 1464 2459 1522 2465
rect 3053 2465 3065 2499
rect 3099 2465 3111 2499
rect 3053 2459 3111 2465
rect 3145 2499 3203 2505
rect 3145 2465 3157 2499
rect 3191 2496 3203 2499
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 3191 2468 4077 2496
rect 3191 2465 3203 2468
rect 3145 2459 3203 2465
rect 4065 2465 4077 2468
rect 4111 2465 4123 2499
rect 4065 2459 4123 2465
rect 4316 2499 4374 2505
rect 4316 2465 4328 2499
rect 4362 2496 4374 2499
rect 4801 2499 4859 2505
rect 4801 2496 4813 2499
rect 4362 2468 4813 2496
rect 4362 2465 4374 2468
rect 4316 2459 4374 2465
rect 4801 2465 4813 2468
rect 4847 2496 4859 2499
rect 6086 2496 6092 2508
rect 4847 2468 6092 2496
rect 4847 2465 4859 2468
rect 4801 2459 4859 2465
rect 6086 2456 6092 2468
rect 6144 2456 6150 2508
rect 7168 2499 7226 2505
rect 7168 2465 7180 2499
rect 7214 2496 7226 2499
rect 7650 2496 7656 2508
rect 7214 2468 7656 2496
rect 7214 2465 7226 2468
rect 7168 2459 7226 2465
rect 7650 2456 7656 2468
rect 7708 2456 7714 2508
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2428 1731 2431
rect 1719 2400 5580 2428
rect 1719 2397 1731 2400
rect 1673 2391 1731 2397
rect 2590 2320 2596 2372
rect 2648 2360 2654 2372
rect 3421 2363 3479 2369
rect 3421 2360 3433 2363
rect 2648 2332 3433 2360
rect 2648 2320 2654 2332
rect 3421 2329 3433 2332
rect 3467 2329 3479 2363
rect 3421 2323 3479 2329
rect 4065 2363 4123 2369
rect 4065 2329 4077 2363
rect 4111 2360 4123 2363
rect 4798 2360 4804 2372
rect 4111 2332 4804 2360
rect 4111 2329 4123 2332
rect 4065 2323 4123 2329
rect 4798 2320 4804 2332
rect 4856 2320 4862 2372
rect 5552 2360 5580 2400
rect 5626 2388 5632 2440
rect 5684 2428 5690 2440
rect 6641 2431 6699 2437
rect 6641 2428 6653 2431
rect 5684 2400 6653 2428
rect 5684 2388 5690 2400
rect 6641 2397 6653 2400
rect 6687 2397 6699 2431
rect 7944 2428 7972 2527
rect 8202 2524 8208 2536
rect 8260 2524 8266 2576
rect 8294 2524 8300 2576
rect 8352 2564 8358 2576
rect 9490 2564 9496 2576
rect 8352 2536 8397 2564
rect 9451 2536 9496 2564
rect 8352 2524 8358 2536
rect 9490 2524 9496 2536
rect 9548 2564 9554 2576
rect 9953 2567 10011 2573
rect 9953 2564 9965 2567
rect 9548 2536 9965 2564
rect 9548 2524 9554 2536
rect 9953 2533 9965 2536
rect 9999 2533 10011 2567
rect 9953 2527 10011 2533
rect 10505 2567 10563 2573
rect 10505 2533 10517 2567
rect 10551 2564 10563 2567
rect 10870 2564 10876 2576
rect 10551 2536 10876 2564
rect 10551 2533 10563 2536
rect 10505 2527 10563 2533
rect 10870 2524 10876 2536
rect 10928 2524 10934 2576
rect 11624 2564 11652 2595
rect 11974 2592 11980 2604
rect 12032 2592 12038 2644
rect 12728 2604 13814 2632
rect 12728 2564 12756 2604
rect 11624 2536 12756 2564
rect 12802 2524 12808 2576
rect 12860 2564 12866 2576
rect 13354 2564 13360 2576
rect 12860 2536 12905 2564
rect 13315 2536 13360 2564
rect 12860 2524 12866 2536
rect 13354 2524 13360 2536
rect 13412 2524 13418 2576
rect 13786 2564 13814 2604
rect 14550 2592 14556 2644
rect 14608 2632 14614 2644
rect 14829 2635 14887 2641
rect 14829 2632 14841 2635
rect 14608 2604 14841 2632
rect 14608 2592 14614 2604
rect 14829 2601 14841 2604
rect 14875 2601 14887 2635
rect 18138 2632 18144 2644
rect 14829 2595 14887 2601
rect 15672 2604 17816 2632
rect 18099 2604 18144 2632
rect 14642 2564 14648 2576
rect 13786 2536 14648 2564
rect 14642 2524 14648 2536
rect 14700 2524 14706 2576
rect 15289 2567 15347 2573
rect 15289 2533 15301 2567
rect 15335 2564 15347 2567
rect 15378 2564 15384 2576
rect 15335 2536 15384 2564
rect 15335 2533 15347 2536
rect 15289 2527 15347 2533
rect 15378 2524 15384 2536
rect 15436 2564 15442 2576
rect 15672 2573 15700 2604
rect 15657 2567 15715 2573
rect 15657 2564 15669 2567
rect 15436 2536 15669 2564
rect 15436 2524 15442 2536
rect 15657 2533 15669 2536
rect 15703 2533 15715 2567
rect 15657 2527 15715 2533
rect 16209 2567 16267 2573
rect 16209 2533 16221 2567
rect 16255 2564 16267 2567
rect 16666 2564 16672 2576
rect 16255 2536 16672 2564
rect 16255 2533 16267 2536
rect 16209 2527 16267 2533
rect 16666 2524 16672 2536
rect 16724 2524 16730 2576
rect 16945 2567 17003 2573
rect 16945 2533 16957 2567
rect 16991 2564 17003 2567
rect 17402 2564 17408 2576
rect 16991 2536 17408 2564
rect 16991 2533 17003 2536
rect 16945 2527 17003 2533
rect 8846 2456 8852 2508
rect 8904 2496 8910 2508
rect 9674 2496 9680 2508
rect 8904 2468 9680 2496
rect 8904 2456 8910 2468
rect 9674 2456 9680 2468
rect 9732 2456 9738 2508
rect 11422 2496 11428 2508
rect 11383 2468 11428 2496
rect 11422 2456 11428 2468
rect 11480 2456 11486 2508
rect 13906 2456 13912 2508
rect 13964 2496 13970 2508
rect 14185 2499 14243 2505
rect 14185 2496 14197 2499
rect 13964 2468 14197 2496
rect 13964 2456 13970 2468
rect 14185 2465 14197 2468
rect 14231 2465 14243 2499
rect 14185 2459 14243 2465
rect 8294 2428 8300 2440
rect 7944 2400 8300 2428
rect 6641 2391 6699 2397
rect 8294 2388 8300 2400
rect 8352 2388 8358 2440
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 8680 2400 9873 2428
rect 8680 2360 8708 2400
rect 9861 2397 9873 2400
rect 9907 2428 9919 2431
rect 12713 2431 12771 2437
rect 9907 2400 12664 2428
rect 9907 2397 9919 2400
rect 9861 2391 9919 2397
rect 5552 2332 8708 2360
rect 12636 2360 12664 2400
rect 12713 2397 12725 2431
rect 12759 2428 12771 2431
rect 13449 2431 13507 2437
rect 13449 2428 13461 2431
rect 12759 2400 13461 2428
rect 12759 2397 12771 2400
rect 12713 2391 12771 2397
rect 13449 2397 13461 2400
rect 13495 2397 13507 2431
rect 13449 2391 13507 2397
rect 14001 2363 14059 2369
rect 14001 2360 14013 2363
rect 12636 2332 14013 2360
rect 14001 2329 14013 2332
rect 14047 2329 14059 2363
rect 14001 2323 14059 2329
rect 3881 2295 3939 2301
rect 3881 2261 3893 2295
rect 3927 2292 3939 2295
rect 4430 2292 4436 2304
rect 3927 2264 4436 2292
rect 3927 2261 3939 2264
rect 3881 2255 3939 2261
rect 4430 2252 4436 2264
rect 4488 2292 4494 2304
rect 5399 2295 5457 2301
rect 5399 2292 5411 2295
rect 4488 2264 5411 2292
rect 4488 2252 4494 2264
rect 5399 2261 5411 2264
rect 5445 2261 5457 2295
rect 5399 2255 5457 2261
rect 5537 2295 5595 2301
rect 5537 2261 5549 2295
rect 5583 2292 5595 2295
rect 6089 2295 6147 2301
rect 6089 2292 6101 2295
rect 5583 2264 6101 2292
rect 5583 2261 5595 2264
rect 5537 2255 5595 2261
rect 6089 2261 6101 2264
rect 6135 2261 6147 2295
rect 7650 2292 7656 2304
rect 7611 2264 7656 2292
rect 6089 2255 6147 2261
rect 7650 2252 7656 2264
rect 7708 2252 7714 2304
rect 12437 2295 12495 2301
rect 12437 2261 12449 2295
rect 12483 2292 12495 2295
rect 12802 2292 12808 2304
rect 12483 2264 12808 2292
rect 12483 2261 12495 2264
rect 12437 2255 12495 2261
rect 12802 2252 12808 2264
rect 12860 2252 12866 2304
rect 13449 2295 13507 2301
rect 13449 2261 13461 2295
rect 13495 2292 13507 2295
rect 13722 2292 13728 2304
rect 13495 2264 13728 2292
rect 13495 2261 13507 2264
rect 13449 2255 13507 2261
rect 13722 2252 13728 2264
rect 13780 2252 13786 2304
rect 14200 2292 14228 2459
rect 16390 2456 16396 2508
rect 16448 2496 16454 2508
rect 16960 2496 16988 2527
rect 17402 2524 17408 2536
rect 17460 2524 17466 2576
rect 16448 2468 16988 2496
rect 16448 2456 16454 2468
rect 17034 2456 17040 2508
rect 17092 2496 17098 2508
rect 17788 2505 17816 2604
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 20533 2635 20591 2641
rect 20533 2601 20545 2635
rect 20579 2632 20591 2635
rect 20990 2632 20996 2644
rect 20579 2604 20996 2632
rect 20579 2601 20591 2604
rect 20533 2595 20591 2601
rect 17862 2524 17868 2576
rect 17920 2564 17926 2576
rect 18325 2567 18383 2573
rect 18325 2564 18337 2567
rect 17920 2536 18337 2564
rect 17920 2524 17926 2536
rect 18325 2533 18337 2536
rect 18371 2533 18383 2567
rect 18325 2527 18383 2533
rect 17773 2499 17831 2505
rect 17092 2468 17137 2496
rect 17092 2456 17098 2468
rect 17773 2465 17785 2499
rect 17819 2496 17831 2499
rect 18417 2499 18475 2505
rect 18417 2496 18429 2499
rect 17819 2468 18429 2496
rect 17819 2465 17831 2468
rect 17773 2459 17831 2465
rect 18417 2465 18429 2468
rect 18463 2465 18475 2499
rect 18417 2459 18475 2465
rect 19889 2499 19947 2505
rect 19889 2465 19901 2499
rect 19935 2496 19947 2499
rect 20548 2496 20576 2595
rect 20990 2592 20996 2604
rect 21048 2592 21054 2644
rect 23382 2632 23388 2644
rect 23343 2604 23388 2632
rect 23382 2592 23388 2604
rect 23440 2592 23446 2644
rect 19935 2468 20576 2496
rect 19935 2465 19947 2468
rect 19889 2459 19947 2465
rect 20714 2456 20720 2508
rect 20772 2496 20778 2508
rect 21212 2499 21270 2505
rect 21212 2496 21224 2499
rect 20772 2468 21224 2496
rect 20772 2456 20778 2468
rect 21212 2465 21224 2468
rect 21258 2496 21270 2499
rect 21637 2499 21695 2505
rect 21637 2496 21649 2499
rect 21258 2468 21649 2496
rect 21258 2465 21270 2468
rect 21212 2459 21270 2465
rect 21637 2465 21649 2468
rect 21683 2465 21695 2499
rect 21637 2459 21695 2465
rect 22741 2499 22799 2505
rect 22741 2465 22753 2499
rect 22787 2496 22799 2499
rect 23400 2496 23428 2592
rect 22787 2468 23428 2496
rect 22787 2465 22799 2468
rect 22741 2459 22799 2465
rect 15554 2431 15612 2437
rect 15554 2397 15566 2431
rect 15600 2428 15612 2431
rect 16022 2428 16028 2440
rect 15600 2400 16028 2428
rect 15600 2397 15612 2400
rect 15554 2391 15612 2397
rect 16022 2388 16028 2400
rect 16080 2428 16086 2440
rect 16485 2431 16543 2437
rect 16485 2428 16497 2431
rect 16080 2400 16497 2428
rect 16080 2388 16086 2400
rect 16485 2397 16497 2400
rect 16531 2397 16543 2431
rect 19705 2431 19763 2437
rect 19705 2428 19717 2431
rect 16485 2391 16543 2397
rect 16592 2400 19717 2428
rect 14369 2363 14427 2369
rect 14369 2329 14381 2363
rect 14415 2360 14427 2363
rect 15378 2360 15384 2372
rect 14415 2332 15384 2360
rect 14415 2329 14427 2332
rect 14369 2323 14427 2329
rect 15378 2320 15384 2332
rect 15436 2320 15442 2372
rect 16592 2292 16620 2400
rect 19705 2397 19717 2400
rect 19751 2397 19763 2431
rect 19705 2391 19763 2397
rect 17221 2363 17279 2369
rect 17221 2329 17233 2363
rect 17267 2360 17279 2363
rect 18138 2360 18144 2372
rect 17267 2332 18144 2360
rect 17267 2329 17279 2332
rect 17221 2323 17279 2329
rect 18138 2320 18144 2332
rect 18196 2320 18202 2372
rect 20073 2363 20131 2369
rect 20073 2329 20085 2363
rect 20119 2360 20131 2363
rect 22738 2360 22744 2372
rect 20119 2332 22744 2360
rect 20119 2329 20131 2332
rect 20073 2323 20131 2329
rect 22738 2320 22744 2332
rect 22796 2320 22802 2372
rect 22925 2363 22983 2369
rect 22925 2329 22937 2363
rect 22971 2360 22983 2363
rect 23658 2360 23664 2372
rect 22971 2332 23664 2360
rect 22971 2329 22983 2332
rect 22925 2323 22983 2329
rect 23658 2320 23664 2332
rect 23716 2320 23722 2372
rect 14200 2264 16620 2292
rect 17034 2252 17040 2304
rect 17092 2292 17098 2304
rect 19337 2295 19395 2301
rect 19337 2292 19349 2295
rect 17092 2264 19349 2292
rect 17092 2252 17098 2264
rect 19337 2261 19349 2264
rect 19383 2261 19395 2295
rect 19337 2255 19395 2261
rect 19794 2252 19800 2304
rect 19852 2292 19858 2304
rect 21315 2295 21373 2301
rect 21315 2292 21327 2295
rect 19852 2264 21327 2292
rect 19852 2252 19858 2264
rect 21315 2261 21327 2264
rect 21361 2261 21373 2295
rect 21315 2255 21373 2261
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 7650 1504 7656 1556
rect 7708 1544 7714 1556
rect 10686 1544 10692 1556
rect 7708 1516 10692 1544
rect 7708 1504 7714 1516
rect 10686 1504 10692 1516
rect 10744 1504 10750 1556
rect 17310 76 17316 128
rect 17368 116 17374 128
rect 19150 116 19156 128
rect 17368 88 19156 116
rect 17368 76 17374 88
rect 19150 76 19156 88
rect 19208 76 19214 128
<< via1 >>
rect 20 27480 72 27532
rect 1032 27480 1084 27532
rect 3148 27480 3200 27532
rect 3976 27480 4028 27532
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 6092 24284 6144 24336
rect 6000 24148 6052 24200
rect 6644 24148 6696 24200
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 5264 23851 5316 23860
rect 5264 23817 5273 23851
rect 5273 23817 5307 23851
rect 5307 23817 5316 23851
rect 5264 23808 5316 23817
rect 6000 23740 6052 23792
rect 1032 23604 1084 23656
rect 5264 23604 5316 23656
rect 9588 23808 9640 23860
rect 18236 23808 18288 23860
rect 20352 23808 20404 23860
rect 22468 23808 22520 23860
rect 25136 23851 25188 23860
rect 25136 23817 25145 23851
rect 25145 23817 25179 23851
rect 25179 23817 25188 23851
rect 25136 23808 25188 23817
rect 13912 23604 13964 23656
rect 16028 23647 16080 23656
rect 16028 23613 16037 23647
rect 16037 23613 16071 23647
rect 16071 23613 16080 23647
rect 16028 23604 16080 23613
rect 18328 23647 18380 23656
rect 18328 23613 18337 23647
rect 18337 23613 18371 23647
rect 18371 23613 18380 23647
rect 18328 23604 18380 23613
rect 24676 23740 24728 23792
rect 3792 23536 3844 23588
rect 19340 23536 19392 23588
rect 25136 23604 25188 23656
rect 6092 23468 6144 23520
rect 7012 23511 7064 23520
rect 7012 23477 7021 23511
rect 7021 23477 7055 23511
rect 7055 23477 7064 23511
rect 7012 23468 7064 23477
rect 8116 23468 8168 23520
rect 13820 23468 13872 23520
rect 19432 23468 19484 23520
rect 22744 23468 22796 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 112 23128 164 23180
rect 1584 23128 1636 23180
rect 5356 23171 5408 23180
rect 5356 23137 5374 23171
rect 5374 23137 5408 23171
rect 7472 23264 7524 23316
rect 11704 23264 11756 23316
rect 16028 23264 16080 23316
rect 6460 23239 6512 23248
rect 6460 23205 6469 23239
rect 6469 23205 6503 23239
rect 6503 23205 6512 23239
rect 6460 23196 6512 23205
rect 8024 23239 8076 23248
rect 8024 23205 8033 23239
rect 8033 23205 8067 23239
rect 8067 23205 8076 23239
rect 8024 23196 8076 23205
rect 5356 23128 5408 23137
rect 11060 23128 11112 23180
rect 15292 23128 15344 23180
rect 6644 23060 6696 23112
rect 7932 23103 7984 23112
rect 7932 23069 7941 23103
rect 7941 23069 7975 23103
rect 7975 23069 7984 23103
rect 7932 23060 7984 23069
rect 8208 23103 8260 23112
rect 8208 23069 8217 23103
rect 8217 23069 8251 23103
rect 8251 23069 8260 23103
rect 8208 23060 8260 23069
rect 2504 22924 2556 22976
rect 5540 22924 5592 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 1584 22763 1636 22772
rect 1584 22729 1593 22763
rect 1593 22729 1627 22763
rect 1627 22729 1636 22763
rect 1584 22720 1636 22729
rect 5356 22763 5408 22772
rect 5356 22729 5365 22763
rect 5365 22729 5399 22763
rect 5399 22729 5408 22763
rect 5356 22720 5408 22729
rect 5540 22720 5592 22772
rect 7932 22720 7984 22772
rect 7012 22584 7064 22636
rect 8208 22584 8260 22636
rect 10876 22516 10928 22568
rect 7380 22491 7432 22500
rect 7380 22457 7389 22491
rect 7389 22457 7423 22491
rect 7423 22457 7432 22491
rect 7380 22448 7432 22457
rect 6000 22380 6052 22432
rect 6460 22380 6512 22432
rect 8024 22380 8076 22432
rect 8208 22423 8260 22432
rect 8208 22389 8217 22423
rect 8217 22389 8251 22423
rect 8251 22389 8260 22423
rect 8208 22380 8260 22389
rect 10968 22423 11020 22432
rect 10968 22389 10977 22423
rect 10977 22389 11011 22423
rect 11011 22389 11020 22423
rect 10968 22380 11020 22389
rect 14004 22380 14056 22432
rect 15292 22423 15344 22432
rect 15292 22389 15301 22423
rect 15301 22389 15335 22423
rect 15335 22389 15344 22423
rect 15292 22380 15344 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 6092 22219 6144 22228
rect 6092 22185 6101 22219
rect 6101 22185 6135 22219
rect 6135 22185 6144 22219
rect 6092 22176 6144 22185
rect 7012 22176 7064 22228
rect 10968 22176 11020 22228
rect 7380 22151 7432 22160
rect 7380 22117 7389 22151
rect 7389 22117 7423 22151
rect 7423 22117 7432 22151
rect 7380 22108 7432 22117
rect 6000 22083 6052 22092
rect 6000 22049 6009 22083
rect 6009 22049 6043 22083
rect 6043 22049 6052 22083
rect 6000 22040 6052 22049
rect 7380 21972 7432 22024
rect 8208 22040 8260 22092
rect 11796 22040 11848 22092
rect 13912 22040 13964 22092
rect 12532 21879 12584 21888
rect 12532 21845 12541 21879
rect 12541 21845 12575 21879
rect 12575 21845 12584 21879
rect 12532 21836 12584 21845
rect 12900 21836 12952 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 11796 21675 11848 21684
rect 11796 21641 11805 21675
rect 11805 21641 11839 21675
rect 11839 21641 11848 21675
rect 11796 21632 11848 21641
rect 13912 21632 13964 21684
rect 15752 21632 15804 21684
rect 12532 21539 12584 21548
rect 12532 21505 12541 21539
rect 12541 21505 12575 21539
rect 12575 21505 12584 21539
rect 12532 21496 12584 21505
rect 1216 21428 1268 21480
rect 11428 21471 11480 21480
rect 11428 21437 11437 21471
rect 11437 21437 11471 21471
rect 11471 21437 11480 21471
rect 11428 21428 11480 21437
rect 11520 21403 11572 21412
rect 5080 21292 5132 21344
rect 6000 21292 6052 21344
rect 7380 21335 7432 21344
rect 7380 21301 7389 21335
rect 7389 21301 7423 21335
rect 7423 21301 7432 21335
rect 7380 21292 7432 21301
rect 11520 21369 11529 21403
rect 11529 21369 11563 21403
rect 11563 21369 11572 21403
rect 11520 21360 11572 21369
rect 11704 21292 11756 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 11520 21020 11572 21072
rect 12900 21063 12952 21072
rect 12900 21029 12909 21063
rect 12909 21029 12943 21063
rect 12943 21029 12952 21063
rect 12900 21020 12952 21029
rect 13084 21020 13136 21072
rect 24676 20952 24728 21004
rect 11336 20927 11388 20936
rect 11336 20893 11345 20927
rect 11345 20893 11379 20927
rect 11379 20893 11388 20927
rect 11336 20884 11388 20893
rect 11796 20927 11848 20936
rect 11796 20893 11805 20927
rect 11805 20893 11839 20927
rect 11839 20893 11848 20927
rect 11796 20884 11848 20893
rect 12532 20816 12584 20868
rect 12992 20816 13044 20868
rect 12716 20791 12768 20800
rect 12716 20757 12725 20791
rect 12725 20757 12759 20791
rect 12759 20757 12768 20791
rect 12716 20748 12768 20757
rect 15660 20748 15712 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 11336 20544 11388 20596
rect 11520 20544 11572 20596
rect 24676 20587 24728 20596
rect 24676 20553 24685 20587
rect 24685 20553 24719 20587
rect 24719 20553 24728 20587
rect 24676 20544 24728 20553
rect 12716 20451 12768 20460
rect 12716 20417 12725 20451
rect 12725 20417 12759 20451
rect 12759 20417 12768 20451
rect 12716 20408 12768 20417
rect 12992 20451 13044 20460
rect 12992 20417 13001 20451
rect 13001 20417 13035 20451
rect 13035 20417 13044 20451
rect 12992 20408 13044 20417
rect 12164 20247 12216 20256
rect 12164 20213 12173 20247
rect 12173 20213 12207 20247
rect 12207 20213 12216 20247
rect 12164 20204 12216 20213
rect 13084 20204 13136 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 12900 20000 12952 20052
rect 13084 19975 13136 19984
rect 13084 19941 13093 19975
rect 13093 19941 13127 19975
rect 13127 19941 13136 19975
rect 13084 19932 13136 19941
rect 12164 19864 12216 19916
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 12164 19116 12216 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 11520 17867 11572 17876
rect 11520 17833 11529 17867
rect 11529 17833 11563 17867
rect 11563 17833 11572 17867
rect 11520 17824 11572 17833
rect 24768 17867 24820 17876
rect 24768 17833 24777 17867
rect 24777 17833 24811 17867
rect 24811 17833 24820 17867
rect 24768 17824 24820 17833
rect 11612 17688 11664 17740
rect 24216 17688 24268 17740
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 11612 16940 11664 16992
rect 24216 16940 24268 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 204 16600 256 16652
rect 6368 16643 6420 16652
rect 6368 16609 6412 16643
rect 6412 16609 6420 16643
rect 8208 16643 8260 16652
rect 6368 16600 6420 16609
rect 8208 16609 8217 16643
rect 8217 16609 8251 16643
rect 8251 16609 8260 16643
rect 8208 16600 8260 16609
rect 7564 16575 7616 16584
rect 7564 16541 7573 16575
rect 7573 16541 7607 16575
rect 7607 16541 7616 16575
rect 7564 16532 7616 16541
rect 7472 16396 7524 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 6368 16235 6420 16244
rect 6368 16201 6377 16235
rect 6377 16201 6411 16235
rect 6411 16201 6420 16235
rect 6368 16192 6420 16201
rect 7932 16124 7984 16176
rect 8484 16056 8536 16108
rect 7104 16031 7156 16040
rect 7104 15997 7113 16031
rect 7113 15997 7147 16031
rect 7147 15997 7156 16031
rect 7104 15988 7156 15997
rect 26424 16192 26476 16244
rect 2412 15852 2464 15904
rect 8208 15920 8260 15972
rect 15660 15852 15712 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 18420 15648 18472 15700
rect 19432 15648 19484 15700
rect 7564 15623 7616 15632
rect 7564 15589 7573 15623
rect 7573 15589 7607 15623
rect 7607 15589 7616 15623
rect 7564 15580 7616 15589
rect 6092 15555 6144 15564
rect 6092 15521 6101 15555
rect 6101 15521 6135 15555
rect 6135 15521 6144 15555
rect 6092 15512 6144 15521
rect 6736 15444 6788 15496
rect 7472 15487 7524 15496
rect 7472 15453 7481 15487
rect 7481 15453 7515 15487
rect 7515 15453 7524 15487
rect 7472 15444 7524 15453
rect 7932 15487 7984 15496
rect 7932 15453 7941 15487
rect 7941 15453 7975 15487
rect 7975 15453 7984 15487
rect 7932 15444 7984 15453
rect 7104 15308 7156 15360
rect 8300 15308 8352 15360
rect 8484 15351 8536 15360
rect 8484 15317 8493 15351
rect 8493 15317 8527 15351
rect 8527 15317 8536 15351
rect 8484 15308 8536 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 6092 15147 6144 15156
rect 6092 15113 6101 15147
rect 6101 15113 6135 15147
rect 6135 15113 6144 15147
rect 6092 15104 6144 15113
rect 7564 15104 7616 15156
rect 14188 15147 14240 15156
rect 14188 15113 14197 15147
rect 14197 15113 14231 15147
rect 14231 15113 14240 15147
rect 14188 15104 14240 15113
rect 24768 15147 24820 15156
rect 24768 15113 24777 15147
rect 24777 15113 24811 15147
rect 24811 15113 24820 15147
rect 24768 15104 24820 15113
rect 8300 15079 8352 15088
rect 8300 15045 8309 15079
rect 8309 15045 8343 15079
rect 8343 15045 8352 15079
rect 8300 15036 8352 15045
rect 7472 14968 7524 15020
rect 24492 15011 24544 15020
rect 24492 14977 24501 15011
rect 24501 14977 24535 15011
rect 24535 14977 24544 15011
rect 24492 14968 24544 14977
rect 9128 14943 9180 14952
rect 9128 14909 9137 14943
rect 9137 14909 9171 14943
rect 9171 14909 9180 14943
rect 9128 14900 9180 14909
rect 8024 14832 8076 14884
rect 6184 14764 6236 14816
rect 6276 14764 6328 14816
rect 7012 14807 7064 14816
rect 7012 14773 7021 14807
rect 7021 14773 7055 14807
rect 7055 14773 7064 14807
rect 7012 14764 7064 14773
rect 15844 14764 15896 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 6184 14560 6236 14612
rect 8576 14560 8628 14612
rect 7012 14492 7064 14544
rect 8392 14492 8444 14544
rect 9128 14492 9180 14544
rect 2412 14424 2464 14476
rect 9680 14467 9732 14476
rect 9680 14433 9689 14467
rect 9689 14433 9723 14467
rect 9723 14433 9732 14467
rect 9680 14424 9732 14433
rect 10140 14467 10192 14476
rect 10140 14433 10149 14467
rect 10149 14433 10183 14467
rect 10183 14433 10192 14467
rect 10140 14424 10192 14433
rect 24676 14424 24728 14476
rect 6552 14356 6604 14408
rect 7472 14356 7524 14408
rect 7932 14399 7984 14408
rect 7932 14365 7941 14399
rect 7941 14365 7975 14399
rect 7975 14365 7984 14399
rect 7932 14356 7984 14365
rect 8300 14399 8352 14408
rect 8300 14365 8309 14399
rect 8309 14365 8343 14399
rect 8343 14365 8352 14399
rect 8300 14356 8352 14365
rect 1584 14331 1636 14340
rect 1584 14297 1593 14331
rect 1593 14297 1627 14331
rect 1627 14297 1636 14331
rect 1584 14288 1636 14297
rect 7380 14288 7432 14340
rect 8024 14288 8076 14340
rect 22008 14220 22060 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 2412 14059 2464 14068
rect 2412 14025 2421 14059
rect 2421 14025 2455 14059
rect 2455 14025 2464 14059
rect 2412 14016 2464 14025
rect 8392 14016 8444 14068
rect 11428 14059 11480 14068
rect 11428 14025 11437 14059
rect 11437 14025 11471 14059
rect 11471 14025 11480 14059
rect 11428 14016 11480 14025
rect 24676 14059 24728 14068
rect 24676 14025 24685 14059
rect 24685 14025 24719 14059
rect 24719 14025 24728 14059
rect 24676 14016 24728 14025
rect 20 13880 72 13932
rect 4252 13880 4304 13932
rect 8760 13923 8812 13932
rect 8760 13889 8769 13923
rect 8769 13889 8803 13923
rect 8803 13889 8812 13923
rect 8760 13880 8812 13889
rect 10968 13880 11020 13932
rect 1676 13812 1728 13864
rect 5356 13855 5408 13864
rect 2964 13787 3016 13796
rect 2964 13753 2973 13787
rect 2973 13753 3007 13787
rect 3007 13753 3016 13787
rect 2964 13744 3016 13753
rect 1584 13719 1636 13728
rect 1584 13685 1593 13719
rect 1593 13685 1627 13719
rect 1627 13685 1636 13719
rect 1584 13676 1636 13685
rect 2688 13676 2740 13728
rect 5356 13821 5365 13855
rect 5365 13821 5399 13855
rect 5399 13821 5408 13855
rect 5356 13812 5408 13821
rect 5724 13855 5776 13864
rect 5724 13821 5733 13855
rect 5733 13821 5767 13855
rect 5767 13821 5776 13855
rect 5724 13812 5776 13821
rect 9220 13812 9272 13864
rect 10692 13812 10744 13864
rect 13728 13880 13780 13932
rect 14740 13923 14792 13932
rect 14740 13889 14749 13923
rect 14749 13889 14783 13923
rect 14783 13889 14792 13923
rect 14740 13880 14792 13889
rect 7932 13744 7984 13796
rect 5264 13719 5316 13728
rect 5264 13685 5273 13719
rect 5273 13685 5307 13719
rect 5307 13685 5316 13719
rect 5264 13676 5316 13685
rect 6184 13719 6236 13728
rect 6184 13685 6193 13719
rect 6193 13685 6227 13719
rect 6227 13685 6236 13719
rect 6184 13676 6236 13685
rect 6552 13719 6604 13728
rect 6552 13685 6561 13719
rect 6561 13685 6595 13719
rect 6595 13685 6604 13719
rect 6552 13676 6604 13685
rect 9036 13676 9088 13728
rect 9312 13676 9364 13728
rect 9680 13744 9732 13796
rect 14188 13676 14240 13728
rect 14464 13719 14516 13728
rect 14464 13685 14473 13719
rect 14473 13685 14507 13719
rect 14507 13685 14516 13719
rect 15936 13744 15988 13796
rect 14464 13676 14516 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1676 13472 1728 13524
rect 5080 13472 5132 13524
rect 7472 13515 7524 13524
rect 7472 13481 7481 13515
rect 7481 13481 7515 13515
rect 7515 13481 7524 13515
rect 7472 13472 7524 13481
rect 7932 13515 7984 13524
rect 7932 13481 7941 13515
rect 7941 13481 7975 13515
rect 7975 13481 7984 13515
rect 7932 13472 7984 13481
rect 8208 13472 8260 13524
rect 8760 13472 8812 13524
rect 11704 13472 11756 13524
rect 12164 13515 12216 13524
rect 12164 13481 12173 13515
rect 12173 13481 12207 13515
rect 12207 13481 12216 13515
rect 12164 13472 12216 13481
rect 14740 13515 14792 13524
rect 14740 13481 14749 13515
rect 14749 13481 14783 13515
rect 14783 13481 14792 13515
rect 14740 13472 14792 13481
rect 2596 13447 2648 13456
rect 2596 13413 2605 13447
rect 2605 13413 2639 13447
rect 2639 13413 2648 13447
rect 2596 13404 2648 13413
rect 6184 13404 6236 13456
rect 14464 13404 14516 13456
rect 15476 13447 15528 13456
rect 15476 13413 15485 13447
rect 15485 13413 15519 13447
rect 15519 13413 15528 13447
rect 15476 13404 15528 13413
rect 9680 13379 9732 13388
rect 9680 13345 9689 13379
rect 9689 13345 9723 13379
rect 9723 13345 9732 13379
rect 9680 13336 9732 13345
rect 10140 13379 10192 13388
rect 10140 13345 10149 13379
rect 10149 13345 10183 13379
rect 10183 13345 10192 13379
rect 10140 13336 10192 13345
rect 13728 13379 13780 13388
rect 13728 13345 13737 13379
rect 13737 13345 13771 13379
rect 13771 13345 13780 13379
rect 13728 13336 13780 13345
rect 2320 13268 2372 13320
rect 2504 13311 2556 13320
rect 2504 13277 2513 13311
rect 2513 13277 2547 13311
rect 2547 13277 2556 13311
rect 2504 13268 2556 13277
rect 2872 13311 2924 13320
rect 2872 13277 2881 13311
rect 2881 13277 2915 13311
rect 2915 13277 2924 13311
rect 2872 13268 2924 13277
rect 4068 13311 4120 13320
rect 4068 13277 4077 13311
rect 4077 13277 4111 13311
rect 4111 13277 4120 13311
rect 4068 13268 4120 13277
rect 5540 13311 5592 13320
rect 5540 13277 5549 13311
rect 5549 13277 5583 13311
rect 5583 13277 5592 13311
rect 5540 13268 5592 13277
rect 8576 13268 8628 13320
rect 9036 13268 9088 13320
rect 11244 13311 11296 13320
rect 11244 13277 11253 13311
rect 11253 13277 11287 13311
rect 11287 13277 11296 13311
rect 11244 13268 11296 13277
rect 15752 13268 15804 13320
rect 22008 13268 22060 13320
rect 5724 13200 5776 13252
rect 15936 13243 15988 13252
rect 15936 13209 15945 13243
rect 15945 13209 15979 13243
rect 15979 13209 15988 13243
rect 15936 13200 15988 13209
rect 3148 13132 3200 13184
rect 7288 13132 7340 13184
rect 7748 13132 7800 13184
rect 9220 13132 9272 13184
rect 10508 13132 10560 13184
rect 10692 13175 10744 13184
rect 10692 13141 10701 13175
rect 10701 13141 10735 13175
rect 10735 13141 10744 13175
rect 10692 13132 10744 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 5356 12928 5408 12980
rect 2688 12860 2740 12912
rect 6184 12928 6236 12980
rect 8576 12928 8628 12980
rect 11612 12928 11664 12980
rect 13728 12928 13780 12980
rect 15476 12928 15528 12980
rect 15752 12971 15804 12980
rect 15752 12937 15761 12971
rect 15761 12937 15795 12971
rect 15795 12937 15804 12971
rect 15752 12928 15804 12937
rect 15844 12928 15896 12980
rect 2596 12792 2648 12844
rect 4988 12792 5040 12844
rect 3332 12767 3384 12776
rect 3332 12733 3341 12767
rect 3341 12733 3375 12767
rect 3375 12733 3384 12767
rect 3332 12724 3384 12733
rect 9496 12860 9548 12912
rect 11704 12860 11756 12912
rect 5540 12792 5592 12844
rect 4436 12656 4488 12708
rect 6368 12724 6420 12776
rect 7656 12792 7708 12844
rect 9680 12792 9732 12844
rect 10508 12835 10560 12844
rect 7288 12767 7340 12776
rect 7288 12733 7297 12767
rect 7297 12733 7331 12767
rect 7331 12733 7340 12767
rect 7288 12724 7340 12733
rect 8760 12767 8812 12776
rect 8760 12733 8769 12767
rect 8769 12733 8803 12767
rect 8803 12733 8812 12767
rect 8760 12724 8812 12733
rect 9404 12724 9456 12776
rect 10508 12801 10517 12835
rect 10517 12801 10551 12835
rect 10551 12801 10560 12835
rect 10508 12792 10560 12801
rect 4160 12588 4212 12640
rect 8024 12656 8076 12708
rect 10140 12724 10192 12776
rect 14096 12767 14148 12776
rect 11060 12656 11112 12708
rect 6184 12631 6236 12640
rect 6184 12597 6193 12631
rect 6193 12597 6227 12631
rect 6227 12597 6236 12631
rect 6184 12588 6236 12597
rect 6920 12631 6972 12640
rect 6920 12597 6929 12631
rect 6929 12597 6963 12631
rect 6963 12597 6972 12631
rect 6920 12588 6972 12597
rect 14096 12733 14105 12767
rect 14105 12733 14139 12767
rect 14139 12733 14148 12767
rect 14096 12724 14148 12733
rect 16028 12724 16080 12776
rect 14372 12656 14424 12708
rect 13360 12588 13412 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 2320 12427 2372 12436
rect 2320 12393 2329 12427
rect 2329 12393 2363 12427
rect 2363 12393 2372 12427
rect 2320 12384 2372 12393
rect 4436 12427 4488 12436
rect 4436 12393 4445 12427
rect 4445 12393 4479 12427
rect 4479 12393 4488 12427
rect 4436 12384 4488 12393
rect 4988 12427 5040 12436
rect 4988 12393 4997 12427
rect 4997 12393 5031 12427
rect 5031 12393 5040 12427
rect 4988 12384 5040 12393
rect 5540 12427 5592 12436
rect 5540 12393 5549 12427
rect 5549 12393 5583 12427
rect 5583 12393 5592 12427
rect 5540 12384 5592 12393
rect 8116 12384 8168 12436
rect 9128 12384 9180 12436
rect 11060 12427 11112 12436
rect 11060 12393 11069 12427
rect 11069 12393 11103 12427
rect 11103 12393 11112 12427
rect 11060 12384 11112 12393
rect 24768 12427 24820 12436
rect 24768 12393 24777 12427
rect 24777 12393 24811 12427
rect 24811 12393 24820 12427
rect 24768 12384 24820 12393
rect 2596 12359 2648 12368
rect 2596 12325 2605 12359
rect 2605 12325 2639 12359
rect 2639 12325 2648 12359
rect 2596 12316 2648 12325
rect 3332 12316 3384 12368
rect 3148 12291 3200 12300
rect 3148 12257 3157 12291
rect 3157 12257 3191 12291
rect 3191 12257 3200 12291
rect 3148 12248 3200 12257
rect 3700 12248 3752 12300
rect 6184 12316 6236 12368
rect 6552 12359 6604 12368
rect 6552 12325 6561 12359
rect 6561 12325 6595 12359
rect 6595 12325 6604 12359
rect 6552 12316 6604 12325
rect 11244 12316 11296 12368
rect 6000 12291 6052 12300
rect 2872 12180 2924 12232
rect 3884 12180 3936 12232
rect 5264 12180 5316 12232
rect 6000 12257 6009 12291
rect 6009 12257 6043 12291
rect 6043 12257 6052 12291
rect 6000 12248 6052 12257
rect 6368 12291 6420 12300
rect 6368 12257 6377 12291
rect 6377 12257 6411 12291
rect 6411 12257 6420 12291
rect 6368 12248 6420 12257
rect 8116 12291 8168 12300
rect 8116 12257 8125 12291
rect 8125 12257 8159 12291
rect 8159 12257 8168 12291
rect 8116 12248 8168 12257
rect 8300 12291 8352 12300
rect 8300 12257 8309 12291
rect 8309 12257 8343 12291
rect 8343 12257 8352 12291
rect 8300 12248 8352 12257
rect 9496 12248 9548 12300
rect 10140 12248 10192 12300
rect 11612 12291 11664 12300
rect 11612 12257 11621 12291
rect 11621 12257 11655 12291
rect 11655 12257 11664 12291
rect 11612 12248 11664 12257
rect 14280 12248 14332 12300
rect 15384 12291 15436 12300
rect 15384 12257 15393 12291
rect 15393 12257 15427 12291
rect 15427 12257 15436 12291
rect 15384 12248 15436 12257
rect 24032 12248 24084 12300
rect 6920 12180 6972 12232
rect 8392 12223 8444 12232
rect 8392 12189 8401 12223
rect 8401 12189 8435 12223
rect 8435 12189 8444 12223
rect 8392 12180 8444 12189
rect 8852 12180 8904 12232
rect 13084 12223 13136 12232
rect 13084 12189 13093 12223
rect 13093 12189 13127 12223
rect 13127 12189 13136 12223
rect 13084 12180 13136 12189
rect 4896 12112 4948 12164
rect 7104 12112 7156 12164
rect 9036 12112 9088 12164
rect 1676 12087 1728 12096
rect 1676 12053 1685 12087
rect 1685 12053 1719 12087
rect 1719 12053 1728 12087
rect 1676 12044 1728 12053
rect 4620 12044 4672 12096
rect 7288 12044 7340 12096
rect 7932 12044 7984 12096
rect 15292 12044 15344 12096
rect 15568 12087 15620 12096
rect 15568 12053 15577 12087
rect 15577 12053 15611 12087
rect 15611 12053 15620 12087
rect 15568 12044 15620 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2964 11840 3016 11892
rect 8116 11840 8168 11892
rect 9220 11840 9272 11892
rect 11612 11883 11664 11892
rect 11612 11849 11621 11883
rect 11621 11849 11655 11883
rect 11655 11849 11664 11883
rect 11612 11840 11664 11849
rect 14280 11840 14332 11892
rect 15384 11883 15436 11892
rect 15384 11849 15393 11883
rect 15393 11849 15427 11883
rect 15427 11849 15436 11883
rect 15384 11840 15436 11849
rect 1676 11772 1728 11824
rect 4160 11772 4212 11824
rect 10968 11772 11020 11824
rect 4068 11704 4120 11756
rect 4896 11747 4948 11756
rect 4896 11713 4905 11747
rect 4905 11713 4939 11747
rect 4939 11713 4948 11747
rect 4896 11704 4948 11713
rect 5540 11704 5592 11756
rect 6000 11704 6052 11756
rect 7472 11704 7524 11756
rect 7748 11747 7800 11756
rect 7748 11713 7757 11747
rect 7757 11713 7791 11747
rect 7791 11713 7800 11747
rect 7748 11704 7800 11713
rect 9128 11747 9180 11756
rect 9128 11713 9137 11747
rect 9137 11713 9171 11747
rect 9171 11713 9180 11747
rect 9128 11704 9180 11713
rect 10784 11704 10836 11756
rect 17224 11772 17276 11824
rect 16028 11747 16080 11756
rect 16028 11713 16037 11747
rect 16037 11713 16071 11747
rect 16071 11713 16080 11747
rect 16028 11704 16080 11713
rect 1952 11679 2004 11688
rect 1952 11645 1961 11679
rect 1961 11645 1995 11679
rect 1995 11645 2004 11679
rect 1952 11636 2004 11645
rect 3700 11679 3752 11688
rect 3700 11645 3709 11679
rect 3709 11645 3743 11679
rect 3743 11645 3752 11679
rect 3700 11636 3752 11645
rect 11336 11636 11388 11688
rect 2136 11611 2188 11620
rect 2136 11577 2145 11611
rect 2145 11577 2179 11611
rect 2179 11577 2188 11611
rect 2136 11568 2188 11577
rect 4620 11611 4672 11620
rect 2964 11500 3016 11552
rect 4620 11577 4629 11611
rect 4629 11577 4663 11611
rect 4663 11577 4672 11611
rect 4620 11568 4672 11577
rect 4988 11568 5040 11620
rect 7380 11611 7432 11620
rect 7380 11577 7389 11611
rect 7389 11577 7423 11611
rect 7423 11577 7432 11611
rect 7380 11568 7432 11577
rect 4436 11500 4488 11552
rect 6368 11500 6420 11552
rect 8024 11568 8076 11620
rect 9220 11611 9272 11620
rect 9220 11577 9229 11611
rect 9229 11577 9263 11611
rect 9263 11577 9272 11611
rect 9220 11568 9272 11577
rect 9772 11611 9824 11620
rect 9772 11577 9781 11611
rect 9781 11577 9815 11611
rect 9815 11577 9824 11611
rect 9772 11568 9824 11577
rect 8300 11543 8352 11552
rect 8300 11509 8309 11543
rect 8309 11509 8343 11543
rect 8343 11509 8352 11543
rect 8300 11500 8352 11509
rect 10140 11543 10192 11552
rect 10140 11509 10149 11543
rect 10149 11509 10183 11543
rect 10183 11509 10192 11543
rect 10140 11500 10192 11509
rect 10784 11611 10836 11620
rect 10784 11577 10793 11611
rect 10793 11577 10827 11611
rect 10827 11577 10836 11611
rect 10784 11568 10836 11577
rect 11060 11500 11112 11552
rect 13176 11500 13228 11552
rect 14280 11500 14332 11552
rect 14464 11543 14516 11552
rect 14464 11509 14473 11543
rect 14473 11509 14507 11543
rect 14507 11509 14516 11543
rect 14464 11500 14516 11509
rect 15384 11500 15436 11552
rect 18604 11500 18656 11552
rect 24032 11568 24084 11620
rect 24768 11500 24820 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 2596 11296 2648 11348
rect 3884 11339 3936 11348
rect 3884 11305 3893 11339
rect 3893 11305 3927 11339
rect 3927 11305 3936 11339
rect 3884 11296 3936 11305
rect 4988 11296 5040 11348
rect 7380 11339 7432 11348
rect 7380 11305 7389 11339
rect 7389 11305 7423 11339
rect 7423 11305 7432 11339
rect 7380 11296 7432 11305
rect 9220 11296 9272 11348
rect 9496 11296 9548 11348
rect 6000 11228 6052 11280
rect 7840 11228 7892 11280
rect 8852 11228 8904 11280
rect 11336 11296 11388 11348
rect 22744 11296 22796 11348
rect 10968 11271 11020 11280
rect 10968 11237 10977 11271
rect 10977 11237 11011 11271
rect 11011 11237 11020 11271
rect 10968 11228 11020 11237
rect 14464 11228 14516 11280
rect 15568 11228 15620 11280
rect 16028 11271 16080 11280
rect 16028 11237 16037 11271
rect 16037 11237 16071 11271
rect 16071 11237 16080 11271
rect 16028 11228 16080 11237
rect 16948 11271 17000 11280
rect 16948 11237 16957 11271
rect 16957 11237 16991 11271
rect 16991 11237 17000 11271
rect 16948 11228 17000 11237
rect 17408 11228 17460 11280
rect 1768 11160 1820 11212
rect 2688 11203 2740 11212
rect 2688 11169 2697 11203
rect 2697 11169 2731 11203
rect 2731 11169 2740 11203
rect 2688 11160 2740 11169
rect 2872 11203 2924 11212
rect 2872 11169 2881 11203
rect 2881 11169 2915 11203
rect 2915 11169 2924 11203
rect 2872 11160 2924 11169
rect 4528 11203 4580 11212
rect 4528 11169 4537 11203
rect 4537 11169 4571 11203
rect 4571 11169 4580 11203
rect 4528 11160 4580 11169
rect 11888 11203 11940 11212
rect 11888 11169 11897 11203
rect 11897 11169 11931 11203
rect 11931 11169 11940 11203
rect 11888 11160 11940 11169
rect 13636 11203 13688 11212
rect 13636 11169 13645 11203
rect 13645 11169 13679 11203
rect 13679 11169 13688 11203
rect 13636 11160 13688 11169
rect 1952 11135 2004 11144
rect 1952 11101 1961 11135
rect 1961 11101 1995 11135
rect 1995 11101 2004 11135
rect 1952 11092 2004 11101
rect 3608 11092 3660 11144
rect 6092 11092 6144 11144
rect 6276 11135 6328 11144
rect 6276 11101 6285 11135
rect 6285 11101 6319 11135
rect 6319 11101 6328 11135
rect 6276 11092 6328 11101
rect 3240 11024 3292 11076
rect 2412 10956 2464 11008
rect 5172 10956 5224 11008
rect 9772 11092 9824 11144
rect 10324 11135 10376 11144
rect 10324 11101 10333 11135
rect 10333 11101 10367 11135
rect 10367 11101 10376 11135
rect 10324 11092 10376 11101
rect 12624 11092 12676 11144
rect 12808 11092 12860 11144
rect 17224 11135 17276 11144
rect 17224 11101 17233 11135
rect 17233 11101 17267 11135
rect 17267 11101 17276 11135
rect 17224 11092 17276 11101
rect 16488 10999 16540 11008
rect 16488 10965 16497 10999
rect 16497 10965 16531 10999
rect 16531 10965 16540 10999
rect 16488 10956 16540 10965
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 2688 10795 2740 10804
rect 2688 10761 2697 10795
rect 2697 10761 2731 10795
rect 2731 10761 2740 10795
rect 2688 10752 2740 10761
rect 3700 10752 3752 10804
rect 4528 10795 4580 10804
rect 4528 10761 4537 10795
rect 4537 10761 4571 10795
rect 4571 10761 4580 10795
rect 4528 10752 4580 10761
rect 6000 10795 6052 10804
rect 6000 10761 6009 10795
rect 6009 10761 6043 10795
rect 6043 10761 6052 10795
rect 6000 10752 6052 10761
rect 7840 10795 7892 10804
rect 7840 10761 7849 10795
rect 7849 10761 7883 10795
rect 7883 10761 7892 10795
rect 7840 10752 7892 10761
rect 9220 10795 9272 10804
rect 9220 10761 9229 10795
rect 9229 10761 9263 10795
rect 9263 10761 9272 10795
rect 9220 10752 9272 10761
rect 10324 10752 10376 10804
rect 11888 10795 11940 10804
rect 11888 10761 11897 10795
rect 11897 10761 11931 10795
rect 11931 10761 11940 10795
rect 11888 10752 11940 10761
rect 13636 10795 13688 10804
rect 13636 10761 13645 10795
rect 13645 10761 13679 10795
rect 13679 10761 13688 10795
rect 13636 10752 13688 10761
rect 14372 10795 14424 10804
rect 14372 10761 14381 10795
rect 14381 10761 14415 10795
rect 14415 10761 14424 10795
rect 14372 10752 14424 10761
rect 15384 10795 15436 10804
rect 15384 10761 15393 10795
rect 15393 10761 15427 10795
rect 15427 10761 15436 10795
rect 15384 10752 15436 10761
rect 15568 10752 15620 10804
rect 25228 10752 25280 10804
rect 5540 10684 5592 10736
rect 11336 10684 11388 10736
rect 1676 10659 1728 10668
rect 1676 10625 1685 10659
rect 1685 10625 1719 10659
rect 1719 10625 1728 10659
rect 1676 10616 1728 10625
rect 6092 10616 6144 10668
rect 7380 10616 7432 10668
rect 8392 10616 8444 10668
rect 12716 10659 12768 10668
rect 12716 10625 12725 10659
rect 12725 10625 12759 10659
rect 12759 10625 12768 10659
rect 12716 10616 12768 10625
rect 13084 10616 13136 10668
rect 14740 10616 14792 10668
rect 16488 10659 16540 10668
rect 16488 10625 16497 10659
rect 16497 10625 16531 10659
rect 16531 10625 16540 10659
rect 16488 10616 16540 10625
rect 17224 10616 17276 10668
rect 10048 10591 10100 10600
rect 10048 10557 10057 10591
rect 10057 10557 10091 10591
rect 10091 10557 10100 10591
rect 10048 10548 10100 10557
rect 2412 10480 2464 10532
rect 4712 10523 4764 10532
rect 4712 10489 4721 10523
rect 4721 10489 4755 10523
rect 4755 10489 4764 10523
rect 4712 10480 4764 10489
rect 2228 10412 2280 10464
rect 2872 10412 2924 10464
rect 4528 10412 4580 10464
rect 6276 10480 6328 10532
rect 8208 10523 8260 10532
rect 8208 10489 8217 10523
rect 8217 10489 8251 10523
rect 8251 10489 8260 10523
rect 8208 10480 8260 10489
rect 9772 10412 9824 10464
rect 12808 10523 12860 10532
rect 12808 10489 12817 10523
rect 12817 10489 12851 10523
rect 12851 10489 12860 10523
rect 13360 10523 13412 10532
rect 12808 10480 12860 10489
rect 13360 10489 13369 10523
rect 13369 10489 13403 10523
rect 13403 10489 13412 10523
rect 13360 10480 13412 10489
rect 14372 10480 14424 10532
rect 15660 10480 15712 10532
rect 17408 10455 17460 10464
rect 17408 10421 17417 10455
rect 17417 10421 17451 10455
rect 17451 10421 17460 10455
rect 17408 10412 17460 10421
rect 24124 10548 24176 10600
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 4712 10208 4764 10260
rect 8392 10251 8444 10260
rect 8392 10217 8401 10251
rect 8401 10217 8435 10251
rect 8435 10217 8444 10251
rect 8392 10208 8444 10217
rect 10048 10208 10100 10260
rect 12716 10251 12768 10260
rect 12716 10217 12725 10251
rect 12725 10217 12759 10251
rect 12759 10217 12768 10251
rect 12716 10208 12768 10217
rect 2780 10140 2832 10192
rect 4436 10183 4488 10192
rect 4436 10149 4439 10183
rect 4439 10149 4473 10183
rect 4473 10149 4488 10183
rect 4436 10140 4488 10149
rect 5540 10140 5592 10192
rect 7196 10183 7248 10192
rect 7196 10149 7205 10183
rect 7205 10149 7239 10183
rect 7239 10149 7248 10183
rect 7196 10140 7248 10149
rect 7748 10183 7800 10192
rect 7748 10149 7757 10183
rect 7757 10149 7791 10183
rect 7791 10149 7800 10183
rect 7748 10140 7800 10149
rect 8024 10140 8076 10192
rect 13636 10208 13688 10260
rect 14464 10208 14516 10260
rect 15660 10251 15712 10260
rect 15660 10217 15669 10251
rect 15669 10217 15703 10251
rect 15703 10217 15712 10251
rect 15660 10208 15712 10217
rect 16488 10208 16540 10260
rect 24216 10208 24268 10260
rect 13360 10140 13412 10192
rect 16948 10183 17000 10192
rect 16948 10149 16957 10183
rect 16957 10149 16991 10183
rect 16991 10149 17000 10183
rect 16948 10140 17000 10149
rect 18420 10183 18472 10192
rect 18420 10149 18429 10183
rect 18429 10149 18463 10183
rect 18463 10149 18472 10183
rect 18420 10140 18472 10149
rect 18604 10140 18656 10192
rect 4528 10072 4580 10124
rect 8576 10115 8628 10124
rect 8576 10081 8585 10115
rect 8585 10081 8619 10115
rect 8619 10081 8628 10115
rect 8576 10072 8628 10081
rect 2228 10004 2280 10056
rect 3148 10047 3200 10056
rect 2412 9936 2464 9988
rect 3148 10013 3157 10047
rect 3157 10013 3191 10047
rect 3191 10013 3200 10047
rect 3148 10004 3200 10013
rect 3976 10004 4028 10056
rect 9956 10072 10008 10124
rect 11612 10115 11664 10124
rect 11612 10081 11621 10115
rect 11621 10081 11655 10115
rect 11655 10081 11664 10115
rect 11612 10072 11664 10081
rect 17316 10115 17368 10124
rect 17316 10081 17325 10115
rect 17325 10081 17359 10115
rect 17359 10081 17368 10115
rect 17316 10072 17368 10081
rect 23848 10072 23900 10124
rect 3332 9936 3384 9988
rect 4712 9936 4764 9988
rect 1768 9868 1820 9920
rect 2320 9911 2372 9920
rect 2320 9877 2329 9911
rect 2329 9877 2363 9911
rect 2363 9877 2372 9911
rect 2320 9868 2372 9877
rect 2596 9868 2648 9920
rect 10876 10004 10928 10056
rect 15844 10004 15896 10056
rect 19064 10047 19116 10056
rect 19064 10013 19073 10047
rect 19073 10013 19107 10047
rect 19107 10013 19116 10047
rect 19064 10004 19116 10013
rect 13728 9936 13780 9988
rect 17408 9936 17460 9988
rect 7380 9868 7432 9920
rect 7656 9868 7708 9920
rect 14740 9868 14792 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 1676 9664 1728 9716
rect 3148 9664 3200 9716
rect 7196 9664 7248 9716
rect 11612 9707 11664 9716
rect 11612 9673 11621 9707
rect 11621 9673 11655 9707
rect 11655 9673 11664 9707
rect 11612 9664 11664 9673
rect 13636 9707 13688 9716
rect 13636 9673 13645 9707
rect 13645 9673 13679 9707
rect 13679 9673 13688 9707
rect 13636 9664 13688 9673
rect 15660 9664 15712 9716
rect 18420 9664 18472 9716
rect 23848 9707 23900 9716
rect 23848 9673 23857 9707
rect 23857 9673 23891 9707
rect 23891 9673 23900 9707
rect 23848 9664 23900 9673
rect 4620 9639 4672 9648
rect 4620 9605 4629 9639
rect 4629 9605 4663 9639
rect 4663 9605 4672 9639
rect 4620 9596 4672 9605
rect 5632 9596 5684 9648
rect 2228 9528 2280 9580
rect 6736 9528 6788 9580
rect 7196 9528 7248 9580
rect 1860 9503 1912 9512
rect 1860 9469 1869 9503
rect 1869 9469 1903 9503
rect 1903 9469 1912 9503
rect 1860 9460 1912 9469
rect 2780 9503 2832 9512
rect 2780 9469 2789 9503
rect 2789 9469 2823 9503
rect 2823 9469 2832 9503
rect 2780 9460 2832 9469
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 2688 9324 2740 9376
rect 4712 9324 4764 9376
rect 6092 9324 6144 9376
rect 8576 9596 8628 9648
rect 9404 9639 9456 9648
rect 8208 9392 8260 9444
rect 9404 9605 9413 9639
rect 9413 9605 9447 9639
rect 9447 9605 9456 9639
rect 9404 9596 9456 9605
rect 9772 9596 9824 9648
rect 13728 9596 13780 9648
rect 19064 9596 19116 9648
rect 14740 9571 14792 9580
rect 9864 9460 9916 9512
rect 12164 9460 12216 9512
rect 14740 9537 14749 9571
rect 14749 9537 14783 9571
rect 14783 9537 14792 9571
rect 14740 9528 14792 9537
rect 13912 9460 13964 9512
rect 14648 9503 14700 9512
rect 14648 9469 14657 9503
rect 14657 9469 14691 9503
rect 14691 9469 14700 9503
rect 19524 9571 19576 9580
rect 19524 9537 19533 9571
rect 19533 9537 19567 9571
rect 19567 9537 19576 9571
rect 19524 9528 19576 9537
rect 14648 9460 14700 9469
rect 12716 9392 12768 9444
rect 13636 9392 13688 9444
rect 16488 9460 16540 9512
rect 18696 9435 18748 9444
rect 18696 9401 18705 9435
rect 18705 9401 18739 9435
rect 18739 9401 18748 9435
rect 18696 9392 18748 9401
rect 7288 9324 7340 9376
rect 7472 9324 7524 9376
rect 10876 9324 10928 9376
rect 11152 9367 11204 9376
rect 11152 9333 11161 9367
rect 11161 9333 11195 9367
rect 11195 9333 11204 9367
rect 11152 9324 11204 9333
rect 13912 9324 13964 9376
rect 15844 9367 15896 9376
rect 15844 9333 15853 9367
rect 15853 9333 15887 9367
rect 15887 9333 15896 9367
rect 15844 9324 15896 9333
rect 17316 9367 17368 9376
rect 17316 9333 17325 9367
rect 17325 9333 17359 9367
rect 17359 9333 17368 9367
rect 17316 9324 17368 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2688 9120 2740 9172
rect 2780 9120 2832 9172
rect 3240 9120 3292 9172
rect 5264 9120 5316 9172
rect 5632 9163 5684 9172
rect 5632 9129 5641 9163
rect 5641 9129 5675 9163
rect 5675 9129 5684 9163
rect 5632 9120 5684 9129
rect 6092 9120 6144 9172
rect 6828 9095 6880 9104
rect 6828 9061 6837 9095
rect 6837 9061 6871 9095
rect 6871 9061 6880 9095
rect 6828 9052 6880 9061
rect 11888 9120 11940 9172
rect 13728 9120 13780 9172
rect 15844 9120 15896 9172
rect 16488 9163 16540 9172
rect 16488 9129 16497 9163
rect 16497 9129 16531 9163
rect 16531 9129 16540 9163
rect 16488 9120 16540 9129
rect 18696 9120 18748 9172
rect 7196 9095 7248 9104
rect 7196 9061 7205 9095
rect 7205 9061 7239 9095
rect 7239 9061 7248 9095
rect 11060 9095 11112 9104
rect 7196 9052 7248 9061
rect 11060 9061 11069 9095
rect 11069 9061 11103 9095
rect 11103 9061 11112 9095
rect 11060 9052 11112 9061
rect 11152 9052 11204 9104
rect 12256 9052 12308 9104
rect 12624 9095 12676 9104
rect 12624 9061 12633 9095
rect 12633 9061 12667 9095
rect 12667 9061 12676 9095
rect 13176 9095 13228 9104
rect 12624 9052 12676 9061
rect 13176 9061 13185 9095
rect 13185 9061 13219 9095
rect 13219 9061 13228 9095
rect 13176 9052 13228 9061
rect 15476 9052 15528 9104
rect 15660 9052 15712 9104
rect 3608 8984 3660 9036
rect 1400 8780 1452 8832
rect 2044 8823 2096 8832
rect 2044 8789 2053 8823
rect 2053 8789 2087 8823
rect 2087 8789 2096 8823
rect 2044 8780 2096 8789
rect 3516 8823 3568 8832
rect 3516 8789 3525 8823
rect 3525 8789 3559 8823
rect 3559 8789 3568 8823
rect 3516 8780 3568 8789
rect 3792 8823 3844 8832
rect 3792 8789 3801 8823
rect 3801 8789 3835 8823
rect 3835 8789 3844 8823
rect 3792 8780 3844 8789
rect 3976 8916 4028 8968
rect 4252 8984 4304 9036
rect 5080 8984 5132 9036
rect 6000 8984 6052 9036
rect 8576 9027 8628 9036
rect 8576 8993 8585 9027
rect 8585 8993 8619 9027
rect 8619 8993 8628 9027
rect 8576 8984 8628 8993
rect 9864 9027 9916 9036
rect 9864 8993 9873 9027
rect 9873 8993 9907 9027
rect 9907 8993 9916 9027
rect 9864 8984 9916 8993
rect 7380 8959 7432 8968
rect 7380 8925 7389 8959
rect 7389 8925 7423 8959
rect 7423 8925 7432 8959
rect 7380 8916 7432 8925
rect 7748 8916 7800 8968
rect 9128 8916 9180 8968
rect 10968 8959 11020 8968
rect 10968 8925 10977 8959
rect 10977 8925 11011 8959
rect 11011 8925 11020 8959
rect 10968 8916 11020 8925
rect 17132 9027 17184 9036
rect 17132 8993 17141 9027
rect 17141 8993 17175 9027
rect 17175 8993 17184 9027
rect 17132 8984 17184 8993
rect 14648 8916 14700 8968
rect 16212 8916 16264 8968
rect 8300 8848 8352 8900
rect 9956 8848 10008 8900
rect 4344 8780 4396 8832
rect 6092 8780 6144 8832
rect 8392 8823 8444 8832
rect 8392 8789 8401 8823
rect 8401 8789 8435 8823
rect 8435 8789 8444 8823
rect 8392 8780 8444 8789
rect 8760 8823 8812 8832
rect 8760 8789 8769 8823
rect 8769 8789 8803 8823
rect 8803 8789 8812 8823
rect 8760 8780 8812 8789
rect 13636 8848 13688 8900
rect 10692 8823 10744 8832
rect 10692 8789 10701 8823
rect 10701 8789 10735 8823
rect 10735 8789 10744 8823
rect 10692 8780 10744 8789
rect 12164 8780 12216 8832
rect 14188 8823 14240 8832
rect 14188 8789 14197 8823
rect 14197 8789 14231 8823
rect 14231 8789 14240 8823
rect 14188 8780 14240 8789
rect 14556 8780 14608 8832
rect 18604 8984 18656 9036
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 3976 8576 4028 8628
rect 5540 8576 5592 8628
rect 6000 8576 6052 8628
rect 7196 8576 7248 8628
rect 8576 8619 8628 8628
rect 8576 8585 8585 8619
rect 8585 8585 8619 8619
rect 8619 8585 8628 8619
rect 8576 8576 8628 8585
rect 9864 8576 9916 8628
rect 11060 8619 11112 8628
rect 11060 8585 11069 8619
rect 11069 8585 11103 8619
rect 11103 8585 11112 8619
rect 11060 8576 11112 8585
rect 12256 8619 12308 8628
rect 12256 8585 12265 8619
rect 12265 8585 12299 8619
rect 12299 8585 12308 8619
rect 12256 8576 12308 8585
rect 12624 8619 12676 8628
rect 12624 8585 12633 8619
rect 12633 8585 12667 8619
rect 12667 8585 12676 8619
rect 12624 8576 12676 8585
rect 14648 8619 14700 8628
rect 14648 8585 14657 8619
rect 14657 8585 14691 8619
rect 14691 8585 14700 8619
rect 14648 8576 14700 8585
rect 17132 8619 17184 8628
rect 17132 8585 17141 8619
rect 17141 8585 17175 8619
rect 17175 8585 17184 8619
rect 17132 8576 17184 8585
rect 18604 8619 18656 8628
rect 18604 8585 18613 8619
rect 18613 8585 18647 8619
rect 18647 8585 18656 8619
rect 18604 8576 18656 8585
rect 19524 8576 19576 8628
rect 3792 8551 3844 8560
rect 3792 8517 3801 8551
rect 3801 8517 3835 8551
rect 3835 8517 3844 8551
rect 3792 8508 3844 8517
rect 7748 8551 7800 8560
rect 7748 8517 7757 8551
rect 7757 8517 7791 8551
rect 7791 8517 7800 8551
rect 7748 8508 7800 8517
rect 7932 8551 7984 8560
rect 7932 8517 7941 8551
rect 7941 8517 7975 8551
rect 7975 8517 7984 8551
rect 7932 8508 7984 8517
rect 1952 8440 2004 8492
rect 2688 8483 2740 8492
rect 2688 8449 2697 8483
rect 2697 8449 2731 8483
rect 2731 8449 2740 8483
rect 2688 8440 2740 8449
rect 4620 8440 4672 8492
rect 5264 8483 5316 8492
rect 5264 8449 5273 8483
rect 5273 8449 5307 8483
rect 5307 8449 5316 8483
rect 5264 8440 5316 8449
rect 7380 8440 7432 8492
rect 7472 8440 7524 8492
rect 8852 8440 8904 8492
rect 14096 8483 14148 8492
rect 1400 8304 1452 8356
rect 1768 8279 1820 8288
rect 1768 8245 1777 8279
rect 1777 8245 1811 8279
rect 1811 8245 1820 8279
rect 1768 8236 1820 8245
rect 3516 8415 3568 8424
rect 2964 8304 3016 8356
rect 3516 8381 3525 8415
rect 3525 8381 3559 8415
rect 3559 8381 3568 8415
rect 3516 8372 3568 8381
rect 3700 8415 3752 8424
rect 3700 8381 3709 8415
rect 3709 8381 3743 8415
rect 3743 8381 3752 8415
rect 3700 8372 3752 8381
rect 9680 8372 9732 8424
rect 10692 8372 10744 8424
rect 13636 8415 13688 8424
rect 13636 8381 13645 8415
rect 13645 8381 13679 8415
rect 13679 8381 13688 8415
rect 13636 8372 13688 8381
rect 14096 8449 14105 8483
rect 14105 8449 14139 8483
rect 14139 8449 14148 8483
rect 14096 8440 14148 8449
rect 15936 8508 15988 8560
rect 16120 8440 16172 8492
rect 15384 8372 15436 8424
rect 2504 8236 2556 8288
rect 4620 8279 4672 8288
rect 4620 8245 4629 8279
rect 4629 8245 4663 8279
rect 4663 8245 4672 8279
rect 4620 8236 4672 8245
rect 5540 8304 5592 8356
rect 6092 8304 6144 8356
rect 7472 8347 7524 8356
rect 7472 8313 7481 8347
rect 7481 8313 7515 8347
rect 7515 8313 7524 8347
rect 7472 8304 7524 8313
rect 9772 8304 9824 8356
rect 10968 8236 11020 8288
rect 12716 8236 12768 8288
rect 15476 8236 15528 8288
rect 15844 8347 15896 8356
rect 15844 8313 15853 8347
rect 15853 8313 15887 8347
rect 15887 8313 15896 8347
rect 16396 8347 16448 8356
rect 15844 8304 15896 8313
rect 16396 8313 16405 8347
rect 16405 8313 16439 8347
rect 16439 8313 16448 8347
rect 16396 8304 16448 8313
rect 21180 8236 21232 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 3700 8032 3752 8084
rect 4344 8075 4396 8084
rect 4344 8041 4353 8075
rect 4353 8041 4387 8075
rect 4387 8041 4396 8075
rect 4344 8032 4396 8041
rect 5540 8075 5592 8084
rect 5540 8041 5549 8075
rect 5549 8041 5583 8075
rect 5583 8041 5592 8075
rect 5540 8032 5592 8041
rect 1952 7964 2004 8016
rect 4436 7964 4488 8016
rect 8300 8007 8352 8016
rect 4160 7939 4212 7948
rect 4160 7905 4169 7939
rect 4169 7905 4203 7939
rect 4203 7905 4212 7939
rect 4620 7939 4672 7948
rect 4160 7896 4212 7905
rect 4620 7905 4629 7939
rect 4629 7905 4663 7939
rect 4663 7905 4672 7939
rect 4620 7896 4672 7905
rect 8300 7973 8309 8007
rect 8309 7973 8343 8007
rect 8343 7973 8352 8007
rect 8300 7964 8352 7973
rect 6184 7939 6236 7948
rect 6184 7905 6193 7939
rect 6193 7905 6227 7939
rect 6227 7905 6236 7939
rect 6184 7896 6236 7905
rect 7748 7896 7800 7948
rect 10876 8032 10928 8084
rect 12164 8075 12216 8084
rect 12164 8041 12173 8075
rect 12173 8041 12207 8075
rect 12207 8041 12216 8075
rect 12164 8032 12216 8041
rect 10692 7964 10744 8016
rect 14648 7964 14700 8016
rect 15476 7964 15528 8016
rect 10048 7896 10100 7948
rect 12348 7939 12400 7948
rect 2044 7828 2096 7880
rect 2780 7828 2832 7880
rect 3700 7871 3752 7880
rect 3700 7837 3709 7871
rect 3709 7837 3743 7871
rect 3743 7837 3752 7871
rect 3700 7828 3752 7837
rect 7012 7828 7064 7880
rect 8116 7760 8168 7812
rect 8760 7828 8812 7880
rect 8392 7760 8444 7812
rect 12348 7905 12357 7939
rect 12357 7905 12391 7939
rect 12391 7905 12400 7939
rect 12348 7896 12400 7905
rect 13636 7939 13688 7948
rect 13636 7905 13645 7939
rect 13645 7905 13679 7939
rect 13679 7905 13688 7939
rect 13636 7896 13688 7905
rect 15292 7939 15344 7948
rect 15292 7905 15301 7939
rect 15301 7905 15335 7939
rect 15335 7905 15344 7939
rect 15292 7896 15344 7905
rect 15384 7896 15436 7948
rect 17040 7896 17092 7948
rect 17500 7939 17552 7948
rect 17500 7905 17509 7939
rect 17509 7905 17543 7939
rect 17543 7905 17552 7939
rect 17500 7896 17552 7905
rect 11980 7760 12032 7812
rect 15844 7760 15896 7812
rect 17132 7760 17184 7812
rect 2228 7692 2280 7744
rect 2964 7735 3016 7744
rect 2964 7701 2973 7735
rect 2973 7701 3007 7735
rect 3007 7701 3016 7735
rect 2964 7692 3016 7701
rect 6000 7692 6052 7744
rect 6276 7735 6328 7744
rect 6276 7701 6285 7735
rect 6285 7701 6319 7735
rect 6319 7701 6328 7735
rect 6276 7692 6328 7701
rect 7472 7735 7524 7744
rect 7472 7701 7481 7735
rect 7481 7701 7515 7735
rect 7515 7701 7524 7735
rect 7472 7692 7524 7701
rect 7840 7735 7892 7744
rect 7840 7701 7849 7735
rect 7849 7701 7883 7735
rect 7883 7701 7892 7735
rect 7840 7692 7892 7701
rect 8576 7735 8628 7744
rect 8576 7701 8585 7735
rect 8585 7701 8619 7735
rect 8619 7701 8628 7735
rect 8576 7692 8628 7701
rect 8944 7735 8996 7744
rect 8944 7701 8953 7735
rect 8953 7701 8987 7735
rect 8987 7701 8996 7735
rect 8944 7692 8996 7701
rect 9036 7692 9088 7744
rect 9864 7692 9916 7744
rect 13912 7692 13964 7744
rect 17040 7692 17092 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 4436 7531 4488 7540
rect 4436 7497 4445 7531
rect 4445 7497 4479 7531
rect 4479 7497 4488 7531
rect 4436 7488 4488 7497
rect 6736 7488 6788 7540
rect 7840 7488 7892 7540
rect 8668 7531 8720 7540
rect 8668 7497 8677 7531
rect 8677 7497 8711 7531
rect 8711 7497 8720 7531
rect 8668 7488 8720 7497
rect 9128 7488 9180 7540
rect 9772 7531 9824 7540
rect 2964 7420 3016 7472
rect 8944 7420 8996 7472
rect 9312 7420 9364 7472
rect 9772 7497 9796 7531
rect 9796 7497 9824 7531
rect 9772 7488 9824 7497
rect 9036 7352 9088 7404
rect 9404 7352 9456 7404
rect 10140 7488 10192 7540
rect 11980 7531 12032 7540
rect 11980 7497 11989 7531
rect 11989 7497 12023 7531
rect 12023 7497 12032 7531
rect 11980 7488 12032 7497
rect 13636 7488 13688 7540
rect 13820 7488 13872 7540
rect 15292 7488 15344 7540
rect 15476 7531 15528 7540
rect 15476 7497 15485 7531
rect 15485 7497 15519 7531
rect 15519 7497 15528 7531
rect 15476 7488 15528 7497
rect 17040 7531 17092 7540
rect 17040 7497 17049 7531
rect 17049 7497 17083 7531
rect 17083 7497 17092 7531
rect 17040 7488 17092 7497
rect 17500 7531 17552 7540
rect 17500 7497 17509 7531
rect 17509 7497 17543 7531
rect 17543 7497 17552 7531
rect 17500 7488 17552 7497
rect 25136 7531 25188 7540
rect 25136 7497 25145 7531
rect 25145 7497 25179 7531
rect 25179 7497 25188 7531
rect 25136 7488 25188 7497
rect 13452 7420 13504 7472
rect 10692 7352 10744 7404
rect 14004 7395 14056 7404
rect 14004 7361 14013 7395
rect 14013 7361 14047 7395
rect 14047 7361 14056 7395
rect 14004 7352 14056 7361
rect 16396 7395 16448 7404
rect 16396 7361 16405 7395
rect 16405 7361 16439 7395
rect 16439 7361 16448 7395
rect 16396 7352 16448 7361
rect 1860 7284 1912 7336
rect 2964 7327 3016 7336
rect 2964 7293 2973 7327
rect 2973 7293 3007 7327
rect 3007 7293 3016 7327
rect 2964 7284 3016 7293
rect 3516 7327 3568 7336
rect 3516 7293 3525 7327
rect 3525 7293 3559 7327
rect 3559 7293 3568 7327
rect 3516 7284 3568 7293
rect 3700 7327 3752 7336
rect 3700 7293 3709 7327
rect 3709 7293 3743 7327
rect 3743 7293 3752 7327
rect 3700 7284 3752 7293
rect 3884 7284 3936 7336
rect 6736 7284 6788 7336
rect 4160 7259 4212 7268
rect 4160 7225 4169 7259
rect 4169 7225 4203 7259
rect 4203 7225 4212 7259
rect 4160 7216 4212 7225
rect 5356 7216 5408 7268
rect 6276 7216 6328 7268
rect 8576 7284 8628 7336
rect 8760 7284 8812 7336
rect 12348 7284 12400 7336
rect 15108 7327 15160 7336
rect 15108 7293 15126 7327
rect 15126 7293 15160 7327
rect 15108 7284 15160 7293
rect 25136 7284 25188 7336
rect 7472 7216 7524 7268
rect 8484 7216 8536 7268
rect 9220 7216 9272 7268
rect 9588 7259 9640 7268
rect 9588 7225 9597 7259
rect 9597 7225 9631 7259
rect 9631 7225 9640 7259
rect 9588 7216 9640 7225
rect 13360 7259 13412 7268
rect 13360 7225 13369 7259
rect 13369 7225 13403 7259
rect 13403 7225 13412 7259
rect 13360 7216 13412 7225
rect 13452 7259 13504 7268
rect 13452 7225 13461 7259
rect 13461 7225 13495 7259
rect 13495 7225 13504 7259
rect 16120 7259 16172 7268
rect 13452 7216 13504 7225
rect 16120 7225 16129 7259
rect 16129 7225 16163 7259
rect 16163 7225 16172 7259
rect 16120 7216 16172 7225
rect 16212 7259 16264 7268
rect 16212 7225 16221 7259
rect 16221 7225 16255 7259
rect 16255 7225 16264 7259
rect 18052 7259 18104 7268
rect 16212 7216 16264 7225
rect 18052 7225 18061 7259
rect 18061 7225 18095 7259
rect 18095 7225 18104 7259
rect 18052 7216 18104 7225
rect 2044 7148 2096 7200
rect 2780 7191 2832 7200
rect 2780 7157 2789 7191
rect 2789 7157 2823 7191
rect 2823 7157 2832 7191
rect 2780 7148 2832 7157
rect 5448 7191 5500 7200
rect 5448 7157 5457 7191
rect 5457 7157 5491 7191
rect 5491 7157 5500 7191
rect 5448 7148 5500 7157
rect 6184 7191 6236 7200
rect 6184 7157 6193 7191
rect 6193 7157 6227 7191
rect 6227 7157 6236 7191
rect 6184 7148 6236 7157
rect 7012 7191 7064 7200
rect 7012 7157 7021 7191
rect 7021 7157 7055 7191
rect 7055 7157 7064 7191
rect 7012 7148 7064 7157
rect 9128 7191 9180 7200
rect 9128 7157 9137 7191
rect 9137 7157 9171 7191
rect 9171 7157 9180 7191
rect 9128 7148 9180 7157
rect 9404 7191 9456 7200
rect 9404 7157 9413 7191
rect 9413 7157 9447 7191
rect 9447 7157 9456 7191
rect 9404 7148 9456 7157
rect 11336 7191 11388 7200
rect 11336 7157 11345 7191
rect 11345 7157 11379 7191
rect 11379 7157 11388 7191
rect 11336 7148 11388 7157
rect 15292 7148 15344 7200
rect 25136 7148 25188 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 2964 6944 3016 6996
rect 3700 6944 3752 6996
rect 4252 6944 4304 6996
rect 8852 6944 8904 6996
rect 8944 6944 8996 6996
rect 13452 6987 13504 6996
rect 13452 6953 13461 6987
rect 13461 6953 13495 6987
rect 13495 6953 13504 6987
rect 13452 6944 13504 6953
rect 15108 6987 15160 6996
rect 15108 6953 15117 6987
rect 15117 6953 15151 6987
rect 15151 6953 15160 6987
rect 15108 6944 15160 6953
rect 16120 6944 16172 6996
rect 16488 6944 16540 6996
rect 3516 6919 3568 6928
rect 3516 6885 3525 6919
rect 3525 6885 3559 6919
rect 3559 6885 3568 6919
rect 3516 6876 3568 6885
rect 2228 6808 2280 6860
rect 3148 6808 3200 6860
rect 3884 6808 3936 6860
rect 1860 6740 1912 6792
rect 5080 6876 5132 6928
rect 6460 6919 6512 6928
rect 6460 6885 6469 6919
rect 6469 6885 6503 6919
rect 6503 6885 6512 6919
rect 6460 6876 6512 6885
rect 8760 6919 8812 6928
rect 8760 6885 8769 6919
rect 8769 6885 8803 6919
rect 8803 6885 8812 6919
rect 8760 6876 8812 6885
rect 12716 6876 12768 6928
rect 14556 6876 14608 6928
rect 18052 6876 18104 6928
rect 4620 6851 4672 6860
rect 4620 6817 4629 6851
rect 4629 6817 4663 6851
rect 4663 6817 4672 6851
rect 4620 6808 4672 6817
rect 4988 6808 5040 6860
rect 7748 6808 7800 6860
rect 8116 6808 8168 6860
rect 9496 6808 9548 6860
rect 9680 6851 9732 6860
rect 9680 6817 9689 6851
rect 9689 6817 9723 6851
rect 9723 6817 9732 6851
rect 9680 6808 9732 6817
rect 11244 6851 11296 6860
rect 7012 6740 7064 6792
rect 7564 6740 7616 6792
rect 6000 6715 6052 6724
rect 6000 6681 6009 6715
rect 6009 6681 6043 6715
rect 6043 6681 6052 6715
rect 6736 6715 6788 6724
rect 6000 6672 6052 6681
rect 1676 6647 1728 6656
rect 1676 6613 1685 6647
rect 1685 6613 1719 6647
rect 1719 6613 1728 6647
rect 1676 6604 1728 6613
rect 5448 6604 5500 6656
rect 5540 6647 5592 6656
rect 5540 6613 5549 6647
rect 5549 6613 5583 6647
rect 5583 6613 5592 6647
rect 6736 6681 6745 6715
rect 6745 6681 6779 6715
rect 6779 6681 6788 6715
rect 6736 6672 6788 6681
rect 10048 6740 10100 6792
rect 11244 6817 11253 6851
rect 11253 6817 11287 6851
rect 11287 6817 11296 6851
rect 11244 6808 11296 6817
rect 11336 6808 11388 6860
rect 12256 6783 12308 6792
rect 12256 6749 12265 6783
rect 12265 6749 12299 6783
rect 12299 6749 12308 6783
rect 12256 6740 12308 6749
rect 14648 6740 14700 6792
rect 16212 6808 16264 6860
rect 18420 6851 18472 6860
rect 18420 6817 18429 6851
rect 18429 6817 18463 6851
rect 18463 6817 18472 6851
rect 18420 6808 18472 6817
rect 18880 6851 18932 6860
rect 18880 6817 18889 6851
rect 18889 6817 18923 6851
rect 18923 6817 18932 6851
rect 18880 6808 18932 6817
rect 23204 6808 23256 6860
rect 15384 6783 15436 6792
rect 15384 6749 15393 6783
rect 15393 6749 15427 6783
rect 15427 6749 15436 6783
rect 15384 6740 15436 6749
rect 13452 6672 13504 6724
rect 14004 6672 14056 6724
rect 17500 6740 17552 6792
rect 5540 6604 5592 6613
rect 7012 6604 7064 6656
rect 7748 6604 7800 6656
rect 8300 6647 8352 6656
rect 8300 6613 8309 6647
rect 8309 6613 8343 6647
rect 8343 6613 8352 6647
rect 8300 6604 8352 6613
rect 8576 6604 8628 6656
rect 9312 6604 9364 6656
rect 9496 6604 9548 6656
rect 10784 6604 10836 6656
rect 16764 6647 16816 6656
rect 16764 6613 16773 6647
rect 16773 6613 16807 6647
rect 16807 6613 16816 6647
rect 16764 6604 16816 6613
rect 16856 6604 16908 6656
rect 17224 6604 17276 6656
rect 23940 6647 23992 6656
rect 23940 6613 23949 6647
rect 23949 6613 23983 6647
rect 23983 6613 23992 6647
rect 23940 6604 23992 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 5540 6400 5592 6452
rect 6368 6400 6420 6452
rect 6736 6400 6788 6452
rect 7564 6443 7616 6452
rect 7564 6409 7573 6443
rect 7573 6409 7607 6443
rect 7607 6409 7616 6443
rect 7564 6400 7616 6409
rect 8300 6443 8352 6452
rect 5448 6375 5500 6384
rect 5448 6341 5457 6375
rect 5457 6341 5491 6375
rect 5491 6341 5500 6375
rect 5448 6332 5500 6341
rect 6920 6332 6972 6384
rect 2412 6264 2464 6316
rect 3240 6239 3292 6248
rect 3240 6205 3249 6239
rect 3249 6205 3283 6239
rect 3283 6205 3292 6239
rect 3240 6196 3292 6205
rect 1584 6171 1636 6180
rect 1584 6137 1593 6171
rect 1593 6137 1627 6171
rect 1627 6137 1636 6171
rect 1584 6128 1636 6137
rect 1676 6171 1728 6180
rect 1676 6137 1685 6171
rect 1685 6137 1719 6171
rect 1719 6137 1728 6171
rect 4712 6264 4764 6316
rect 8300 6409 8309 6443
rect 8309 6409 8343 6443
rect 8343 6409 8352 6443
rect 9128 6443 9180 6452
rect 8300 6400 8352 6409
rect 9128 6409 9137 6443
rect 9137 6409 9171 6443
rect 9171 6409 9180 6443
rect 9128 6400 9180 6409
rect 9312 6400 9364 6452
rect 9956 6400 10008 6452
rect 10692 6443 10744 6452
rect 10692 6409 10701 6443
rect 10701 6409 10735 6443
rect 10735 6409 10744 6443
rect 10692 6400 10744 6409
rect 12716 6400 12768 6452
rect 14556 6443 14608 6452
rect 14556 6409 14565 6443
rect 14565 6409 14599 6443
rect 14599 6409 14608 6443
rect 14556 6400 14608 6409
rect 16856 6400 16908 6452
rect 17224 6443 17276 6452
rect 17224 6409 17233 6443
rect 17233 6409 17267 6443
rect 17267 6409 17276 6443
rect 17224 6400 17276 6409
rect 18420 6400 18472 6452
rect 23940 6443 23992 6452
rect 23940 6409 23949 6443
rect 23949 6409 23983 6443
rect 23983 6409 23992 6443
rect 23940 6400 23992 6409
rect 25136 6443 25188 6452
rect 25136 6409 25145 6443
rect 25145 6409 25179 6443
rect 25179 6409 25188 6443
rect 25136 6400 25188 6409
rect 8116 6332 8168 6384
rect 8484 6332 8536 6384
rect 9680 6332 9732 6384
rect 9404 6307 9456 6316
rect 3700 6239 3752 6248
rect 3700 6205 3709 6239
rect 3709 6205 3743 6239
rect 3743 6205 3752 6239
rect 3700 6196 3752 6205
rect 3976 6196 4028 6248
rect 5356 6196 5408 6248
rect 9404 6273 9413 6307
rect 9413 6273 9447 6307
rect 9447 6273 9456 6307
rect 9404 6264 9456 6273
rect 10048 6264 10100 6316
rect 15108 6264 15160 6316
rect 5632 6196 5684 6248
rect 9588 6239 9640 6248
rect 9588 6205 9597 6239
rect 9597 6205 9631 6239
rect 9631 6205 9640 6239
rect 9588 6196 9640 6205
rect 9772 6239 9824 6248
rect 9772 6205 9778 6239
rect 9778 6205 9824 6239
rect 9772 6196 9824 6205
rect 10692 6196 10744 6248
rect 11152 6239 11204 6248
rect 11152 6205 11161 6239
rect 11161 6205 11195 6239
rect 11195 6205 11204 6239
rect 11152 6196 11204 6205
rect 16488 6196 16540 6248
rect 16764 6196 16816 6248
rect 17132 6196 17184 6248
rect 1676 6128 1728 6137
rect 3516 6128 3568 6180
rect 7748 6128 7800 6180
rect 8024 6171 8076 6180
rect 8024 6137 8033 6171
rect 8033 6137 8067 6171
rect 8067 6137 8076 6171
rect 8024 6128 8076 6137
rect 8576 6128 8628 6180
rect 8760 6171 8812 6180
rect 8760 6137 8769 6171
rect 8769 6137 8803 6171
rect 8803 6137 8812 6171
rect 8760 6128 8812 6137
rect 9312 6128 9364 6180
rect 11244 6128 11296 6180
rect 3976 6060 4028 6112
rect 4068 6060 4120 6112
rect 4620 6060 4672 6112
rect 4896 6060 4948 6112
rect 6184 6060 6236 6112
rect 7012 6103 7064 6112
rect 7012 6069 7021 6103
rect 7021 6069 7055 6103
rect 7055 6069 7064 6103
rect 7012 6060 7064 6069
rect 8116 6060 8168 6112
rect 8208 6060 8260 6112
rect 12716 6060 12768 6112
rect 14740 6128 14792 6180
rect 15476 6128 15528 6180
rect 13360 6103 13412 6112
rect 13360 6069 13369 6103
rect 13369 6069 13403 6103
rect 13403 6069 13412 6103
rect 13360 6060 13412 6069
rect 14004 6103 14056 6112
rect 14004 6069 14013 6103
rect 14013 6069 14047 6103
rect 14047 6069 14056 6103
rect 14004 6060 14056 6069
rect 15936 6103 15988 6112
rect 15936 6069 15945 6103
rect 15945 6069 15979 6103
rect 15979 6069 15988 6103
rect 15936 6060 15988 6069
rect 16212 6103 16264 6112
rect 16212 6069 16221 6103
rect 16221 6069 16255 6103
rect 16255 6069 16264 6103
rect 16212 6060 16264 6069
rect 17040 6060 17092 6112
rect 18880 6196 18932 6248
rect 24860 6171 24912 6180
rect 23204 6060 23256 6112
rect 23940 6060 23992 6112
rect 24860 6137 24869 6171
rect 24869 6137 24903 6171
rect 24903 6137 24912 6171
rect 24860 6128 24912 6137
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1676 5856 1728 5908
rect 2228 5899 2280 5908
rect 2228 5865 2237 5899
rect 2237 5865 2271 5899
rect 2271 5865 2280 5899
rect 2228 5856 2280 5865
rect 3516 5856 3568 5908
rect 3884 5899 3936 5908
rect 3884 5865 3893 5899
rect 3893 5865 3927 5899
rect 3927 5865 3936 5899
rect 3884 5856 3936 5865
rect 6000 5856 6052 5908
rect 6460 5856 6512 5908
rect 8024 5856 8076 5908
rect 8760 5856 8812 5908
rect 11244 5856 11296 5908
rect 11612 5856 11664 5908
rect 12716 5856 12768 5908
rect 15108 5899 15160 5908
rect 15108 5865 15117 5899
rect 15117 5865 15151 5899
rect 15151 5865 15160 5899
rect 15108 5856 15160 5865
rect 15384 5856 15436 5908
rect 2872 5788 2924 5840
rect 1768 5720 1820 5772
rect 3424 5788 3476 5840
rect 4344 5788 4396 5840
rect 4528 5720 4580 5772
rect 6368 5763 6420 5772
rect 6368 5729 6377 5763
rect 6377 5729 6411 5763
rect 6411 5729 6420 5763
rect 6368 5720 6420 5729
rect 6460 5720 6512 5772
rect 8208 5788 8260 5840
rect 9496 5831 9548 5840
rect 9496 5797 9505 5831
rect 9505 5797 9539 5831
rect 9539 5797 9548 5831
rect 9496 5788 9548 5797
rect 7748 5720 7800 5772
rect 7932 5720 7984 5772
rect 8116 5720 8168 5772
rect 9680 5763 9732 5772
rect 9680 5729 9689 5763
rect 9689 5729 9723 5763
rect 9723 5729 9732 5763
rect 9680 5720 9732 5729
rect 9772 5720 9824 5772
rect 12256 5788 12308 5840
rect 16672 5831 16724 5840
rect 16672 5797 16681 5831
rect 16681 5797 16715 5831
rect 16715 5797 16724 5831
rect 16672 5788 16724 5797
rect 17776 5788 17828 5840
rect 23204 5788 23256 5840
rect 13912 5763 13964 5772
rect 2596 5652 2648 5704
rect 3332 5652 3384 5704
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 6828 5695 6880 5704
rect 6828 5661 6837 5695
rect 6837 5661 6871 5695
rect 6871 5661 6880 5695
rect 6828 5652 6880 5661
rect 8208 5695 8260 5704
rect 8208 5661 8217 5695
rect 8217 5661 8251 5695
rect 8251 5661 8260 5695
rect 8208 5652 8260 5661
rect 9128 5652 9180 5704
rect 10048 5695 10100 5704
rect 3240 5584 3292 5636
rect 5540 5584 5592 5636
rect 6184 5584 6236 5636
rect 9680 5584 9732 5636
rect 10048 5661 10057 5695
rect 10057 5661 10091 5695
rect 10091 5661 10100 5695
rect 10048 5652 10100 5661
rect 13912 5729 13921 5763
rect 13921 5729 13955 5763
rect 13955 5729 13964 5763
rect 13912 5720 13964 5729
rect 11980 5652 12032 5704
rect 13636 5652 13688 5704
rect 15476 5720 15528 5772
rect 17500 5763 17552 5772
rect 17500 5729 17509 5763
rect 17509 5729 17543 5763
rect 17543 5729 17552 5763
rect 17500 5720 17552 5729
rect 23112 5720 23164 5772
rect 14372 5695 14424 5704
rect 14372 5661 14381 5695
rect 14381 5661 14415 5695
rect 14415 5661 14424 5695
rect 14372 5652 14424 5661
rect 14648 5652 14700 5704
rect 16948 5652 17000 5704
rect 18144 5695 18196 5704
rect 18144 5661 18153 5695
rect 18153 5661 18187 5695
rect 18187 5661 18196 5695
rect 18144 5652 18196 5661
rect 10692 5584 10744 5636
rect 10876 5627 10928 5636
rect 10876 5593 10885 5627
rect 10885 5593 10919 5627
rect 10919 5593 10928 5627
rect 10876 5584 10928 5593
rect 13820 5584 13872 5636
rect 16764 5584 16816 5636
rect 17132 5627 17184 5636
rect 17132 5593 17141 5627
rect 17141 5593 17175 5627
rect 17175 5593 17184 5627
rect 25044 5652 25096 5704
rect 17132 5584 17184 5593
rect 24032 5584 24084 5636
rect 24860 5584 24912 5636
rect 3148 5516 3200 5568
rect 5356 5559 5408 5568
rect 5356 5525 5365 5559
rect 5365 5525 5399 5559
rect 5399 5525 5408 5559
rect 5356 5516 5408 5525
rect 6000 5516 6052 5568
rect 7104 5516 7156 5568
rect 7748 5559 7800 5568
rect 7748 5525 7757 5559
rect 7757 5525 7791 5559
rect 7791 5525 7800 5559
rect 7748 5516 7800 5525
rect 8116 5559 8168 5568
rect 8116 5525 8125 5559
rect 8125 5525 8159 5559
rect 8159 5525 8168 5559
rect 8116 5516 8168 5525
rect 8484 5559 8536 5568
rect 8484 5525 8493 5559
rect 8493 5525 8527 5559
rect 8527 5525 8536 5559
rect 8484 5516 8536 5525
rect 9956 5559 10008 5568
rect 9956 5525 9965 5559
rect 9965 5525 9999 5559
rect 9999 5525 10008 5559
rect 9956 5516 10008 5525
rect 10140 5559 10192 5568
rect 10140 5525 10149 5559
rect 10149 5525 10183 5559
rect 10183 5525 10192 5559
rect 10140 5516 10192 5525
rect 13728 5516 13780 5568
rect 23848 5516 23900 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 1768 5312 1820 5364
rect 4344 5244 4396 5296
rect 5816 5244 5868 5296
rect 6092 5244 6144 5296
rect 112 4972 164 5024
rect 2596 5108 2648 5160
rect 3884 5176 3936 5228
rect 3056 5040 3108 5092
rect 4528 5151 4580 5160
rect 4528 5117 4537 5151
rect 4537 5117 4571 5151
rect 4571 5117 4580 5151
rect 4528 5108 4580 5117
rect 6736 5244 6788 5296
rect 7932 5244 7984 5296
rect 8116 5287 8168 5296
rect 8116 5253 8125 5287
rect 8125 5253 8159 5287
rect 8159 5253 8168 5287
rect 8116 5244 8168 5253
rect 7012 5176 7064 5228
rect 8208 5219 8260 5228
rect 8208 5185 8217 5219
rect 8217 5185 8251 5219
rect 8251 5185 8260 5219
rect 8208 5176 8260 5185
rect 6920 5108 6972 5160
rect 7380 5108 7432 5160
rect 8024 5108 8076 5160
rect 4620 5083 4672 5092
rect 4620 5049 4629 5083
rect 4629 5049 4663 5083
rect 4663 5049 4672 5083
rect 4620 5040 4672 5049
rect 6460 5040 6512 5092
rect 7196 5040 7248 5092
rect 9312 5312 9364 5364
rect 11796 5312 11848 5364
rect 12532 5312 12584 5364
rect 16212 5312 16264 5364
rect 16948 5355 17000 5364
rect 16948 5321 16957 5355
rect 16957 5321 16991 5355
rect 16991 5321 17000 5355
rect 16948 5312 17000 5321
rect 18144 5312 18196 5364
rect 23112 5355 23164 5364
rect 23112 5321 23121 5355
rect 23121 5321 23155 5355
rect 23155 5321 23164 5355
rect 23112 5312 23164 5321
rect 23204 5312 23256 5364
rect 25044 5355 25096 5364
rect 25044 5321 25053 5355
rect 25053 5321 25087 5355
rect 25087 5321 25096 5355
rect 25044 5312 25096 5321
rect 11980 5244 12032 5296
rect 16028 5244 16080 5296
rect 11060 5176 11112 5228
rect 17040 5176 17092 5228
rect 9680 5108 9732 5160
rect 10876 5151 10928 5160
rect 10876 5117 10885 5151
rect 10885 5117 10919 5151
rect 10919 5117 10928 5151
rect 10876 5108 10928 5117
rect 11244 5151 11296 5160
rect 11244 5117 11253 5151
rect 11253 5117 11287 5151
rect 11287 5117 11296 5151
rect 11244 5108 11296 5117
rect 12440 5108 12492 5160
rect 11336 5040 11388 5092
rect 11520 5083 11572 5092
rect 11520 5049 11529 5083
rect 11529 5049 11563 5083
rect 11563 5049 11572 5083
rect 11520 5040 11572 5049
rect 11980 5040 12032 5092
rect 13912 5108 13964 5160
rect 14280 5151 14332 5160
rect 14280 5117 14289 5151
rect 14289 5117 14323 5151
rect 14323 5117 14332 5151
rect 14280 5108 14332 5117
rect 14556 5151 14608 5160
rect 14556 5117 14565 5151
rect 14565 5117 14599 5151
rect 14599 5117 14608 5151
rect 14556 5108 14608 5117
rect 14740 5108 14792 5160
rect 15200 5151 15252 5160
rect 15200 5117 15209 5151
rect 15209 5117 15243 5151
rect 15243 5117 15252 5151
rect 15200 5108 15252 5117
rect 15384 5151 15436 5160
rect 15384 5117 15393 5151
rect 15393 5117 15427 5151
rect 15427 5117 15436 5151
rect 15384 5108 15436 5117
rect 16856 5108 16908 5160
rect 18696 5151 18748 5160
rect 18696 5117 18705 5151
rect 18705 5117 18739 5151
rect 18739 5117 18748 5151
rect 18696 5108 18748 5117
rect 24124 5108 24176 5160
rect 17960 5040 18012 5092
rect 3976 4972 4028 5024
rect 5264 4972 5316 5024
rect 6368 4972 6420 5024
rect 7012 5015 7064 5024
rect 7012 4981 7021 5015
rect 7021 4981 7055 5015
rect 7055 4981 7064 5015
rect 7012 4972 7064 4981
rect 8760 4972 8812 5024
rect 9772 4972 9824 5024
rect 10692 5015 10744 5024
rect 10692 4981 10701 5015
rect 10701 4981 10735 5015
rect 10735 4981 10744 5015
rect 10692 4972 10744 4981
rect 16672 5015 16724 5024
rect 16672 4981 16681 5015
rect 16681 4981 16715 5015
rect 16715 4981 16724 5015
rect 16672 4972 16724 4981
rect 17776 5015 17828 5024
rect 17776 4981 17785 5015
rect 17785 4981 17819 5015
rect 17819 4981 17828 5015
rect 17776 4972 17828 4981
rect 22284 5015 22336 5024
rect 22284 4981 22293 5015
rect 22293 4981 22327 5015
rect 22327 4981 22336 5015
rect 22284 4972 22336 4981
rect 23940 5015 23992 5024
rect 23940 4981 23949 5015
rect 23949 4981 23983 5015
rect 23983 4981 23992 5015
rect 23940 4972 23992 4981
rect 27068 4972 27120 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 2872 4811 2924 4820
rect 2872 4777 2881 4811
rect 2881 4777 2915 4811
rect 2915 4777 2924 4811
rect 2872 4768 2924 4777
rect 4068 4768 4120 4820
rect 5816 4768 5868 4820
rect 6736 4768 6788 4820
rect 7380 4811 7432 4820
rect 7380 4777 7389 4811
rect 7389 4777 7423 4811
rect 7423 4777 7432 4811
rect 7380 4768 7432 4777
rect 1400 4743 1452 4752
rect 1400 4709 1409 4743
rect 1409 4709 1443 4743
rect 1443 4709 1452 4743
rect 1400 4700 1452 4709
rect 2688 4700 2740 4752
rect 4620 4700 4672 4752
rect 7564 4768 7616 4820
rect 7748 4768 7800 4820
rect 10048 4768 10100 4820
rect 11428 4768 11480 4820
rect 13636 4768 13688 4820
rect 14740 4768 14792 4820
rect 14832 4768 14884 4820
rect 15384 4768 15436 4820
rect 15936 4768 15988 4820
rect 7656 4743 7708 4752
rect 7656 4709 7665 4743
rect 7665 4709 7699 4743
rect 7699 4709 7708 4743
rect 7656 4700 7708 4709
rect 7932 4700 7984 4752
rect 10416 4700 10468 4752
rect 11612 4700 11664 4752
rect 12900 4700 12952 4752
rect 15200 4700 15252 4752
rect 16672 4700 16724 4752
rect 1768 4675 1820 4684
rect 1768 4641 1777 4675
rect 1777 4641 1811 4675
rect 1811 4641 1820 4675
rect 1768 4632 1820 4641
rect 2964 4675 3016 4684
rect 2964 4641 2973 4675
rect 2973 4641 3007 4675
rect 3007 4641 3016 4675
rect 2964 4632 3016 4641
rect 6184 4675 6236 4684
rect 6184 4641 6193 4675
rect 6193 4641 6227 4675
rect 6227 4641 6236 4675
rect 6184 4632 6236 4641
rect 6460 4675 6512 4684
rect 6460 4641 6469 4675
rect 6469 4641 6503 4675
rect 6503 4641 6512 4675
rect 6460 4632 6512 4641
rect 8300 4632 8352 4684
rect 4436 4607 4488 4616
rect 4436 4573 4445 4607
rect 4445 4573 4479 4607
rect 4479 4573 4488 4607
rect 4436 4564 4488 4573
rect 6644 4607 6696 4616
rect 3332 4496 3384 4548
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 6644 4564 6696 4573
rect 7564 4607 7616 4616
rect 7564 4573 7573 4607
rect 7573 4573 7607 4607
rect 7607 4573 7616 4607
rect 7564 4564 7616 4573
rect 10508 4607 10560 4616
rect 10508 4573 10517 4607
rect 10517 4573 10551 4607
rect 10551 4573 10560 4607
rect 10508 4564 10560 4573
rect 12348 4632 12400 4684
rect 13268 4632 13320 4684
rect 13820 4675 13872 4684
rect 13820 4641 13829 4675
rect 13829 4641 13863 4675
rect 13863 4641 13872 4675
rect 13820 4632 13872 4641
rect 14280 4632 14332 4684
rect 17776 4768 17828 4820
rect 22560 4743 22612 4752
rect 22560 4709 22569 4743
rect 22569 4709 22603 4743
rect 22603 4709 22612 4743
rect 22560 4700 22612 4709
rect 24124 4743 24176 4752
rect 24124 4709 24133 4743
rect 24133 4709 24167 4743
rect 24167 4709 24176 4743
rect 24124 4700 24176 4709
rect 18788 4675 18840 4684
rect 18788 4641 18797 4675
rect 18797 4641 18831 4675
rect 18831 4641 18840 4675
rect 18788 4632 18840 4641
rect 13912 4564 13964 4616
rect 14188 4607 14240 4616
rect 14188 4573 14197 4607
rect 14197 4573 14231 4607
rect 14231 4573 14240 4607
rect 14188 4564 14240 4573
rect 14372 4564 14424 4616
rect 16672 4564 16724 4616
rect 3884 4428 3936 4480
rect 7012 4496 7064 4548
rect 8668 4496 8720 4548
rect 9956 4496 10008 4548
rect 11888 4496 11940 4548
rect 12624 4496 12676 4548
rect 22468 4607 22520 4616
rect 22468 4573 22477 4607
rect 22477 4573 22511 4607
rect 22511 4573 22520 4607
rect 22468 4564 22520 4573
rect 22744 4607 22796 4616
rect 22744 4573 22753 4607
rect 22753 4573 22787 4607
rect 22787 4573 22796 4607
rect 22744 4564 22796 4573
rect 23848 4564 23900 4616
rect 24032 4607 24084 4616
rect 24032 4573 24041 4607
rect 24041 4573 24075 4607
rect 24075 4573 24084 4607
rect 24032 4564 24084 4573
rect 24216 4564 24268 4616
rect 5448 4471 5500 4480
rect 5448 4437 5457 4471
rect 5457 4437 5491 4471
rect 5491 4437 5500 4471
rect 5448 4428 5500 4437
rect 6920 4471 6972 4480
rect 6920 4437 6929 4471
rect 6929 4437 6963 4471
rect 6963 4437 6972 4471
rect 6920 4428 6972 4437
rect 11336 4428 11388 4480
rect 16304 4471 16356 4480
rect 16304 4437 16313 4471
rect 16313 4437 16347 4471
rect 16347 4437 16356 4471
rect 16304 4428 16356 4437
rect 18696 4428 18748 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 1860 4267 1912 4276
rect 1860 4233 1869 4267
rect 1869 4233 1903 4267
rect 1903 4233 1912 4267
rect 1860 4224 1912 4233
rect 2964 4267 3016 4276
rect 2964 4233 2973 4267
rect 2973 4233 3007 4267
rect 3007 4233 3016 4267
rect 2964 4224 3016 4233
rect 3700 4224 3752 4276
rect 3884 4267 3936 4276
rect 3884 4233 3893 4267
rect 3893 4233 3927 4267
rect 3927 4233 3936 4267
rect 3884 4224 3936 4233
rect 4252 4267 4304 4276
rect 4252 4233 4261 4267
rect 4261 4233 4295 4267
rect 4295 4233 4304 4267
rect 4252 4224 4304 4233
rect 4620 4267 4672 4276
rect 4620 4233 4629 4267
rect 4629 4233 4663 4267
rect 4663 4233 4672 4267
rect 4620 4224 4672 4233
rect 5172 4224 5224 4276
rect 4528 4156 4580 4208
rect 6184 4199 6236 4208
rect 6184 4165 6193 4199
rect 6193 4165 6227 4199
rect 6227 4165 6236 4199
rect 6184 4156 6236 4165
rect 3976 4131 4028 4140
rect 3976 4097 3985 4131
rect 3985 4097 4019 4131
rect 4019 4097 4028 4131
rect 3976 4088 4028 4097
rect 4804 4088 4856 4140
rect 5724 4088 5776 4140
rect 1768 4063 1820 4072
rect 1768 4029 1777 4063
rect 1777 4029 1811 4063
rect 1811 4029 1820 4063
rect 1768 4020 1820 4029
rect 2504 4063 2556 4072
rect 2504 4029 2513 4063
rect 2513 4029 2547 4063
rect 2547 4029 2556 4063
rect 2504 4020 2556 4029
rect 3240 4020 3292 4072
rect 3608 4063 3660 4072
rect 3608 4029 3617 4063
rect 3617 4029 3651 4063
rect 3651 4029 3660 4063
rect 3608 4020 3660 4029
rect 5264 4063 5316 4072
rect 5264 4029 5273 4063
rect 5273 4029 5307 4063
rect 5307 4029 5316 4063
rect 5264 4020 5316 4029
rect 5448 4020 5500 4072
rect 8116 4224 8168 4276
rect 8208 4224 8260 4276
rect 10508 4224 10560 4276
rect 10876 4224 10928 4276
rect 13268 4224 13320 4276
rect 14004 4224 14056 4276
rect 16856 4267 16908 4276
rect 16856 4233 16865 4267
rect 16865 4233 16899 4267
rect 16899 4233 16908 4267
rect 16856 4224 16908 4233
rect 22468 4224 22520 4276
rect 23940 4267 23992 4276
rect 23940 4233 23949 4267
rect 23949 4233 23983 4267
rect 23983 4233 23992 4267
rect 23940 4224 23992 4233
rect 6736 4156 6788 4208
rect 7380 4199 7432 4208
rect 7380 4165 7389 4199
rect 7389 4165 7423 4199
rect 7423 4165 7432 4199
rect 7380 4156 7432 4165
rect 8668 4199 8720 4208
rect 8668 4165 8677 4199
rect 8677 4165 8711 4199
rect 8711 4165 8720 4199
rect 8668 4156 8720 4165
rect 11428 4156 11480 4208
rect 13544 4156 13596 4208
rect 17040 4156 17092 4208
rect 17224 4156 17276 4208
rect 18788 4156 18840 4208
rect 24124 4156 24176 4208
rect 4804 3952 4856 4004
rect 8208 4088 8260 4140
rect 6644 4020 6696 4072
rect 9680 4063 9732 4072
rect 9680 4029 9698 4063
rect 9698 4029 9732 4063
rect 11888 4088 11940 4140
rect 12532 4131 12584 4140
rect 12532 4097 12541 4131
rect 12541 4097 12575 4131
rect 12575 4097 12584 4131
rect 12532 4088 12584 4097
rect 13820 4088 13872 4140
rect 14832 4131 14884 4140
rect 10416 4063 10468 4072
rect 9680 4020 9732 4029
rect 10416 4029 10425 4063
rect 10425 4029 10459 4063
rect 10459 4029 10468 4063
rect 10416 4020 10468 4029
rect 10692 4020 10744 4072
rect 11980 4020 12032 4072
rect 14832 4097 14841 4131
rect 14841 4097 14875 4131
rect 14875 4097 14884 4131
rect 14832 4088 14884 4097
rect 15292 4088 15344 4140
rect 18972 4088 19024 4140
rect 22284 4088 22336 4140
rect 22744 4131 22796 4140
rect 22744 4097 22753 4131
rect 22753 4097 22787 4131
rect 22787 4097 22796 4131
rect 22744 4088 22796 4097
rect 24216 4088 24268 4140
rect 14740 4063 14792 4072
rect 14740 4029 14749 4063
rect 14749 4029 14783 4063
rect 14783 4029 14792 4063
rect 14740 4020 14792 4029
rect 16672 4020 16724 4072
rect 17224 4020 17276 4072
rect 21088 4063 21140 4072
rect 21088 4029 21097 4063
rect 21097 4029 21131 4063
rect 21131 4029 21140 4063
rect 21088 4020 21140 4029
rect 7656 3952 7708 4004
rect 9128 3952 9180 4004
rect 12624 3995 12676 4004
rect 12624 3961 12633 3995
rect 12633 3961 12667 3995
rect 12667 3961 12676 3995
rect 12624 3952 12676 3961
rect 13820 3952 13872 4004
rect 15844 3995 15896 4004
rect 7380 3884 7432 3936
rect 9312 3884 9364 3936
rect 9404 3884 9456 3936
rect 12348 3884 12400 3936
rect 13544 3884 13596 3936
rect 15844 3961 15853 3995
rect 15853 3961 15887 3995
rect 15887 3961 15896 3995
rect 15844 3952 15896 3961
rect 16856 3952 16908 4004
rect 17776 3952 17828 4004
rect 18052 3995 18104 4004
rect 18052 3961 18061 3995
rect 18061 3961 18095 3995
rect 18095 3961 18104 3995
rect 18052 3952 18104 3961
rect 22192 3995 22244 4004
rect 22192 3961 22201 3995
rect 22201 3961 22235 3995
rect 22235 3961 22244 3995
rect 22192 3952 22244 3961
rect 24216 3995 24268 4004
rect 24216 3961 24225 3995
rect 24225 3961 24259 3995
rect 24259 3961 24268 3995
rect 24216 3952 24268 3961
rect 18144 3884 18196 3936
rect 19984 3884 20036 3936
rect 22560 3884 22612 3936
rect 23940 3884 23992 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1584 3680 1636 3732
rect 3608 3723 3660 3732
rect 3608 3689 3617 3723
rect 3617 3689 3651 3723
rect 3651 3689 3660 3723
rect 3608 3680 3660 3689
rect 3976 3680 4028 3732
rect 4988 3680 5040 3732
rect 6460 3680 6512 3732
rect 6644 3680 6696 3732
rect 7932 3723 7984 3732
rect 2596 3612 2648 3664
rect 3148 3655 3200 3664
rect 3148 3621 3157 3655
rect 3157 3621 3191 3655
rect 3191 3621 3200 3655
rect 3148 3612 3200 3621
rect 3240 3612 3292 3664
rect 1308 3544 1360 3596
rect 1860 3544 1912 3596
rect 4712 3544 4764 3596
rect 6736 3612 6788 3664
rect 7932 3689 7941 3723
rect 7941 3689 7975 3723
rect 7975 3689 7984 3723
rect 7932 3680 7984 3689
rect 9312 3723 9364 3732
rect 9312 3689 9321 3723
rect 9321 3689 9355 3723
rect 9355 3689 9364 3723
rect 9312 3680 9364 3689
rect 10876 3723 10928 3732
rect 10876 3689 10885 3723
rect 10885 3689 10919 3723
rect 10919 3689 10928 3723
rect 10876 3680 10928 3689
rect 14280 3680 14332 3732
rect 14740 3680 14792 3732
rect 15844 3680 15896 3732
rect 17960 3680 18012 3732
rect 22284 3680 22336 3732
rect 24032 3680 24084 3732
rect 9864 3587 9916 3596
rect 9864 3553 9873 3587
rect 9873 3553 9907 3587
rect 9907 3553 9916 3587
rect 9864 3544 9916 3553
rect 10324 3587 10376 3596
rect 10324 3553 10333 3587
rect 10333 3553 10367 3587
rect 10367 3553 10376 3587
rect 10324 3544 10376 3553
rect 10692 3612 10744 3664
rect 11612 3612 11664 3664
rect 13544 3612 13596 3664
rect 15292 3612 15344 3664
rect 17224 3655 17276 3664
rect 17224 3621 17233 3655
rect 17233 3621 17267 3655
rect 17267 3621 17276 3655
rect 17224 3612 17276 3621
rect 17776 3612 17828 3664
rect 18696 3612 18748 3664
rect 19064 3612 19116 3664
rect 22192 3655 22244 3664
rect 22192 3621 22201 3655
rect 22201 3621 22235 3655
rect 22235 3621 22244 3655
rect 22192 3612 22244 3621
rect 1952 3476 2004 3528
rect 3792 3476 3844 3528
rect 3056 3408 3108 3460
rect 4252 3408 4304 3460
rect 4436 3408 4488 3460
rect 5540 3408 5592 3460
rect 6092 3476 6144 3528
rect 5724 3408 5776 3460
rect 6644 3408 6696 3460
rect 8208 3476 8260 3528
rect 11520 3476 11572 3528
rect 11980 3476 12032 3528
rect 13636 3476 13688 3528
rect 13820 3519 13872 3528
rect 13820 3485 13829 3519
rect 13829 3485 13863 3519
rect 13863 3485 13872 3519
rect 13820 3476 13872 3485
rect 14556 3476 14608 3528
rect 6828 3408 6880 3460
rect 12532 3408 12584 3460
rect 848 3340 900 3392
rect 1768 3340 1820 3392
rect 3424 3340 3476 3392
rect 4620 3383 4672 3392
rect 4620 3349 4629 3383
rect 4629 3349 4663 3383
rect 4663 3349 4672 3383
rect 4620 3340 4672 3349
rect 4988 3383 5040 3392
rect 4988 3349 4997 3383
rect 4997 3349 5031 3383
rect 5031 3349 5040 3383
rect 4988 3340 5040 3349
rect 6276 3340 6328 3392
rect 8760 3340 8812 3392
rect 12808 3340 12860 3392
rect 16672 3340 16724 3392
rect 18420 3476 18472 3528
rect 20904 3544 20956 3596
rect 22560 3587 22612 3596
rect 22560 3553 22569 3587
rect 22569 3553 22603 3587
rect 22603 3553 22612 3587
rect 22560 3544 22612 3553
rect 22744 3544 22796 3596
rect 23480 3544 23532 3596
rect 24216 3544 24268 3596
rect 24952 3544 25004 3596
rect 18972 3519 19024 3528
rect 18972 3485 18981 3519
rect 18981 3485 19015 3519
rect 19015 3485 19024 3519
rect 18972 3476 19024 3485
rect 17408 3340 17460 3392
rect 23388 3340 23440 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1952 3179 2004 3188
rect 1952 3145 1961 3179
rect 1961 3145 1995 3179
rect 1995 3145 2004 3179
rect 1952 3136 2004 3145
rect 3056 3179 3108 3188
rect 3056 3145 3065 3179
rect 3065 3145 3099 3179
rect 3099 3145 3108 3179
rect 3056 3136 3108 3145
rect 3424 3179 3476 3188
rect 3424 3145 3433 3179
rect 3433 3145 3467 3179
rect 3467 3145 3476 3179
rect 3424 3136 3476 3145
rect 5172 3136 5224 3188
rect 6000 3136 6052 3188
rect 6276 3179 6328 3188
rect 6276 3145 6285 3179
rect 6285 3145 6319 3179
rect 6319 3145 6328 3179
rect 6276 3136 6328 3145
rect 6736 3136 6788 3188
rect 3608 3068 3660 3120
rect 2688 2975 2740 2984
rect 2688 2941 2697 2975
rect 2697 2941 2731 2975
rect 2731 2941 2740 2975
rect 2688 2932 2740 2941
rect 4620 3000 4672 3052
rect 4988 3000 5040 3052
rect 6092 3000 6144 3052
rect 8300 3136 8352 3188
rect 9588 3136 9640 3188
rect 9864 3136 9916 3188
rect 10324 3179 10376 3188
rect 10324 3145 10333 3179
rect 10333 3145 10367 3179
rect 10367 3145 10376 3179
rect 10324 3136 10376 3145
rect 11612 3136 11664 3188
rect 13544 3179 13596 3188
rect 10692 3068 10744 3120
rect 13544 3145 13553 3179
rect 13553 3145 13587 3179
rect 13587 3145 13596 3179
rect 13544 3136 13596 3145
rect 14188 3136 14240 3188
rect 8944 3000 8996 3052
rect 10876 3043 10928 3052
rect 10876 3009 10885 3043
rect 10885 3009 10919 3043
rect 10919 3009 10928 3043
rect 10876 3000 10928 3009
rect 13360 3000 13412 3052
rect 8116 2932 8168 2984
rect 2780 2907 2832 2916
rect 2780 2873 2789 2907
rect 2789 2873 2823 2907
rect 2823 2873 2832 2907
rect 2780 2864 2832 2873
rect 3424 2864 3476 2916
rect 4344 2907 4396 2916
rect 4344 2873 4353 2907
rect 4353 2873 4387 2907
rect 4387 2873 4396 2907
rect 4344 2864 4396 2873
rect 4896 2864 4948 2916
rect 7380 2907 7432 2916
rect 4712 2839 4764 2848
rect 4712 2805 4721 2839
rect 4721 2805 4755 2839
rect 4755 2805 4764 2839
rect 7380 2873 7389 2907
rect 7389 2873 7423 2907
rect 7423 2873 7432 2907
rect 7380 2864 7432 2873
rect 8852 2864 8904 2916
rect 4712 2796 4764 2805
rect 8392 2796 8444 2848
rect 9128 2839 9180 2848
rect 9128 2805 9137 2839
rect 9137 2805 9171 2839
rect 9171 2805 9180 2839
rect 9128 2796 9180 2805
rect 10692 2907 10744 2916
rect 10692 2873 10701 2907
rect 10701 2873 10735 2907
rect 10735 2873 10744 2907
rect 12532 2907 12584 2916
rect 10692 2864 10744 2873
rect 12532 2873 12541 2907
rect 12541 2873 12575 2907
rect 12575 2873 12584 2907
rect 12532 2864 12584 2873
rect 15384 3136 15436 3188
rect 17040 3136 17092 3188
rect 17224 3136 17276 3188
rect 18052 3136 18104 3188
rect 19064 3179 19116 3188
rect 19064 3145 19073 3179
rect 19073 3145 19107 3179
rect 19107 3145 19116 3179
rect 19064 3136 19116 3145
rect 22560 3136 22612 3188
rect 23480 3179 23532 3188
rect 23480 3145 23489 3179
rect 23489 3145 23523 3179
rect 23523 3145 23532 3179
rect 23480 3136 23532 3145
rect 24952 3136 25004 3188
rect 26976 3136 27028 3188
rect 15292 3068 15344 3120
rect 16672 3043 16724 3052
rect 16672 3009 16681 3043
rect 16681 3009 16715 3043
rect 16715 3009 16724 3043
rect 16672 3000 16724 3009
rect 18144 3043 18196 3052
rect 18144 3009 18153 3043
rect 18153 3009 18187 3043
rect 18187 3009 18196 3043
rect 18144 3000 18196 3009
rect 18420 3043 18472 3052
rect 18420 3009 18429 3043
rect 18429 3009 18463 3043
rect 18463 3009 18472 3043
rect 18420 3000 18472 3009
rect 22652 3043 22704 3052
rect 22652 3009 22661 3043
rect 22661 3009 22695 3043
rect 22695 3009 22704 3043
rect 22652 3000 22704 3009
rect 11152 2796 11204 2848
rect 16396 2907 16448 2916
rect 16396 2873 16405 2907
rect 16405 2873 16439 2907
rect 16439 2873 16448 2907
rect 16396 2864 16448 2873
rect 15292 2796 15344 2848
rect 15384 2796 15436 2848
rect 17868 2864 17920 2916
rect 18052 2796 18104 2848
rect 25780 2932 25832 2984
rect 19432 2839 19484 2848
rect 19432 2805 19441 2839
rect 19441 2805 19475 2839
rect 19475 2805 19484 2839
rect 19432 2796 19484 2805
rect 20904 2839 20956 2848
rect 20904 2805 20913 2839
rect 20913 2805 20947 2839
rect 20947 2805 20956 2839
rect 20904 2796 20956 2805
rect 20996 2796 21048 2848
rect 21456 2796 21508 2848
rect 23112 2796 23164 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 1860 2635 1912 2644
rect 1860 2601 1869 2635
rect 1869 2601 1903 2635
rect 1903 2601 1912 2635
rect 1860 2592 1912 2601
rect 2780 2592 2832 2644
rect 2228 2567 2280 2576
rect 2228 2533 2237 2567
rect 2237 2533 2271 2567
rect 2271 2533 2280 2567
rect 2228 2524 2280 2533
rect 3240 2524 3292 2576
rect 4528 2592 4580 2644
rect 5080 2635 5132 2644
rect 5080 2601 5089 2635
rect 5089 2601 5123 2635
rect 5123 2601 5132 2635
rect 5908 2635 5960 2644
rect 5080 2592 5132 2601
rect 5172 2524 5224 2576
rect 5908 2601 5917 2635
rect 5917 2601 5951 2635
rect 5951 2601 5960 2635
rect 5908 2592 5960 2601
rect 6920 2592 6972 2644
rect 8116 2592 8168 2644
rect 10692 2592 10744 2644
rect 11152 2635 11204 2644
rect 11152 2601 11161 2635
rect 11161 2601 11195 2635
rect 11195 2601 11204 2635
rect 11152 2592 11204 2601
rect 11980 2635 12032 2644
rect 5356 2524 5408 2576
rect 8208 2567 8260 2576
rect 6092 2456 6144 2508
rect 7656 2456 7708 2508
rect 2596 2320 2648 2372
rect 4804 2320 4856 2372
rect 5632 2431 5684 2440
rect 5632 2397 5641 2431
rect 5641 2397 5675 2431
rect 5675 2397 5684 2431
rect 5632 2388 5684 2397
rect 8208 2533 8217 2567
rect 8217 2533 8251 2567
rect 8251 2533 8260 2567
rect 8208 2524 8260 2533
rect 8300 2567 8352 2576
rect 8300 2533 8309 2567
rect 8309 2533 8343 2567
rect 8343 2533 8352 2567
rect 9496 2567 9548 2576
rect 8300 2524 8352 2533
rect 9496 2533 9505 2567
rect 9505 2533 9539 2567
rect 9539 2533 9548 2567
rect 9496 2524 9548 2533
rect 10876 2524 10928 2576
rect 11980 2601 11989 2635
rect 11989 2601 12023 2635
rect 12023 2601 12032 2635
rect 11980 2592 12032 2601
rect 12808 2567 12860 2576
rect 12808 2533 12817 2567
rect 12817 2533 12851 2567
rect 12851 2533 12860 2567
rect 13360 2567 13412 2576
rect 12808 2524 12860 2533
rect 13360 2533 13369 2567
rect 13369 2533 13403 2567
rect 13403 2533 13412 2567
rect 13360 2524 13412 2533
rect 14556 2592 14608 2644
rect 18144 2635 18196 2644
rect 14648 2524 14700 2576
rect 15384 2524 15436 2576
rect 16672 2524 16724 2576
rect 8852 2499 8904 2508
rect 8852 2465 8861 2499
rect 8861 2465 8895 2499
rect 8895 2465 8904 2499
rect 8852 2456 8904 2465
rect 9680 2456 9732 2508
rect 11428 2499 11480 2508
rect 11428 2465 11437 2499
rect 11437 2465 11471 2499
rect 11471 2465 11480 2499
rect 11428 2456 11480 2465
rect 13912 2456 13964 2508
rect 8300 2388 8352 2440
rect 4436 2252 4488 2304
rect 7656 2295 7708 2304
rect 7656 2261 7665 2295
rect 7665 2261 7699 2295
rect 7699 2261 7708 2295
rect 7656 2252 7708 2261
rect 12808 2252 12860 2304
rect 13728 2295 13780 2304
rect 13728 2261 13737 2295
rect 13737 2261 13771 2295
rect 13771 2261 13780 2295
rect 13728 2252 13780 2261
rect 16396 2456 16448 2508
rect 17408 2524 17460 2576
rect 17040 2499 17092 2508
rect 17040 2465 17049 2499
rect 17049 2465 17083 2499
rect 17083 2465 17092 2499
rect 18144 2601 18153 2635
rect 18153 2601 18187 2635
rect 18187 2601 18196 2635
rect 18144 2592 18196 2601
rect 17868 2524 17920 2576
rect 17040 2456 17092 2465
rect 20996 2592 21048 2644
rect 23388 2635 23440 2644
rect 23388 2601 23397 2635
rect 23397 2601 23431 2635
rect 23431 2601 23440 2635
rect 23388 2592 23440 2601
rect 20720 2456 20772 2508
rect 16028 2388 16080 2440
rect 15384 2320 15436 2372
rect 18144 2320 18196 2372
rect 22744 2320 22796 2372
rect 23664 2320 23716 2372
rect 17040 2252 17092 2304
rect 19800 2252 19852 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 7656 1504 7708 1556
rect 10692 1504 10744 1556
rect 17316 76 17368 128
rect 19156 76 19208 128
<< metal2 >>
rect 20 27532 72 27538
rect 1030 27532 1086 28000
rect 1030 27520 1032 27532
rect 20 27474 72 27480
rect 1084 27520 1086 27532
rect 3146 27532 3202 28000
rect 3146 27520 3148 27532
rect 1032 27474 1084 27480
rect 3200 27520 3202 27532
rect 3976 27532 4028 27538
rect 3148 27474 3200 27480
rect 5262 27520 5318 28000
rect 7470 27520 7526 28000
rect 9586 27520 9642 28000
rect 11702 27520 11758 28000
rect 13910 27520 13966 28000
rect 16026 27554 16082 28000
rect 15764 27526 16082 27554
rect 3976 27474 4028 27480
rect 32 13938 60 27474
rect 1044 27443 1072 27474
rect 3160 27443 3188 27474
rect 1030 26480 1086 26489
rect 1030 26415 1086 26424
rect 110 24984 166 24993
rect 110 24919 166 24928
rect 124 23186 152 24919
rect 1044 23662 1072 26415
rect 1032 23656 1084 23662
rect 1032 23598 1084 23604
rect 3792 23588 3844 23594
rect 3792 23530 3844 23536
rect 112 23180 164 23186
rect 112 23122 164 23128
rect 1584 23180 1636 23186
rect 1584 23122 1636 23128
rect 1596 22778 1624 23122
rect 2504 22976 2556 22982
rect 2504 22918 2556 22924
rect 1584 22772 1636 22778
rect 1584 22714 1636 22720
rect 1214 22400 1270 22409
rect 1214 22335 1270 22344
rect 1228 21486 1256 22335
rect 1216 21480 1268 21486
rect 1216 21422 1268 21428
rect 110 21040 166 21049
rect 166 20998 244 21026
rect 110 20975 166 20984
rect 110 16960 166 16969
rect 110 16895 166 16904
rect 124 15609 152 16895
rect 216 16658 244 20998
rect 204 16652 256 16658
rect 204 16594 256 16600
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 110 15600 166 15609
rect 110 15535 166 15544
rect 1582 14648 1638 14657
rect 1582 14583 1638 14592
rect 1596 14346 1624 14583
rect 2424 14482 2452 15846
rect 2412 14476 2464 14482
rect 2412 14418 2464 14424
rect 1584 14340 1636 14346
rect 1584 14282 1636 14288
rect 2424 14074 2452 14418
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 20 13932 72 13938
rect 20 13874 72 13880
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1584 13728 1636 13734
rect 1584 13670 1636 13676
rect 1596 13569 1624 13670
rect 1582 13560 1638 13569
rect 1688 13530 1716 13806
rect 1582 13495 1638 13504
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 2516 13326 2544 22918
rect 2964 13796 3016 13802
rect 2964 13738 3016 13744
rect 2688 13728 2740 13734
rect 2688 13670 2740 13676
rect 2596 13456 2648 13462
rect 2596 13398 2648 13404
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2332 12442 2360 13262
rect 2608 12850 2636 13398
rect 2700 12918 2728 13670
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 2688 12912 2740 12918
rect 2688 12854 2740 12860
rect 2596 12844 2648 12850
rect 2596 12786 2648 12792
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2596 12368 2648 12374
rect 2700 12356 2728 12854
rect 2648 12328 2728 12356
rect 2596 12310 2648 12316
rect 1676 12096 1728 12102
rect 1676 12038 1728 12044
rect 1688 11830 1716 12038
rect 1676 11824 1728 11830
rect 1676 11766 1728 11772
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1676 10668 1728 10674
rect 1676 10610 1728 10616
rect 1688 9722 1716 10610
rect 1780 9926 1808 11154
rect 1964 11150 1992 11630
rect 2136 11620 2188 11626
rect 2136 11562 2188 11568
rect 1952 11144 2004 11150
rect 1952 11086 2004 11092
rect 1858 10432 1914 10441
rect 1858 10367 1914 10376
rect 1768 9920 1820 9926
rect 1768 9862 1820 9868
rect 1676 9716 1728 9722
rect 1676 9658 1728 9664
rect 1780 9489 1808 9862
rect 1872 9518 1900 10367
rect 1860 9512 1912 9518
rect 1766 9480 1822 9489
rect 1860 9454 1912 9460
rect 1766 9415 1822 9424
rect 2148 9217 2176 11562
rect 2608 11354 2636 12310
rect 2884 12238 2912 13262
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2976 11898 3004 13738
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3160 12306 3188 13126
rect 3332 12776 3384 12782
rect 3332 12718 3384 12724
rect 3344 12374 3372 12718
rect 3332 12368 3384 12374
rect 3332 12310 3384 12316
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 3700 12300 3752 12306
rect 3700 12242 3752 12248
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2976 11558 3004 11834
rect 3712 11694 3740 12242
rect 3700 11688 3752 11694
rect 3700 11630 3752 11636
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2596 11348 2648 11354
rect 2596 11290 2648 11296
rect 2688 11212 2740 11218
rect 2688 11154 2740 11160
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2424 10538 2452 10950
rect 2700 10810 2728 11154
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 2412 10532 2464 10538
rect 2412 10474 2464 10480
rect 2228 10464 2280 10470
rect 2280 10424 2360 10452
rect 2228 10406 2280 10412
rect 2228 10056 2280 10062
rect 2228 9998 2280 10004
rect 2240 9586 2268 9998
rect 2332 9926 2360 10424
rect 2424 9994 2452 10474
rect 2884 10470 2912 11154
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 2872 10464 2924 10470
rect 2872 10406 2924 10412
rect 2780 10192 2832 10198
rect 2780 10134 2832 10140
rect 2412 9988 2464 9994
rect 2412 9930 2464 9936
rect 2320 9920 2372 9926
rect 2320 9862 2372 9868
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2134 9208 2190 9217
rect 2332 9160 2360 9862
rect 2134 9143 2190 9152
rect 2240 9132 2360 9160
rect 1400 8832 1452 8838
rect 1400 8774 1452 8780
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 1412 8362 1440 8774
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1400 8356 1452 8362
rect 1400 8298 1452 8304
rect 112 5024 164 5030
rect 112 4966 164 4972
rect 124 1057 152 4966
rect 1412 4758 1440 8298
rect 1768 8288 1820 8294
rect 1768 8230 1820 8236
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 1688 6186 1716 6598
rect 1584 6180 1636 6186
rect 1584 6122 1636 6128
rect 1676 6180 1728 6186
rect 1676 6122 1728 6128
rect 1400 4752 1452 4758
rect 1400 4694 1452 4700
rect 1306 4584 1362 4593
rect 1306 4519 1362 4528
rect 1320 3602 1348 4519
rect 1596 3738 1624 6122
rect 1688 5914 1716 6122
rect 1676 5908 1728 5914
rect 1676 5850 1728 5856
rect 1780 5778 1808 8230
rect 1964 8022 1992 8434
rect 1952 8016 2004 8022
rect 1952 7958 2004 7964
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1872 6798 1900 7278
rect 1964 7188 1992 7958
rect 2056 7886 2084 8774
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2240 7750 2268 9132
rect 2228 7744 2280 7750
rect 2228 7686 2280 7692
rect 2044 7200 2096 7206
rect 1964 7160 2044 7188
rect 2044 7142 2096 7148
rect 1860 6792 1912 6798
rect 1860 6734 1912 6740
rect 1768 5772 1820 5778
rect 1768 5714 1820 5720
rect 1780 5370 1808 5714
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 1768 4684 1820 4690
rect 1768 4626 1820 4632
rect 1780 4078 1808 4626
rect 1872 4282 1900 6734
rect 2056 5953 2084 7142
rect 2240 6866 2268 7686
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 2042 5944 2098 5953
rect 2240 5914 2268 6802
rect 2424 6322 2452 9930
rect 2596 9920 2648 9926
rect 2596 9862 2648 9868
rect 2504 8288 2556 8294
rect 2504 8230 2556 8236
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2042 5879 2098 5888
rect 2228 5908 2280 5914
rect 1860 4276 1912 4282
rect 1860 4218 1912 4224
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 1308 3596 1360 3602
rect 1308 3538 1360 3544
rect 1780 3398 1808 4014
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 848 3392 900 3398
rect 848 3334 900 3340
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 110 1048 166 1057
rect 110 983 166 992
rect 570 82 626 480
rect 860 82 888 3334
rect 1872 2650 1900 3538
rect 1952 3528 2004 3534
rect 1952 3470 2004 3476
rect 1964 3194 1992 3470
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 1860 2644 1912 2650
rect 1860 2586 1912 2592
rect 570 54 888 82
rect 1674 82 1730 480
rect 2056 82 2084 5879
rect 2228 5850 2280 5856
rect 2516 4078 2544 8230
rect 2608 5710 2636 9862
rect 2792 9518 2820 10134
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2700 9178 2728 9318
rect 2792 9178 2820 9454
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2700 8498 2728 9114
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2792 7206 2820 7822
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2884 7018 2912 10406
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3160 9722 3188 9998
rect 3148 9716 3200 9722
rect 3148 9658 3200 9664
rect 3252 9178 3280 11018
rect 3332 9988 3384 9994
rect 3332 9930 3384 9936
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 2964 8356 3016 8362
rect 2964 8298 3016 8304
rect 2976 7750 3004 8298
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2976 7478 3004 7686
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 2976 7342 3004 7414
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 2792 6990 2912 7018
rect 2976 7002 3004 7278
rect 3238 7168 3294 7177
rect 3238 7103 3294 7112
rect 2964 6996 3016 7002
rect 2596 5704 2648 5710
rect 2648 5664 2728 5692
rect 2596 5646 2648 5652
rect 2596 5160 2648 5166
rect 2596 5102 2648 5108
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 2226 2680 2282 2689
rect 2226 2615 2282 2624
rect 2240 2582 2268 2615
rect 2228 2576 2280 2582
rect 2228 2518 2280 2524
rect 1674 54 2084 82
rect 2516 82 2544 4014
rect 2608 3670 2636 5102
rect 2700 4758 2728 5664
rect 2688 4752 2740 4758
rect 2688 4694 2740 4700
rect 2792 4154 2820 6990
rect 2964 6938 3016 6944
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 2962 6488 3018 6497
rect 2962 6423 3018 6432
rect 2872 5840 2924 5846
rect 2872 5782 2924 5788
rect 2884 4826 2912 5782
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2976 4690 3004 6423
rect 3160 5574 3188 6802
rect 3252 6254 3280 7103
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3252 5642 3280 6190
rect 3344 5710 3372 9930
rect 3620 9625 3648 11086
rect 3700 10804 3752 10810
rect 3700 10746 3752 10752
rect 3606 9616 3662 9625
rect 3606 9551 3662 9560
rect 3606 9072 3662 9081
rect 3606 9007 3608 9016
rect 3660 9007 3662 9016
rect 3608 8978 3660 8984
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3528 8430 3556 8774
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3516 7336 3568 7342
rect 3620 7324 3648 8978
rect 3712 8430 3740 10746
rect 3804 8945 3832 23530
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3896 11354 3924 12174
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3988 11234 4016 27474
rect 5276 23866 5304 27520
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6092 24336 6144 24342
rect 6092 24278 6144 24284
rect 6000 24200 6052 24206
rect 6000 24142 6052 24148
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5264 23860 5316 23866
rect 5264 23802 5316 23808
rect 5276 23662 5304 23802
rect 6012 23798 6040 24142
rect 6000 23792 6052 23798
rect 6000 23734 6052 23740
rect 5264 23656 5316 23662
rect 5264 23598 5316 23604
rect 6104 23526 6132 24278
rect 6644 24200 6696 24206
rect 6644 24142 6696 24148
rect 6092 23520 6144 23526
rect 6092 23462 6144 23468
rect 5356 23180 5408 23186
rect 5356 23122 5408 23128
rect 5368 22778 5396 23122
rect 5540 22976 5592 22982
rect 5540 22918 5592 22924
rect 5552 22778 5580 22918
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5356 22772 5408 22778
rect 5356 22714 5408 22720
rect 5540 22772 5592 22778
rect 5540 22714 5592 22720
rect 6000 22432 6052 22438
rect 6000 22374 6052 22380
rect 6012 22098 6040 22374
rect 6104 22234 6132 23462
rect 6460 23248 6512 23254
rect 6460 23190 6512 23196
rect 6472 22438 6500 23190
rect 6656 23118 6684 24142
rect 7012 23520 7064 23526
rect 7012 23462 7064 23468
rect 6644 23112 6696 23118
rect 6644 23054 6696 23060
rect 7024 22642 7052 23462
rect 7484 23322 7512 27520
rect 9600 23866 9628 27520
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 9588 23860 9640 23866
rect 9588 23802 9640 23808
rect 8116 23520 8168 23526
rect 8116 23462 8168 23468
rect 7472 23316 7524 23322
rect 7472 23258 7524 23264
rect 8024 23248 8076 23254
rect 8024 23190 8076 23196
rect 7932 23112 7984 23118
rect 7932 23054 7984 23060
rect 7944 22778 7972 23054
rect 7932 22772 7984 22778
rect 7932 22714 7984 22720
rect 7012 22636 7064 22642
rect 7012 22578 7064 22584
rect 6460 22432 6512 22438
rect 6460 22374 6512 22380
rect 7024 22234 7052 22578
rect 7380 22500 7432 22506
rect 7380 22442 7432 22448
rect 6092 22228 6144 22234
rect 6092 22170 6144 22176
rect 7012 22228 7064 22234
rect 7012 22170 7064 22176
rect 7392 22166 7420 22442
rect 8036 22438 8064 23190
rect 8024 22432 8076 22438
rect 8024 22374 8076 22380
rect 7380 22160 7432 22166
rect 7380 22102 7432 22108
rect 6000 22092 6052 22098
rect 6000 22034 6052 22040
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 6012 21350 6040 22034
rect 7380 22024 7432 22030
rect 7380 21966 7432 21972
rect 7392 21350 7420 21966
rect 5080 21344 5132 21350
rect 5080 21286 5132 21292
rect 6000 21344 6052 21350
rect 6000 21286 6052 21292
rect 7380 21344 7432 21350
rect 7380 21286 7432 21292
rect 4252 13932 4304 13938
rect 4252 13874 4304 13880
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 4080 11762 4108 13262
rect 4264 12889 4292 13874
rect 5092 13530 5120 21286
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6380 16250 6408 16594
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 6092 15564 6144 15570
rect 6092 15506 6144 15512
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6104 15162 6132 15506
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 5080 13524 5132 13530
rect 5080 13466 5132 13472
rect 4250 12880 4306 12889
rect 4250 12815 4306 12824
rect 4988 12844 5040 12850
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4172 11830 4200 12582
rect 4160 11824 4212 11830
rect 4160 11766 4212 11772
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 3896 11206 4016 11234
rect 3790 8936 3846 8945
rect 3790 8871 3846 8880
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3804 8566 3832 8774
rect 3792 8560 3844 8566
rect 3792 8502 3844 8508
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3712 8090 3740 8366
rect 3700 8084 3752 8090
rect 3700 8026 3752 8032
rect 3700 7880 3752 7886
rect 3700 7822 3752 7828
rect 3712 7342 3740 7822
rect 3896 7342 3924 11206
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 3988 9674 4016 9998
rect 3988 9646 4108 9674
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3988 8634 4016 8910
rect 4080 8820 4108 9646
rect 4172 9081 4200 11766
rect 4158 9072 4214 9081
rect 4264 9042 4292 12815
rect 4988 12786 5040 12792
rect 4436 12708 4488 12714
rect 4436 12650 4488 12656
rect 4448 12442 4476 12650
rect 5000 12442 5028 12786
rect 4436 12436 4488 12442
rect 4436 12378 4488 12384
rect 4988 12436 5040 12442
rect 4988 12378 5040 12384
rect 4448 11558 4476 12378
rect 4896 12164 4948 12170
rect 4896 12106 4948 12112
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4632 11626 4660 12038
rect 4908 11762 4936 12106
rect 4896 11756 4948 11762
rect 4896 11698 4948 11704
rect 5000 11626 5028 12378
rect 5276 12238 5304 13670
rect 5368 12986 5396 13806
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5264 12232 5316 12238
rect 5264 12174 5316 12180
rect 4620 11620 4672 11626
rect 4620 11562 4672 11568
rect 4988 11620 5040 11626
rect 4988 11562 5040 11568
rect 4436 11552 4488 11558
rect 4436 11494 4488 11500
rect 4448 10198 4476 11494
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 4540 10810 4568 11154
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4540 10470 4568 10746
rect 4632 10713 4660 11562
rect 5000 11354 5028 11562
rect 4988 11348 5040 11354
rect 4988 11290 5040 11296
rect 5172 11008 5224 11014
rect 5172 10950 5224 10956
rect 4618 10704 4674 10713
rect 4618 10639 4674 10648
rect 4712 10532 4764 10538
rect 4712 10474 4764 10480
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4436 10192 4488 10198
rect 4436 10134 4488 10140
rect 4540 10130 4568 10406
rect 4724 10266 4752 10474
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 4618 10024 4674 10033
rect 4724 9994 4752 10202
rect 4618 9959 4674 9968
rect 4712 9988 4764 9994
rect 4632 9654 4660 9959
rect 4712 9930 4764 9936
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4158 9007 4214 9016
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 4344 8832 4396 8838
rect 4080 8792 4344 8820
rect 4344 8774 4396 8780
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 4356 8090 4384 8774
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4632 8294 4660 8434
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 4436 8016 4488 8022
rect 4436 7958 4488 7964
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 3568 7296 3648 7324
rect 3700 7336 3752 7342
rect 3516 7278 3568 7284
rect 3700 7278 3752 7284
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3528 7041 3556 7278
rect 3514 7032 3570 7041
rect 3712 7002 3740 7278
rect 4172 7274 4200 7890
rect 4448 7546 4476 7958
rect 4632 7954 4660 8230
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4160 7268 4212 7274
rect 4160 7210 4212 7216
rect 4172 7177 4200 7210
rect 4158 7168 4214 7177
rect 4158 7103 4214 7112
rect 3974 7032 4030 7041
rect 3514 6967 3570 6976
rect 3700 6996 3752 7002
rect 3528 6934 3556 6967
rect 3974 6967 4030 6976
rect 4252 6996 4304 7002
rect 3700 6938 3752 6944
rect 3516 6928 3568 6934
rect 3516 6870 3568 6876
rect 3712 6254 3740 6938
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 3700 6248 3752 6254
rect 3700 6190 3752 6196
rect 3516 6180 3568 6186
rect 3516 6122 3568 6128
rect 3422 5944 3478 5953
rect 3528 5914 3556 6122
rect 3896 5914 3924 6802
rect 3988 6254 4016 6967
rect 4252 6938 4304 6944
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3988 6118 4016 6190
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 3422 5879 3478 5888
rect 3516 5908 3568 5914
rect 3436 5846 3464 5879
rect 3516 5850 3568 5856
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3424 5840 3476 5846
rect 3424 5782 3476 5788
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3240 5636 3292 5642
rect 3240 5578 3292 5584
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 3056 5092 3108 5098
rect 3056 5034 3108 5040
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 2976 4282 3004 4626
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 2792 4126 3004 4154
rect 2596 3664 2648 3670
rect 2596 3606 2648 3612
rect 2608 2378 2636 3606
rect 2686 3088 2742 3097
rect 2686 3023 2742 3032
rect 2700 2990 2728 3023
rect 2688 2984 2740 2990
rect 2976 2961 3004 4126
rect 3068 3466 3096 5034
rect 3160 3670 3188 5510
rect 3252 4078 3280 5578
rect 3344 4554 3372 5646
rect 3698 5264 3754 5273
rect 3896 5234 3924 5850
rect 4080 5710 4108 6054
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 3698 5199 3754 5208
rect 3884 5228 3936 5234
rect 3332 4548 3384 4554
rect 3332 4490 3384 4496
rect 3712 4282 3740 5199
rect 3884 5170 3936 5176
rect 3976 5024 4028 5030
rect 3790 4992 3846 5001
rect 3976 4966 4028 4972
rect 3790 4927 3846 4936
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 3608 4072 3660 4078
rect 3608 4014 3660 4020
rect 3620 3738 3648 4014
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3148 3664 3200 3670
rect 3148 3606 3200 3612
rect 3240 3664 3292 3670
rect 3240 3606 3292 3612
rect 3056 3460 3108 3466
rect 3056 3402 3108 3408
rect 3068 3194 3096 3402
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 2688 2926 2740 2932
rect 2962 2952 3018 2961
rect 2780 2916 2832 2922
rect 2962 2887 3018 2896
rect 2780 2858 2832 2864
rect 2792 2650 2820 2858
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 3252 2582 3280 3606
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 3436 3194 3464 3334
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 3436 2922 3464 3130
rect 3620 3126 3648 3674
rect 3804 3534 3832 4927
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 3896 4282 3924 4422
rect 3884 4276 3936 4282
rect 3884 4218 3936 4224
rect 3988 4146 4016 4966
rect 4080 4826 4108 5646
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4264 4282 4292 6938
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4632 6118 4660 6802
rect 4724 6322 4752 9318
rect 5078 9208 5134 9217
rect 5078 9143 5134 9152
rect 5092 9042 5120 9143
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 4802 8936 4858 8945
rect 4802 8871 4858 8880
rect 4712 6316 4764 6322
rect 4712 6258 4764 6264
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4344 5840 4396 5846
rect 4344 5782 4396 5788
rect 4356 5302 4384 5782
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4344 5296 4396 5302
rect 4344 5238 4396 5244
rect 4540 5166 4568 5714
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 4620 5092 4672 5098
rect 4620 5034 4672 5040
rect 4632 4758 4660 5034
rect 4620 4752 4672 4758
rect 4620 4694 4672 4700
rect 4436 4616 4488 4622
rect 4436 4558 4488 4564
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3988 3738 4016 4082
rect 4448 4049 4476 4558
rect 4632 4282 4660 4694
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4528 4208 4580 4214
rect 4528 4150 4580 4156
rect 4434 4040 4490 4049
rect 4264 3998 4434 4026
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 3608 3120 3660 3126
rect 3608 3062 3660 3068
rect 3424 2916 3476 2922
rect 3424 2858 3476 2864
rect 3240 2576 3292 2582
rect 3240 2518 3292 2524
rect 2596 2372 2648 2378
rect 2596 2314 2648 2320
rect 2870 82 2926 480
rect 2516 54 2926 82
rect 3804 82 3832 3470
rect 4264 3466 4292 3998
rect 4434 3975 4490 3984
rect 4252 3460 4304 3466
rect 4252 3402 4304 3408
rect 4436 3460 4488 3466
rect 4436 3402 4488 3408
rect 4344 2916 4396 2922
rect 4344 2858 4396 2864
rect 4356 2689 4384 2858
rect 4342 2680 4398 2689
rect 4342 2615 4398 2624
rect 4448 2310 4476 3402
rect 4540 2650 4568 4150
rect 4816 4146 4844 8871
rect 5080 6928 5132 6934
rect 5080 6870 5132 6876
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4804 4004 4856 4010
rect 4804 3946 4856 3952
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4618 3496 4674 3505
rect 4618 3431 4674 3440
rect 4632 3398 4660 3431
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4632 3058 4660 3334
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4724 2854 4752 3538
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4528 2644 4580 2650
rect 4528 2586 4580 2592
rect 4816 2378 4844 3946
rect 4908 2922 4936 6054
rect 5000 3738 5028 6802
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 5000 3398 5028 3674
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 5000 3058 5028 3334
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 4896 2916 4948 2922
rect 4896 2858 4948 2864
rect 4804 2372 4856 2378
rect 4804 2314 4856 2320
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 4066 82 4122 480
rect 3804 54 4122 82
rect 4908 82 4936 2858
rect 5092 2650 5120 6870
rect 5184 4282 5212 10950
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5276 8498 5304 9114
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5368 8378 5396 12922
rect 5552 12850 5580 13262
rect 5736 13258 5764 13806
rect 5724 13252 5776 13258
rect 5724 13194 5776 13200
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5552 12442 5580 12786
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6012 11762 6040 12242
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 5552 10742 5580 11698
rect 6000 11280 6052 11286
rect 6000 11222 6052 11228
rect 6104 11234 6132 15098
rect 6182 14920 6238 14929
rect 6182 14855 6238 14864
rect 6196 14822 6224 14855
rect 6184 14816 6236 14822
rect 6184 14758 6236 14764
rect 6276 14816 6328 14822
rect 6276 14758 6328 14764
rect 6184 14612 6236 14618
rect 6184 14554 6236 14560
rect 6196 13734 6224 14554
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6196 13462 6224 13670
rect 6184 13456 6236 13462
rect 6184 13398 6236 13404
rect 6196 12986 6224 13398
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 6196 12646 6224 12922
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 6196 12374 6224 12582
rect 6184 12368 6236 12374
rect 6184 12310 6236 12316
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 6012 10810 6040 11222
rect 6104 11206 6224 11234
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 6104 10674 6132 11086
rect 6092 10668 6144 10674
rect 6092 10610 6144 10616
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5552 9636 5580 10134
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5632 9648 5684 9654
rect 5552 9608 5632 9636
rect 5632 9590 5684 9596
rect 5644 9178 5672 9590
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 6104 9178 6132 9318
rect 5632 9172 5684 9178
rect 5552 9132 5632 9160
rect 5552 8634 5580 9132
rect 5632 9114 5684 9120
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 6196 9058 6224 11206
rect 6288 11150 6316 14758
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 6564 13734 6592 14350
rect 6552 13728 6604 13734
rect 6552 13670 6604 13676
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6380 12306 6408 12718
rect 6564 12374 6592 13670
rect 6552 12368 6604 12374
rect 6552 12310 6604 12316
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6380 11558 6408 12242
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6288 10538 6316 11086
rect 6276 10532 6328 10538
rect 6276 10474 6328 10480
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 6104 9030 6224 9058
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6012 8634 6040 8978
rect 6104 8838 6132 9030
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5276 8350 5396 8378
rect 6104 8362 6132 8774
rect 5540 8356 5592 8362
rect 5276 5030 5304 8350
rect 5540 8298 5592 8304
rect 6092 8356 6144 8362
rect 6092 8298 6144 8304
rect 5552 8090 5580 8298
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5356 7268 5408 7274
rect 5356 7210 5408 7216
rect 5368 6254 5396 7210
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5460 6662 5488 7142
rect 6012 6730 6040 7686
rect 6196 7206 6224 7890
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6288 7274 6316 7686
rect 6276 7268 6328 7274
rect 6276 7210 6328 7216
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 6000 6724 6052 6730
rect 6000 6666 6052 6672
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5460 6390 5488 6598
rect 5552 6458 5580 6598
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5552 6236 5580 6394
rect 5632 6248 5684 6254
rect 5552 6208 5632 6236
rect 5368 5574 5396 6190
rect 5552 5642 5580 6208
rect 5632 6190 5684 6196
rect 6012 5914 6040 6666
rect 6090 6352 6146 6361
rect 6090 6287 6146 6296
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 5540 5636 5592 5642
rect 5540 5578 5592 5584
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5170 4176 5226 4185
rect 5170 4111 5226 4120
rect 5184 3194 5212 4111
rect 5276 4078 5304 4966
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5368 2972 5396 5510
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5460 4078 5488 4422
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5552 3466 5580 5578
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5816 5296 5868 5302
rect 5816 5238 5868 5244
rect 5828 4826 5856 5238
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5736 3466 5764 4082
rect 5540 3460 5592 3466
rect 5540 3402 5592 3408
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6012 3194 6040 5510
rect 6104 5302 6132 6287
rect 6196 6202 6224 7142
rect 6380 6458 6408 11494
rect 6748 9586 6776 15438
rect 7116 15366 7144 15982
rect 7104 15360 7156 15366
rect 7104 15302 7156 15308
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 7024 14550 7052 14758
rect 7012 14544 7064 14550
rect 7012 14486 7064 14492
rect 7392 14346 7420 21286
rect 7564 16584 7616 16590
rect 7564 16526 7616 16532
rect 7472 16448 7524 16454
rect 7472 16390 7524 16396
rect 7484 15502 7512 16390
rect 7576 15638 7604 16526
rect 7932 16176 7984 16182
rect 7932 16118 7984 16124
rect 7564 15632 7616 15638
rect 7564 15574 7616 15580
rect 7472 15496 7524 15502
rect 7472 15438 7524 15444
rect 7484 15026 7512 15438
rect 7576 15162 7604 15574
rect 7944 15502 7972 16118
rect 7932 15496 7984 15502
rect 7932 15438 7984 15444
rect 7564 15156 7616 15162
rect 7564 15098 7616 15104
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7944 14414 7972 15438
rect 8024 14884 8076 14890
rect 8024 14826 8076 14832
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 7380 14340 7432 14346
rect 7380 14282 7432 14288
rect 7484 13530 7512 14350
rect 8036 14346 8064 14826
rect 8024 14340 8076 14346
rect 8024 14282 8076 14288
rect 7932 13796 7984 13802
rect 7932 13738 7984 13744
rect 7944 13530 7972 13738
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7932 13524 7984 13530
rect 7932 13466 7984 13472
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7300 12782 7328 13126
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6932 12238 6960 12582
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 6826 9616 6882 9625
rect 6736 9580 6788 9586
rect 6826 9551 6882 9560
rect 6736 9522 6788 9528
rect 6840 9518 6868 9551
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6840 9110 6868 9454
rect 6828 9104 6880 9110
rect 6828 9046 6880 9052
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6748 7342 6776 7482
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6460 6928 6512 6934
rect 6460 6870 6512 6876
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 6196 6174 6316 6202
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6196 5642 6224 6054
rect 6184 5636 6236 5642
rect 6184 5578 6236 5584
rect 6092 5296 6144 5302
rect 6092 5238 6144 5244
rect 6104 4185 6132 5238
rect 6288 5001 6316 6174
rect 6472 5914 6500 6870
rect 6748 6730 6776 7278
rect 7024 7206 7052 7822
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 7024 6798 7052 7142
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 6736 6724 6788 6730
rect 6736 6666 6788 6672
rect 6748 6458 6776 6666
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 6368 5772 6420 5778
rect 6368 5714 6420 5720
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6380 5030 6408 5714
rect 6472 5098 6500 5714
rect 6748 5302 6776 6394
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 6460 5092 6512 5098
rect 6460 5034 6512 5040
rect 6368 5024 6420 5030
rect 6274 4992 6330 5001
rect 6368 4966 6420 4972
rect 6274 4927 6330 4936
rect 6472 4690 6500 5034
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6196 4214 6224 4626
rect 6184 4208 6236 4214
rect 6090 4176 6146 4185
rect 6184 4150 6236 4156
rect 6090 4111 6146 4120
rect 6196 3913 6224 4150
rect 6182 3904 6238 3913
rect 6182 3839 6238 3848
rect 6472 3738 6500 4626
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6656 4078 6684 4558
rect 6748 4214 6776 4762
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 6104 3058 6132 3470
rect 6656 3466 6684 3674
rect 6748 3670 6776 4150
rect 6736 3664 6788 3670
rect 6736 3606 6788 3612
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 6288 3194 6316 3334
rect 6748 3194 6776 3606
rect 6840 3466 6868 5646
rect 6932 5166 6960 6326
rect 7024 6118 7052 6598
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 7116 5574 7144 12106
rect 7300 12102 7328 12718
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7380 11620 7432 11626
rect 7380 11562 7432 11568
rect 7392 11354 7420 11562
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7392 10674 7420 11290
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7196 10192 7248 10198
rect 7196 10134 7248 10140
rect 7208 9722 7236 10134
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7208 9110 7236 9522
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7196 9104 7248 9110
rect 7196 9046 7248 9052
rect 7208 8634 7236 9046
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6932 4486 6960 5102
rect 7024 5030 7052 5170
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 7012 5024 7064 5030
rect 7208 5001 7236 5034
rect 7012 4966 7064 4972
rect 7194 4992 7250 5001
rect 7024 4554 7052 4966
rect 7194 4927 7250 4936
rect 7012 4548 7064 4554
rect 7012 4490 7064 4496
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 5368 2944 5672 2972
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 5172 2576 5224 2582
rect 5356 2576 5408 2582
rect 5224 2536 5356 2564
rect 5172 2518 5224 2524
rect 5356 2518 5408 2524
rect 5644 2446 5672 2944
rect 5906 2952 5962 2961
rect 5906 2887 5962 2896
rect 5920 2650 5948 2887
rect 6932 2650 6960 4422
rect 5908 2644 5960 2650
rect 5908 2586 5960 2592
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 6092 2508 6144 2514
rect 6092 2450 6144 2456
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5170 82 5226 480
rect 4908 54 5226 82
rect 6104 82 6132 2450
rect 6366 82 6422 480
rect 6104 54 6422 82
rect 7300 82 7328 9318
rect 7392 8974 7420 9862
rect 7484 9382 7512 11698
rect 7668 9926 7696 12786
rect 7760 11762 7788 13126
rect 8024 12708 8076 12714
rect 8024 12650 8076 12656
rect 8036 12288 8064 12650
rect 8128 12442 8156 23462
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 11716 23322 11744 27520
rect 13924 23662 13952 27520
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 13912 23656 13964 23662
rect 13912 23598 13964 23604
rect 13820 23520 13872 23526
rect 13820 23462 13872 23468
rect 11704 23316 11756 23322
rect 11704 23258 11756 23264
rect 11060 23180 11112 23186
rect 11060 23122 11112 23128
rect 8208 23112 8260 23118
rect 8208 23054 8260 23060
rect 8220 22642 8248 23054
rect 8208 22636 8260 22642
rect 8208 22578 8260 22584
rect 10876 22568 10928 22574
rect 10966 22536 11022 22545
rect 10928 22516 10966 22522
rect 10876 22510 10966 22516
rect 10888 22494 10966 22510
rect 10966 22471 11022 22480
rect 8208 22432 8260 22438
rect 8208 22374 8260 22380
rect 10968 22432 11020 22438
rect 11072 22420 11100 23122
rect 11020 22392 11100 22420
rect 10968 22374 11020 22380
rect 8220 22098 8248 22374
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10980 22234 11008 22374
rect 10968 22228 11020 22234
rect 10968 22170 11020 22176
rect 8208 22092 8260 22098
rect 8208 22034 8260 22040
rect 11796 22092 11848 22098
rect 11796 22034 11848 22040
rect 11808 21690 11836 22034
rect 12532 21888 12584 21894
rect 12532 21830 12584 21836
rect 12900 21888 12952 21894
rect 12900 21830 12952 21836
rect 11796 21684 11848 21690
rect 11796 21626 11848 21632
rect 11428 21480 11480 21486
rect 11428 21422 11480 21428
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 11336 20936 11388 20942
rect 11336 20878 11388 20884
rect 11348 20602 11376 20878
rect 11336 20596 11388 20602
rect 11336 20538 11388 20544
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8220 15978 8248 16594
rect 8484 16108 8536 16114
rect 8484 16050 8536 16056
rect 8208 15972 8260 15978
rect 8208 15914 8260 15920
rect 8220 13530 8248 15914
rect 8496 15366 8524 16050
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 8312 15094 8340 15302
rect 8300 15088 8352 15094
rect 8300 15030 8352 15036
rect 8312 14414 8340 15030
rect 8392 14544 8444 14550
rect 8496 14521 8524 15302
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 8392 14486 8444 14492
rect 8482 14512 8538 14521
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 8404 14074 8432 14486
rect 8482 14447 8538 14456
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 8588 13326 8616 14554
rect 9140 14550 9168 14894
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 9128 14544 9180 14550
rect 9128 14486 9180 14492
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 10140 14476 10192 14482
rect 10140 14418 10192 14424
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8772 13530 8800 13874
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 9310 13832 9366 13841
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 9048 13326 9076 13670
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 8588 12986 8616 13262
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8758 12880 8814 12889
rect 8758 12815 8814 12824
rect 8772 12782 8800 12815
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8116 12436 8168 12442
rect 8116 12378 8168 12384
rect 8116 12300 8168 12306
rect 8036 12260 8116 12288
rect 8116 12242 8168 12248
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7760 10198 7788 11698
rect 7840 11280 7892 11286
rect 7840 11222 7892 11228
rect 7852 10810 7880 11222
rect 7840 10804 7892 10810
rect 7840 10746 7892 10752
rect 7748 10192 7800 10198
rect 7748 10134 7800 10140
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7392 8498 7420 8910
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7472 8492 7524 8498
rect 7524 8452 7604 8480
rect 7472 8434 7524 8440
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 7484 7750 7512 8298
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7484 7274 7512 7686
rect 7472 7268 7524 7274
rect 7472 7210 7524 7216
rect 7576 6798 7604 8452
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7576 6458 7604 6734
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7668 6338 7696 9862
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7760 8566 7788 8910
rect 7944 8566 7972 12038
rect 8128 11898 8156 12242
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 8024 11620 8076 11626
rect 8024 11562 8076 11568
rect 8036 10198 8064 11562
rect 8312 11558 8340 12242
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8208 10532 8260 10538
rect 8208 10474 8260 10480
rect 8024 10192 8076 10198
rect 8024 10134 8076 10140
rect 8220 9450 8248 10474
rect 8208 9444 8260 9450
rect 8208 9386 8260 9392
rect 8312 8906 8340 11494
rect 8404 10674 8432 12174
rect 8864 11286 8892 12174
rect 9048 12170 9076 13262
rect 9232 13190 9260 13806
rect 9692 13814 9720 14418
rect 9310 13767 9366 13776
rect 9508 13802 9720 13814
rect 9508 13796 9732 13802
rect 9508 13786 9680 13796
rect 9324 13734 9352 13767
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 9508 12918 9536 13786
rect 9680 13738 9732 13744
rect 10152 13394 10180 14418
rect 11440 14074 11468 21422
rect 11520 21412 11572 21418
rect 11520 21354 11572 21360
rect 11532 21078 11560 21354
rect 11704 21344 11756 21350
rect 11704 21286 11756 21292
rect 11520 21072 11572 21078
rect 11520 21014 11572 21020
rect 11532 20602 11560 21014
rect 11520 20596 11572 20602
rect 11520 20538 11572 20544
rect 11518 18184 11574 18193
rect 11518 18119 11574 18128
rect 11532 17882 11560 18119
rect 11520 17876 11572 17882
rect 11520 17818 11572 17824
rect 11612 17740 11664 17746
rect 11612 17682 11664 17688
rect 11624 16998 11652 17682
rect 11612 16992 11664 16998
rect 11612 16934 11664 16940
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 9496 12912 9548 12918
rect 9496 12854 9548 12860
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9128 12436 9180 12442
rect 9128 12378 9180 12384
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 9140 11762 9168 12378
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 9232 11626 9260 11834
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 9232 11354 9260 11562
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 8852 11280 8904 11286
rect 8852 11222 8904 11228
rect 9232 10810 9260 11290
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 8404 10266 8432 10610
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8576 10124 8628 10130
rect 8576 10066 8628 10072
rect 8588 9654 8616 10066
rect 9416 9654 9444 12718
rect 9508 12306 9536 12854
rect 9692 12850 9720 13330
rect 10704 13190 10732 13806
rect 10508 13184 10560 13190
rect 10508 13126 10560 13132
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10520 12850 10548 13126
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 10152 12306 10180 12718
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 9508 11354 9536 12242
rect 9772 11620 9824 11626
rect 9772 11562 9824 11568
rect 9496 11348 9548 11354
rect 9496 11290 9548 11296
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 9404 9648 9456 9654
rect 9404 9590 9456 9596
rect 8588 9042 8616 9590
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 7748 8560 7800 8566
rect 7748 8502 7800 8508
rect 7932 8560 7984 8566
rect 7932 8502 7984 8508
rect 8312 8022 8340 8842
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7760 6866 7788 7890
rect 8404 7818 8432 8774
rect 8588 8634 8616 8978
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8666 8392 8722 8401
rect 8666 8327 8722 8336
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 7852 7546 7880 7686
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 8128 6866 8156 7754
rect 8576 7744 8628 7750
rect 8576 7686 8628 7692
rect 8588 7342 8616 7686
rect 8680 7546 8708 8327
rect 8772 7886 8800 8774
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8484 7268 8536 7274
rect 8484 7210 8536 7216
rect 7748 6860 7800 6866
rect 7748 6802 7800 6808
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 7760 6662 7788 6802
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7576 6310 7696 6338
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 7392 4826 7420 5102
rect 7576 4826 7604 6310
rect 7760 6186 7788 6598
rect 8128 6390 8156 6802
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8312 6458 8340 6598
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8116 6384 8168 6390
rect 8312 6361 8340 6394
rect 8496 6390 8524 7210
rect 8772 6934 8800 7278
rect 8864 7002 8892 8434
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 8956 7478 8984 7686
rect 8944 7472 8996 7478
rect 8944 7414 8996 7420
rect 9048 7410 9076 7686
rect 9140 7546 9168 8910
rect 9508 7857 9536 11290
rect 9784 11150 9812 11562
rect 10152 11558 10180 12242
rect 10980 11830 11008 13874
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11060 12708 11112 12714
rect 11060 12650 11112 12656
rect 11072 12442 11100 12650
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 10968 11824 11020 11830
rect 10968 11766 11020 11772
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10796 11626 10824 11698
rect 10784 11620 10836 11626
rect 10784 11562 10836 11568
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9784 9654 9812 10406
rect 10060 10266 10088 10542
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9772 9648 9824 9654
rect 9772 9590 9824 9596
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9494 7848 9550 7857
rect 9494 7783 9550 7792
rect 9692 7698 9720 8366
rect 9784 8362 9812 9590
rect 9864 9512 9916 9518
rect 9864 9454 9916 9460
rect 9876 9042 9904 9454
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 9876 8634 9904 8978
rect 9968 8906 9996 10066
rect 9956 8900 10008 8906
rect 9956 8842 10008 8848
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9772 8356 9824 8362
rect 9772 8298 9824 8304
rect 10048 7948 10100 7954
rect 10048 7890 10100 7896
rect 9864 7744 9916 7750
rect 9692 7670 9812 7698
rect 9864 7686 9916 7692
rect 9784 7546 9812 7670
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9140 7206 9168 7482
rect 9312 7472 9364 7478
rect 9312 7414 9364 7420
rect 9220 7268 9272 7274
rect 9220 7210 9272 7216
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 8852 6996 8904 7002
rect 8852 6938 8904 6944
rect 8944 6996 8996 7002
rect 8944 6938 8996 6944
rect 8760 6928 8812 6934
rect 8760 6870 8812 6876
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8484 6384 8536 6390
rect 8116 6326 8168 6332
rect 8298 6352 8354 6361
rect 7748 6180 7800 6186
rect 7748 6122 7800 6128
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 7760 5778 7788 6122
rect 8036 5914 8064 6122
rect 8128 6118 8156 6326
rect 8484 6326 8536 6332
rect 8298 6287 8354 6296
rect 8588 6186 8616 6598
rect 8576 6180 8628 6186
rect 8576 6122 8628 6128
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 7760 5574 7788 5714
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7760 4826 7788 5510
rect 7944 5302 7972 5714
rect 7932 5296 7984 5302
rect 7932 5238 7984 5244
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7944 4758 7972 5238
rect 8036 5166 8064 5850
rect 8128 5778 8156 6054
rect 8220 5846 8248 6054
rect 8772 5914 8800 6122
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8116 5568 8168 5574
rect 8220 5545 8248 5646
rect 8484 5568 8536 5574
rect 8116 5510 8168 5516
rect 8206 5536 8262 5545
rect 8128 5302 8156 5510
rect 8484 5510 8536 5516
rect 8206 5471 8262 5480
rect 8116 5296 8168 5302
rect 8116 5238 8168 5244
rect 8220 5234 8248 5471
rect 8496 5409 8524 5510
rect 8482 5400 8538 5409
rect 8482 5335 8538 5344
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 7656 4752 7708 4758
rect 7656 4694 7708 4700
rect 7932 4752 7984 4758
rect 7932 4694 7984 4700
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 7378 4312 7434 4321
rect 7378 4247 7434 4256
rect 7392 4214 7420 4247
rect 7380 4208 7432 4214
rect 7380 4150 7432 4156
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7392 3097 7420 3878
rect 7576 3369 7604 4558
rect 7668 4010 7696 4694
rect 7656 4004 7708 4010
rect 7656 3946 7708 3952
rect 7944 3738 7972 4694
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8128 4185 8156 4218
rect 8114 4176 8170 4185
rect 8220 4146 8248 4218
rect 8114 4111 8170 4120
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 7562 3360 7618 3369
rect 7562 3295 7618 3304
rect 7378 3088 7434 3097
rect 7378 3023 7434 3032
rect 7392 2922 7420 3023
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 7380 2916 7432 2922
rect 7380 2858 7432 2864
rect 8128 2650 8156 2926
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 8220 2582 8248 3470
rect 8312 3194 8340 4626
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 8680 4214 8708 4490
rect 8668 4208 8720 4214
rect 8668 4150 8720 4156
rect 8772 3398 8800 4966
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8956 3058 8984 6938
rect 9140 6458 9168 7142
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 9140 6361 9168 6394
rect 9126 6352 9182 6361
rect 9126 6287 9182 6296
rect 9140 5710 9168 6287
rect 9232 6168 9260 7210
rect 9324 6662 9352 7414
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9416 7206 9444 7346
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 9404 7200 9456 7206
rect 9600 7177 9628 7210
rect 9404 7142 9456 7148
rect 9586 7168 9642 7177
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9324 6458 9352 6598
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9416 6322 9444 7142
rect 9586 7103 9642 7112
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9508 6662 9536 6802
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 9600 6254 9628 7103
rect 9678 7032 9734 7041
rect 9678 6967 9734 6976
rect 9692 6866 9720 6967
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9588 6248 9640 6254
rect 9508 6208 9588 6236
rect 9312 6180 9364 6186
rect 9232 6140 9312 6168
rect 9312 6122 9364 6128
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9324 5370 9352 6122
rect 9508 5846 9536 6208
rect 9588 6190 9640 6196
rect 9496 5840 9548 5846
rect 9496 5782 9548 5788
rect 9692 5778 9720 6326
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9784 5778 9812 6190
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 9324 5273 9352 5306
rect 9310 5264 9366 5273
rect 9310 5199 9366 5208
rect 9692 5166 9720 5578
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9784 5030 9812 5714
rect 9876 5681 9904 7686
rect 10060 6798 10088 7890
rect 10152 7546 10180 11494
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10980 11286 11008 11766
rect 11072 11558 11100 12378
rect 11256 12374 11284 13262
rect 11624 12986 11652 16934
rect 11716 13814 11744 21286
rect 11808 20942 11836 21626
rect 12544 21554 12572 21830
rect 12532 21548 12584 21554
rect 12532 21490 12584 21496
rect 11796 20936 11848 20942
rect 11796 20878 11848 20884
rect 12544 20874 12572 21490
rect 12912 21078 12940 21830
rect 13832 21434 13860 23462
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15304 22438 15332 23122
rect 14004 22432 14056 22438
rect 14004 22374 14056 22380
rect 15292 22432 15344 22438
rect 15292 22374 15344 22380
rect 13912 22092 13964 22098
rect 13912 22034 13964 22040
rect 13924 21690 13952 22034
rect 13912 21684 13964 21690
rect 13912 21626 13964 21632
rect 13740 21406 13860 21434
rect 12900 21072 12952 21078
rect 12900 21014 12952 21020
rect 13084 21072 13136 21078
rect 13084 21014 13136 21020
rect 12532 20868 12584 20874
rect 12532 20810 12584 20816
rect 12716 20800 12768 20806
rect 12716 20742 12768 20748
rect 12728 20466 12756 20742
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12728 20369 12756 20402
rect 12714 20360 12770 20369
rect 12714 20295 12770 20304
rect 12164 20256 12216 20262
rect 12164 20198 12216 20204
rect 12176 19922 12204 20198
rect 12912 20058 12940 21014
rect 12992 20868 13044 20874
rect 12992 20810 13044 20816
rect 13004 20466 13032 20810
rect 12992 20460 13044 20466
rect 12992 20402 13044 20408
rect 13096 20262 13124 21014
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 13096 19990 13124 20198
rect 13084 19984 13136 19990
rect 13084 19926 13136 19932
rect 12164 19916 12216 19922
rect 12164 19858 12216 19864
rect 12176 19174 12204 19858
rect 12164 19168 12216 19174
rect 12164 19110 12216 19116
rect 11716 13786 11836 13814
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11716 12918 11744 13466
rect 11704 12912 11756 12918
rect 11704 12854 11756 12860
rect 11244 12368 11296 12374
rect 11244 12310 11296 12316
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11624 11898 11652 12242
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 11348 11354 11376 11630
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 10968 11280 11020 11286
rect 10968 11222 11020 11228
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 10336 10810 10364 11086
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 11348 10742 11376 11290
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10888 9382 10916 9998
rect 11624 9722 11652 10066
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10704 8430 10732 8774
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10704 8022 10732 8366
rect 10888 8090 10916 9318
rect 11164 9110 11192 9318
rect 11060 9104 11112 9110
rect 11060 9046 11112 9052
rect 11152 9104 11204 9110
rect 11152 9046 11204 9052
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 10980 8294 11008 8910
rect 11072 8634 11100 9046
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10692 8016 10744 8022
rect 10692 7958 10744 7964
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10704 6644 10732 7346
rect 10784 6656 10836 6662
rect 10704 6616 10784 6644
rect 10704 6458 10732 6616
rect 10784 6598 10836 6604
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 9862 5672 9918 5681
rect 9862 5607 9918 5616
rect 9968 5574 9996 6394
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10060 5710 10088 6258
rect 10704 6254 10732 6394
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9968 4554 9996 5510
rect 10060 4826 10088 5646
rect 10692 5636 10744 5642
rect 10692 5578 10744 5584
rect 10876 5636 10928 5642
rect 10876 5578 10928 5584
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 9956 4548 10008 4554
rect 9956 4490 10008 4496
rect 10152 4185 10180 5510
rect 10704 5030 10732 5578
rect 10888 5166 10916 5578
rect 10876 5160 10928 5166
rect 10876 5102 10928 5108
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10416 4752 10468 4758
rect 10416 4694 10468 4700
rect 10428 4321 10456 4694
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10414 4312 10470 4321
rect 10520 4282 10548 4558
rect 10414 4247 10470 4256
rect 10508 4276 10560 4282
rect 10138 4176 10194 4185
rect 10138 4111 10194 4120
rect 9680 4072 9732 4078
rect 9402 4040 9458 4049
rect 9128 4004 9180 4010
rect 9680 4014 9732 4020
rect 9862 4040 9918 4049
rect 9402 3975 9458 3984
rect 9128 3946 9180 3952
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 8852 2916 8904 2922
rect 8852 2858 8904 2864
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 8208 2576 8260 2582
rect 8208 2518 8260 2524
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 7656 2508 7708 2514
rect 7656 2450 7708 2456
rect 7668 2310 7696 2450
rect 8312 2446 8340 2518
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 7668 1562 7696 2246
rect 7656 1556 7708 1562
rect 7656 1498 7708 1504
rect 7562 82 7618 480
rect 7300 54 7618 82
rect 8404 82 8432 2790
rect 8864 2514 8892 2858
rect 9140 2854 9168 3946
rect 9416 3942 9444 3975
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9324 3738 9352 3878
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9586 3496 9642 3505
rect 9586 3431 9642 3440
rect 9600 3194 9628 3431
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 9494 2680 9550 2689
rect 9494 2615 9550 2624
rect 9508 2582 9536 2615
rect 9496 2576 9548 2582
rect 9496 2518 9548 2524
rect 9692 2514 9720 4014
rect 9862 3975 9918 3984
rect 9876 3602 9904 3975
rect 9864 3596 9916 3602
rect 10152 3584 10180 4111
rect 10428 4078 10456 4247
rect 10508 4218 10560 4224
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10704 3670 10732 4014
rect 10888 3738 10916 4218
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10692 3664 10744 3670
rect 10692 3606 10744 3612
rect 10324 3596 10376 3602
rect 10152 3556 10324 3584
rect 9864 3538 9916 3544
rect 10324 3538 10376 3544
rect 9876 3194 9904 3538
rect 10336 3194 10364 3538
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 10692 3120 10744 3126
rect 10692 3062 10744 3068
rect 10704 2922 10732 3062
rect 10876 3052 10928 3058
rect 10980 3040 11008 8230
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11348 6866 11376 7142
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 11164 5545 11192 6190
rect 11256 6186 11284 6802
rect 11244 6180 11296 6186
rect 11244 6122 11296 6128
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11150 5536 11206 5545
rect 11150 5471 11206 5480
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 11072 4049 11100 5170
rect 11256 5166 11284 5850
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 11336 5092 11388 5098
rect 11336 5034 11388 5040
rect 11520 5092 11572 5098
rect 11520 5034 11572 5040
rect 11348 4486 11376 5034
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11440 4214 11468 4762
rect 11428 4208 11480 4214
rect 11428 4150 11480 4156
rect 11058 4040 11114 4049
rect 11058 3975 11114 3984
rect 10928 3012 11008 3040
rect 10876 2994 10928 3000
rect 10692 2916 10744 2922
rect 10692 2858 10744 2864
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10704 2650 10732 2858
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 10888 2582 10916 2994
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 11164 2650 11192 2790
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 10876 2576 10928 2582
rect 10876 2518 10928 2524
rect 11440 2514 11468 4150
rect 11532 3534 11560 5034
rect 11624 4758 11652 5850
rect 11808 5370 11836 13786
rect 12176 13530 12204 19110
rect 13740 13938 13768 21406
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13740 12986 13768 13330
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13360 12640 13412 12646
rect 13360 12582 13412 12588
rect 13084 12232 13136 12238
rect 13084 12174 13136 12180
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11900 10810 11928 11154
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11900 9178 11928 10746
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 12176 8838 12204 9454
rect 12636 9110 12664 11086
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12728 10266 12756 10610
rect 12820 10538 12848 11086
rect 13096 10674 13124 12174
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 12808 10532 12860 10538
rect 12808 10474 12860 10480
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12716 9444 12768 9450
rect 12716 9386 12768 9392
rect 12256 9104 12308 9110
rect 12256 9046 12308 9052
rect 12624 9104 12676 9110
rect 12624 9046 12676 9052
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12176 8090 12204 8774
rect 12268 8634 12296 9046
rect 12636 8634 12664 9046
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12728 8294 12756 9386
rect 13188 9110 13216 11494
rect 13372 10538 13400 12582
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13648 10810 13676 11154
rect 13636 10804 13688 10810
rect 13636 10746 13688 10752
rect 13360 10532 13412 10538
rect 13360 10474 13412 10480
rect 13372 10198 13400 10474
rect 13648 10266 13676 10746
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13360 10192 13412 10198
rect 13360 10134 13412 10140
rect 13648 9722 13676 10202
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13636 9716 13688 9722
rect 13636 9658 13688 9664
rect 13740 9654 13768 9930
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13636 9444 13688 9450
rect 13636 9386 13688 9392
rect 13176 9104 13228 9110
rect 13176 9046 13228 9052
rect 13648 8906 13676 9386
rect 13740 9178 13768 9590
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 13924 9382 13952 9454
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13636 8900 13688 8906
rect 13636 8842 13688 8848
rect 13648 8430 13676 8842
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 11980 7812 12032 7818
rect 11980 7754 12032 7760
rect 11992 7546 12020 7754
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 11992 5710 12020 7482
rect 12360 7342 12388 7890
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12728 6934 12756 8230
rect 13648 7954 13676 8366
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13648 7546 13676 7890
rect 13924 7750 13952 9318
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 13452 7472 13504 7478
rect 13452 7414 13504 7420
rect 13464 7274 13492 7414
rect 13360 7268 13412 7274
rect 13360 7210 13412 7216
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 12716 6928 12768 6934
rect 12716 6870 12768 6876
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 12268 5846 12296 6734
rect 12728 6458 12756 6870
rect 13372 6712 13400 7210
rect 13464 7002 13492 7210
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13452 6724 13504 6730
rect 13372 6684 13452 6712
rect 13452 6666 13504 6672
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12728 6118 12756 6394
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 12728 5914 12756 6054
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12256 5840 12308 5846
rect 12256 5782 12308 5788
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11992 5302 12020 5646
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 11980 5296 12032 5302
rect 11980 5238 12032 5244
rect 11992 5098 12020 5238
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 11980 5092 12032 5098
rect 11980 5034 12032 5040
rect 11612 4752 11664 4758
rect 11612 4694 11664 4700
rect 11624 3670 11652 4694
rect 12348 4684 12400 4690
rect 12348 4626 12400 4632
rect 11888 4548 11940 4554
rect 11888 4490 11940 4496
rect 11900 4146 11928 4490
rect 11978 4176 12034 4185
rect 11888 4140 11940 4146
rect 11978 4111 12034 4120
rect 11888 4082 11940 4088
rect 11992 4078 12020 4111
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 12360 3942 12388 4626
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 11624 3194 11652 3606
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 11992 2650 12020 3470
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 8852 2508 8904 2514
rect 8852 2450 8904 2456
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 11428 2508 11480 2514
rect 11428 2450 11480 2456
rect 9770 1864 9826 1873
rect 9770 1799 9826 1808
rect 8666 82 8722 480
rect 8404 54 8722 82
rect 9784 82 9812 1799
rect 10692 1556 10744 1562
rect 10692 1498 10744 1504
rect 9862 82 9918 480
rect 9784 54 9918 82
rect 10704 82 10732 1498
rect 11058 82 11114 480
rect 10704 54 11114 82
rect 570 0 626 54
rect 1674 0 1730 54
rect 2870 0 2926 54
rect 4066 0 4122 54
rect 5170 0 5226 54
rect 6366 0 6422 54
rect 7562 0 7618 54
rect 8666 0 8722 54
rect 9862 0 9918 54
rect 11058 0 11114 54
rect 12162 82 12218 480
rect 12452 82 12480 5102
rect 12544 4146 12572 5306
rect 13372 5273 13400 6054
rect 13358 5264 13414 5273
rect 13358 5199 13414 5208
rect 13464 5148 13492 6666
rect 13636 5704 13688 5710
rect 13636 5646 13688 5652
rect 13372 5120 13492 5148
rect 12900 4752 12952 4758
rect 12900 4694 12952 4700
rect 12624 4548 12676 4554
rect 12624 4490 12676 4496
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12636 4010 12664 4490
rect 12624 4004 12676 4010
rect 12624 3946 12676 3952
rect 12532 3460 12584 3466
rect 12532 3402 12584 3408
rect 12544 2922 12572 3402
rect 12808 3392 12860 3398
rect 12912 3369 12940 4694
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13280 4282 13308 4626
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 12808 3334 12860 3340
rect 12898 3360 12954 3369
rect 12532 2916 12584 2922
rect 12532 2858 12584 2864
rect 12544 2825 12572 2858
rect 12530 2816 12586 2825
rect 12530 2751 12586 2760
rect 12820 2689 12848 3334
rect 12898 3295 12954 3304
rect 12806 2680 12862 2689
rect 12806 2615 12862 2624
rect 12820 2582 12848 2615
rect 12808 2576 12860 2582
rect 12808 2518 12860 2524
rect 12820 2310 12848 2518
rect 12808 2304 12860 2310
rect 12808 2246 12860 2252
rect 12912 1737 12940 3295
rect 13372 3058 13400 5120
rect 13648 4826 13676 5646
rect 13832 5642 13860 7482
rect 13924 5778 13952 7686
rect 14016 7410 14044 22374
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15764 21690 15792 27526
rect 16026 27520 16082 27526
rect 18234 27520 18290 28000
rect 20350 27520 20406 28000
rect 22466 27520 22522 28000
rect 24674 27520 24730 28000
rect 26790 27554 26846 28000
rect 26436 27526 26846 27554
rect 18248 23866 18276 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20364 23866 20392 27520
rect 22480 23866 22508 27520
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 18236 23860 18288 23866
rect 18236 23802 18288 23808
rect 20352 23860 20404 23866
rect 20352 23802 20404 23808
rect 22468 23860 22520 23866
rect 22468 23802 22520 23808
rect 24688 23798 24716 27520
rect 25134 26208 25190 26217
rect 25134 26143 25190 26152
rect 25148 23866 25176 26143
rect 25136 23860 25188 23866
rect 25136 23802 25188 23808
rect 24676 23792 24728 23798
rect 24676 23734 24728 23740
rect 25148 23662 25176 23802
rect 16028 23656 16080 23662
rect 16028 23598 16080 23604
rect 18328 23656 18380 23662
rect 18328 23598 18380 23604
rect 25136 23656 25188 23662
rect 25136 23598 25188 23604
rect 16040 23322 16068 23598
rect 16028 23316 16080 23322
rect 16028 23258 16080 23264
rect 18340 22545 18368 23598
rect 19340 23588 19392 23594
rect 19340 23530 19392 23536
rect 18326 22536 18382 22545
rect 18326 22471 18382 22480
rect 15752 21684 15804 21690
rect 15752 21626 15804 21632
rect 15660 20800 15712 20806
rect 15660 20742 15712 20748
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15672 20369 15700 20742
rect 15658 20360 15714 20369
rect 15658 20295 15714 20304
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 14186 15600 14242 15609
rect 14186 15535 14242 15544
rect 14200 15162 14228 15535
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14188 15156 14240 15162
rect 14188 15098 14240 15104
rect 15672 14521 15700 15846
rect 18420 15700 18472 15706
rect 18420 15642 18472 15648
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 15658 14512 15714 14521
rect 15658 14447 15714 14456
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 14188 13728 14240 13734
rect 14188 13670 14240 13676
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14108 8498 14136 12718
rect 14200 11665 14228 13670
rect 14476 13462 14504 13670
rect 14752 13530 14780 13874
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14464 13456 14516 13462
rect 14464 13398 14516 13404
rect 15476 13456 15528 13462
rect 15476 13398 15528 13404
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15488 12986 15516 13398
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15764 12986 15792 13262
rect 15856 12986 15884 14758
rect 15936 13796 15988 13802
rect 15936 13738 15988 13744
rect 15948 13258 15976 13738
rect 15936 13252 15988 13258
rect 15936 13194 15988 13200
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 14372 12708 14424 12714
rect 14372 12650 14424 12656
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 14292 11898 14320 12242
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14186 11656 14242 11665
rect 14186 11591 14242 11600
rect 14292 11558 14320 11834
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14384 10810 14412 12650
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14464 11552 14516 11558
rect 14464 11494 14516 11500
rect 14476 11286 14504 11494
rect 14464 11280 14516 11286
rect 14464 11222 14516 11228
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14384 10538 14412 10746
rect 14372 10532 14424 10538
rect 14372 10474 14424 10480
rect 14476 10266 14504 11222
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14752 9926 14780 10610
rect 15304 10577 15332 12038
rect 15396 11898 15424 12242
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15396 11558 15424 11834
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15396 10810 15424 11494
rect 15580 11286 15608 12038
rect 15568 11280 15620 11286
rect 15568 11222 15620 11228
rect 15580 10810 15608 11222
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15290 10568 15346 10577
rect 15290 10503 15346 10512
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15672 10266 15700 10474
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14752 9586 14780 9862
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15672 9722 15700 10202
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14648 9512 14700 9518
rect 14568 9472 14648 9500
rect 14568 8838 14596 9472
rect 14648 9454 14700 9460
rect 15672 9110 15700 9658
rect 15856 9382 15884 9998
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 15856 9178 15884 9318
rect 15844 9172 15896 9178
rect 15844 9114 15896 9120
rect 15476 9104 15528 9110
rect 15476 9046 15528 9052
rect 15660 9104 15712 9110
rect 15660 9046 15712 9052
rect 14648 8968 14700 8974
rect 14648 8910 14700 8916
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14200 8401 14228 8774
rect 14660 8634 14688 8910
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14186 8392 14242 8401
rect 14186 8327 14242 8336
rect 14660 8022 14688 8570
rect 15384 8424 15436 8430
rect 15384 8366 15436 8372
rect 14648 8016 14700 8022
rect 14648 7958 14700 7964
rect 15396 7954 15424 8366
rect 15488 8294 15516 9046
rect 15948 8566 15976 13194
rect 16028 12776 16080 12782
rect 16028 12718 16080 12724
rect 16040 11762 16068 12718
rect 17224 11824 17276 11830
rect 17224 11766 17276 11772
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 16040 11286 16068 11698
rect 16028 11280 16080 11286
rect 16028 11222 16080 11228
rect 16948 11280 17000 11286
rect 16948 11222 17000 11228
rect 16488 11008 16540 11014
rect 16488 10950 16540 10956
rect 16500 10674 16528 10950
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 16500 10266 16528 10610
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16960 10198 16988 11222
rect 17236 11150 17264 11766
rect 17408 11280 17460 11286
rect 17408 11222 17460 11228
rect 17224 11144 17276 11150
rect 17224 11086 17276 11092
rect 17236 10674 17264 11086
rect 17224 10668 17276 10674
rect 17224 10610 17276 10616
rect 17420 10470 17448 11222
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 16948 10192 17000 10198
rect 16948 10134 17000 10140
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 16500 9178 16528 9454
rect 17328 9382 17356 10066
rect 17420 9994 17448 10406
rect 18432 10198 18460 15642
rect 19352 13841 19380 23530
rect 19432 23520 19484 23526
rect 19432 23462 19484 23468
rect 22744 23520 22796 23526
rect 22744 23462 22796 23468
rect 24766 23488 24822 23497
rect 19444 15706 19472 23462
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19432 15700 19484 15706
rect 19432 15642 19484 15648
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 22008 14272 22060 14278
rect 22008 14214 22060 14220
rect 19338 13832 19394 13841
rect 19338 13767 19394 13776
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 22020 13326 22048 14214
rect 22008 13320 22060 13326
rect 22008 13262 22060 13268
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 18604 11552 18656 11558
rect 18604 11494 18656 11500
rect 18616 10713 18644 11494
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 22756 11354 22784 23462
rect 24766 23423 24822 23432
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24674 21040 24730 21049
rect 24674 20975 24676 20984
rect 24728 20975 24730 20984
rect 24676 20946 24728 20952
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24688 20602 24716 20946
rect 24676 20596 24728 20602
rect 24676 20538 24728 20544
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24780 18714 24808 23423
rect 24688 18686 24808 18714
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24216 17740 24268 17746
rect 24216 17682 24268 17688
rect 24228 16998 24256 17682
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24216 16992 24268 16998
rect 24216 16934 24268 16940
rect 24032 12300 24084 12306
rect 24032 12242 24084 12248
rect 24044 11626 24072 12242
rect 24122 11656 24178 11665
rect 24032 11620 24084 11626
rect 24122 11591 24178 11600
rect 24032 11562 24084 11568
rect 22744 11348 22796 11354
rect 22744 11290 22796 11296
rect 18602 10704 18658 10713
rect 18602 10639 18658 10648
rect 24044 10577 24072 11562
rect 24136 10606 24164 11591
rect 24124 10600 24176 10606
rect 24030 10568 24086 10577
rect 24124 10542 24176 10548
rect 24030 10503 24086 10512
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 24228 10266 24256 16934
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24492 15020 24544 15026
rect 24492 14962 24544 14968
rect 24504 14929 24532 14962
rect 24490 14920 24546 14929
rect 24490 14855 24546 14864
rect 24688 14482 24716 18686
rect 24766 18592 24822 18601
rect 24766 18527 24822 18536
rect 24780 17882 24808 18527
rect 24768 17876 24820 17882
rect 24768 17818 24820 17824
rect 26436 16250 26464 27526
rect 26790 27520 26846 27526
rect 26424 16244 26476 16250
rect 26424 16186 26476 16192
rect 24766 16008 24822 16017
rect 24766 15943 24822 15952
rect 24780 15162 24808 15943
rect 24768 15156 24820 15162
rect 24768 15098 24820 15104
rect 24676 14476 24728 14482
rect 24676 14418 24728 14424
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24688 14074 24716 14418
rect 24676 14068 24728 14074
rect 24676 14010 24728 14016
rect 24766 13696 24822 13705
rect 24766 13631 24822 13640
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24780 12442 24808 13631
rect 24768 12436 24820 12442
rect 24768 12378 24820 12384
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24768 11552 24820 11558
rect 24768 11494 24820 11500
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24216 10260 24268 10266
rect 24216 10202 24268 10208
rect 18420 10192 18472 10198
rect 18420 10134 18472 10140
rect 18604 10192 18656 10198
rect 18604 10134 18656 10140
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 18432 9722 18460 10134
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 17132 9036 17184 9042
rect 17132 8978 17184 8984
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 15936 8560 15988 8566
rect 15936 8502 15988 8508
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 15844 8356 15896 8362
rect 15844 8298 15896 8304
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 15488 8022 15516 8230
rect 15476 8016 15528 8022
rect 15476 7958 15528 7964
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 15384 7948 15436 7954
rect 15384 7890 15436 7896
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15304 7546 15332 7890
rect 15488 7546 15516 7958
rect 15856 7818 15884 8298
rect 15844 7812 15896 7818
rect 15844 7754 15896 7760
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 14016 6730 14044 7346
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 15120 7002 15148 7278
rect 16132 7274 16160 8434
rect 16224 7274 16252 8910
rect 17144 8634 17172 8978
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 16396 8356 16448 8362
rect 16396 8298 16448 8304
rect 16408 7410 16436 8298
rect 17040 7948 17092 7954
rect 17040 7890 17092 7896
rect 17052 7750 17080 7890
rect 17144 7818 17172 8570
rect 17132 7812 17184 7818
rect 17132 7754 17184 7760
rect 17040 7744 17092 7750
rect 17040 7686 17092 7692
rect 17052 7546 17080 7686
rect 17040 7540 17092 7546
rect 17040 7482 17092 7488
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 16120 7268 16172 7274
rect 16120 7210 16172 7216
rect 16212 7268 16264 7274
rect 16212 7210 16264 7216
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 14556 6928 14608 6934
rect 14556 6870 14608 6876
rect 14004 6724 14056 6730
rect 14004 6666 14056 6672
rect 14568 6458 14596 6870
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13544 4208 13596 4214
rect 13544 4150 13596 4156
rect 13556 3942 13584 4150
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13556 3670 13584 3878
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 13556 3194 13584 3606
rect 13636 3528 13688 3534
rect 13740 3516 13768 5510
rect 13832 4690 13860 5578
rect 13924 5166 13952 5714
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 13832 4146 13860 4626
rect 13912 4616 13964 4622
rect 13912 4558 13964 4564
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13832 3534 13860 3946
rect 13688 3488 13768 3516
rect 13636 3470 13688 3476
rect 13544 3188 13596 3194
rect 13544 3130 13596 3136
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 13266 2952 13322 2961
rect 13266 2887 13322 2896
rect 12898 1728 12954 1737
rect 12898 1663 12954 1672
rect 12162 54 12480 82
rect 13280 82 13308 2887
rect 13372 2582 13400 2994
rect 13360 2576 13412 2582
rect 13360 2518 13412 2524
rect 13740 2417 13768 3488
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13924 2514 13952 4558
rect 14016 4282 14044 6054
rect 14660 5710 14688 6734
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 14740 6180 14792 6186
rect 14740 6122 14792 6128
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 14648 5704 14700 5710
rect 14648 5646 14700 5652
rect 14278 5400 14334 5409
rect 14278 5335 14334 5344
rect 14292 5166 14320 5335
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 14292 4690 14320 5102
rect 14280 4684 14332 4690
rect 14280 4626 14332 4632
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 14200 3194 14228 4558
rect 14292 3738 14320 4626
rect 14384 4622 14412 5646
rect 14752 5166 14780 6122
rect 15120 5914 15148 6258
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14556 5160 14608 5166
rect 14556 5102 14608 5108
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 14568 3534 14596 5102
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 14752 4078 14780 4762
rect 14844 4146 14872 4762
rect 15212 4758 15240 5102
rect 15200 4752 15252 4758
rect 15200 4694 15252 4700
rect 15304 4706 15332 7142
rect 16132 7002 16160 7210
rect 16120 6996 16172 7002
rect 16120 6938 16172 6944
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 15384 6792 15436 6798
rect 15384 6734 15436 6740
rect 15396 5914 15424 6734
rect 15476 6180 15528 6186
rect 15476 6122 15528 6128
rect 15384 5908 15436 5914
rect 15384 5850 15436 5856
rect 15488 5778 15516 6122
rect 16224 6118 16252 6802
rect 16500 6254 16528 6938
rect 16764 6656 16816 6662
rect 16764 6598 16816 6604
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 16776 6254 16804 6598
rect 16868 6458 16896 6598
rect 17236 6458 17264 6598
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 17224 6452 17276 6458
rect 17224 6394 17276 6400
rect 17236 6361 17264 6394
rect 17222 6352 17278 6361
rect 17222 6287 17278 6296
rect 16488 6248 16540 6254
rect 16488 6190 16540 6196
rect 16764 6248 16816 6254
rect 16764 6190 16816 6196
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15396 4826 15424 5102
rect 15948 4826 15976 6054
rect 16224 5370 16252 6054
rect 16672 5840 16724 5846
rect 16672 5782 16724 5788
rect 16212 5364 16264 5370
rect 16212 5306 16264 5312
rect 16028 5296 16080 5302
rect 16028 5238 16080 5244
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 15212 4468 15240 4694
rect 15304 4678 15424 4706
rect 15212 4440 15332 4468
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15304 4146 15332 4440
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 14752 3738 14780 4014
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 15304 3670 15332 4082
rect 15292 3664 15344 3670
rect 15292 3606 15344 3612
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14568 2650 14596 3470
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15396 3194 15424 4678
rect 15844 4004 15896 4010
rect 15844 3946 15896 3952
rect 15856 3738 15884 3946
rect 15844 3732 15896 3738
rect 15844 3674 15896 3680
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15292 3120 15344 3126
rect 15292 3062 15344 3068
rect 15304 2854 15332 3062
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 15384 2848 15436 2854
rect 15384 2790 15436 2796
rect 14556 2644 14608 2650
rect 14556 2586 14608 2592
rect 15396 2582 15424 2790
rect 14648 2576 14700 2582
rect 14648 2518 14700 2524
rect 15384 2576 15436 2582
rect 15384 2518 15436 2524
rect 13912 2508 13964 2514
rect 13912 2450 13964 2456
rect 13726 2408 13782 2417
rect 13726 2343 13782 2352
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 13740 2009 13768 2246
rect 13726 2000 13782 2009
rect 13726 1935 13782 1944
rect 13358 82 13414 480
rect 13280 54 13414 82
rect 12162 0 12218 54
rect 13358 0 13414 54
rect 14554 82 14610 480
rect 14660 82 14688 2518
rect 16040 2446 16068 5238
rect 16684 5030 16712 5782
rect 16948 5704 17000 5710
rect 16948 5646 17000 5652
rect 16764 5636 16816 5642
rect 16764 5578 16816 5584
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 16684 4758 16712 4966
rect 16672 4752 16724 4758
rect 16672 4694 16724 4700
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16316 4049 16344 4422
rect 16684 4078 16712 4558
rect 16672 4072 16724 4078
rect 16302 4040 16358 4049
rect 16672 4014 16724 4020
rect 16302 3975 16358 3984
rect 16672 3392 16724 3398
rect 16672 3334 16724 3340
rect 16684 3058 16712 3334
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 16396 2916 16448 2922
rect 16396 2858 16448 2864
rect 16408 2514 16436 2858
rect 16684 2582 16712 2994
rect 16672 2576 16724 2582
rect 16672 2518 16724 2524
rect 16396 2508 16448 2514
rect 16396 2450 16448 2456
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 15384 2372 15436 2378
rect 15384 2314 15436 2320
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14554 54 14688 82
rect 15396 82 15424 2314
rect 15658 82 15714 480
rect 15396 54 15714 82
rect 16776 82 16804 5578
rect 16960 5370 16988 5646
rect 16948 5364 17000 5370
rect 16948 5306 17000 5312
rect 17052 5234 17080 6054
rect 17144 5642 17172 6190
rect 17132 5636 17184 5642
rect 17132 5578 17184 5584
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16868 4282 16896 5102
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 16868 4010 16896 4218
rect 17040 4208 17092 4214
rect 17224 4208 17276 4214
rect 17092 4168 17224 4196
rect 17040 4150 17092 4156
rect 17224 4150 17276 4156
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 16856 4004 16908 4010
rect 16856 3946 16908 3952
rect 17236 3670 17264 4014
rect 17224 3664 17276 3670
rect 17224 3606 17276 3612
rect 17236 3194 17264 3606
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 17052 2514 17080 3130
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 17052 2310 17080 2450
rect 17040 2304 17092 2310
rect 17040 2246 17092 2252
rect 16854 82 16910 480
rect 17328 134 17356 9318
rect 18616 9042 18644 10134
rect 23848 10124 23900 10130
rect 23848 10066 23900 10072
rect 19064 10056 19116 10062
rect 23860 10033 23888 10066
rect 19064 9998 19116 10004
rect 23846 10024 23902 10033
rect 19076 9654 19104 9998
rect 23846 9959 23902 9968
rect 23860 9722 23888 9959
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 23848 9716 23900 9722
rect 23848 9658 23900 9664
rect 19064 9648 19116 9654
rect 19064 9590 19116 9596
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 18696 9444 18748 9450
rect 18696 9386 18748 9392
rect 18708 9178 18736 9386
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18604 9036 18656 9042
rect 18604 8978 18656 8984
rect 18616 8634 18644 8978
rect 19536 8634 19564 9522
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 19524 8628 19576 8634
rect 19524 8570 19576 8576
rect 21180 8288 21232 8294
rect 21180 8230 21232 8236
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 17500 7948 17552 7954
rect 17500 7890 17552 7896
rect 17512 7546 17540 7890
rect 18418 7848 18474 7857
rect 18418 7783 18474 7792
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 18052 7268 18104 7274
rect 18052 7210 18104 7216
rect 18064 6934 18092 7210
rect 18052 6928 18104 6934
rect 18052 6870 18104 6876
rect 18432 6866 18460 7783
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 18880 6860 18932 6866
rect 18880 6802 18932 6808
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17512 5778 17540 6734
rect 18432 6458 18460 6802
rect 18420 6452 18472 6458
rect 18420 6394 18472 6400
rect 18892 6254 18920 6802
rect 18880 6248 18932 6254
rect 18880 6190 18932 6196
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 17776 5840 17828 5846
rect 17776 5782 17828 5788
rect 17500 5772 17552 5778
rect 17500 5714 17552 5720
rect 17512 5681 17540 5714
rect 17498 5672 17554 5681
rect 17498 5607 17554 5616
rect 17788 5030 17816 5782
rect 18144 5704 18196 5710
rect 18144 5646 18196 5652
rect 18156 5545 18184 5646
rect 18142 5536 18198 5545
rect 18142 5471 18198 5480
rect 18156 5370 18184 5471
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 18696 5160 18748 5166
rect 18696 5102 18748 5108
rect 17960 5092 18012 5098
rect 17960 5034 18012 5040
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 17788 4826 17816 4966
rect 17776 4820 17828 4826
rect 17776 4762 17828 4768
rect 17776 4004 17828 4010
rect 17776 3946 17828 3952
rect 17788 3670 17816 3946
rect 17972 3738 18000 5034
rect 18708 4486 18736 5102
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 18788 4684 18840 4690
rect 18788 4626 18840 4632
rect 18696 4480 18748 4486
rect 18696 4422 18748 4428
rect 18708 4185 18736 4422
rect 18800 4214 18828 4626
rect 18788 4208 18840 4214
rect 18694 4176 18750 4185
rect 18788 4150 18840 4156
rect 18694 4111 18750 4120
rect 18972 4140 19024 4146
rect 18052 4004 18104 4010
rect 18052 3946 18104 3952
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 17776 3664 17828 3670
rect 17776 3606 17828 3612
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 17420 2582 17448 3334
rect 18064 3194 18092 3946
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 18052 3188 18104 3194
rect 18052 3130 18104 3136
rect 17868 2916 17920 2922
rect 17868 2858 17920 2864
rect 17880 2582 17908 2858
rect 18064 2854 18092 3130
rect 18156 3058 18184 3878
rect 18708 3670 18736 4111
rect 18972 4082 19024 4088
rect 18696 3664 18748 3670
rect 18696 3606 18748 3612
rect 18984 3534 19012 4082
rect 21088 4072 21140 4078
rect 21088 4014 21140 4020
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19064 3664 19116 3670
rect 19064 3606 19116 3612
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18972 3528 19024 3534
rect 18972 3470 19024 3476
rect 18432 3058 18460 3470
rect 19076 3194 19104 3606
rect 19064 3188 19116 3194
rect 19064 3130 19116 3136
rect 19996 3097 20024 3878
rect 20904 3596 20956 3602
rect 20904 3538 20956 3544
rect 19982 3088 20038 3097
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18420 3052 18472 3058
rect 19982 3023 20038 3032
rect 18420 2994 18472 3000
rect 18052 2848 18104 2854
rect 18052 2790 18104 2796
rect 18156 2650 18184 2994
rect 20916 2854 20944 3538
rect 19432 2848 19484 2854
rect 19432 2790 19484 2796
rect 20904 2848 20956 2854
rect 20904 2790 20956 2796
rect 20996 2848 21048 2854
rect 20996 2790 21048 2796
rect 19444 2689 19472 2790
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19430 2680 19486 2689
rect 18144 2644 18196 2650
rect 19622 2672 19918 2692
rect 19430 2615 19486 2624
rect 18144 2586 18196 2592
rect 17408 2576 17460 2582
rect 17408 2518 17460 2524
rect 17868 2576 17920 2582
rect 17868 2518 17920 2524
rect 20720 2508 20772 2514
rect 20720 2450 20772 2456
rect 18144 2372 18196 2378
rect 18144 2314 18196 2320
rect 16776 54 16910 82
rect 17316 128 17368 134
rect 17316 70 17368 76
rect 18050 82 18106 480
rect 18156 82 18184 2314
rect 19800 2304 19852 2310
rect 19800 2246 19852 2252
rect 19812 1737 19840 2246
rect 19798 1728 19854 1737
rect 19798 1663 19854 1672
rect 14554 0 14610 54
rect 15658 0 15714 54
rect 16854 0 16910 54
rect 18050 54 18184 82
rect 19154 128 19210 480
rect 19154 76 19156 128
rect 19208 76 19210 128
rect 18050 0 18106 54
rect 19154 0 19210 76
rect 20350 82 20406 480
rect 20732 82 20760 2450
rect 20916 1737 20944 2790
rect 21008 2650 21036 2790
rect 20996 2644 21048 2650
rect 20996 2586 21048 2592
rect 21100 1873 21128 4014
rect 21086 1864 21142 1873
rect 21086 1799 21142 1808
rect 20902 1728 20958 1737
rect 20902 1663 20958 1672
rect 20350 54 20760 82
rect 21192 82 21220 8230
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 23204 6860 23256 6866
rect 23204 6802 23256 6808
rect 23216 6118 23244 6802
rect 23940 6656 23992 6662
rect 23940 6598 23992 6604
rect 23952 6458 23980 6598
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 23940 6452 23992 6458
rect 23940 6394 23992 6400
rect 23952 6118 23980 6394
rect 23204 6112 23256 6118
rect 23204 6054 23256 6060
rect 23940 6112 23992 6118
rect 23940 6054 23992 6060
rect 23216 5846 23244 6054
rect 23204 5840 23256 5846
rect 23110 5808 23166 5817
rect 23204 5782 23256 5788
rect 23110 5743 23112 5752
rect 23164 5743 23166 5752
rect 23112 5714 23164 5720
rect 23124 5370 23152 5714
rect 23216 5370 23244 5782
rect 24032 5636 24084 5642
rect 24032 5578 24084 5584
rect 23848 5568 23900 5574
rect 24044 5545 24072 5578
rect 23848 5510 23900 5516
rect 24030 5536 24086 5545
rect 23112 5364 23164 5370
rect 23112 5306 23164 5312
rect 23204 5364 23256 5370
rect 23204 5306 23256 5312
rect 23216 5273 23244 5306
rect 23202 5264 23258 5273
rect 23202 5199 23258 5208
rect 22284 5024 22336 5030
rect 22284 4966 22336 4972
rect 22296 4146 22324 4966
rect 22560 4752 22612 4758
rect 22560 4694 22612 4700
rect 22468 4616 22520 4622
rect 22468 4558 22520 4564
rect 22480 4282 22508 4558
rect 22468 4276 22520 4282
rect 22468 4218 22520 4224
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 22192 4004 22244 4010
rect 22192 3946 22244 3952
rect 22204 3670 22232 3946
rect 22296 3738 22324 4082
rect 22572 4049 22600 4694
rect 23860 4622 23888 5510
rect 24030 5471 24086 5480
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24124 5160 24176 5166
rect 24124 5102 24176 5108
rect 23940 5024 23992 5030
rect 23940 4966 23992 4972
rect 22744 4616 22796 4622
rect 22744 4558 22796 4564
rect 23848 4616 23900 4622
rect 23848 4558 23900 4564
rect 22756 4146 22784 4558
rect 23952 4282 23980 4966
rect 24136 4758 24164 5102
rect 24124 4752 24176 4758
rect 24124 4694 24176 4700
rect 24032 4616 24084 4622
rect 24032 4558 24084 4564
rect 23940 4276 23992 4282
rect 23940 4218 23992 4224
rect 22744 4140 22796 4146
rect 22744 4082 22796 4088
rect 22558 4040 22614 4049
rect 22558 3975 22614 3984
rect 22572 3942 22600 3975
rect 22560 3936 22612 3942
rect 22560 3878 22612 3884
rect 22284 3732 22336 3738
rect 22284 3674 22336 3680
rect 22192 3664 22244 3670
rect 22192 3606 22244 3612
rect 22572 3602 22600 3878
rect 22756 3602 22784 4082
rect 23952 3942 23980 4218
rect 23940 3936 23992 3942
rect 23940 3878 23992 3884
rect 24044 3738 24072 4558
rect 24136 4214 24164 4694
rect 24216 4616 24268 4622
rect 24216 4558 24268 4564
rect 24124 4208 24176 4214
rect 24124 4150 24176 4156
rect 24228 4146 24256 4558
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24780 4154 24808 11494
rect 25226 10976 25282 10985
rect 25226 10911 25282 10920
rect 25240 10810 25268 10911
rect 25228 10804 25280 10810
rect 25228 10746 25280 10752
rect 25134 8392 25190 8401
rect 25134 8327 25190 8336
rect 25148 7546 25176 8327
rect 25136 7540 25188 7546
rect 25136 7482 25188 7488
rect 25148 7342 25176 7482
rect 25136 7336 25188 7342
rect 25136 7278 25188 7284
rect 25136 7200 25188 7206
rect 25136 7142 25188 7148
rect 25148 6458 25176 7142
rect 25136 6452 25188 6458
rect 25136 6394 25188 6400
rect 24860 6180 24912 6186
rect 24860 6122 24912 6128
rect 24872 5642 24900 6122
rect 25044 5704 25096 5710
rect 25044 5646 25096 5652
rect 24860 5636 24912 5642
rect 24860 5578 24912 5584
rect 25056 5370 25084 5646
rect 25044 5364 25096 5370
rect 25044 5306 25096 5312
rect 27068 5024 27120 5030
rect 27068 4966 27120 4972
rect 24216 4140 24268 4146
rect 24780 4126 24900 4154
rect 24216 4082 24268 4088
rect 24216 4004 24268 4010
rect 24216 3946 24268 3952
rect 24032 3732 24084 3738
rect 24032 3674 24084 3680
rect 24228 3602 24256 3946
rect 22560 3596 22612 3602
rect 22560 3538 22612 3544
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 23480 3596 23532 3602
rect 23480 3538 23532 3544
rect 24216 3596 24268 3602
rect 24216 3538 24268 3544
rect 22572 3194 22600 3538
rect 23388 3392 23440 3398
rect 23388 3334 23440 3340
rect 22560 3188 22612 3194
rect 22560 3130 22612 3136
rect 22652 3052 22704 3058
rect 22652 2994 22704 3000
rect 22664 2961 22692 2994
rect 22650 2952 22706 2961
rect 22650 2887 22706 2896
rect 21456 2848 21508 2854
rect 21456 2790 21508 2796
rect 23112 2848 23164 2854
rect 23112 2790 23164 2796
rect 21468 2009 21496 2790
rect 23124 2417 23152 2790
rect 23400 2650 23428 3334
rect 23492 3194 23520 3538
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 23480 3188 23532 3194
rect 23480 3130 23532 3136
rect 23388 2644 23440 2650
rect 23388 2586 23440 2592
rect 23110 2408 23166 2417
rect 22744 2372 22796 2378
rect 23110 2343 23166 2352
rect 23664 2372 23716 2378
rect 22744 2314 22796 2320
rect 23664 2314 23716 2320
rect 21454 2000 21510 2009
rect 21454 1935 21510 1944
rect 21546 82 21602 480
rect 21192 54 21602 82
rect 20350 0 20406 54
rect 21546 0 21602 54
rect 22650 82 22706 480
rect 22756 82 22784 2314
rect 22650 54 22784 82
rect 23676 82 23704 2314
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 23846 82 23902 480
rect 23676 54 23902 82
rect 24872 82 24900 4126
rect 24952 3596 25004 3602
rect 24952 3538 25004 3544
rect 24964 3194 24992 3538
rect 26974 3496 27030 3505
rect 26974 3431 27030 3440
rect 26988 3194 27016 3431
rect 24952 3188 25004 3194
rect 24952 3130 25004 3136
rect 26976 3188 27028 3194
rect 26976 3130 27028 3136
rect 25780 2984 25832 2990
rect 25780 2926 25832 2932
rect 25042 82 25098 480
rect 24872 54 25098 82
rect 25792 82 25820 2926
rect 26146 82 26202 480
rect 25792 54 26202 82
rect 27080 82 27108 4966
rect 27342 82 27398 480
rect 27080 54 27398 82
rect 22650 0 22706 54
rect 23846 0 23902 54
rect 25042 0 25098 54
rect 26146 0 26202 54
rect 27342 0 27398 54
<< via2 >>
rect 1030 26424 1086 26480
rect 110 24928 166 24984
rect 1214 22344 1270 22400
rect 110 20984 166 21040
rect 110 16904 166 16960
rect 110 15544 166 15600
rect 1582 14592 1638 14648
rect 1582 13504 1638 13560
rect 1858 10376 1914 10432
rect 1766 9424 1822 9480
rect 2134 9152 2190 9208
rect 1306 4528 1362 4584
rect 2042 5888 2098 5944
rect 110 992 166 1048
rect 3238 7112 3294 7168
rect 2226 2624 2282 2680
rect 2962 6432 3018 6488
rect 3606 9560 3662 9616
rect 3606 9036 3662 9072
rect 3606 9016 3608 9036
rect 3608 9016 3660 9036
rect 3660 9016 3662 9036
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 4250 12824 4306 12880
rect 3790 8880 3846 8936
rect 4158 9016 4214 9072
rect 4618 10648 4674 10704
rect 4618 9968 4674 10024
rect 3514 6976 3570 7032
rect 4158 7112 4214 7168
rect 3974 6976 4030 7032
rect 3422 5888 3478 5944
rect 2686 3032 2742 3088
rect 3698 5208 3754 5264
rect 3790 4936 3846 4992
rect 2962 2896 3018 2952
rect 5078 9152 5134 9208
rect 4802 8880 4858 8936
rect 4434 3984 4490 4040
rect 4342 2624 4398 2680
rect 4618 3440 4674 3496
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 6182 14864 6238 14920
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 6090 6296 6146 6352
rect 5170 4120 5226 4176
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 6826 9560 6882 9616
rect 6274 4936 6330 4992
rect 6090 4120 6146 4176
rect 6182 3848 6238 3904
rect 7194 4936 7250 4992
rect 5906 2896 5962 2952
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 10966 22480 11022 22536
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 8482 14456 8538 14512
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 8758 12824 8814 12880
rect 9310 13776 9366 13832
rect 11518 18128 11574 18184
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 8666 8336 8722 8392
rect 9494 7792 9550 7848
rect 8298 6296 8354 6352
rect 8206 5480 8262 5536
rect 8482 5344 8538 5400
rect 7378 4256 7434 4312
rect 8114 4120 8170 4176
rect 7562 3304 7618 3360
rect 7378 3032 7434 3088
rect 9126 6296 9182 6352
rect 9586 7112 9642 7168
rect 9678 6976 9734 7032
rect 9310 5208 9366 5264
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 12714 20304 12770 20360
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 9862 5616 9918 5672
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10414 4256 10470 4312
rect 10138 4120 10194 4176
rect 9402 3984 9458 4040
rect 9586 3440 9642 3496
rect 9494 2624 9550 2680
rect 9862 3984 9918 4040
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 11150 5480 11206 5536
rect 11058 3984 11114 4040
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 11978 4120 12034 4176
rect 9770 1808 9826 1864
rect 13358 5208 13414 5264
rect 12530 2760 12586 2816
rect 12898 3304 12954 3360
rect 12806 2624 12862 2680
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 25134 26152 25190 26208
rect 18326 22480 18382 22536
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 15658 20304 15714 20360
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14186 15544 14242 15600
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 15658 14456 15714 14512
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14186 11600 14242 11656
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 15290 10512 15346 10568
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14186 8336 14242 8392
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19338 13776 19394 13832
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 24766 23432 24822 23488
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24674 21004 24730 21040
rect 24674 20984 24676 21004
rect 24676 20984 24728 21004
rect 24728 20984 24730 21004
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24122 11600 24178 11656
rect 18602 10648 18658 10704
rect 24030 10512 24086 10568
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24490 14864 24546 14920
rect 24766 18536 24822 18592
rect 24766 15952 24822 16008
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24766 13640 24822 13696
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 13266 2896 13322 2952
rect 12898 1672 12954 1728
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14278 5344 14334 5400
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 17222 6296 17278 6352
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 13726 2352 13782 2408
rect 13726 1944 13782 2000
rect 16302 3984 16358 4040
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 23846 9968 23902 10024
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 18418 7792 18474 7848
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 17498 5616 17554 5672
rect 18142 5480 18198 5536
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 18694 4120 18750 4176
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19982 3032 20038 3088
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 19430 2624 19486 2680
rect 19798 1672 19854 1728
rect 21086 1808 21142 1864
rect 20902 1672 20958 1728
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 23110 5772 23166 5808
rect 23110 5752 23112 5772
rect 23112 5752 23164 5772
rect 23164 5752 23166 5772
rect 23202 5208 23258 5264
rect 24030 5480 24086 5536
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 22558 3984 22614 4040
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 25226 10920 25282 10976
rect 25134 8336 25190 8392
rect 22650 2896 22706 2952
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 23110 2352 23166 2408
rect 21454 1944 21510 2000
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 26974 3440 27030 3496
<< metal3 >>
rect 0 26936 480 27056
rect 62 26482 122 26936
rect 27520 26664 28000 26784
rect 1025 26482 1091 26485
rect 62 26480 1091 26482
rect 62 26424 1030 26480
rect 1086 26424 1091 26480
rect 62 26422 1091 26424
rect 1025 26419 1091 26422
rect 25129 26210 25195 26213
rect 27662 26210 27722 26664
rect 25129 26208 27722 26210
rect 25129 26152 25134 26208
rect 25190 26152 27722 26208
rect 25129 26150 27722 26152
rect 25129 26147 25195 26150
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 5610 25056 5930 25057
rect 0 24984 480 25016
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 0 24928 110 24984
rect 166 24928 480 24984
rect 0 24896 480 24928
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 27520 24172 28000 24200
rect 27520 24108 27660 24172
rect 27724 24108 28000 24172
rect 27520 24080 28000 24108
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 24761 23490 24827 23493
rect 27654 23490 27660 23492
rect 24761 23488 27660 23490
rect 24761 23432 24766 23488
rect 24822 23432 27660 23488
rect 24761 23430 27660 23432
rect 24761 23427 24827 23430
rect 27654 23428 27660 23430
rect 27724 23428 27730 23492
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 0 22856 480 22976
rect 5610 22880 5930 22881
rect 62 22402 122 22856
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 10961 22538 11027 22541
rect 18321 22538 18387 22541
rect 10961 22536 18387 22538
rect 10961 22480 10966 22536
rect 11022 22480 18326 22536
rect 18382 22480 18387 22536
rect 10961 22478 18387 22480
rect 10961 22475 11027 22478
rect 18321 22475 18387 22478
rect 1209 22402 1275 22405
rect 62 22400 1275 22402
rect 62 22344 1214 22400
rect 1270 22344 1275 22400
rect 62 22342 1275 22344
rect 1209 22339 1275 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 27520 21496 28000 21616
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 0 21040 480 21072
rect 0 20984 110 21040
rect 166 20984 480 21040
rect 0 20952 480 20984
rect 24669 21042 24735 21045
rect 27662 21042 27722 21496
rect 24669 21040 27722 21042
rect 24669 20984 24674 21040
rect 24730 20984 27722 21040
rect 24669 20982 27722 20984
rect 24669 20979 24735 20982
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 12709 20362 12775 20365
rect 15653 20362 15719 20365
rect 12709 20360 15719 20362
rect 12709 20304 12714 20360
rect 12770 20304 15658 20360
rect 15714 20304 15719 20360
rect 12709 20302 15719 20304
rect 12709 20299 12775 20302
rect 15653 20299 15719 20302
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 10277 19072 10597 19073
rect 0 18912 480 19032
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 27520 19048 28000 19168
rect 19610 19007 19930 19008
rect 62 18186 122 18912
rect 24761 18594 24827 18597
rect 27662 18594 27722 19048
rect 24761 18592 27722 18594
rect 24761 18536 24766 18592
rect 24822 18536 27722 18592
rect 24761 18534 27722 18536
rect 24761 18531 24827 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 11513 18186 11579 18189
rect 62 18184 11579 18186
rect 62 18128 11518 18184
rect 11574 18128 11579 18184
rect 62 18126 11579 18128
rect 11513 18123 11579 18126
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 0 16960 480 16992
rect 0 16904 110 16960
rect 166 16904 480 16960
rect 0 16872 480 16904
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 27520 16464 28000 16584
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 24761 16010 24827 16013
rect 27662 16010 27722 16464
rect 24761 16008 27722 16010
rect 24761 15952 24766 16008
rect 24822 15952 27722 16008
rect 24761 15950 27722 15952
rect 24761 15947 24827 15950
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 105 15602 171 15605
rect 14181 15602 14247 15605
rect 105 15600 14247 15602
rect 105 15544 110 15600
rect 166 15544 14186 15600
rect 14242 15544 14247 15600
rect 105 15542 14247 15544
rect 105 15539 171 15542
rect 14181 15539 14247 15542
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 0 14968 480 15088
rect 62 14650 122 14968
rect 6177 14922 6243 14925
rect 24485 14922 24551 14925
rect 6177 14920 24551 14922
rect 6177 14864 6182 14920
rect 6238 14864 24490 14920
rect 24546 14864 24551 14920
rect 6177 14862 24551 14864
rect 6177 14859 6243 14862
rect 24485 14859 24551 14862
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 1577 14650 1643 14653
rect 62 14648 1643 14650
rect 62 14592 1582 14648
rect 1638 14592 1643 14648
rect 62 14590 1643 14592
rect 1577 14587 1643 14590
rect 8477 14514 8543 14517
rect 15653 14514 15719 14517
rect 8477 14512 15719 14514
rect 8477 14456 8482 14512
rect 8538 14456 15658 14512
rect 15714 14456 15719 14512
rect 8477 14454 15719 14456
rect 8477 14451 8543 14454
rect 15653 14451 15719 14454
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 27520 13880 28000 14000
rect 9305 13834 9371 13837
rect 19333 13834 19399 13837
rect 9305 13832 19399 13834
rect 9305 13776 9310 13832
rect 9366 13776 19338 13832
rect 19394 13776 19399 13832
rect 9305 13774 19399 13776
rect 9305 13771 9371 13774
rect 19333 13771 19399 13774
rect 24761 13698 24827 13701
rect 27662 13698 27722 13880
rect 24761 13696 27722 13698
rect 24761 13640 24766 13696
rect 24822 13640 27722 13696
rect 24761 13638 27722 13640
rect 24761 13635 24827 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 1577 13562 1643 13565
rect 62 13560 1643 13562
rect 62 13504 1582 13560
rect 1638 13504 1643 13560
rect 62 13502 1643 13504
rect 62 13048 122 13502
rect 1577 13499 1643 13502
rect 5610 13088 5930 13089
rect 0 12928 480 13048
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 4245 12882 4311 12885
rect 8753 12882 8819 12885
rect 4245 12880 8819 12882
rect 4245 12824 4250 12880
rect 4306 12824 8758 12880
rect 8814 12824 8819 12880
rect 4245 12822 8819 12824
rect 4245 12819 4311 12822
rect 8753 12819 8819 12822
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 14181 11658 14247 11661
rect 24117 11658 24183 11661
rect 14181 11656 24183 11658
rect 14181 11600 14186 11656
rect 14242 11600 24122 11656
rect 24178 11600 24183 11656
rect 14181 11598 24183 11600
rect 14181 11595 14247 11598
rect 24117 11595 24183 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 27520 11296 28000 11416
rect 0 10888 480 11008
rect 25221 10978 25287 10981
rect 27662 10978 27722 11296
rect 25221 10976 27722 10978
rect 25221 10920 25226 10976
rect 25282 10920 27722 10976
rect 25221 10918 27722 10920
rect 25221 10915 25287 10918
rect 5610 10912 5930 10913
rect 62 10434 122 10888
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 4613 10706 4679 10709
rect 18597 10706 18663 10709
rect 4613 10704 18663 10706
rect 4613 10648 4618 10704
rect 4674 10648 18602 10704
rect 18658 10648 18663 10704
rect 4613 10646 18663 10648
rect 4613 10643 4679 10646
rect 18597 10643 18663 10646
rect 15285 10570 15351 10573
rect 24025 10570 24091 10573
rect 15285 10568 24091 10570
rect 15285 10512 15290 10568
rect 15346 10512 24030 10568
rect 24086 10512 24091 10568
rect 15285 10510 24091 10512
rect 15285 10507 15351 10510
rect 24025 10507 24091 10510
rect 1853 10434 1919 10437
rect 62 10432 1919 10434
rect 62 10376 1858 10432
rect 1914 10376 1919 10432
rect 62 10374 1919 10376
rect 1853 10371 1919 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 4613 10026 4679 10029
rect 23841 10026 23907 10029
rect 4613 10024 23907 10026
rect 4613 9968 4618 10024
rect 4674 9968 23846 10024
rect 23902 9968 23907 10024
rect 4613 9966 23907 9968
rect 4613 9963 4679 9966
rect 23841 9963 23907 9966
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 3601 9618 3667 9621
rect 6821 9618 6887 9621
rect 3601 9616 6887 9618
rect 3601 9560 3606 9616
rect 3662 9560 6826 9616
rect 6882 9560 6887 9616
rect 3601 9558 6887 9560
rect 3601 9555 3667 9558
rect 6821 9555 6887 9558
rect 1761 9482 1827 9485
rect 62 9480 1827 9482
rect 62 9424 1766 9480
rect 1822 9424 1827 9480
rect 62 9422 1827 9424
rect 62 8968 122 9422
rect 1761 9419 1827 9422
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 2129 9210 2195 9213
rect 5073 9210 5139 9213
rect 2129 9208 5139 9210
rect 2129 9152 2134 9208
rect 2190 9152 5078 9208
rect 5134 9152 5139 9208
rect 2129 9150 5139 9152
rect 2129 9147 2195 9150
rect 5073 9147 5139 9150
rect 3601 9074 3667 9077
rect 4153 9074 4219 9077
rect 3601 9072 4219 9074
rect 3601 9016 3606 9072
rect 3662 9016 4158 9072
rect 4214 9016 4219 9072
rect 3601 9014 4219 9016
rect 3601 9011 3667 9014
rect 4153 9011 4219 9014
rect 0 8848 480 8968
rect 3785 8938 3851 8941
rect 4797 8938 4863 8941
rect 3785 8936 4863 8938
rect 3785 8880 3790 8936
rect 3846 8880 4802 8936
rect 4858 8880 4863 8936
rect 3785 8878 4863 8880
rect 3785 8875 3851 8878
rect 4797 8875 4863 8878
rect 27520 8848 28000 8968
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 8661 8394 8727 8397
rect 14181 8394 14247 8397
rect 8661 8392 14247 8394
rect 8661 8336 8666 8392
rect 8722 8336 14186 8392
rect 14242 8336 14247 8392
rect 8661 8334 14247 8336
rect 8661 8331 8727 8334
rect 14181 8331 14247 8334
rect 25129 8394 25195 8397
rect 27662 8394 27722 8848
rect 25129 8392 27722 8394
rect 25129 8336 25134 8392
rect 25190 8336 27722 8392
rect 25129 8334 27722 8336
rect 25129 8331 25195 8334
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 9489 7850 9555 7853
rect 18413 7850 18479 7853
rect 9489 7848 18479 7850
rect 9489 7792 9494 7848
rect 9550 7792 18418 7848
rect 18474 7792 18479 7848
rect 9489 7790 18479 7792
rect 9489 7787 9555 7790
rect 18413 7787 18479 7790
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 3233 7170 3299 7173
rect 4153 7170 4219 7173
rect 9581 7170 9647 7173
rect 3233 7168 9647 7170
rect 3233 7112 3238 7168
rect 3294 7112 4158 7168
rect 4214 7112 9586 7168
rect 9642 7112 9647 7168
rect 3233 7110 9647 7112
rect 3233 7107 3299 7110
rect 4153 7107 4219 7110
rect 9581 7107 9647 7110
rect 10277 7104 10597 7105
rect 0 6944 480 7064
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 3509 7034 3575 7037
rect 3969 7034 4035 7037
rect 9673 7034 9739 7037
rect 3509 7032 9739 7034
rect 3509 6976 3514 7032
rect 3570 6976 3974 7032
rect 4030 6976 9678 7032
rect 9734 6976 9739 7032
rect 3509 6974 9739 6976
rect 3509 6971 3575 6974
rect 3969 6971 4035 6974
rect 9673 6971 9739 6974
rect 62 6490 122 6944
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 2957 6490 3023 6493
rect 62 6488 3023 6490
rect 62 6432 2962 6488
rect 3018 6432 3023 6488
rect 62 6430 3023 6432
rect 2957 6427 3023 6430
rect 6085 6354 6151 6357
rect 8293 6354 8359 6357
rect 6085 6352 8359 6354
rect 6085 6296 6090 6352
rect 6146 6296 8298 6352
rect 8354 6296 8359 6352
rect 6085 6294 8359 6296
rect 6085 6291 6151 6294
rect 8293 6291 8359 6294
rect 9121 6354 9187 6357
rect 17217 6354 17283 6357
rect 9121 6352 17283 6354
rect 9121 6296 9126 6352
rect 9182 6296 17222 6352
rect 17278 6296 17283 6352
rect 9121 6294 17283 6296
rect 9121 6291 9187 6294
rect 17217 6291 17283 6294
rect 27520 6264 28000 6384
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 2037 5946 2103 5949
rect 3417 5946 3483 5949
rect 2037 5944 3483 5946
rect 2037 5888 2042 5944
rect 2098 5888 3422 5944
rect 3478 5888 3483 5944
rect 2037 5886 3483 5888
rect 2037 5883 2103 5886
rect 3417 5883 3483 5886
rect 23105 5810 23171 5813
rect 27662 5810 27722 6264
rect 23105 5808 27722 5810
rect 23105 5752 23110 5808
rect 23166 5752 27722 5808
rect 23105 5750 27722 5752
rect 23105 5747 23171 5750
rect 9857 5674 9923 5677
rect 17493 5674 17559 5677
rect 9857 5672 17559 5674
rect 9857 5616 9862 5672
rect 9918 5616 17498 5672
rect 17554 5616 17559 5672
rect 9857 5614 17559 5616
rect 9857 5611 9923 5614
rect 17493 5611 17559 5614
rect 8201 5538 8267 5541
rect 11145 5538 11211 5541
rect 8201 5536 11211 5538
rect 8201 5480 8206 5536
rect 8262 5480 11150 5536
rect 11206 5480 11211 5536
rect 8201 5478 11211 5480
rect 8201 5475 8267 5478
rect 11145 5475 11211 5478
rect 18137 5538 18203 5541
rect 24025 5538 24091 5541
rect 18137 5536 24091 5538
rect 18137 5480 18142 5536
rect 18198 5480 24030 5536
rect 24086 5480 24091 5536
rect 18137 5478 24091 5480
rect 18137 5475 18203 5478
rect 24025 5475 24091 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 8477 5402 8543 5405
rect 14273 5402 14339 5405
rect 8477 5400 14339 5402
rect 8477 5344 8482 5400
rect 8538 5344 14278 5400
rect 14334 5344 14339 5400
rect 8477 5342 14339 5344
rect 8477 5339 8543 5342
rect 14273 5339 14339 5342
rect 3693 5266 3759 5269
rect 9305 5266 9371 5269
rect 3693 5264 9371 5266
rect 3693 5208 3698 5264
rect 3754 5208 9310 5264
rect 9366 5208 9371 5264
rect 3693 5206 9371 5208
rect 3693 5203 3759 5206
rect 9305 5203 9371 5206
rect 13353 5266 13419 5269
rect 23197 5266 23263 5269
rect 13353 5264 23263 5266
rect 13353 5208 13358 5264
rect 13414 5208 23202 5264
rect 23258 5208 23263 5264
rect 13353 5206 23263 5208
rect 13353 5203 13419 5206
rect 23197 5203 23263 5206
rect 0 4904 480 5024
rect 3785 4994 3851 4997
rect 6269 4994 6335 4997
rect 7189 4994 7255 4997
rect 3785 4992 7255 4994
rect 3785 4936 3790 4992
rect 3846 4936 6274 4992
rect 6330 4936 7194 4992
rect 7250 4936 7255 4992
rect 3785 4934 7255 4936
rect 3785 4931 3851 4934
rect 6269 4931 6335 4934
rect 7189 4931 7255 4934
rect 10277 4928 10597 4929
rect 62 4586 122 4904
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 1301 4586 1367 4589
rect 62 4584 1367 4586
rect 62 4528 1306 4584
rect 1362 4528 1367 4584
rect 62 4526 1367 4528
rect 1301 4523 1367 4526
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 7373 4314 7439 4317
rect 10409 4314 10475 4317
rect 7373 4312 10475 4314
rect 7373 4256 7378 4312
rect 7434 4256 10414 4312
rect 10470 4256 10475 4312
rect 7373 4254 10475 4256
rect 7373 4251 7439 4254
rect 10409 4251 10475 4254
rect 5165 4178 5231 4181
rect 6085 4178 6151 4181
rect 5165 4176 6151 4178
rect 5165 4120 5170 4176
rect 5226 4120 6090 4176
rect 6146 4120 6151 4176
rect 5165 4118 6151 4120
rect 5165 4115 5231 4118
rect 6085 4115 6151 4118
rect 8109 4178 8175 4181
rect 10133 4178 10199 4181
rect 8109 4176 10199 4178
rect 8109 4120 8114 4176
rect 8170 4120 10138 4176
rect 10194 4120 10199 4176
rect 8109 4118 10199 4120
rect 8109 4115 8175 4118
rect 10133 4115 10199 4118
rect 11973 4178 12039 4181
rect 18689 4178 18755 4181
rect 11973 4176 18755 4178
rect 11973 4120 11978 4176
rect 12034 4120 18694 4176
rect 18750 4120 18755 4176
rect 11973 4118 18755 4120
rect 11973 4115 12039 4118
rect 18689 4115 18755 4118
rect 4429 4042 4495 4045
rect 9397 4042 9463 4045
rect 9857 4042 9923 4045
rect 11053 4042 11119 4045
rect 4429 4040 9463 4042
rect 4429 3984 4434 4040
rect 4490 3984 9402 4040
rect 9458 3984 9463 4040
rect 4429 3982 9463 3984
rect 4429 3979 4495 3982
rect 9397 3979 9463 3982
rect 9630 4040 11119 4042
rect 9630 3984 9862 4040
rect 9918 3984 11058 4040
rect 11114 3984 11119 4040
rect 9630 3982 11119 3984
rect 6177 3906 6243 3909
rect 9630 3906 9690 3982
rect 9857 3979 9923 3982
rect 11053 3979 11119 3982
rect 16297 4042 16363 4045
rect 22553 4042 22619 4045
rect 16297 4040 22619 4042
rect 16297 3984 16302 4040
rect 16358 3984 22558 4040
rect 22614 3984 22619 4040
rect 16297 3982 22619 3984
rect 16297 3979 16363 3982
rect 22553 3979 22619 3982
rect 6177 3904 9690 3906
rect 6177 3848 6182 3904
rect 6238 3848 9690 3904
rect 6177 3846 9690 3848
rect 6177 3843 6243 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 27520 3680 28000 3800
rect 4613 3498 4679 3501
rect 9581 3498 9647 3501
rect 4613 3496 9647 3498
rect 4613 3440 4618 3496
rect 4674 3440 9586 3496
rect 9642 3440 9647 3496
rect 4613 3438 9647 3440
rect 4613 3435 4679 3438
rect 9581 3435 9647 3438
rect 26969 3498 27035 3501
rect 27662 3498 27722 3680
rect 26969 3496 27722 3498
rect 26969 3440 26974 3496
rect 27030 3440 27722 3496
rect 26969 3438 27722 3440
rect 26969 3435 27035 3438
rect 7557 3362 7623 3365
rect 12893 3362 12959 3365
rect 7557 3360 12959 3362
rect 7557 3304 7562 3360
rect 7618 3304 12898 3360
rect 12954 3304 12959 3360
rect 7557 3302 12959 3304
rect 7557 3299 7623 3302
rect 12893 3299 12959 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 2681 3090 2747 3093
rect 7373 3090 7439 3093
rect 2681 3088 7439 3090
rect 2681 3032 2686 3088
rect 2742 3032 7378 3088
rect 7434 3032 7439 3088
rect 2681 3030 7439 3032
rect 2681 3027 2747 3030
rect 7373 3027 7439 3030
rect 16246 3028 16252 3092
rect 16316 3090 16322 3092
rect 19977 3090 20043 3093
rect 16316 3088 20043 3090
rect 16316 3032 19982 3088
rect 20038 3032 20043 3088
rect 16316 3030 20043 3032
rect 16316 3028 16322 3030
rect 19977 3027 20043 3030
rect 0 2864 480 2984
rect 2957 2954 3023 2957
rect 5901 2954 5967 2957
rect 2957 2952 5967 2954
rect 2957 2896 2962 2952
rect 3018 2896 5906 2952
rect 5962 2896 5967 2952
rect 2957 2894 5967 2896
rect 2957 2891 3023 2894
rect 5901 2891 5967 2894
rect 13261 2954 13327 2957
rect 22645 2954 22711 2957
rect 13261 2952 22711 2954
rect 13261 2896 13266 2952
rect 13322 2896 22650 2952
rect 22706 2896 22711 2952
rect 13261 2894 22711 2896
rect 13261 2891 13327 2894
rect 22645 2891 22711 2894
rect 62 2682 122 2864
rect 12525 2818 12591 2821
rect 12934 2818 12940 2820
rect 12525 2816 12940 2818
rect 12525 2760 12530 2816
rect 12586 2760 12940 2816
rect 12525 2758 12940 2760
rect 12525 2755 12591 2758
rect 12934 2756 12940 2758
rect 13004 2756 13010 2820
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 2221 2682 2287 2685
rect 62 2680 2287 2682
rect 62 2624 2226 2680
rect 2282 2624 2287 2680
rect 62 2622 2287 2624
rect 2221 2619 2287 2622
rect 4337 2682 4403 2685
rect 9489 2682 9555 2685
rect 4337 2680 9555 2682
rect 4337 2624 4342 2680
rect 4398 2624 9494 2680
rect 9550 2624 9555 2680
rect 4337 2622 9555 2624
rect 4337 2619 4403 2622
rect 9489 2619 9555 2622
rect 12801 2682 12867 2685
rect 19425 2682 19491 2685
rect 12801 2680 19491 2682
rect 12801 2624 12806 2680
rect 12862 2624 19430 2680
rect 19486 2624 19491 2680
rect 12801 2622 19491 2624
rect 12801 2619 12867 2622
rect 19425 2619 19491 2622
rect 13721 2410 13787 2413
rect 23105 2410 23171 2413
rect 13721 2408 23171 2410
rect 13721 2352 13726 2408
rect 13782 2352 23110 2408
rect 23166 2352 23171 2408
rect 13721 2350 23171 2352
rect 13721 2347 13787 2350
rect 23105 2347 23171 2350
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 13721 2002 13787 2005
rect 21449 2002 21515 2005
rect 13721 2000 21515 2002
rect 13721 1944 13726 2000
rect 13782 1944 21454 2000
rect 21510 1944 21515 2000
rect 13721 1942 21515 1944
rect 13721 1939 13787 1942
rect 21449 1939 21515 1942
rect 9765 1866 9831 1869
rect 21081 1866 21147 1869
rect 9765 1864 21147 1866
rect 9765 1808 9770 1864
rect 9826 1808 21086 1864
rect 21142 1808 21147 1864
rect 9765 1806 21147 1808
rect 9765 1803 9831 1806
rect 21081 1803 21147 1806
rect 12893 1730 12959 1733
rect 19793 1730 19859 1733
rect 12893 1728 19859 1730
rect 12893 1672 12898 1728
rect 12954 1672 19798 1728
rect 19854 1672 19859 1728
rect 12893 1670 19859 1672
rect 12893 1667 12959 1670
rect 19793 1667 19859 1670
rect 20897 1730 20963 1733
rect 20897 1728 27722 1730
rect 20897 1672 20902 1728
rect 20958 1672 27722 1728
rect 20897 1670 27722 1672
rect 20897 1667 20963 1670
rect 27662 1352 27722 1670
rect 27520 1232 28000 1352
rect 0 1048 480 1080
rect 0 992 110 1048
rect 166 992 480 1048
rect 0 960 480 992
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 27660 24108 27724 24172
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 27660 23428 27724 23492
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 16252 3028 16316 3092
rect 12940 2756 13004 2820
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 12939 2820 13005 2821
rect 12939 2756 12940 2820
rect 13004 2756 13005 2820
rect 12939 2755 13005 2756
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 12942 1818 13002 2755
rect 14944 2208 15264 3232
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 16251 3092 16317 3093
rect 16251 3028 16252 3092
rect 16316 3028 16317 3092
rect 16251 3027 16317 3028
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 16254 1818 16314 3027
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 27659 24172 27725 24173
rect 27659 24108 27660 24172
rect 27724 24108 27725 24172
rect 27659 24107 27725 24108
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 27662 23493 27722 24107
rect 27659 23492 27725 23493
rect 27659 23428 27660 23492
rect 27724 23428 27725 23492
rect 27659 23427 27725 23428
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 12854 1582 13090 1818
rect 16166 1582 16402 1818
<< metal5 >>
rect 12812 1818 16444 1860
rect 12812 1582 12854 1818
rect 13090 1582 16166 1818
rect 16402 1582 16444 1818
rect 12812 1540 16444 1582
use scs8hd_decap_4  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _176_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 866 592
use scs8hd_inv_8  _177_
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _199_
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_19
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_23
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_36
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_37
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_40
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_41
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_or4_4  _123_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use scs8hd_or4_4  _163_
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__C
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__D
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_68
timestamp 1586364061
transform 1 0 7360 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6992 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7084 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7176 0 1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8740 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_75
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_79
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_94
timestamp 1586364061
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_107
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_117
timestamp 1586364061
transform 1 0 11868 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_111
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_111
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _232_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_136
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _231_
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14536 0 1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_146
timestamp 1586364061
transform 1 0 14536 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_142
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_165
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_157
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_161
timestamp 1586364061
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _228_
timestamp 1586364061
transform 1 0 17020 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17296 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_169
timestamp 1586364061
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_177
timestamp 1586364061
transform 1 0 17388 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_174
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_178
timestamp 1586364061
transform 1 0 17480 0 1 2720
box -38 -48 314 592
use scs8hd_inv_8  _193_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _191_
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _242_
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_197
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_210
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_212
timestamp 1586364061
transform 1 0 20608 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 20424 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_217
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_214
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_216
timestamp 1586364061
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_221
timestamp 1586364061
transform 1 0 21436 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_221
timestamp 1586364061
transform 1 0 21436 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _241_
timestamp 1586364061
transform 1 0 22724 0 -1 2720
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22632 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_225 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21804 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_233
timestamp 1586364061
transform 1 0 22540 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_225
timestamp 1586364061
transform 1 0 21804 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_239
timestamp 1586364061
transform 1 0 23092 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 23276 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_247
timestamp 1586364061
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_243
timestamp 1586364061
transform 1 0 23460 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24012 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_249 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24196 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_1_254
timestamp 1586364061
transform 1 0 24472 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_259
timestamp 1586364061
transform 1 0 24932 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_6  FILLER_1_271 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 26036 0 1 2720
box -38 -48 590 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 1840 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_10
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use scs8hd_or4_4  _166_
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__D
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 4600 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_29
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_36
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_40
timestamp 1586364061
transform 1 0 4784 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 6164 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 4968 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_53
timestamp 1586364061
transform 1 0 5980 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6716 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_57
timestamp 1586364061
transform 1 0 6348 0 -1 3808
box -38 -48 222 592
use scs8hd_conb_1  _223_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__146__C
timestamp 1586364061
transform 1 0 7912 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 8280 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_72
timestamp 1586364061
transform 1 0 7728 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_76
timestamp 1586364061
transform 1 0 8096 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_83
timestamp 1586364061
transform 1 0 8740 0 -1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _119_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9844 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_87
timestamp 1586364061
transform 1 0 9108 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_91
timestamp 1586364061
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_104
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_108
timestamp 1586364061
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11684 0 -1 3808
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_2_112
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_126
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_130
timestamp 1586364061
transform 1 0 13064 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_143
timestamp 1586364061
transform 1 0 14260 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_147
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_151
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_165
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_169
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_182
timestamp 1586364061
transform 1 0 17848 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_12  FILLER_2_199
timestamp 1586364061
transform 1 0 19412 0 -1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_211
timestamp 1586364061
transform 1 0 20516 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_218
timestamp 1586364061
transform 1 0 21160 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_8  _194_
timestamp 1586364061
transform 1 0 22172 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_226
timestamp 1586364061
transform 1 0 21896 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23736 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_238
timestamp 1586364061
transform 1 0 23000 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_2_249
timestamp 1586364061
transform 1 0 24012 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24748 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24564 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_253
timestamp 1586364061
transform 1 0 24380 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_260
timestamp 1586364061
transform 1 0 25024 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_272
timestamp 1586364061
transform 1 0 26128 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_nand2_4  _108_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_or4_4  _130_
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_16
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  FILLER_3_22
timestamp 1586364061
transform 1 0 3128 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_36
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_40
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7452 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7268 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_66
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 8648 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_80
timestamp 1586364061
transform 1 0 8464 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_84
timestamp 1586364061
transform 1 0 8832 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_88
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_99
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_138
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_151
timestamp 1586364061
transform 1 0 14996 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_157
timestamp 1586364061
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16744 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_168
timestamp 1586364061
transform 1 0 16560 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_172
timestamp 1586364061
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_176
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 406 592
use scs8hd_inv_8  _192_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_180
timestamp 1586364061
transform 1 0 17664 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_conb_1  _213_
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_197
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_3_204
timestamp 1586364061
transform 1 0 19872 0 1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_215
timestamp 1586364061
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_219
timestamp 1586364061
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_223
timestamp 1586364061
transform 1 0 21620 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23920 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_236
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_240
timestamp 1586364061
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 1 3808
box -38 -48 866 592
use scs8hd_decap_12  FILLER_3_259
timestamp 1586364061
transform 1 0 24932 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_3_271
timestamp 1586364061
transform 1 0 26036 0 1 3808
box -38 -48 590 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_inv_8  _101_
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_12
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 2760 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_16
timestamp 1586364061
transform 1 0 2576 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4324 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_29
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 314 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 5336 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_48
timestamp 1586364061
transform 1 0 5520 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__D
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_61
timestamp 1586364061
transform 1 0 6716 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_65
timestamp 1586364061
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__D
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_78
timestamp 1586364061
transform 1 0 8280 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_82
timestamp 1586364061
transform 1 0 8648 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 9844 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_86
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_90
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 10212 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_97
timestamp 1586364061
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_101
timestamp 1586364061
transform 1 0 10396 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_113
timestamp 1586364061
transform 1 0 11500 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_121
timestamp 1586364061
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_128
timestamp 1586364061
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_132
timestamp 1586364061
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15364 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 590 592
use scs8hd_inv_8  _182_
timestamp 1586364061
transform 1 0 17112 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 16928 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_8  _179_
timestamp 1586364061
transform 1 0 18676 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 18124 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_183
timestamp 1586364061
transform 1 0 17940 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_187
timestamp 1586364061
transform 1 0 18308 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_200
timestamp 1586364061
transform 1 0 19504 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_212
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22356 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_4  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23920 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_240
timestamp 1586364061
transform 1 0 23184 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_4_257
timestamp 1586364061
transform 1 0 24748 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_4_269
timestamp 1586364061
transform 1 0 25852 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_inv_8  _137_
timestamp 1586364061
transform 1 0 2300 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 1564 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_22
timestamp 1586364061
transform 1 0 3128 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_26
timestamp 1586364061
transform 1 0 3496 0 1 4896
box -38 -48 130 592
use scs8hd_inv_8  _205_
timestamp 1586364061
transform 1 0 3864 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_29
timestamp 1586364061
transform 1 0 3772 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _098_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_43
timestamp 1586364061
transform 1 0 5060 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_47
timestamp 1586364061
transform 1 0 5428 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _114_
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 7268 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_65
timestamp 1586364061
transform 1 0 7084 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_69
timestamp 1586364061
transform 1 0 7452 0 1 4896
box -38 -48 222 592
use scs8hd_or4_4  _149_
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_82
timestamp 1586364061
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use scs8hd_or2_4  _099_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__C
timestamp 1586364061
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__D
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_97
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_101
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_130
timestamp 1586364061
transform 1 0 13064 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_134
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 14812 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_151
timestamp 1586364061
transform 1 0 14996 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15364 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_166
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16560 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_170
timestamp 1586364061
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_174
timestamp 1586364061
transform 1 0 17112 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _178_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 774 592
use scs8hd_conb_1  _224_
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_204
timestamp 1586364061
transform 1 0 19872 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_216
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 1142 592
use scs8hd_conb_1  _214_
timestamp 1586364061
transform 1 0 22264 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_228
timestamp 1586364061
transform 1 0 22080 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_233
timestamp 1586364061
transform 1 0 22540 0 1 4896
box -38 -48 406 592
use scs8hd_inv_8  _195_
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_237
timestamp 1586364061
transform 1 0 22908 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_265
timestamp 1586364061
transform 1 0 25484 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_6
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_1  _103_
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_13
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_10
timestamp 1586364061
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 1 5984
box -38 -48 866 592
use scs8hd_nor3_4  _169_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3036 0 1 5984
box -38 -48 1234 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__C
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_17
timestamp 1586364061
transform 1 0 2668 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_34
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_38
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 406 592
use scs8hd_or4_4  _160_
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__160__D
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 6072 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__C
timestamp 1586364061
transform 1 0 5704 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_43
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_47
timestamp 1586364061
transform 1 0 5428 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_52
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_60
timestamp 1586364061
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 6440 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_buf_1  _139_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_65
timestamp 1586364061
transform 1 0 7084 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_69
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_65
timestamp 1586364061
transform 1 0 7084 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__D
timestamp 1586364061
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 866 592
use scs8hd_or4_4  _143_
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 866 592
use scs8hd_or4_4  _146_
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__D
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_82
timestamp 1586364061
transform 1 0 8648 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_88
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_84
timestamp 1586364061
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_86
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__D
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_or4_4  _118_
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_or4_4  _115_
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 866 592
use scs8hd_buf_1  _097_
timestamp 1586364061
transform 1 0 11132 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_107
timestamp 1586364061
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_101
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_105
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_116
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_112
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_111
timestamp 1586364061
transform 1 0 11316 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_121
timestamp 1586364061
transform 1 0 12236 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1050 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 11408 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_125
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_133
timestamp 1586364061
transform 1 0 13340 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_134
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_142
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14812 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 1050 592
use scs8hd_buf_2  _229_
timestamp 1586364061
transform 1 0 15364 0 -1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__126__D
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15916 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_159
timestamp 1586364061
transform 1 0 15732 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_162
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_166
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__C
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_176
timestamp 1586364061
transform 1 0 17296 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_173
timestamp 1586364061
transform 1 0 17020 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_177
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 406 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_180
timestamp 1586364061
transform 1 0 17664 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_193
timestamp 1586364061
transform 1 0 18860 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_205
timestamp 1586364061
transform 1 0 19964 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_197
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_201
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_213
timestamp 1586364061
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_213
timestamp 1586364061
transform 1 0 20700 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_235
timestamp 1586364061
transform 1 0 22724 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_225
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23000 0 -1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24012 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23920 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_241
timestamp 1586364061
transform 1 0 23276 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_4  FILLER_7_237
timestamp 1586364061
transform 1 0 22908 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_241
timestamp 1586364061
transform 1 0 23276 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25116 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_258
timestamp 1586364061
transform 1 0 24840 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_259
timestamp 1586364061
transform 1 0 24932 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_270
timestamp 1586364061
transform 1 0 25944 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_274
timestamp 1586364061
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_263
timestamp 1586364061
transform 1 0 25300 0 1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_275
timestamp 1586364061
transform 1 0 26404 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_inv_8  _207_
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_8_12
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 406 592
use scs8hd_buf_1  _167_
timestamp 1586364061
transform 1 0 2944 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 2668 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__C
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_16
timestamp 1586364061
transform 1 0 2576 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_19
timestamp 1586364061
transform 1 0 2852 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_nand2_4  _138_
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__C
timestamp 1586364061
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 5888 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_46
timestamp 1586364061
transform 1 0 5336 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_50
timestamp 1586364061
transform 1 0 5704 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_54
timestamp 1586364061
transform 1 0 6072 0 -1 7072
box -38 -48 222 592
use scs8hd_or4_4  _157_
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_67
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 314 592
use scs8hd_or4_4  _140_
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__D
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_72
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 314 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__D
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__143__C
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_106
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12236 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 11684 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_113
timestamp 1586364061
transform 1 0 11500 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_132
timestamp 1586364061
transform 1 0 13248 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_136
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 222 592
use scs8hd_conb_1  _218_
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_140
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_163
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use scs8hd_or4_4  _126_
timestamp 1586364061
transform 1 0 16836 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16652 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_167
timestamp 1586364061
transform 1 0 16468 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 18400 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_180
timestamp 1586364061
transform 1 0 17664 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_186
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_197
timestamp 1586364061
transform 1 0 19228 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_209
timestamp 1586364061
transform 1 0 20332 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_inv_8  _183_
timestamp 1586364061
transform 1 0 23644 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_6  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_8_254
timestamp 1586364061
transform 1 0 24472 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_266
timestamp 1586364061
transform 1 0 25576 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_274
timestamp 1586364061
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_buf_1  _109_
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_9
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_13
timestamp 1586364061
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use scs8hd_nor3_4  _171_
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_30
timestamp 1586364061
transform 1 0 3864 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_34
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_38
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 406 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _122_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_65
timestamp 1586364061
transform 1 0 7084 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_69
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 130 592
use scs8hd_or4_4  _134_
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 7544 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_72
timestamp 1586364061
transform 1 0 7728 0 1 7072
box -38 -48 314 592
use scs8hd_or4_4  _104_
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_84
timestamp 1586364061
transform 1 0 8832 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_88
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__D
timestamp 1586364061
transform 1 0 10948 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_101
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_105
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_109
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _208_
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 11868 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_119
timestamp 1586364061
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 12604 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_127
timestamp 1586364061
transform 1 0 12788 0 1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14996 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_141
timestamp 1586364061
transform 1 0 14076 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_145
timestamp 1586364061
transform 1 0 14444 0 1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_154
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_158
timestamp 1586364061
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _190_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_205
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_217
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_229
timestamp 1586364061
transform 1 0 22172 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_241
timestamp 1586364061
transform 1 0 23276 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_253
timestamp 1586364061
transform 1 0 24380 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_262
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_9_274
timestamp 1586364061
transform 1 0 26312 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1472 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 2852 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_21
timestamp 1586364061
transform 1 0 3036 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_25
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_nor3_4  _168_
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_29
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_8  _121_
timestamp 1586364061
transform 1 0 5980 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 5796 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_45
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_49
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__D
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__D
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_62
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_66
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use scs8hd_or4_4  _153_
timestamp 1586364061
transform 1 0 7544 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__C
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_79
timestamp 1586364061
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_83
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 8924 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 9292 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_87
timestamp 1586364061
transform 1 0 9108 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 11040 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_106
timestamp 1586364061
transform 1 0 10856 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_110
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 590 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 866 592
use scs8hd_fill_1  FILLER_10_116
timestamp 1586364061
transform 1 0 11776 0 -1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 13524 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_126
timestamp 1586364061
transform 1 0 12696 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_132
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_144
timestamp 1586364061
transform 1 0 14352 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_152
timestamp 1586364061
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_165
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 774 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 17020 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_12  FILLER_10_182
timestamp 1586364061
transform 1 0 17848 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_194
timestamp 1586364061
transform 1 0 18952 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_or2_4  _102_
timestamp 1586364061
transform 1 0 1472 0 1 8160
box -38 -48 682 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_11
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use scs8hd_nor3_4  _170_
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_32
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_36
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_40
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_or4_4  _110_
timestamp 1586364061
transform 1 0 7452 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_66
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_78
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_83
timestamp 1586364061
transform 1 0 8740 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 8924 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_87
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_91
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_106
timestamp 1586364061
transform 1 0 10856 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 13340 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 13156 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_127
timestamp 1586364061
transform 1 0 12788 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_142
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_148
timestamp 1586364061
transform 1 0 14720 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_152
timestamp 1586364061
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_156
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_167
timestamp 1586364061
transform 1 0 16468 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 774 592
use scs8hd_conb_1  _219_
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 18584 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_187
timestamp 1586364061
transform 1 0 18308 0 1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_11_192
timestamp 1586364061
transform 1 0 18768 0 1 8160
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19320 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19780 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_201
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_205
timestamp 1586364061
transform 1 0 19964 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_217
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_229
timestamp 1586364061
transform 1 0 22172 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_11_241
timestamp 1586364061
transform 1 0 23276 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1932 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_11
timestamp 1586364061
transform 1 0 2116 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4508 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_35
timestamp 1586364061
transform 1 0 4324 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_39
timestamp 1586364061
transform 1 0 4692 0 -1 9248
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5244 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_60
timestamp 1586364061
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  _129_
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_73
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_77
timestamp 1586364061
transform 1 0 8188 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  _132_
timestamp 1586364061
transform 1 0 9844 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 10304 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_98
timestamp 1586364061
transform 1 0 10120 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12236 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_115
timestamp 1586364061
transform 1 0 11684 0 -1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_132
timestamp 1586364061
transform 1 0 13248 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_136
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_144
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_150
timestamp 1586364061
transform 1 0 14904 0 -1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_165
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_8  _184_
timestamp 1586364061
transform 1 0 17020 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 16468 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_169
timestamp 1586364061
transform 1 0 16652 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_8  _189_
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_182
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_189
timestamp 1586364061
transform 1 0 18492 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_199
timestamp 1586364061
transform 1 0 19412 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_211
timestamp 1586364061
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use scs8hd_conb_1  _212_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_6
timestamp 1586364061
transform 1 0 1656 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_10
timestamp 1586364061
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_10
timestamp 1586364061
transform 1 0 2024 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_8  _206_
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_23
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_40
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_43
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_48
timestamp 1586364061
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_44
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_47
timestamp 1586364061
transform 1 0 5428 0 -1 10336
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_59
timestamp 1586364061
transform 1 0 6532 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_73
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_73
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_77
timestamp 1586364061
transform 1 0 8188 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_77
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8280 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _152_
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 314 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_8  _095_
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 9384 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_84
timestamp 1586364061
transform 1 0 8832 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_88
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_8  _202_
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 866 592
use scs8hd_conb_1  _216_
timestamp 1586364061
transform 1 0 11132 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_101
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_105
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_106
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_112
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_116
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 406 592
use scs8hd_decap_6  FILLER_14_119
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_134
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_138
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_127
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_138
timestamp 1586364061
transform 1 0 13800 0 -1 10336
box -38 -48 590 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_151
timestamp 1586364061
transform 1 0 14996 0 1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_144
timestamp 1586364061
transform 1 0 14352 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_147
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_156
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_14_165
timestamp 1586364061
transform 1 0 16284 0 -1 10336
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17296 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_168
timestamp 1586364061
transform 1 0 16560 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_172
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_13_178
timestamp 1586364061
transform 1 0 17480 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_173
timestamp 1586364061
transform 1 0 17020 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_179
timestamp 1586364061
transform 1 0 17572 0 -1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19504 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_198
timestamp 1586364061
transform 1 0 19320 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_202
timestamp 1586364061
transform 1 0 19688 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_196
timestamp 1586364061
transform 1 0 19136 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_214
timestamp 1586364061
transform 1 0 20792 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_14_208
timestamp 1586364061
transform 1 0 20240 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_226
timestamp 1586364061
transform 1 0 21896 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_238
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_249
timestamp 1586364061
transform 1 0 24012 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_243
timestamp 1586364061
transform 1 0 23460 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_247
timestamp 1586364061
transform 1 0 23828 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_261
timestamp 1586364061
transform 1 0 25116 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_259
timestamp 1586364061
transform 1 0 24932 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_273
timestamp 1586364061
transform 1 0 26220 0 1 9248
box -38 -48 406 592
use scs8hd_decap_4  FILLER_14_271
timestamp 1586364061
transform 1 0 26036 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_conb_1  _211_
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_14
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_18
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_22
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_26
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_30
timestamp 1586364061
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_34
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5888 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_47
timestamp 1586364061
transform 1 0 5428 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_54
timestamp 1586364061
transform 1 0 6072 0 1 10336
box -38 -48 222 592
use scs8hd_conb_1  _210_
timestamp 1586364061
transform 1 0 7084 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_58
timestamp 1586364061
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_68
timestamp 1586364061
transform 1 0 7360 0 1 10336
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8280 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8096 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7728 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_89
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_93
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_108
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_112
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_134
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_138
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14444 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_142
timestamp 1586364061
transform 1 0 14168 0 1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_156
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_160
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _187_
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_205
timestamp 1586364061
transform 1 0 19964 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_217
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_229
timestamp 1586364061
transform 1 0 22172 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_241
timestamp 1586364061
transform 1 0 23276 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 774 592
use scs8hd_buf_2  _240_
timestamp 1586364061
transform 1 0 24564 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 25116 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_253
timestamp 1586364061
transform 1 0 24380 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_259
timestamp 1586364061
transform 1 0 24932 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_263
timestamp 1586364061
transform 1 0 25300 0 1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_15_275
timestamp 1586364061
transform 1 0 26404 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_10
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _164_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_8  _204_
timestamp 1586364061
transform 1 0 4324 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5888 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_48
timestamp 1586364061
transform 1 0 5520 0 -1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_61
timestamp 1586364061
transform 1 0 6716 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_4  FILLER_16_69
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 9936 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_88
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 -1 11424
box -38 -48 866 592
use scs8hd_fill_1  FILLER_16_98
timestamp 1586364061
transform 1 0 10120 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_108
timestamp 1586364061
transform 1 0 11040 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_8  _198_
timestamp 1586364061
transform 1 0 11776 0 -1 11424
box -38 -48 866 592
use scs8hd_inv_8  _188_
timestamp 1586364061
transform 1 0 13340 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_8  FILLER_16_142
timestamp 1586364061
transform 1 0 14168 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_150
timestamp 1586364061
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  FILLER_16_168
timestamp 1586364061
transform 1 0 16560 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_180
timestamp 1586364061
transform 1 0 17664 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_192
timestamp 1586364061
transform 1 0 18768 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_204
timestamp 1586364061
transform 1 0 19872 0 -1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_212
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_12
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_16
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4508 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_29
timestamp 1586364061
transform 1 0 3772 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_34
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_46
timestamp 1586364061
transform 1 0 5336 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_50
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_76
timestamp 1586364061
transform 1 0 8096 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_80
timestamp 1586364061
transform 1 0 8464 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 866 592
use scs8hd_fill_2  FILLER_17_84
timestamp 1586364061
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_95
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_99
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _196_
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_112
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_116
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 774 592
use scs8hd_conb_1  _220_
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 14904 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_140
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_143
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_148
timestamp 1586364061
transform 1 0 14720 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_152
timestamp 1586364061
transform 1 0 15088 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_165
timestamp 1586364061
transform 1 0 16284 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_169
timestamp 1586364061
transform 1 0 16652 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_181
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_248
timestamp 1586364061
transform 1 0 23920 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 24564 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_252
timestamp 1586364061
transform 1 0 24288 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_7
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_11
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 5796 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_43
timestamp 1586364061
transform 1 0 5060 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_47
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_50
timestamp 1586364061
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_60
timestamp 1586364061
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 774 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 7820 0 -1 12512
box -38 -48 866 592
use scs8hd_fill_1  FILLER_18_72
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_82
timestamp 1586364061
transform 1 0 8648 0 -1 12512
box -38 -48 406 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 9936 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_109
timestamp 1586364061
transform 1 0 11132 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_8  _197_
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11316 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_122
timestamp 1586364061
transform 1 0 12328 0 -1 12512
box -38 -48 774 592
use scs8hd_conb_1  _221_
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_133
timestamp 1586364061
transform 1 0 13340 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_144
timestamp 1586364061
transform 1 0 14352 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_152
timestamp 1586364061
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use scs8hd_inv_8  _186_
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_175
timestamp 1586364061
transform 1 0 17204 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_187
timestamp 1586364061
transform 1 0 18308 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_199
timestamp 1586364061
transform 1 0 19412 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_211
timestamp 1586364061
transform 1 0 20516 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_buf_2  _239_
timestamp 1586364061
transform 1 0 24564 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_4  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_259
timestamp 1586364061
transform 1 0 24932 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_271
timestamp 1586364061
transform 1 0 26036 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_6
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 1564 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_10
timestamp 1586364061
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_8  _175_
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 3312 0 1 12512
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 3128 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_16
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_20
timestamp 1586364061
transform 1 0 2944 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 774 592
use scs8hd_conb_1  _222_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_35
timestamp 1586364061
transform 1 0 4324 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_35
timestamp 1586364061
transform 1 0 4324 0 -1 13600
box -38 -48 774 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5520 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_43
timestamp 1586364061
transform 1 0 5060 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_46
timestamp 1586364061
transform 1 0 5336 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_59
timestamp 1586364061
transform 1 0 6532 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_67
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7544 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_75
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_79
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_81
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 774 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9292 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_90
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_91
timestamp 1586364061
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11224 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_103
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_107
timestamp 1586364061
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 406 592
use scs8hd_conb_1  _215_
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_121
timestamp 1586364061
transform 1 0 12236 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_8  _185_
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13156 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_126
timestamp 1586364061
transform 1 0 12696 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_130
timestamp 1586364061
transform 1 0 13064 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_133
timestamp 1586364061
transform 1 0 13340 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_137
timestamp 1586364061
transform 1 0 13708 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_133
timestamp 1586364061
transform 1 0 13340 0 -1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14076 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13892 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_152
timestamp 1586364061
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16284 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_156
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_163
timestamp 1586364061
transform 1 0 16100 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_163
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_167
timestamp 1586364061
transform 1 0 16468 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_175
timestamp 1586364061
transform 1 0 17204 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_263
timestamp 1586364061
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_buf_2  _233_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_11
timestamp 1586364061
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use scs8hd_inv_8  _174_
timestamp 1586364061
transform 1 0 2944 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_29
timestamp 1586364061
transform 1 0 3772 0 1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_21_41
timestamp 1586364061
transform 1 0 4876 0 1 13600
box -38 -48 130 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7360 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_66
timestamp 1586364061
transform 1 0 7176 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7544 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_81
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9292 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 9752 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_85
timestamp 1586364061
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_92
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_96
timestamp 1586364061
transform 1 0 9936 0 1 13600
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10488 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_21_113
timestamp 1586364061
transform 1 0 11500 0 1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_21_121
timestamp 1586364061
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_126
timestamp 1586364061
transform 1 0 12696 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_130
timestamp 1586364061
transform 1 0 13064 0 1 13600
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_142
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_156
timestamp 1586364061
transform 1 0 15456 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_168
timestamp 1586364061
transform 1 0 16560 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_21_180
timestamp 1586364061
transform 1 0 17664 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_253
timestamp 1586364061
transform 1 0 24380 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_buf_2  _230_
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_19
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_22_40
timestamp 1586364061
transform 1 0 4784 0 -1 14688
box -38 -48 314 592
use scs8hd_conb_1  _225_
timestamp 1586364061
transform 1 0 5060 0 -1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6072 0 -1 14688
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_22_46
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_6  FILLER_22_65
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_82
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_90
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_102
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_114
timestamp 1586364061
transform 1 0 11592 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_126
timestamp 1586364061
transform 1 0 12696 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_138
timestamp 1586364061
transform 1 0 13800 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_22_150
timestamp 1586364061
transform 1 0 14904 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_178
timestamp 1586364061
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_190
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_202
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_258
timestamp 1586364061
transform 1 0 24840 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_270
timestamp 1586364061
transform 1 0 25944 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_274
timestamp 1586364061
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 6072 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_47
timestamp 1586364061
transform 1 0 5428 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_52
timestamp 1586364061
transform 1 0 5888 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6440 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_56
timestamp 1586364061
transform 1 0 6256 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_60
timestamp 1586364061
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_66
timestamp 1586364061
transform 1 0 7176 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_70
timestamp 1586364061
transform 1 0 7544 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_80
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use scs8hd_inv_8  _180_
timestamp 1586364061
transform 1 0 9200 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_84
timestamp 1586364061
transform 1 0 8832 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_97
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_109
timestamp 1586364061
transform 1 0 11132 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_23_121
timestamp 1586364061
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 406 592
use scs8hd_buf_2  _227_
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_139
timestamp 1586364061
transform 1 0 13892 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_144
timestamp 1586364061
transform 1 0 14352 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_148
timestamp 1586364061
transform 1 0 14720 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_160
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_172
timestamp 1586364061
transform 1 0 16928 0 1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_23_180
timestamp 1586364061
transform 1 0 17664 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_232
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 774 592
use scs8hd_buf_2  _236_
timestamp 1586364061
transform 1 0 24564 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 25116 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_253
timestamp 1586364061
transform 1 0 24380 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_259
timestamp 1586364061
transform 1 0 24932 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_263
timestamp 1586364061
transform 1 0 25300 0 1 14688
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_23_275
timestamp 1586364061
transform 1 0 26404 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_inv_8  _203_
timestamp 1586364061
transform 1 0 5796 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_6  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_50
timestamp 1586364061
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_60
timestamp 1586364061
transform 1 0 6624 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_64
timestamp 1586364061
transform 1 0 6992 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_67
timestamp 1586364061
transform 1 0 7268 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_77
timestamp 1586364061
transform 1 0 8188 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_81
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_89
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_178
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7084 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_68
timestamp 1586364061
transform 1 0 7360 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8096 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 7544 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_72
timestamp 1586364061
transform 1 0 7728 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_85
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_97
timestamp 1586364061
transform 1 0 10028 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_109
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_121
timestamp 1586364061
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_147
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_171
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_220
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_253
timestamp 1586364061
transform 1 0 24380 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_258
timestamp 1586364061
transform 1 0 24840 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_262
timestamp 1586364061
transform 1 0 25208 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_25_274
timestamp 1586364061
transform 1 0 26312 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6348 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_60
timestamp 1586364061
transform 1 0 6624 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_inv_8  _181_
timestamp 1586364061
transform 1 0 7544 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_12  FILLER_26_79
timestamp 1586364061
transform 1 0 8372 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_91
timestamp 1586364061
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_27_110
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_117
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_113
timestamp 1586364061
transform 1 0 11500 0 1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_121
timestamp 1586364061
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 24564 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_253
timestamp 1586364061
transform 1 0 24380 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 590 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 11316 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_115
timestamp 1586364061
transform 1 0 11684 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_127
timestamp 1586364061
transform 1 0 12788 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_139
timestamp 1586364061
transform 1 0 13892 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_28_151
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_buf_2  _235_
timestamp 1586364061
transform 1 0 24564 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_4  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_259
timestamp 1586364061
transform 1 0 24932 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_271
timestamp 1586364061
transform 1 0 26036 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 12604 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_127
timestamp 1586364061
transform 1 0 12788 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_139
timestamp 1586364061
transform 1 0 13892 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_151
timestamp 1586364061
transform 1 0 14996 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_163
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_8  _173_
timestamp 1586364061
transform 1 0 12328 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_4  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_121
timestamp 1586364061
transform 1 0 12236 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_131
timestamp 1586364061
transform 1 0 13156 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_135
timestamp 1586364061
transform 1 0 13524 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_32_147
timestamp 1586364061
transform 1 0 14628 0 -1 20128
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_33_106
timestamp 1586364061
transform 1 0 10856 0 1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_109
timestamp 1586364061
transform 1 0 11132 0 -1 21216
box -38 -48 130 592
use scs8hd_conb_1  _217_
timestamp 1586364061
transform 1 0 11316 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_114
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_119
timestamp 1586364061
transform 1 0 12052 0 -1 21216
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_134
timestamp 1586364061
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_138
timestamp 1586364061
transform 1 0 13800 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_136
timestamp 1586364061
transform 1 0 13616 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_150
timestamp 1586364061
transform 1 0 14904 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_148
timestamp 1586364061
transform 1 0 14720 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_152
timestamp 1586364061
transform 1 0 15088 0 -1 21216
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_162
timestamp 1586364061
transform 1 0 16008 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_174
timestamp 1586364061
transform 1 0 17112 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_182
timestamp 1586364061
transform 1 0 17848 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_253
timestamp 1586364061
transform 1 0 24380 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_258
timestamp 1586364061
transform 1 0 24840 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_4  FILLER_34_270
timestamp 1586364061
transform 1 0 25944 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_274
timestamp 1586364061
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_6
timestamp 1586364061
transform 1 0 1656 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_10
timestamp 1586364061
transform 1 0 2024 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_22
timestamp 1586364061
transform 1 0 3128 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_34
timestamp 1586364061
transform 1 0 4232 0 1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_46
timestamp 1586364061
transform 1 0 5336 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_50
timestamp 1586364061
transform 1 0 5704 0 1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 7360 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_70
timestamp 1586364061
transform 1 0 7544 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_82
timestamp 1586364061
transform 1 0 8648 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_94
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 774 592
use scs8hd_inv_8  _172_
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 10580 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_102
timestamp 1586364061
transform 1 0 10488 0 1 21216
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_114
timestamp 1586364061
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13708 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_132
timestamp 1586364061
transform 1 0 13248 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_136
timestamp 1586364061
transform 1 0 13616 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_139
timestamp 1586364061
transform 1 0 13892 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_151
timestamp 1586364061
transform 1 0 14996 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_163
timestamp 1586364061
transform 1 0 16100 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_175
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_inv_8  _201_
timestamp 1586364061
transform 1 0 5796 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_6  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_50
timestamp 1586364061
transform 1 0 5704 0 -1 22304
box -38 -48 130 592
use scs8hd_inv_8  _200_
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_60
timestamp 1586364061
transform 1 0 6624 0 -1 22304
box -38 -48 590 592
use scs8hd_decap_12  FILLER_36_77
timestamp 1586364061
transform 1 0 8188 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_36_89
timestamp 1586364061
transform 1 0 9292 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_114
timestamp 1586364061
transform 1 0 11592 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_36_122
timestamp 1586364061
transform 1 0 12328 0 -1 22304
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13708 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_140
timestamp 1586364061
transform 1 0 13984 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_152
timestamp 1586364061
transform 1 0 15088 0 -1 22304
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_19
timestamp 1586364061
transform 1 0 2852 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_31
timestamp 1586364061
transform 1 0 3956 0 1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5244 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_43
timestamp 1586364061
transform 1 0 5060 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_47
timestamp 1586364061
transform 1 0 5428 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_54
timestamp 1586364061
transform 1 0 6072 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6256 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_58
timestamp 1586364061
transform 1 0 6440 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8740 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_75
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_79
timestamp 1586364061
transform 1 0 8372 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9200 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_90
timestamp 1586364061
transform 1 0 9384 0 1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 10856 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_102
timestamp 1586364061
transform 1 0 10488 0 1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_37_108
timestamp 1586364061
transform 1 0 11040 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_120
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_153
timestamp 1586364061
transform 1 0 15180 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_156
timestamp 1586364061
transform 1 0 15456 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_168
timestamp 1586364061
transform 1 0 16560 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_180
timestamp 1586364061
transform 1 0 17664 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_6
timestamp 1586364061
transform 1 0 1656 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_18
timestamp 1586364061
transform 1 0 2760 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_30
timestamp 1586364061
transform 1 0 3864 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5244 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_48
timestamp 1586364061
transform 1 0 5520 0 -1 23392
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_8  FILLER_38_65
timestamp 1586364061
transform 1 0 7084 0 -1 23392
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_8  FILLER_38_82
timestamp 1586364061
transform 1 0 8648 0 -1 23392
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_90
timestamp 1586364061
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_2  _234_
timestamp 1586364061
transform 1 0 10856 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_110
timestamp 1586364061
transform 1 0 11224 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_122
timestamp 1586364061
transform 1 0 12328 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_134
timestamp 1586364061
transform 1 0 13432 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_38_146
timestamp 1586364061
transform 1 0 14536 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_38_152
timestamp 1586364061
transform 1 0 15088 0 -1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_157
timestamp 1586364061
transform 1 0 15548 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_169
timestamp 1586364061
transform 1 0 16652 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_181
timestamp 1586364061
transform 1 0 17756 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_193
timestamp 1586364061
transform 1 0 18860 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_205
timestamp 1586364061
transform 1 0 19964 0 -1 23392
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_213
timestamp 1586364061
transform 1 0 20700 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_22
timestamp 1586364061
transform 1 0 3128 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4784 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_6  FILLER_39_34
timestamp 1586364061
transform 1 0 4232 0 1 23392
box -38 -48 590 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5244 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_43
timestamp 1586364061
transform 1 0 5060 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_47
timestamp 1586364061
transform 1 0 5428 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_53
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_40_50
timestamp 1586364061
transform 1 0 5704 0 -1 24480
box -38 -48 130 592
use scs8hd_conb_1  _209_
timestamp 1586364061
transform 1 0 6992 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_57
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_67
timestamp 1586364061
transform 1 0 7268 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_60
timestamp 1586364061
transform 1 0 6624 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_79
timestamp 1586364061
transform 1 0 8372 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_72
timestamp 1586364061
transform 1 0 7728 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_84
timestamp 1586364061
transform 1 0 8832 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_88
timestamp 1586364061
transform 1 0 9200 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_84
timestamp 1586364061
transform 1 0 8832 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_100
timestamp 1586364061
transform 1 0 10304 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_112
timestamp 1586364061
transform 1 0 11408 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_120
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_138
timestamp 1586364061
transform 1 0 13800 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_142
timestamp 1586364061
transform 1 0 14168 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _243_
timestamp 1586364061
transform 1 0 16008 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_154
timestamp 1586364061
transform 1 0 15272 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_166
timestamp 1586364061
transform 1 0 16376 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 16560 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_170
timestamp 1586364061
transform 1 0 16744 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _238_
timestamp 1586364061
transform 1 0 18308 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 18860 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_182
timestamp 1586364061
transform 1 0 17848 0 1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_191
timestamp 1586364061
transform 1 0 18676 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19872 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_195
timestamp 1586364061
transform 1 0 19044 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_202
timestamp 1586364061
transform 1 0 19688 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_206
timestamp 1586364061
transform 1 0 20056 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _237_
timestamp 1586364061
transform 1 0 20424 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 20976 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_214
timestamp 1586364061
transform 1 0 20792 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_218
timestamp 1586364061
transform 1 0 21160 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_230
timestamp 1586364061
transform 1 0 22264 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_242
timestamp 1586364061
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_253
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_258
timestamp 1586364061
transform 1 0 24840 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_262
timestamp 1586364061
transform 1 0 25208 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_274
timestamp 1586364061
transform 1 0 26312 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
<< labels >>
rlabel metal2 s 1030 27520 1086 28000 6 address[0]
port 0 nsew default input
rlabel metal2 s 2870 0 2926 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 3146 27520 3202 28000 6 address[2]
port 2 nsew default input
rlabel metal2 s 4066 0 4122 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 5170 0 5226 480 6 address[4]
port 4 nsew default input
rlabel metal3 s 0 960 480 1080 6 address[5]
port 5 nsew default input
rlabel metal2 s 7562 0 7618 480 6 bottom_left_grid_pin_11_
port 6 nsew default input
rlabel metal2 s 8666 0 8722 480 6 bottom_left_grid_pin_13_
port 7 nsew default input
rlabel metal3 s 0 4904 480 5024 6 bottom_left_grid_pin_15_
port 8 nsew default input
rlabel metal3 s 27520 1232 28000 1352 6 bottom_left_grid_pin_1_
port 9 nsew default input
rlabel metal3 s 27520 3680 28000 3800 6 bottom_left_grid_pin_3_
port 10 nsew default input
rlabel metal2 s 6366 0 6422 480 6 bottom_left_grid_pin_5_
port 11 nsew default input
rlabel metal3 s 0 2864 480 2984 6 bottom_left_grid_pin_7_
port 12 nsew default input
rlabel metal2 s 5262 27520 5318 28000 6 bottom_left_grid_pin_9_
port 13 nsew default input
rlabel metal2 s 9862 0 9918 480 6 bottom_right_grid_pin_11_
port 14 nsew default input
rlabel metal3 s 0 6944 480 7064 6 chanx_right_in[0]
port 15 nsew default input
rlabel metal3 s 0 8848 480 8968 6 chanx_right_in[1]
port 16 nsew default input
rlabel metal2 s 7470 27520 7526 28000 6 chanx_right_in[2]
port 17 nsew default input
rlabel metal2 s 11058 0 11114 480 6 chanx_right_in[3]
port 18 nsew default input
rlabel metal2 s 9586 27520 9642 28000 6 chanx_right_in[4]
port 19 nsew default input
rlabel metal3 s 27520 6264 28000 6384 6 chanx_right_in[5]
port 20 nsew default input
rlabel metal2 s 12162 0 12218 480 6 chanx_right_in[6]
port 21 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chanx_right_in[7]
port 22 nsew default input
rlabel metal3 s 0 10888 480 11008 6 chanx_right_in[8]
port 23 nsew default input
rlabel metal2 s 11702 27520 11758 28000 6 chanx_right_out[0]
port 24 nsew default tristate
rlabel metal3 s 0 12928 480 13048 6 chanx_right_out[1]
port 25 nsew default tristate
rlabel metal2 s 14554 0 14610 480 6 chanx_right_out[2]
port 26 nsew default tristate
rlabel metal2 s 15658 0 15714 480 6 chanx_right_out[3]
port 27 nsew default tristate
rlabel metal3 s 0 14968 480 15088 6 chanx_right_out[4]
port 28 nsew default tristate
rlabel metal2 s 16854 0 16910 480 6 chanx_right_out[5]
port 29 nsew default tristate
rlabel metal2 s 18050 0 18106 480 6 chanx_right_out[6]
port 30 nsew default tristate
rlabel metal3 s 0 16872 480 16992 6 chanx_right_out[7]
port 31 nsew default tristate
rlabel metal3 s 0 18912 480 19032 6 chanx_right_out[8]
port 32 nsew default tristate
rlabel metal2 s 19154 0 19210 480 6 chany_bottom_in[0]
port 33 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chany_bottom_in[1]
port 34 nsew default input
rlabel metal3 s 27520 8848 28000 8968 6 chany_bottom_in[2]
port 35 nsew default input
rlabel metal3 s 0 20952 480 21072 6 chany_bottom_in[3]
port 36 nsew default input
rlabel metal3 s 0 22856 480 22976 6 chany_bottom_in[4]
port 37 nsew default input
rlabel metal2 s 20350 0 20406 480 6 chany_bottom_in[5]
port 38 nsew default input
rlabel metal3 s 0 24896 480 25016 6 chany_bottom_in[6]
port 39 nsew default input
rlabel metal2 s 16026 27520 16082 28000 6 chany_bottom_in[7]
port 40 nsew default input
rlabel metal2 s 21546 0 21602 480 6 chany_bottom_in[8]
port 41 nsew default input
rlabel metal2 s 18234 27520 18290 28000 6 chany_bottom_out[0]
port 42 nsew default tristate
rlabel metal2 s 22650 0 22706 480 6 chany_bottom_out[1]
port 43 nsew default tristate
rlabel metal2 s 23846 0 23902 480 6 chany_bottom_out[2]
port 44 nsew default tristate
rlabel metal3 s 27520 11296 28000 11416 6 chany_bottom_out[3]
port 45 nsew default tristate
rlabel metal3 s 27520 13880 28000 14000 6 chany_bottom_out[4]
port 46 nsew default tristate
rlabel metal2 s 20350 27520 20406 28000 6 chany_bottom_out[5]
port 47 nsew default tristate
rlabel metal2 s 22466 27520 22522 28000 6 chany_bottom_out[6]
port 48 nsew default tristate
rlabel metal3 s 27520 16464 28000 16584 6 chany_bottom_out[7]
port 49 nsew default tristate
rlabel metal3 s 27520 19048 28000 19168 6 chany_bottom_out[8]
port 50 nsew default tristate
rlabel metal2 s 1674 0 1730 480 6 data_in
port 51 nsew default input
rlabel metal2 s 570 0 626 480 6 enable
port 52 nsew default input
rlabel metal2 s 24674 27520 24730 28000 6 right_bottom_grid_pin_12_
port 53 nsew default input
rlabel metal2 s 27342 0 27398 480 6 right_top_grid_pin_11_
port 54 nsew default input
rlabel metal3 s 27520 24080 28000 24200 6 right_top_grid_pin_13_
port 55 nsew default input
rlabel metal3 s 27520 26664 28000 26784 6 right_top_grid_pin_15_
port 56 nsew default input
rlabel metal3 s 27520 21496 28000 21616 6 right_top_grid_pin_1_
port 57 nsew default input
rlabel metal2 s 25042 0 25098 480 6 right_top_grid_pin_3_
port 58 nsew default input
rlabel metal3 s 0 26936 480 27056 6 right_top_grid_pin_5_
port 59 nsew default input
rlabel metal2 s 26146 0 26202 480 6 right_top_grid_pin_7_
port 60 nsew default input
rlabel metal2 s 26790 27520 26846 28000 6 right_top_grid_pin_9_
port 61 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 62 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 63 nsew default input
<< end >>
