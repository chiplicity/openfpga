* NGSPICE file created from grid_io_left.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_1 abstract view
.subckt scs8hd_ebufn_1 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_and4_4 abstract view
.subckt scs8hd_and4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

.subckt grid_io_left address[0] address[1] address[2] address[3] data_in enable gfpga_pad_GPIO_PAD[0]
+ gfpga_pad_GPIO_PAD[1] gfpga_pad_GPIO_PAD[2] gfpga_pad_GPIO_PAD[3] gfpga_pad_GPIO_PAD[4]
+ gfpga_pad_GPIO_PAD[5] gfpga_pad_GPIO_PAD[6] gfpga_pad_GPIO_PAD[7] right_width_0_height_0__pin_0_
+ right_width_0_height_0__pin_10_ right_width_0_height_0__pin_11_ right_width_0_height_0__pin_12_
+ right_width_0_height_0__pin_13_ right_width_0_height_0__pin_14_ right_width_0_height_0__pin_15_
+ right_width_0_height_0__pin_1_ right_width_0_height_0__pin_2_ right_width_0_height_0__pin_3_
+ right_width_0_height_0__pin_4_ right_width_0_height_0__pin_5_ right_width_0_height_0__pin_6_
+ right_width_0_height_0__pin_7_ right_width_0_height_0__pin_8_ right_width_0_height_0__pin_9_
+ vpwr vgnd
XFILLER_596_56 vgnd vpwr scs8hd_decap_12
XFILLER_379_80 vgnd vpwr scs8hd_fill_1
XFILLER_449_39 vgnd vpwr scs8hd_decap_12
XPHY_1707 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1718 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1729 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_465_27 vgnd vpwr scs8hd_decap_12
XFILLER_481_15 vgnd vpwr scs8hd_decap_12
XFILLER_77_15 vgnd vpwr scs8hd_decap_12
XFILLER_481_59 vpwr vgnd scs8hd_fill_2
XFILLER_77_59 vpwr vgnd scs8hd_fill_2
XFILLER_172_3 vgnd vpwr scs8hd_decap_12
XFILLER_289_80 vgnd vpwr scs8hd_fill_1
XFILLER_359_39 vgnd vpwr scs8hd_decap_12
XFILLER_437_3 vgnd vpwr scs8hd_decap_12
XFILLER_375_27 vgnd vpwr scs8hd_decap_12
XFILLER_308_32 vgnd vpwr scs8hd_decap_12
XFILLER_391_15 vgnd vpwr scs8hd_decap_12
XFILLER_391_59 vpwr vgnd scs8hd_fill_2
XFILLER_83_80 vgnd vpwr scs8hd_fill_1
XFILLER_199_80 vgnd vpwr scs8hd_fill_1
XFILLER_269_39 vgnd vpwr scs8hd_decap_12
XFILLER_566_15 vgnd vpwr scs8hd_decap_12
XFILLER_285_27 vgnd vpwr scs8hd_decap_12
XFILLER_218_32 vgnd vpwr scs8hd_decap_12
XFILLER_515_74 vgnd vpwr scs8hd_decap_6
XFILLER_531_62 vgnd vpwr scs8hd_decap_12
XFILLER_531_51 vgnd vpwr scs8hd_decap_8
XFILLER_63_39 vgnd vpwr scs8hd_decap_12
XFILLER_179_39 vgnd vpwr scs8hd_decap_12
XFILLER_400_44 vgnd vpwr scs8hd_decap_12
XPHY_905 vgnd vpwr scs8hd_decap_3
XPHY_916 vgnd vpwr scs8hd_decap_3
XPHY_927 vgnd vpwr scs8hd_decap_3
XPHY_1504 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1515 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_938 vgnd vpwr scs8hd_decap_3
XPHY_949 vgnd vpwr scs8hd_decap_3
XPHY_1526 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1537 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1548 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_476_15 vgnd vpwr scs8hd_decap_12
XFILLER_195_27 vpwr vgnd scs8hd_fill_2
XPHY_1559 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
XFILLER_128_32 vgnd vpwr scs8hd_decap_12
XFILLER_572_80 vgnd vpwr scs8hd_fill_1
XFILLER_425_74 vgnd vpwr scs8hd_decap_6
XFILLER_387_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_51 vgnd vpwr scs8hd_decap_8
XFILLER_441_51 vgnd vpwr scs8hd_decap_8
XFILLER_441_62 vgnd vpwr scs8hd_decap_12
XFILLER_554_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_310_44 vgnd vpwr scs8hd_decap_12
XFILLER_386_15 vgnd vpwr scs8hd_decap_12
XFILLER_335_74 vgnd vpwr scs8hd_decap_6
XFILLER_482_80 vgnd vpwr scs8hd_fill_1
XFILLER_78_80 vgnd vpwr scs8hd_fill_1
XFILLER_204_56 vgnd vpwr scs8hd_decap_12
XFILLER_351_51 vgnd vpwr scs8hd_decap_8
XFILLER_351_62 vgnd vpwr scs8hd_decap_12
XFILLER_220_22 vgnd vpwr scs8hd_decap_8
XFILLER_220_44 vgnd vpwr scs8hd_decap_12
XFILLER_296_15 vgnd vpwr scs8hd_decap_12
XFILLER_245_74 vgnd vpwr scs8hd_decap_6
XFILLER_392_80 vgnd vpwr scs8hd_fill_1
XFILLER_114_56 vgnd vpwr scs8hd_decap_12
XFILLER_261_51 vgnd vpwr scs8hd_decap_8
XFILLER_261_62 vgnd vpwr scs8hd_decap_12
XFILLER_74_27 vgnd vpwr scs8hd_decap_4
XFILLER_130_44 vgnd vpwr scs8hd_decap_12
XPHY_702 vgnd vpwr scs8hd_decap_3
XFILLER_90_15 vgnd vpwr scs8hd_decap_12
XPHY_713 vgnd vpwr scs8hd_decap_3
XPHY_724 vgnd vpwr scs8hd_decap_3
XPHY_735 vgnd vpwr scs8hd_decap_3
XPHY_1323 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1312 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1301 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_746 vgnd vpwr scs8hd_decap_3
XPHY_757 vgnd vpwr scs8hd_decap_3
XPHY_768 vgnd vpwr scs8hd_decap_3
XFILLER_567_80 vgnd vpwr scs8hd_fill_1
XPHY_1334 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_135_3 vgnd vpwr scs8hd_decap_12
XPHY_1345 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1356 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_779 vgnd vpwr scs8hd_decap_3
XPHY_1367 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1378 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1389 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_302_3 vgnd vpwr scs8hd_decap_12
XFILLER_155_74 vgnd vpwr scs8hd_decap_6
XFILLER_171_51 vgnd vpwr scs8hd_decap_8
XFILLER_171_62 vgnd vpwr scs8hd_decap_12
XFILLER_0_79 vpwr vgnd scs8hd_fill_2
XFILLER_547_39 vgnd vpwr scs8hd_decap_12
XFILLER_477_80 vgnd vpwr scs8hd_fill_1
XFILLER_563_27 vgnd vpwr scs8hd_decap_12
XFILLER_50_3 vgnd vpwr scs8hd_decap_12
XFILLER_588_68 vgnd vpwr scs8hd_decap_12
XFILLER_387_80 vgnd vpwr scs8hd_fill_1
XFILLER_457_39 vgnd vpwr scs8hd_decap_12
XFILLER_473_27 vgnd vpwr scs8hd_decap_12
XFILLER_69_27 vgnd vpwr scs8hd_decap_12
XFILLER_406_32 vgnd vpwr scs8hd_decap_12
XFILLER_85_15 vgnd vpwr scs8hd_decap_12
XFILLER_85_59 vpwr vgnd scs8hd_fill_2
XFILLER_252_3 vgnd vpwr scs8hd_decap_12
XPHY_510 vgnd vpwr scs8hd_decap_3
XFILLER_498_68 vgnd vpwr scs8hd_decap_12
XPHY_521 vgnd vpwr scs8hd_decap_3
XPHY_532 vgnd vpwr scs8hd_decap_3
XPHY_543 vgnd vpwr scs8hd_decap_3
XPHY_1131 vgnd vpwr scs8hd_decap_3
XPHY_1120 vgnd vpwr scs8hd_decap_3
XPHY_554 vgnd vpwr scs8hd_decap_3
XPHY_565 vgnd vpwr scs8hd_decap_3
XPHY_576 vgnd vpwr scs8hd_decap_3
XPHY_587 vgnd vpwr scs8hd_decap_3
XFILLER_367_39 vgnd vpwr scs8hd_decap_8
XFILLER_517_3 vgnd vpwr scs8hd_decap_12
XPHY_1175 vgnd vpwr scs8hd_decap_3
XPHY_1164 vgnd vpwr scs8hd_decap_3
XPHY_1153 vgnd vpwr scs8hd_decap_3
XPHY_1142 vgnd vpwr scs8hd_decap_3
XFILLER_297_80 vgnd vpwr scs8hd_fill_1
XPHY_598 vgnd vpwr scs8hd_decap_3
XPHY_1197 vgnd vpwr scs8hd_decap_3
XPHY_1186 vgnd vpwr scs8hd_decap_3
XFILLER_166_73 vgnd vpwr scs8hd_decap_8
XFILLER_383_27 vgnd vpwr scs8hd_decap_12
XFILLER_316_32 vgnd vpwr scs8hd_decap_12
XFILLER_201_35 vgnd vpwr scs8hd_decap_12
XFILLER_558_27 vgnd vpwr scs8hd_decap_4
XFILLER_98_3 vgnd vpwr scs8hd_decap_12
XFILLER_91_80 vgnd vpwr scs8hd_fill_1
XFILLER_277_39 vgnd vpwr scs8hd_decap_12
XFILLER_574_15 vgnd vpwr scs8hd_decap_12
XFILLER_293_27 vgnd vpwr scs8hd_decap_12
XFILLER_226_32 vgnd vpwr scs8hd_decap_12
XFILLER_523_74 vgnd vpwr scs8hd_decap_6
XFILLER_468_27 vgnd vpwr scs8hd_decap_4
XFILLER_71_39 vgnd vpwr scs8hd_decap_12
XFILLER_187_39 vgnd vpwr scs8hd_decap_12
XFILLER_484_15 vgnd vpwr scs8hd_decap_12
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
XFILLER_136_32 vgnd vpwr scs8hd_decap_12
XFILLER_580_80 vgnd vpwr scs8hd_fill_1
XFILLER_433_74 vgnd vpwr scs8hd_decap_6
XFILLER_29_74 vgnd vpwr scs8hd_decap_6
XFILLER_467_3 vgnd vpwr scs8hd_decap_12
XFILLER_302_56 vgnd vpwr scs8hd_decap_12
XFILLER_45_62 vgnd vpwr scs8hd_decap_12
XFILLER_45_51 vgnd vpwr scs8hd_decap_8
XFILLER_378_27 vgnd vpwr scs8hd_decap_4
XPHY_340 vgnd vpwr scs8hd_decap_3
XPHY_351 vgnd vpwr scs8hd_decap_3
XPHY_362 vgnd vpwr scs8hd_decap_3
XPHY_373 vgnd vpwr scs8hd_decap_3
XPHY_384 vgnd vpwr scs8hd_decap_3
XPHY_395 vgnd vpwr scs8hd_decap_3
XFILLER_394_15 vgnd vpwr scs8hd_decap_12
XFILLER_6_56 vgnd vpwr scs8hd_decap_12
XFILLER_343_74 vgnd vpwr scs8hd_decap_6
XFILLER_490_80 vgnd vpwr scs8hd_fill_1
XFILLER_86_80 vgnd vpwr scs8hd_fill_1
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
XFILLER_212_12 vpwr vgnd scs8hd_fill_2
XFILLER_569_15 vgnd vpwr scs8hd_decap_12
XFILLER_569_59 vpwr vgnd scs8hd_fill_2
XFILLER_288_27 vgnd vpwr scs8hd_decap_4
XFILLER_106_68 vgnd vpwr scs8hd_decap_12
XFILLER_253_74 vgnd vpwr scs8hd_decap_6
XFILLER_122_56 vgnd vpwr scs8hd_decap_12
XFILLER_479_15 vgnd vpwr scs8hd_decap_12
XFILLER_82_27 vgnd vpwr scs8hd_decap_4
XFILLER_479_59 vpwr vgnd scs8hd_fill_2
XFILLER_198_27 vgnd vpwr scs8hd_decap_4
XFILLER_215_3 vgnd vpwr scs8hd_decap_12
XFILLER_575_80 vgnd vpwr scs8hd_fill_1
XFILLER_584_3 vgnd vpwr scs8hd_decap_12
XFILLER_163_74 vgnd vpwr scs8hd_decap_6
XFILLER_389_15 vgnd vpwr scs8hd_decap_12
XFILLER_389_59 vpwr vgnd scs8hd_fill_2
XPHY_170 vgnd vpwr scs8hd_decap_3
XPHY_192 vgnd vpwr scs8hd_decap_3
XPHY_181 vgnd vpwr scs8hd_decap_3
XFILLER_555_39 vgnd vpwr scs8hd_decap_12
XFILLER_485_80 vgnd vpwr scs8hd_fill_1
XFILLER_571_27 vgnd vpwr scs8hd_decap_12
XFILLER_504_32 vgnd vpwr scs8hd_decap_12
XFILLER_299_15 vgnd vpwr scs8hd_decap_12
XFILLER_299_59 vpwr vgnd scs8hd_fill_2
XFILLER_596_68 vgnd vpwr scs8hd_decap_12
XPHY_1708 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1719 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_529_62 vgnd vpwr scs8hd_decap_12
XFILLER_529_51 vgnd vpwr scs8hd_decap_8
XFILLER_395_80 vgnd vpwr scs8hd_fill_1
XFILLER_465_39 vgnd vpwr scs8hd_decap_12
XFILLER_77_27 vgnd vpwr scs8hd_decap_12
XFILLER_481_27 vgnd vpwr scs8hd_decap_12
XFILLER_414_32 vgnd vpwr scs8hd_decap_12
XFILLER_93_15 vgnd vpwr scs8hd_decap_12
XFILLER_93_59 vpwr vgnd scs8hd_fill_2
XFILLER_165_3 vgnd vpwr scs8hd_decap_12
XFILLER_332_3 vgnd vpwr scs8hd_decap_12
XFILLER_439_51 vgnd vpwr scs8hd_decap_8
XFILLER_439_62 vgnd vpwr scs8hd_decap_12
XFILLER_375_39 vgnd vpwr scs8hd_decap_12
XFILLER_308_44 vgnd vpwr scs8hd_decap_12
XFILLER_391_27 vgnd vpwr scs8hd_decap_12
XFILLER_324_32 vgnd vpwr scs8hd_decap_12
XFILLER_566_27 vgnd vpwr scs8hd_decap_4
XFILLER_80_3 vgnd vpwr scs8hd_decap_12
XFILLER_349_51 vgnd vpwr scs8hd_decap_8
XFILLER_349_62 vgnd vpwr scs8hd_decap_12
XFILLER_285_39 vgnd vpwr scs8hd_decap_12
XFILLER_582_15 vgnd vpwr scs8hd_decap_12
XFILLER_218_44 vgnd vpwr scs8hd_decap_12
XFILLER_234_32 vgnd vpwr scs8hd_decap_12
XFILLER_531_74 vgnd vpwr scs8hd_decap_6
XFILLER_400_56 vgnd vpwr scs8hd_decap_12
XPHY_906 vgnd vpwr scs8hd_decap_3
XPHY_917 vgnd vpwr scs8hd_decap_3
XPHY_1505 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_928 vgnd vpwr scs8hd_decap_3
XPHY_939 vgnd vpwr scs8hd_decap_3
XFILLER_259_51 vgnd vpwr scs8hd_decap_8
XFILLER_259_62 vgnd vpwr scs8hd_decap_12
XPHY_1516 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1527 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1538 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1549 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_476_27 vgnd vpwr scs8hd_decap_4
XFILLER_12_44 vgnd vpwr scs8hd_decap_12
XFILLER_128_44 vgnd vpwr scs8hd_decap_12
XFILLER_492_15 vgnd vpwr scs8hd_decap_12
XFILLER_88_15 vgnd vpwr scs8hd_decap_12
XFILLER_144_32 vgnd vpwr scs8hd_decap_12
XFILLER_282_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_74 vgnd vpwr scs8hd_decap_6
XFILLER_441_74 vgnd vpwr scs8hd_decap_6
XFILLER_547_3 vgnd vpwr scs8hd_decap_12
XFILLER_53_62 vgnd vpwr scs8hd_decap_12
XFILLER_53_51 vgnd vpwr scs8hd_decap_8
XFILLER_310_56 vgnd vpwr scs8hd_decap_12
XFILLER_169_51 vgnd vpwr scs8hd_decap_8
XFILLER_169_62 vgnd vpwr scs8hd_decap_12
XFILLER_386_27 vgnd vpwr scs8hd_decap_4
XFILLER_204_24 vgnd vpwr scs8hd_decap_6
XFILLER_204_68 vgnd vpwr scs8hd_decap_12
XFILLER_94_80 vgnd vpwr scs8hd_fill_1
XFILLER_351_74 vgnd vpwr scs8hd_decap_6
XFILLER_577_15 vgnd vpwr scs8hd_decap_12
XFILLER_220_56 vgnd vpwr scs8hd_decap_12
XFILLER_296_27 vgnd vpwr scs8hd_decap_4
XFILLER_114_68 vgnd vpwr scs8hd_decap_12
XFILLER_261_74 vgnd vpwr scs8hd_decap_6
XFILLER_487_15 vgnd vpwr scs8hd_decap_12
XFILLER_130_56 vgnd vpwr scs8hd_decap_12
XFILLER_90_27 vgnd vpwr scs8hd_decap_4
XPHY_703 vgnd vpwr scs8hd_decap_3
XPHY_714 vgnd vpwr scs8hd_decap_3
XPHY_725 vgnd vpwr scs8hd_decap_3
XPHY_736 vgnd vpwr scs8hd_decap_3
XPHY_1324 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1313 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1302 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_747 vgnd vpwr scs8hd_decap_3
XPHY_758 vgnd vpwr scs8hd_decap_3
XPHY_769 vgnd vpwr scs8hd_decap_3
XFILLER_487_59 vpwr vgnd scs8hd_fill_2
XPHY_1335 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1346 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1357 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_128_3 vgnd vpwr scs8hd_decap_12
XPHY_1368 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1379 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_583_80 vgnd vpwr scs8hd_fill_1
XFILLER_497_3 vgnd vpwr scs8hd_decap_12
XFILLER_602_32 vgnd vpwr scs8hd_decap_12
XFILLER_171_74 vgnd vpwr scs8hd_decap_6
XFILLER_0_47 vgnd vpwr scs8hd_decap_12
XFILLER_0_36 vgnd vpwr scs8hd_fill_1
XFILLER_397_15 vgnd vpwr scs8hd_decap_12
XFILLER_397_59 vpwr vgnd scs8hd_fill_2
XFILLER_563_39 vgnd vpwr scs8hd_decap_12
XFILLER_493_80 vgnd vpwr scs8hd_fill_1
XFILLER_89_80 vgnd vpwr scs8hd_fill_1
XFILLER_43_3 vgnd vpwr scs8hd_decap_12
XFILLER_512_32 vgnd vpwr scs8hd_decap_12
XFILLER_100_15 vgnd vpwr scs8hd_decap_12
XFILLER_537_62 vgnd vpwr scs8hd_decap_12
XFILLER_537_51 vgnd vpwr scs8hd_decap_8
XFILLER_69_39 vgnd vpwr scs8hd_decap_12
XFILLER_473_39 vgnd vpwr scs8hd_decap_12
XFILLER_406_44 vgnd vpwr scs8hd_decap_12
XFILLER_85_27 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _10_/X vgnd vpwr scs8hd_diode_2
XFILLER_422_32 vgnd vpwr scs8hd_decap_12
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
XPHY_500 vgnd vpwr scs8hd_decap_3
XFILLER_578_80 vgnd vpwr scs8hd_fill_1
XFILLER_245_3 vgnd vpwr scs8hd_decap_12
XPHY_511 vgnd vpwr scs8hd_decap_3
XPHY_522 vgnd vpwr scs8hd_decap_3
XPHY_533 vgnd vpwr scs8hd_decap_3
XPHY_544 vgnd vpwr scs8hd_decap_3
XPHY_1132 vgnd vpwr scs8hd_decap_3
XPHY_1121 vgnd vpwr scs8hd_decap_3
XPHY_1110 vgnd vpwr scs8hd_decap_3
XPHY_555 vgnd vpwr scs8hd_decap_3
XPHY_566 vgnd vpwr scs8hd_decap_3
XPHY_577 vgnd vpwr scs8hd_decap_3
XPHY_1165 vgnd vpwr scs8hd_decap_3
XPHY_1154 vgnd vpwr scs8hd_decap_3
XPHY_1143 vgnd vpwr scs8hd_decap_3
XPHY_588 vgnd vpwr scs8hd_decap_3
XPHY_599 vgnd vpwr scs8hd_decap_3
XFILLER_412_3 vgnd vpwr scs8hd_decap_12
XPHY_1198 vgnd vpwr scs8hd_decap_3
XPHY_1187 vgnd vpwr scs8hd_decap_3
XPHY_1176 vgnd vpwr scs8hd_decap_3
XFILLER_447_51 vgnd vpwr scs8hd_decap_8
XFILLER_447_62 vgnd vpwr scs8hd_decap_12
XFILLER_383_39 vgnd vpwr scs8hd_decap_12
XFILLER_316_44 vgnd vpwr scs8hd_decap_12
XFILLER_332_32 vgnd vpwr scs8hd_decap_12
XFILLER_201_47 vgnd vpwr scs8hd_decap_12
XFILLER_488_80 vgnd vpwr scs8hd_fill_1
XFILLER_574_27 vgnd vpwr scs8hd_decap_4
XFILLER_357_51 vgnd vpwr scs8hd_decap_8
XFILLER_357_62 vgnd vpwr scs8hd_decap_12
XFILLER_226_11 vgnd vpwr scs8hd_decap_3
XFILLER_293_39 vgnd vpwr scs8hd_decap_12
XFILLER_590_15 vgnd vpwr scs8hd_decap_12
XFILLER_226_22 vgnd vpwr scs8hd_decap_8
XFILLER_226_44 vgnd vpwr scs8hd_decap_12
XFILLER_242_32 vgnd vpwr scs8hd_decap_12
XFILLER_398_80 vgnd vpwr scs8hd_fill_1
XFILLER_267_51 vgnd vpwr scs8hd_decap_8
XFILLER_267_62 vgnd vpwr scs8hd_decap_12
XFILLER_484_27 vgnd vpwr scs8hd_decap_4
XFILLER_217_7 vgnd vpwr scs8hd_decap_4
XFILLER_20_44 vgnd vpwr scs8hd_decap_12
XFILLER_136_44 vgnd vpwr scs8hd_decap_12
XFILLER_96_15 vgnd vpwr scs8hd_decap_12
XFILLER_195_3 vgnd vpwr scs8hd_decap_4
XFILLER_152_32 vgnd vpwr scs8hd_decap_12
XFILLER_362_3 vgnd vpwr scs8hd_decap_12
XFILLER_45_74 vgnd vpwr scs8hd_decap_6
XFILLER_302_68 vgnd vpwr scs8hd_decap_12
XPHY_330 vgnd vpwr scs8hd_decap_3
XPHY_341 vgnd vpwr scs8hd_decap_3
XPHY_352 vgnd vpwr scs8hd_decap_3
XFILLER_101_80 vgnd vpwr scs8hd_fill_1
XFILLER_61_51 vgnd vpwr scs8hd_decap_8
XPHY_363 vgnd vpwr scs8hd_decap_3
XPHY_374 vgnd vpwr scs8hd_decap_3
XPHY_385 vgnd vpwr scs8hd_decap_3
XFILLER_61_62 vgnd vpwr scs8hd_decap_12
XFILLER_177_51 vgnd vpwr scs8hd_decap_8
XPHY_396 vgnd vpwr scs8hd_decap_3
XFILLER_394_27 vgnd vpwr scs8hd_decap_4
XFILLER_177_62 vgnd vpwr scs8hd_decap_12
XFILLER_6_68 vgnd vpwr scs8hd_decap_12
XFILLER_212_24 vgnd vpwr scs8hd_decap_3
XFILLER_212_57 vgnd vpwr scs8hd_decap_12
XFILLER_569_27 vgnd vpwr scs8hd_decap_12
XFILLER_585_15 vgnd vpwr scs8hd_decap_12
XFILLER_585_59 vpwr vgnd scs8hd_fill_2
XFILLER_122_68 vgnd vpwr scs8hd_decap_12
XFILLER_479_27 vgnd vpwr scs8hd_decap_12
XFILLER_495_15 vgnd vpwr scs8hd_decap_12
XFILLER_495_59 vpwr vgnd scs8hd_fill_2
XFILLER_110_3 vgnd vpwr scs8hd_decap_12
XFILLER_591_80 vgnd vpwr scs8hd_fill_1
XFILLER_577_3 vgnd vpwr scs8hd_decap_12
XFILLER_389_27 vgnd vpwr scs8hd_decap_12
XPHY_160 vgnd vpwr scs8hd_decap_3
XPHY_193 vgnd vpwr scs8hd_decap_3
XPHY_182 vgnd vpwr scs8hd_decap_3
XPHY_171 vgnd vpwr scs8hd_decap_3
XFILLER_207_35 vgnd vpwr scs8hd_decap_12
XFILLER_571_39 vgnd vpwr scs8hd_decap_12
XFILLER_97_80 vgnd vpwr scs8hd_fill_1
XFILLER_504_44 vgnd vpwr scs8hd_decap_12
XFILLER_299_27 vgnd vpwr scs8hd_decap_12
XFILLER_520_32 vgnd vpwr scs8hd_decap_12
XPHY_1709 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_529_74 vgnd vpwr scs8hd_decap_6
XFILLER_545_51 vgnd vpwr scs8hd_decap_8
XFILLER_184_19 vgnd vpwr scs8hd_fill_1
XFILLER_545_62 vgnd vpwr scs8hd_decap_12
XFILLER_481_39 vgnd vpwr scs8hd_decap_12
XFILLER_77_39 vgnd vpwr scs8hd_decap_12
XFILLER_414_44 vgnd vpwr scs8hd_decap_12
XFILLER_93_27 vgnd vpwr scs8hd_decap_12
XFILLER_26_32 vgnd vpwr scs8hd_decap_12
XFILLER_430_32 vgnd vpwr scs8hd_decap_12
XFILLER_158_3 vgnd vpwr scs8hd_decap_12
XFILLER_325_3 vgnd vpwr scs8hd_decap_12
XFILLER_439_74 vgnd vpwr scs8hd_decap_6
XFILLER_586_80 vgnd vpwr scs8hd_fill_1
XFILLER_308_56 vgnd vpwr scs8hd_decap_12
XFILLER_455_51 vgnd vpwr scs8hd_decap_8
XFILLER_455_62 vgnd vpwr scs8hd_decap_12
XFILLER_391_39 vgnd vpwr scs8hd_decap_12
XFILLER_324_44 vgnd vpwr scs8hd_decap_12
XFILLER_340_32 vgnd vpwr scs8hd_decap_12
XFILLER_349_74 vgnd vpwr scs8hd_decap_6
XFILLER_496_80 vgnd vpwr scs8hd_fill_1
XFILLER_73_3 vgnd vpwr scs8hd_decap_12
XFILLER_365_51 vgnd vpwr scs8hd_decap_8
XFILLER_582_27 vgnd vpwr scs8hd_decap_4
XFILLER_218_56 vgnd vpwr scs8hd_decap_12
XFILLER_365_62 vgnd vpwr scs8hd_decap_12
XFILLER_234_44 vgnd vpwr scs8hd_decap_12
XFILLER_103_15 vgnd vpwr scs8hd_decap_12
XFILLER_250_32 vgnd vpwr scs8hd_decap_12
XFILLER_103_59 vpwr vgnd scs8hd_fill_2
XPHY_907 vgnd vpwr scs8hd_decap_3
XPHY_918 vgnd vpwr scs8hd_decap_3
XPHY_1506 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_400_68 vgnd vpwr scs8hd_decap_12
XPHY_929 vgnd vpwr scs8hd_decap_3
XPHY_1517 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1528 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1539 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_259_74 vgnd vpwr scs8hd_decap_6
XFILLER_12_56 vgnd vpwr scs8hd_decap_12
XFILLER_275_51 vgnd vpwr scs8hd_decap_8
XFILLER_128_56 vgnd vpwr scs8hd_decap_12
XFILLER_88_27 vgnd vpwr scs8hd_decap_4
XFILLER_275_62 vgnd vpwr scs8hd_decap_12
XFILLER_492_27 vgnd vpwr scs8hd_decap_4
XFILLER_144_44 vgnd vpwr scs8hd_decap_12
XFILLER_160_32 vgnd vpwr scs8hd_decap_12
XFILLER_275_3 vgnd vpwr scs8hd_decap_12
XFILLER_442_3 vgnd vpwr scs8hd_decap_12
XFILLER_310_68 vgnd vpwr scs8hd_decap_12
XFILLER_53_74 vgnd vpwr scs8hd_decap_6
XFILLER_169_74 vgnd vpwr scs8hd_decap_6
XFILLER_185_62 vgnd vpwr scs8hd_decap_12
XFILLER_577_27 vgnd vpwr scs8hd_decap_8
XFILLER_220_68 vgnd vpwr scs8hd_decap_12
XFILLER_593_15 vgnd vpwr scs8hd_decap_12
XFILLER_593_59 vpwr vgnd scs8hd_fill_2
XFILLER_130_68 vgnd vpwr scs8hd_decap_12
XPHY_704 vgnd vpwr scs8hd_decap_3
XPHY_715 vgnd vpwr scs8hd_decap_3
XPHY_726 vgnd vpwr scs8hd_decap_3
XFILLER_487_27 vgnd vpwr scs8hd_decap_12
XPHY_1314 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1303 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_737 vgnd vpwr scs8hd_decap_3
XPHY_748 vgnd vpwr scs8hd_decap_3
XPHY_759 vgnd vpwr scs8hd_decap_3
XPHY_1336 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1325 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1347 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1358 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1369 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_99_15 vgnd vpwr scs8hd_decap_12
XFILLER_99_59 vpwr vgnd scs8hd_fill_2
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_392_3 vgnd vpwr scs8hd_decap_12
XFILLER_602_44 vgnd vpwr scs8hd_decap_12
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XFILLER_104_80 vgnd vpwr scs8hd_fill_1
XFILLER_0_59 vgnd vpwr scs8hd_decap_3
XFILLER_397_27 vgnd vpwr scs8hd_decap_12
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XFILLER_512_44 vgnd vpwr scs8hd_decap_12
XFILLER_588_15 vgnd vpwr scs8hd_decap_12
XFILLER_100_27 vgnd vpwr scs8hd_decap_4
XFILLER_537_74 vgnd vpwr scs8hd_decap_6
XFILLER_553_62 vgnd vpwr scs8hd_decap_12
XFILLER_553_51 vgnd vpwr scs8hd_decap_8
XFILLER_406_56 vgnd vpwr scs8hd_decap_12
XFILLER_85_39 vgnd vpwr scs8hd_decap_12
XFILLER_18_44 vgnd vpwr scs8hd_decap_12
XFILLER_422_44 vgnd vpwr scs8hd_decap_12
XFILLER_498_15 vgnd vpwr scs8hd_decap_12
XPHY_501 vgnd vpwr scs8hd_decap_3
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XPHY_512 vgnd vpwr scs8hd_decap_3
XPHY_523 vgnd vpwr scs8hd_decap_3
XPHY_534 vgnd vpwr scs8hd_decap_3
XPHY_1122 vgnd vpwr scs8hd_decap_3
XPHY_1111 vgnd vpwr scs8hd_decap_3
XPHY_1100 vgnd vpwr scs8hd_decap_3
XFILLER_140_3 vgnd vpwr scs8hd_decap_12
XFILLER_238_3 vgnd vpwr scs8hd_decap_12
XPHY_545 vgnd vpwr scs8hd_decap_3
XPHY_556 vgnd vpwr scs8hd_decap_3
XPHY_567 vgnd vpwr scs8hd_decap_3
XPHY_578 vgnd vpwr scs8hd_decap_3
XPHY_1166 vgnd vpwr scs8hd_decap_3
XPHY_1155 vgnd vpwr scs8hd_decap_3
XPHY_1144 vgnd vpwr scs8hd_decap_3
XPHY_1133 vgnd vpwr scs8hd_decap_3
XPHY_589 vgnd vpwr scs8hd_decap_3
XPHY_1199 vgnd vpwr scs8hd_decap_3
XPHY_1188 vgnd vpwr scs8hd_decap_3
XPHY_1177 vgnd vpwr scs8hd_decap_3
XFILLER_594_80 vgnd vpwr scs8hd_fill_1
XFILLER_405_3 vgnd vpwr scs8hd_decap_12
XFILLER_447_74 vgnd vpwr scs8hd_decap_6
XFILLER_59_62 vgnd vpwr scs8hd_decap_12
XFILLER_59_51 vgnd vpwr scs8hd_decap_8
XFILLER_316_56 vgnd vpwr scs8hd_decap_12
XFILLER_463_51 vgnd vpwr scs8hd_decap_8
XFILLER_463_62 vgnd vpwr scs8hd_decap_12
XFILLER_332_44 vgnd vpwr scs8hd_decap_12
XFILLER_201_59 vpwr vgnd scs8hd_fill_2
XFILLER_357_74 vgnd vpwr scs8hd_decap_6
XFILLER_590_27 vgnd vpwr scs8hd_decap_4
XFILLER_226_56 vgnd vpwr scs8hd_decap_12
XFILLER_373_51 vgnd vpwr scs8hd_decap_8
XFILLER_373_62 vgnd vpwr scs8hd_decap_12
XFILLER_242_44 vgnd vpwr scs8hd_decap_12
XFILLER_1_80 vgnd vpwr scs8hd_fill_1
XFILLER_111_15 vgnd vpwr scs8hd_decap_12
XFILLER_111_59 vpwr vgnd scs8hd_fill_2
XFILLER_267_74 vgnd vpwr scs8hd_decap_6
XFILLER_20_56 vgnd vpwr scs8hd_decap_12
XFILLER_136_56 vgnd vpwr scs8hd_decap_12
XFILLER_283_51 vgnd vpwr scs8hd_decap_8
XFILLER_283_62 vgnd vpwr scs8hd_decap_12
XFILLER_96_27 vgnd vpwr scs8hd_decap_4
XFILLER_152_44 vgnd vpwr scs8hd_decap_12
XFILLER_188_3 vgnd vpwr scs8hd_decap_12
XFILLER_589_80 vgnd vpwr scs8hd_fill_1
XFILLER_355_3 vgnd vpwr scs8hd_decap_12
XFILLER_522_3 vgnd vpwr scs8hd_decap_12
XPHY_320 vgnd vpwr scs8hd_decap_3
XPHY_331 vgnd vpwr scs8hd_decap_3
XPHY_342 vgnd vpwr scs8hd_decap_3
XPHY_353 vgnd vpwr scs8hd_decap_3
XPHY_364 vgnd vpwr scs8hd_decap_3
XPHY_375 vgnd vpwr scs8hd_decap_3
XPHY_386 vgnd vpwr scs8hd_decap_3
XFILLER_61_74 vgnd vpwr scs8hd_decap_6
XPHY_397 vgnd vpwr scs8hd_decap_3
XFILLER_177_74 vgnd vpwr scs8hd_decap_6
XFILLER_193_62 vgnd vpwr scs8hd_decap_12
XFILLER_569_39 vgnd vpwr scs8hd_decap_12
XFILLER_212_69 vgnd vpwr scs8hd_decap_12
XFILLER_499_80 vgnd vpwr scs8hd_fill_1
XFILLER_585_27 vgnd vpwr scs8hd_decap_12
XFILLER_518_32 vgnd vpwr scs8hd_decap_12
XFILLER_106_15 vgnd vpwr scs8hd_decap_12
XFILLER_479_39 vgnd vpwr scs8hd_decap_12
XFILLER_202_80 vgnd vpwr scs8hd_fill_1
XFILLER_495_27 vgnd vpwr scs8hd_decap_12
XANTENNA__04__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_428_32 vgnd vpwr scs8hd_decap_12
XFILLER_103_3 vgnd vpwr scs8hd_decap_12
XFILLER_472_3 vgnd vpwr scs8hd_decap_12
XFILLER_389_39 vgnd vpwr scs8hd_decap_12
XFILLER_112_80 vgnd vpwr scs8hd_fill_1
XPHY_161 vgnd vpwr scs8hd_decap_3
XPHY_150 vgnd vpwr scs8hd_decap_3
XPHY_194 vgnd vpwr scs8hd_decap_3
XPHY_183 vgnd vpwr scs8hd_decap_3
XPHY_172 vgnd vpwr scs8hd_decap_3
XFILLER_338_32 vgnd vpwr scs8hd_decap_12
XFILLER_207_47 vgnd vpwr scs8hd_decap_12
XFILLER_504_56 vgnd vpwr scs8hd_decap_12
XFILLER_299_39 vgnd vpwr scs8hd_decap_12
XFILLER_520_44 vgnd vpwr scs8hd_decap_12
XFILLER_596_15 vgnd vpwr scs8hd_decap_12
XFILLER_248_32 vgnd vpwr scs8hd_decap_12
XFILLER_545_74 vgnd vpwr scs8hd_decap_6
XFILLER_561_62 vgnd vpwr scs8hd_decap_12
XFILLER_561_51 vgnd vpwr scs8hd_decap_8
XFILLER_414_56 vgnd vpwr scs8hd_decap_12
XFILLER_93_39 vgnd vpwr scs8hd_decap_12
XFILLER_430_44 vgnd vpwr scs8hd_decap_12
XFILLER_26_44 vgnd vpwr scs8hd_decap_12
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_158_32 vgnd vpwr scs8hd_decap_12
XFILLER_220_3 vgnd vpwr scs8hd_decap_8
XFILLER_318_3 vgnd vpwr scs8hd_decap_12
XFILLER_308_68 vgnd vpwr scs8hd_decap_12
XFILLER_455_74 vgnd vpwr scs8hd_decap_6
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
XFILLER_107_80 vgnd vpwr scs8hd_fill_1
XFILLER_67_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_59 vpwr vgnd scs8hd_fill_2
XFILLER_324_56 vgnd vpwr scs8hd_decap_12
XFILLER_471_51 vgnd vpwr scs8hd_decap_8
XFILLER_471_62 vgnd vpwr scs8hd_decap_12
XFILLER_67_62 vgnd vpwr scs8hd_decap_12
XFILLER_340_44 vgnd vpwr scs8hd_decap_12
XFILLER_66_3 vgnd vpwr scs8hd_decap_12
XFILLER_218_68 vgnd vpwr scs8hd_decap_12
XFILLER_365_74 vgnd vpwr scs8hd_decap_6
XFILLER_234_56 vgnd vpwr scs8hd_decap_12
XFILLER_381_51 vgnd vpwr scs8hd_decap_8
XFILLER_381_62 vgnd vpwr scs8hd_decap_12
XFILLER_103_27 vgnd vpwr scs8hd_decap_12
XFILLER_250_44 vgnd vpwr scs8hd_decap_12
XPHY_908 vgnd vpwr scs8hd_decap_3
XPHY_919 vgnd vpwr scs8hd_decap_3
XPHY_1507 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1518 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1529 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_68 vgnd vpwr scs8hd_decap_12
XFILLER_128_68 vgnd vpwr scs8hd_decap_12
XFILLER_275_74 vgnd vpwr scs8hd_decap_6
XFILLER_144_56 vgnd vpwr scs8hd_decap_12
XFILLER_291_51 vgnd vpwr scs8hd_decap_8
XFILLER_291_62 vgnd vpwr scs8hd_decap_12
XFILLER_160_44 vgnd vpwr scs8hd_decap_12
XFILLER_170_3 vgnd vpwr scs8hd_decap_12
XFILLER_268_3 vgnd vpwr scs8hd_decap_12
XFILLER_597_80 vgnd vpwr scs8hd_fill_1
XFILLER_435_3 vgnd vpwr scs8hd_decap_12
XFILLER_602_3 vgnd vpwr scs8hd_decap_12
XFILLER_185_74 vgnd vpwr scs8hd_decap_6
Xlogical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ right_width_0_height_0__pin_8_ logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[4] vgnd vpwr scs8hd_ebufn_1
XFILLER_577_39 vpwr vgnd scs8hd_fill_2
XFILLER_300_80 vgnd vpwr scs8hd_fill_1
XFILLER_593_27 vgnd vpwr scs8hd_decap_12
XFILLER_526_32 vgnd vpwr scs8hd_decap_12
XFILLER_114_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_80 vgnd vpwr scs8hd_fill_1
XPHY_705 vgnd vpwr scs8hd_decap_3
XPHY_716 vgnd vpwr scs8hd_decap_3
XPHY_727 vgnd vpwr scs8hd_decap_3
XFILLER_487_39 vgnd vpwr scs8hd_decap_12
XPHY_1315 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1304 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_738 vgnd vpwr scs8hd_decap_3
XPHY_749 vgnd vpwr scs8hd_decap_3
XPHY_1337 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1326 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1348 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_210_80 vgnd vpwr scs8hd_fill_1
XPHY_1359 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_99_27 vgnd vpwr scs8hd_decap_12
XANTENNA__12__A _07_/C vgnd vpwr scs8hd_diode_2
XFILLER_436_32 vgnd vpwr scs8hd_decap_12
XFILLER_385_3 vgnd vpwr scs8hd_decap_12
XFILLER_602_56 vgnd vpwr scs8hd_decap_12
XFILLER_552_3 vgnd vpwr scs8hd_decap_12
XFILLER_0_27 vpwr vgnd scs8hd_fill_2
XFILLER_397_39 vgnd vpwr scs8hd_decap_12
XFILLER_120_80 vgnd vpwr scs8hd_fill_1
XFILLER_346_32 vgnd vpwr scs8hd_decap_12
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
XFILLER_512_56 vgnd vpwr scs8hd_decap_12
XFILLER_588_27 vgnd vpwr scs8hd_decap_4
XFILLER_231_68 vgnd vpwr scs8hd_fill_1
XFILLER_231_79 vpwr vgnd scs8hd_fill_2
XFILLER_109_15 vgnd vpwr scs8hd_decap_12
XFILLER_256_32 vgnd vpwr scs8hd_decap_12
XFILLER_109_59 vpwr vgnd scs8hd_fill_2
XFILLER_553_74 vgnd vpwr scs8hd_decap_6
XFILLER_406_68 vgnd vpwr scs8hd_decap_12
XFILLER_205_80 vgnd vpwr scs8hd_fill_1
XFILLER_422_56 vgnd vpwr scs8hd_decap_12
XFILLER_18_56 vgnd vpwr scs8hd_decap_12
XFILLER_498_27 vgnd vpwr scs8hd_decap_4
XANTENNA__07__A _07_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XPHY_502 vgnd vpwr scs8hd_decap_3
XPHY_513 vgnd vpwr scs8hd_decap_3
XPHY_524 vgnd vpwr scs8hd_decap_3
XPHY_535 vgnd vpwr scs8hd_decap_3
XPHY_1123 vgnd vpwr scs8hd_decap_3
XPHY_1112 vgnd vpwr scs8hd_decap_3
XPHY_1101 vgnd vpwr scs8hd_decap_3
XPHY_546 vgnd vpwr scs8hd_decap_3
XPHY_557 vgnd vpwr scs8hd_decap_3
XPHY_568 vgnd vpwr scs8hd_decap_3
XPHY_1156 vgnd vpwr scs8hd_decap_3
XPHY_1145 vgnd vpwr scs8hd_decap_3
XPHY_1134 vgnd vpwr scs8hd_decap_3
XFILLER_133_3 vgnd vpwr scs8hd_decap_12
XPHY_579 vgnd vpwr scs8hd_decap_3
XPHY_1189 vgnd vpwr scs8hd_decap_3
XPHY_1178 vgnd vpwr scs8hd_decap_3
XPHY_1167 vgnd vpwr scs8hd_decap_3
XFILLER_50_32 vgnd vpwr scs8hd_decap_12
XFILLER_166_32 vgnd vpwr scs8hd_decap_12
XFILLER_300_3 vgnd vpwr scs8hd_decap_12
XFILLER_316_68 vgnd vpwr scs8hd_decap_12
XFILLER_463_74 vgnd vpwr scs8hd_decap_6
XFILLER_59_74 vgnd vpwr scs8hd_decap_6
XFILLER_115_80 vgnd vpwr scs8hd_fill_1
XFILLER_332_56 vgnd vpwr scs8hd_decap_12
XFILLER_75_62 vgnd vpwr scs8hd_decap_12
XFILLER_75_51 vgnd vpwr scs8hd_decap_8
XPHY_1690 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_226_68 vgnd vpwr scs8hd_decap_12
XFILLER_373_74 vgnd vpwr scs8hd_decap_6
XFILLER_599_15 vgnd vpwr scs8hd_decap_12
XFILLER_242_56 vgnd vpwr scs8hd_decap_12
XFILLER_599_59 vpwr vgnd scs8hd_fill_2
XFILLER_111_27 vgnd vpwr scs8hd_decap_12
XFILLER_20_68 vgnd vpwr scs8hd_decap_12
XFILLER_136_68 vgnd vpwr scs8hd_decap_12
XFILLER_283_74 vgnd vpwr scs8hd_decap_6
XFILLER_152_56 vgnd vpwr scs8hd_decap_12
XFILLER_302_15 vgnd vpwr scs8hd_decap_12
XPHY_310 vgnd vpwr scs8hd_decap_3
XFILLER_250_3 vgnd vpwr scs8hd_decap_12
XFILLER_348_3 vgnd vpwr scs8hd_decap_12
XPHY_321 vgnd vpwr scs8hd_decap_3
XPHY_332 vgnd vpwr scs8hd_decap_3
XPHY_343 vgnd vpwr scs8hd_decap_3
XPHY_354 vgnd vpwr scs8hd_decap_3
XPHY_365 vgnd vpwr scs8hd_decap_3
XPHY_376 vgnd vpwr scs8hd_decap_3
XFILLER_515_3 vgnd vpwr scs8hd_decap_12
XPHY_387 vgnd vpwr scs8hd_decap_3
XPHY_398 vgnd vpwr scs8hd_decap_3
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XFILLER_193_74 vgnd vpwr scs8hd_decap_6
XFILLER_212_48 vgnd vpwr scs8hd_fill_1
XFILLER_96_3 vgnd vpwr scs8hd_decap_12
XFILLER_585_39 vgnd vpwr scs8hd_decap_12
XFILLER_518_44 vgnd vpwr scs8hd_decap_12
XFILLER_534_32 vgnd vpwr scs8hd_decap_12
XFILLER_106_27 vgnd vpwr scs8hd_decap_4
XFILLER_122_15 vgnd vpwr scs8hd_decap_12
XFILLER_559_62 vgnd vpwr scs8hd_decap_12
XFILLER_559_51 vgnd vpwr scs8hd_decap_8
XFILLER_495_39 vgnd vpwr scs8hd_decap_12
XFILLER_428_44 vgnd vpwr scs8hd_decap_12
XANTENNA__20__A gfpga_pad_GPIO_PAD[1] vgnd vpwr scs8hd_diode_2
XFILLER_444_32 vgnd vpwr scs8hd_decap_12
XFILLER_298_3 vgnd vpwr scs8hd_decap_12
XFILLER_465_3 vgnd vpwr scs8hd_decap_12
XFILLER_469_51 vgnd vpwr scs8hd_decap_8
XFILLER_469_62 vgnd vpwr scs8hd_decap_12
XPHY_151 vgnd vpwr scs8hd_decap_3
XPHY_140 vgnd vpwr scs8hd_decap_3
XPHY_184 vgnd vpwr scs8hd_decap_3
XPHY_173 vgnd vpwr scs8hd_decap_3
XPHY_162 vgnd vpwr scs8hd_decap_3
XPHY_195 vgnd vpwr scs8hd_decap_3
XFILLER_338_44 vgnd vpwr scs8hd_decap_12
XFILLER_207_15 vgnd vpwr scs8hd_decap_3
XFILLER_354_32 vgnd vpwr scs8hd_decap_12
XFILLER_207_59 vpwr vgnd scs8hd_fill_2
XFILLER_504_68 vgnd vpwr scs8hd_decap_12
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XFILLER_303_80 vgnd vpwr scs8hd_fill_1
XFILLER_520_56 vgnd vpwr scs8hd_decap_12
XFILLER_596_27 vgnd vpwr scs8hd_decap_4
XFILLER_379_51 vgnd vpwr scs8hd_decap_8
XFILLER_379_62 vgnd vpwr scs8hd_decap_12
XFILLER_248_44 vgnd vpwr scs8hd_decap_12
XFILLER_7_80 vgnd vpwr scs8hd_fill_1
XFILLER_117_15 vgnd vpwr scs8hd_decap_12
XFILLER_264_32 vgnd vpwr scs8hd_decap_12
XFILLER_117_59 vpwr vgnd scs8hd_fill_2
XFILLER_414_68 vgnd vpwr scs8hd_decap_12
XFILLER_561_74 vgnd vpwr scs8hd_decap_6
XFILLER_213_80 vgnd vpwr scs8hd_fill_1
XFILLER_26_56 vgnd vpwr scs8hd_decap_12
XFILLER_430_56 vgnd vpwr scs8hd_decap_12
XFILLER_289_51 vgnd vpwr scs8hd_decap_8
XFILLER_289_62 vgnd vpwr scs8hd_decap_12
XANTENNA__15__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_158_44 vgnd vpwr scs8hd_decap_12
XFILLER_213_3 vgnd vpwr scs8hd_decap_12
XFILLER_174_32 vgnd vpwr scs8hd_decap_12
XFILLER_582_3 vgnd vpwr scs8hd_decap_12
XFILLER_3_27 vgnd vpwr scs8hd_decap_12
XFILLER_67_74 vgnd vpwr scs8hd_decap_6
XFILLER_324_68 vgnd vpwr scs8hd_decap_12
XFILLER_471_74 vgnd vpwr scs8hd_decap_6
XFILLER_123_80 vgnd vpwr scs8hd_fill_1
XFILLER_83_62 vgnd vpwr scs8hd_decap_12
XFILLER_83_51 vgnd vpwr scs8hd_decap_8
XFILLER_340_56 vgnd vpwr scs8hd_decap_12
XFILLER_199_62 vgnd vpwr scs8hd_decap_12
XFILLER_59_3 vgnd vpwr scs8hd_decap_12
XFILLER_234_68 vgnd vpwr scs8hd_decap_12
XFILLER_381_74 vgnd vpwr scs8hd_decap_6
XFILLER_103_39 vgnd vpwr scs8hd_decap_12
XFILLER_250_56 vgnd vpwr scs8hd_decap_12
XFILLER_400_15 vgnd vpwr scs8hd_decap_12
XPHY_909 vgnd vpwr scs8hd_decap_3
XPHY_1508 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1519 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_144_68 vgnd vpwr scs8hd_decap_12
XFILLER_291_74 vgnd vpwr scs8hd_decap_6
XFILLER_160_56 vgnd vpwr scs8hd_decap_12
XFILLER_163_3 vgnd vpwr scs8hd_decap_12
XFILLER_310_15 vgnd vpwr scs8hd_decap_12
XFILLER_330_3 vgnd vpwr scs8hd_decap_12
XFILLER_428_3 vgnd vpwr scs8hd_decap_12
XFILLER_185_31 vgnd vpwr scs8hd_decap_12
XFILLER_118_80 vgnd vpwr scs8hd_fill_1
XFILLER_593_39 vgnd vpwr scs8hd_decap_12
XFILLER_229_68 vgnd vpwr scs8hd_fill_1
XFILLER_229_79 vpwr vgnd scs8hd_fill_2
XFILLER_526_44 vgnd vpwr scs8hd_decap_12
XFILLER_542_32 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _12_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_114_27 vgnd vpwr scs8hd_decap_4
XFILLER_130_15 vgnd vpwr scs8hd_decap_12
XPHY_706 vgnd vpwr scs8hd_decap_3
XPHY_717 vgnd vpwr scs8hd_decap_3
XPHY_1305 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_728 vgnd vpwr scs8hd_decap_3
XPHY_739 vgnd vpwr scs8hd_decap_3
XFILLER_567_62 vgnd vpwr scs8hd_decap_12
XFILLER_567_51 vgnd vpwr scs8hd_decap_8
XPHY_1338 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1327 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1316 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1349 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_99_39 vgnd vpwr scs8hd_decap_12
XANTENNA__12__B _14_/B vgnd vpwr scs8hd_diode_2
XFILLER_436_44 vgnd vpwr scs8hd_decap_12
XFILLER_305_15 vgnd vpwr scs8hd_decap_12
XFILLER_48_32 vgnd vpwr scs8hd_decap_12
XFILLER_305_59 vpwr vgnd scs8hd_fill_2
XFILLER_452_32 vgnd vpwr scs8hd_decap_12
XFILLER_280_3 vgnd vpwr scs8hd_decap_12
XFILLER_378_3 vgnd vpwr scs8hd_decap_12
XFILLER_602_68 vgnd vpwr scs8hd_decap_12
XFILLER_545_3 vgnd vpwr scs8hd_decap_12
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
XFILLER_401_80 vgnd vpwr scs8hd_fill_1
XFILLER_9_59 vpwr vgnd scs8hd_fill_2
XFILLER_477_51 vgnd vpwr scs8hd_decap_8
XFILLER_477_62 vgnd vpwr scs8hd_decap_12
XFILLER_196_30 vgnd vpwr scs8hd_fill_1
XFILLER_346_44 vgnd vpwr scs8hd_decap_12
XFILLER_215_15 vgnd vpwr scs8hd_decap_12
XFILLER_215_59 vpwr vgnd scs8hd_fill_2
XFILLER_362_32 vgnd vpwr scs8hd_decap_12
XFILLER_512_68 vgnd vpwr scs8hd_decap_12
XFILLER_311_80 vgnd vpwr scs8hd_fill_1
XFILLER_387_51 vgnd vpwr scs8hd_decap_8
XFILLER_387_62 vgnd vpwr scs8hd_decap_12
XFILLER_109_27 vgnd vpwr scs8hd_decap_12
XFILLER_256_44 vgnd vpwr scs8hd_decap_12
XFILLER_125_15 vgnd vpwr scs8hd_decap_12
XFILLER_125_59 vpwr vgnd scs8hd_fill_2
XFILLER_272_32 vgnd vpwr scs8hd_decap_12
XFILLER_18_68 vgnd vpwr scs8hd_decap_12
XFILLER_422_68 vgnd vpwr scs8hd_decap_12
XANTENNA__07__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_221_80 vgnd vpwr scs8hd_fill_1
XPHY_503 vgnd vpwr scs8hd_decap_3
XPHY_514 vgnd vpwr scs8hd_decap_3
XPHY_525 vgnd vpwr scs8hd_decap_3
XPHY_1113 vgnd vpwr scs8hd_decap_3
XPHY_1102 vgnd vpwr scs8hd_decap_3
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
XPHY_536 vgnd vpwr scs8hd_decap_3
XPHY_547 vgnd vpwr scs8hd_decap_3
XPHY_558 vgnd vpwr scs8hd_decap_3
XPHY_569 vgnd vpwr scs8hd_decap_3
XFILLER_297_51 vgnd vpwr scs8hd_decap_8
XPHY_1157 vgnd vpwr scs8hd_decap_3
XPHY_1146 vgnd vpwr scs8hd_decap_3
XPHY_1135 vgnd vpwr scs8hd_decap_3
XPHY_1124 vgnd vpwr scs8hd_decap_3
XFILLER_297_62 vgnd vpwr scs8hd_decap_12
XPHY_1179 vgnd vpwr scs8hd_decap_3
XPHY_1168 vgnd vpwr scs8hd_decap_3
XFILLER_126_3 vgnd vpwr scs8hd_decap_12
XANTENNA__23__A gfpga_pad_GPIO_PAD[4] vgnd vpwr scs8hd_diode_2
XFILLER_50_44 vgnd vpwr scs8hd_decap_12
XFILLER_166_44 vgnd vpwr scs8hd_decap_12
XFILLER_495_3 vgnd vpwr scs8hd_decap_12
XFILLER_182_32 vgnd vpwr scs8hd_decap_12
XFILLER_332_68 vgnd vpwr scs8hd_decap_12
XFILLER_75_74 vgnd vpwr scs8hd_decap_6
XFILLER_131_80 vgnd vpwr scs8hd_fill_1
XFILLER_91_51 vgnd vpwr scs8hd_decap_8
XFILLER_91_62 vgnd vpwr scs8hd_decap_12
XPHY_1680 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1691 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XFILLER_306_80 vgnd vpwr scs8hd_fill_1
XFILLER_599_27 vgnd vpwr scs8hd_decap_12
XFILLER_242_68 vgnd vpwr scs8hd_decap_12
XFILLER_111_39 vgnd vpwr scs8hd_decap_12
XFILLER_216_80 vgnd vpwr scs8hd_fill_1
XFILLER_152_68 vgnd vpwr scs8hd_decap_12
XANTENNA__18__A gfpga_pad_GPIO_PAD[7] vgnd vpwr scs8hd_diode_2
XFILLER_302_27 vgnd vpwr scs8hd_decap_4
XPHY_300 vgnd vpwr scs8hd_decap_3
XPHY_311 vgnd vpwr scs8hd_decap_3
XPHY_322 vgnd vpwr scs8hd_decap_3
XPHY_333 vgnd vpwr scs8hd_decap_3
XFILLER_243_3 vgnd vpwr scs8hd_decap_12
XPHY_344 vgnd vpwr scs8hd_decap_3
XPHY_355 vgnd vpwr scs8hd_decap_3
XPHY_366 vgnd vpwr scs8hd_decap_3
XPHY_377 vgnd vpwr scs8hd_decap_3
XPHY_388 vgnd vpwr scs8hd_decap_3
XPHY_399 vgnd vpwr scs8hd_decap_3
XFILLER_410_3 vgnd vpwr scs8hd_decap_12
XFILLER_508_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_193_31 vgnd vpwr scs8hd_decap_12
XFILLER_10_80 vgnd vpwr scs8hd_fill_1
XFILLER_126_80 vgnd vpwr scs8hd_fill_1
XFILLER_212_16 vgnd vpwr scs8hd_decap_8
XFILLER_89_3 vgnd vpwr scs8hd_decap_12
XFILLER_518_56 vgnd vpwr scs8hd_decap_12
XFILLER_534_44 vgnd vpwr scs8hd_decap_12
XFILLER_403_15 vgnd vpwr scs8hd_decap_12
XFILLER_550_32 vgnd vpwr scs8hd_decap_12
XFILLER_122_27 vgnd vpwr scs8hd_decap_4
XFILLER_403_59 vpwr vgnd scs8hd_fill_2
XFILLER_559_74 vgnd vpwr scs8hd_decap_6
XFILLER_575_51 vgnd vpwr scs8hd_decap_8
XFILLER_575_62 vgnd vpwr scs8hd_decap_12
XFILLER_428_56 vgnd vpwr scs8hd_decap_12
XFILLER_444_44 vgnd vpwr scs8hd_decap_12
XFILLER_193_3 vpwr vgnd scs8hd_fill_2
XFILLER_313_15 vgnd vpwr scs8hd_decap_12
XFILLER_56_32 vgnd vpwr scs8hd_decap_12
XFILLER_460_32 vgnd vpwr scs8hd_decap_12
XFILLER_313_59 vpwr vgnd scs8hd_fill_2
XFILLER_360_3 vgnd vpwr scs8hd_decap_12
XFILLER_458_3 vgnd vpwr scs8hd_decap_12
XPHY_152 vgnd vpwr scs8hd_decap_3
XPHY_141 vgnd vpwr scs8hd_decap_3
XPHY_130 vgnd vpwr scs8hd_decap_3
XFILLER_469_74 vgnd vpwr scs8hd_decap_6
XPHY_185 vgnd vpwr scs8hd_decap_3
XPHY_174 vgnd vpwr scs8hd_decap_3
XPHY_163 vgnd vpwr scs8hd_decap_3
XPHY_196 vgnd vpwr scs8hd_decap_3
XFILLER_485_51 vgnd vpwr scs8hd_decap_8
XFILLER_338_56 vgnd vpwr scs8hd_decap_12
XFILLER_485_62 vgnd vpwr scs8hd_decap_12
XFILLER_354_44 vgnd vpwr scs8hd_decap_12
XFILLER_223_15 vgnd vpwr scs8hd_decap_12
XFILLER_370_32 vgnd vpwr scs8hd_decap_12
XFILLER_223_59 vpwr vgnd scs8hd_fill_2
XFILLER_520_68 vgnd vpwr scs8hd_decap_12
XFILLER_379_74 vgnd vpwr scs8hd_decap_6
XFILLER_395_51 vgnd vpwr scs8hd_decap_8
XFILLER_248_56 vgnd vpwr scs8hd_decap_12
XFILLER_395_62 vgnd vpwr scs8hd_decap_12
XFILLER_117_27 vgnd vpwr scs8hd_decap_12
XFILLER_264_44 vgnd vpwr scs8hd_decap_12
XFILLER_133_15 vgnd vpwr scs8hd_decap_12
XFILLER_280_32 vgnd vpwr scs8hd_decap_12
XFILLER_133_59 vpwr vgnd scs8hd_fill_2
XFILLER_430_68 vgnd vpwr scs8hd_decap_12
XFILLER_26_68 vgnd vpwr scs8hd_decap_12
XFILLER_289_74 vgnd vpwr scs8hd_decap_6
XANTENNA__15__B _14_/B vgnd vpwr scs8hd_diode_2
XFILLER_42_56 vgnd vpwr scs8hd_decap_12
XFILLER_158_56 vgnd vpwr scs8hd_decap_12
XFILLER_308_15 vgnd vpwr scs8hd_decap_12
XFILLER_206_3 vpwr vgnd scs8hd_fill_2
XFILLER_174_44 vgnd vpwr scs8hd_decap_12
XFILLER_3_39 vgnd vpwr scs8hd_decap_12
XFILLER_575_3 vgnd vpwr scs8hd_decap_12
XFILLER_190_21 vgnd vpwr scs8hd_decap_8
XFILLER_190_32 vgnd vpwr scs8hd_decap_12
XFILLER_404_80 vgnd vpwr scs8hd_fill_1
XFILLER_340_68 vgnd vpwr scs8hd_decap_12
XFILLER_83_74 vgnd vpwr scs8hd_decap_6
XFILLER_199_74 vgnd vpwr scs8hd_decap_6
XFILLER_314_80 vgnd vpwr scs8hd_fill_1
XFILLER_250_68 vgnd vpwr scs8hd_decap_12
XFILLER_400_27 vgnd vpwr scs8hd_decap_4
XPHY_1509 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
XFILLER_128_15 vgnd vpwr scs8hd_decap_12
XFILLER_224_80 vgnd vpwr scs8hd_fill_1
XFILLER_160_68 vgnd vpwr scs8hd_decap_12
XFILLER_310_27 vgnd vpwr scs8hd_decap_4
XFILLER_156_3 vgnd vpwr scs8hd_decap_12
XFILLER_323_3 vgnd vpwr scs8hd_decap_12
XFILLER_185_43 vgnd vpwr scs8hd_decap_12
XFILLER_134_80 vgnd vpwr scs8hd_fill_1
XFILLER_501_15 vgnd vpwr scs8hd_decap_12
XFILLER_501_59 vpwr vgnd scs8hd_fill_2
XFILLER_71_3 vgnd vpwr scs8hd_decap_12
XFILLER_526_56 vgnd vpwr scs8hd_decap_12
XFILLER_309_80 vgnd vpwr scs8hd_fill_1
XFILLER_542_44 vgnd vpwr scs8hd_decap_12
XFILLER_411_15 vgnd vpwr scs8hd_decap_12
XFILLER_130_27 vgnd vpwr scs8hd_decap_4
XFILLER_411_59 vpwr vgnd scs8hd_fill_2
XPHY_707 vgnd vpwr scs8hd_decap_3
XPHY_718 vgnd vpwr scs8hd_decap_3
XPHY_1306 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_729 vgnd vpwr scs8hd_decap_3
XPHY_1339 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1328 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1317 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_567_74 vgnd vpwr scs8hd_decap_6
XANTENNA__12__C _07_/A vgnd vpwr scs8hd_diode_2
XFILLER_583_62 vgnd vpwr scs8hd_decap_12
XFILLER_583_51 vgnd vpwr scs8hd_decap_8
XFILLER_219_80 vgnd vpwr scs8hd_fill_1
XFILLER_436_56 vgnd vpwr scs8hd_decap_12
XFILLER_305_27 vgnd vpwr scs8hd_decap_12
XFILLER_452_44 vgnd vpwr scs8hd_decap_12
XFILLER_48_44 vgnd vpwr scs8hd_decap_12
XFILLER_273_3 vgnd vpwr scs8hd_decap_12
XFILLER_321_15 vgnd vpwr scs8hd_decap_12
XFILLER_64_32 vgnd vpwr scs8hd_decap_12
XFILLER_321_59 vpwr vgnd scs8hd_fill_2
XFILLER_538_3 vgnd vpwr scs8hd_decap_12
XFILLER_440_3 vgnd vpwr scs8hd_decap_12
XFILLER_9_27 vgnd vpwr scs8hd_decap_12
XFILLER_477_74 vgnd vpwr scs8hd_decap_6
XFILLER_13_80 vgnd vpwr scs8hd_fill_1
XFILLER_129_80 vgnd vpwr scs8hd_fill_1
XFILLER_89_51 vgnd vpwr scs8hd_decap_8
XFILLER_346_56 vgnd vpwr scs8hd_decap_12
XFILLER_493_51 vgnd vpwr scs8hd_decap_8
XFILLER_493_62 vgnd vpwr scs8hd_decap_12
XFILLER_89_62 vgnd vpwr scs8hd_decap_12
XFILLER_215_27 vgnd vpwr scs8hd_decap_12
XFILLER_362_44 vgnd vpwr scs8hd_decap_12
XFILLER_231_15 vgnd vpwr scs8hd_decap_12
XFILLER_231_59 vpwr vgnd scs8hd_fill_2
XFILLER_387_74 vgnd vpwr scs8hd_decap_6
XFILLER_109_39 vgnd vpwr scs8hd_decap_12
XFILLER_256_56 vgnd vpwr scs8hd_decap_12
XFILLER_406_15 vgnd vpwr scs8hd_decap_12
XFILLER_125_27 vgnd vpwr scs8hd_decap_12
XFILLER_272_44 vgnd vpwr scs8hd_decap_12
XFILLER_205_60 vgnd vpwr scs8hd_fill_1
XFILLER_141_15 vgnd vpwr scs8hd_decap_12
XFILLER_141_59 vpwr vgnd scs8hd_fill_2
XFILLER_502_80 vgnd vpwr scs8hd_fill_1
XANTENNA__07__C _07_/C vgnd vpwr scs8hd_diode_2
XPHY_504 vgnd vpwr scs8hd_decap_3
XPHY_515 vgnd vpwr scs8hd_decap_3
XPHY_526 vgnd vpwr scs8hd_decap_3
XPHY_1114 vgnd vpwr scs8hd_decap_3
XPHY_1103 vgnd vpwr scs8hd_decap_3
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XPHY_537 vgnd vpwr scs8hd_decap_3
XPHY_548 vgnd vpwr scs8hd_decap_3
XPHY_559 vgnd vpwr scs8hd_decap_3
XPHY_1147 vgnd vpwr scs8hd_decap_3
XPHY_1136 vgnd vpwr scs8hd_decap_3
XPHY_1125 vgnd vpwr scs8hd_decap_3
XFILLER_297_74 vgnd vpwr scs8hd_decap_6
XPHY_1169 vgnd vpwr scs8hd_decap_3
XPHY_1158 vgnd vpwr scs8hd_decap_3
XFILLER_50_56 vgnd vpwr scs8hd_decap_12
XFILLER_119_3 vgnd vpwr scs8hd_decap_12
XFILLER_166_56 vgnd vpwr scs8hd_decap_12
XFILLER_316_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
XFILLER_182_44 vgnd vpwr scs8hd_decap_12
XFILLER_390_3 vgnd vpwr scs8hd_decap_12
XFILLER_488_3 vgnd vpwr scs8hd_decap_12
XFILLER_412_80 vgnd vpwr scs8hd_fill_1
XFILLER_91_74 vgnd vpwr scs8hd_decap_6
XPHY_1670 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1681 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1692 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XFILLER_599_39 vgnd vpwr scs8hd_decap_12
XFILLER_322_80 vgnd vpwr scs8hd_fill_1
XFILLER_548_32 vgnd vpwr scs8hd_decap_12
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XFILLER_136_15 vgnd vpwr scs8hd_decap_12
XFILLER_195_7 vgnd vpwr scs8hd_fill_1
XPHY_301 vgnd vpwr scs8hd_decap_3
XFILLER_101_51 vgnd vpwr scs8hd_decap_8
XPHY_312 vgnd vpwr scs8hd_decap_3
XPHY_323 vgnd vpwr scs8hd_decap_3
XPHY_334 vgnd vpwr scs8hd_decap_3
XFILLER_101_62 vgnd vpwr scs8hd_decap_12
XPHY_345 vgnd vpwr scs8hd_decap_3
XPHY_356 vgnd vpwr scs8hd_decap_3
XPHY_367 vgnd vpwr scs8hd_decap_3
XFILLER_236_3 vgnd vpwr scs8hd_decap_12
XFILLER_458_32 vgnd vpwr scs8hd_decap_12
XPHY_378 vgnd vpwr scs8hd_decap_3
XPHY_389 vgnd vpwr scs8hd_decap_3
XFILLER_403_3 vgnd vpwr scs8hd_decap_12
XFILLER_193_43 vgnd vpwr scs8hd_decap_12
XFILLER_407_80 vgnd vpwr scs8hd_fill_1
XFILLER_142_80 vgnd vpwr scs8hd_fill_1
XFILLER_368_32 vgnd vpwr scs8hd_decap_12
XPHY_890 vgnd vpwr scs8hd_decap_3
XFILLER_518_68 vgnd vpwr scs8hd_decap_12
XFILLER_534_56 vgnd vpwr scs8hd_decap_12
XFILLER_317_80 vgnd vpwr scs8hd_fill_1
XFILLER_550_44 vgnd vpwr scs8hd_decap_12
XFILLER_403_27 vgnd vpwr scs8hd_decap_12
XFILLER_15_15 vgnd vpwr scs8hd_decap_12
XFILLER_15_59 vpwr vgnd scs8hd_fill_2
XFILLER_278_32 vgnd vpwr scs8hd_decap_12
XFILLER_575_74 vgnd vpwr scs8hd_decap_6
XFILLER_428_68 vgnd vpwr scs8hd_decap_12
XFILLER_591_62 vgnd vpwr scs8hd_decap_12
XFILLER_591_51 vgnd vpwr scs8hd_decap_8
XFILLER_227_80 vgnd vpwr scs8hd_fill_1
XFILLER_444_56 vgnd vpwr scs8hd_decap_12
XFILLER_313_27 vgnd vpwr scs8hd_decap_12
XFILLER_460_44 vgnd vpwr scs8hd_decap_12
XFILLER_56_44 vgnd vpwr scs8hd_decap_12
XFILLER_186_3 vgnd vpwr scs8hd_decap_12
XFILLER_353_3 vgnd vpwr scs8hd_decap_12
XFILLER_72_32 vgnd vpwr scs8hd_decap_12
XPHY_142 vgnd vpwr scs8hd_decap_3
XPHY_131 vgnd vpwr scs8hd_decap_3
XPHY_120 vgnd vpwr scs8hd_decap_3
XFILLER_188_21 vgnd vpwr scs8hd_decap_8
XFILLER_188_32 vgnd vpwr scs8hd_decap_12
XFILLER_520_3 vgnd vpwr scs8hd_decap_12
XPHY_175 vgnd vpwr scs8hd_decap_3
XPHY_164 vgnd vpwr scs8hd_decap_3
XPHY_153 vgnd vpwr scs8hd_decap_3
XPHY_197 vgnd vpwr scs8hd_decap_3
XPHY_186 vgnd vpwr scs8hd_decap_3
XFILLER_338_68 vgnd vpwr scs8hd_decap_12
XFILLER_485_74 vgnd vpwr scs8hd_decap_6
XFILLER_21_80 vgnd vpwr scs8hd_fill_1
XFILLER_137_80 vgnd vpwr scs8hd_fill_1
XFILLER_354_56 vgnd vpwr scs8hd_decap_12
XFILLER_97_62 vgnd vpwr scs8hd_decap_12
XFILLER_97_51 vgnd vpwr scs8hd_decap_8
XFILLER_504_15 vgnd vpwr scs8hd_decap_12
XFILLER_223_27 vgnd vpwr scs8hd_decap_12
XFILLER_370_44 vgnd vpwr scs8hd_decap_12
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_600_80 vgnd vpwr scs8hd_fill_1
XFILLER_248_68 vgnd vpwr scs8hd_decap_12
XFILLER_395_74 vgnd vpwr scs8hd_decap_6
XFILLER_117_39 vgnd vpwr scs8hd_decap_12
XFILLER_264_56 vgnd vpwr scs8hd_decap_12
XFILLER_414_15 vgnd vpwr scs8hd_decap_12
XFILLER_133_27 vgnd vpwr scs8hd_decap_12
XFILLER_280_44 vgnd vpwr scs8hd_decap_12
XFILLER_510_80 vgnd vpwr scs8hd_fill_1
XANTENNA__15__C _07_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_68 vgnd vpwr scs8hd_decap_12
XFILLER_158_68 vgnd vpwr scs8hd_decap_12
XFILLER_308_27 vgnd vpwr scs8hd_decap_4
XFILLER_101_3 vgnd vpwr scs8hd_decap_12
XFILLER_174_56 vgnd vpwr scs8hd_decap_12
XFILLER_324_15 vgnd vpwr scs8hd_decap_12
XFILLER_568_3 vgnd vpwr scs8hd_decap_12
XFILLER_190_44 vgnd vpwr scs8hd_decap_12
XFILLER_470_3 vgnd vpwr scs8hd_decap_12
XFILLER_199_31 vgnd vpwr scs8hd_decap_12
XFILLER_16_80 vgnd vpwr scs8hd_fill_1
XFILLER_420_80 vgnd vpwr scs8hd_fill_1
XFILLER_234_15 vgnd vpwr scs8hd_decap_12
XFILLER_330_80 vgnd vpwr scs8hd_fill_1
XFILLER_556_32 vgnd vpwr scs8hd_decap_12
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
XFILLER_409_15 vgnd vpwr scs8hd_decap_12
XFILLER_128_27 vgnd vpwr scs8hd_decap_4
XFILLER_409_59 vpwr vgnd scs8hd_fill_2
XFILLER_144_15 vgnd vpwr scs8hd_decap_12
XFILLER_505_80 vgnd vpwr scs8hd_fill_1
XFILLER_240_80 vgnd vpwr scs8hd_fill_1
XFILLER_149_3 vgnd vpwr scs8hd_decap_12
XFILLER_319_15 vgnd vpwr scs8hd_decap_12
XFILLER_466_32 vgnd vpwr scs8hd_decap_12
XFILLER_316_3 vgnd vpwr scs8hd_decap_12
XFILLER_319_59 vpwr vgnd scs8hd_fill_2
XFILLER_185_55 vgnd vpwr scs8hd_decap_6
XFILLER_415_80 vgnd vpwr scs8hd_fill_1
XFILLER_501_27 vgnd vpwr scs8hd_decap_12
XFILLER_150_80 vgnd vpwr scs8hd_fill_1
XFILLER_229_15 vgnd vpwr scs8hd_decap_12
XFILLER_376_32 vgnd vpwr scs8hd_decap_12
XFILLER_229_59 vpwr vgnd scs8hd_fill_2
XFILLER_64_3 vgnd vpwr scs8hd_decap_12
XFILLER_526_68 vgnd vpwr scs8hd_decap_12
XFILLER_542_56 vgnd vpwr scs8hd_decap_12
XFILLER_325_80 vgnd vpwr scs8hd_fill_1
XFILLER_411_27 vgnd vpwr scs8hd_decap_12
XPHY_708 vgnd vpwr scs8hd_decap_3
XPHY_719 vgnd vpwr scs8hd_decap_3
XPHY_1329 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1318 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1307 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_15 vgnd vpwr scs8hd_decap_12
XFILLER_23_59 vpwr vgnd scs8hd_fill_2
XFILLER_139_15 vgnd vpwr scs8hd_decap_12
XFILLER_286_32 vgnd vpwr scs8hd_decap_12
XFILLER_139_59 vpwr vgnd scs8hd_fill_2
XANTENNA__12__D _08_/Y vgnd vpwr scs8hd_diode_2
XFILLER_583_74 vgnd vpwr scs8hd_decap_6
XFILLER_436_68 vgnd vpwr scs8hd_decap_12
XFILLER_235_80 vgnd vpwr scs8hd_fill_1
XFILLER_305_39 vgnd vpwr scs8hd_decap_12
XFILLER_452_56 vgnd vpwr scs8hd_decap_12
XFILLER_602_15 vgnd vpwr scs8hd_decap_12
XFILLER_48_56 vgnd vpwr scs8hd_decap_12
XFILLER_321_27 vgnd vpwr scs8hd_decap_12
XFILLER_64_44 vgnd vpwr scs8hd_decap_12
XFILLER_266_3 vgnd vpwr scs8hd_decap_12
XFILLER_433_3 vgnd vpwr scs8hd_decap_12
XFILLER_80_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_39 vgnd vpwr scs8hd_decap_12
XFILLER_196_32 vgnd vpwr scs8hd_decap_12
XFILLER_600_3 vgnd vpwr scs8hd_decap_12
XFILLER_346_68 vgnd vpwr scs8hd_decap_12
XFILLER_493_74 vgnd vpwr scs8hd_decap_6
XFILLER_89_74 vgnd vpwr scs8hd_decap_6
XFILLER_145_80 vgnd vpwr scs8hd_fill_1
XFILLER_215_39 vgnd vpwr scs8hd_decap_12
XFILLER_362_56 vgnd vpwr scs8hd_decap_12
XFILLER_512_15 vgnd vpwr scs8hd_decap_12
XFILLER_231_27 vgnd vpwr scs8hd_decap_12
XFILLER_256_68 vgnd vpwr scs8hd_decap_12
XFILLER_406_27 vgnd vpwr scs8hd_decap_4
XFILLER_125_39 vgnd vpwr scs8hd_decap_12
XFILLER_272_56 vgnd vpwr scs8hd_decap_12
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
XFILLER_422_15 vgnd vpwr scs8hd_decap_12
XFILLER_141_27 vgnd vpwr scs8hd_decap_12
XANTENNA__07__D enable vgnd vpwr scs8hd_diode_2
XPHY_505 vgnd vpwr scs8hd_decap_3
XPHY_516 vgnd vpwr scs8hd_decap_3
XPHY_1104 vgnd vpwr scs8hd_decap_3
XPHY_527 vgnd vpwr scs8hd_decap_3
XPHY_538 vgnd vpwr scs8hd_decap_3
XPHY_549 vgnd vpwr scs8hd_decap_3
XPHY_1148 vgnd vpwr scs8hd_decap_3
XPHY_1137 vgnd vpwr scs8hd_decap_3
XPHY_1126 vgnd vpwr scs8hd_decap_3
XPHY_1115 vgnd vpwr scs8hd_decap_3
XPHY_1159 vgnd vpwr scs8hd_decap_3
XFILLER_50_68 vgnd vpwr scs8hd_decap_12
XFILLER_166_68 vgnd vpwr scs8hd_fill_1
XFILLER_316_27 vgnd vpwr scs8hd_decap_4
XFILLER_182_56 vgnd vpwr scs8hd_decap_12
XFILLER_332_15 vgnd vpwr scs8hd_decap_12
XFILLER_383_3 vgnd vpwr scs8hd_decap_12
XFILLER_550_3 vgnd vpwr scs8hd_decap_12
XFILLER_201_19 vpwr vgnd scs8hd_fill_2
XFILLER_24_80 vgnd vpwr scs8hd_fill_1
XPHY_1660 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1671 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1682 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1693 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_507_15 vgnd vpwr scs8hd_decap_12
XFILLER_507_59 vpwr vgnd scs8hd_fill_2
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
XFILLER_242_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
XFILLER_548_44 vgnd vpwr scs8hd_decap_12
XFILLER_564_32 vgnd vpwr scs8hd_decap_12
XFILLER_417_15 vgnd vpwr scs8hd_decap_12
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XFILLER_417_59 vpwr vgnd scs8hd_fill_2
XFILLER_136_27 vgnd vpwr scs8hd_decap_4
XFILLER_152_15 vgnd vpwr scs8hd_decap_12
XFILLER_513_80 vgnd vpwr scs8hd_fill_1
XFILLER_589_62 vgnd vpwr scs8hd_decap_12
XFILLER_589_51 vgnd vpwr scs8hd_decap_8
XPHY_302 vgnd vpwr scs8hd_decap_3
XPHY_313 vgnd vpwr scs8hd_decap_3
XPHY_324 vgnd vpwr scs8hd_decap_3
XFILLER_101_74 vgnd vpwr scs8hd_decap_6
XPHY_335 vgnd vpwr scs8hd_decap_3
XPHY_346 vgnd vpwr scs8hd_decap_3
XPHY_357 vgnd vpwr scs8hd_decap_3
XPHY_368 vgnd vpwr scs8hd_decap_3
XFILLER_458_44 vgnd vpwr scs8hd_decap_12
XFILLER_131_3 vgnd vpwr scs8hd_decap_12
XPHY_379 vgnd vpwr scs8hd_decap_3
XFILLER_229_3 vgnd vpwr scs8hd_decap_12
XFILLER_327_15 vgnd vpwr scs8hd_decap_12
XFILLER_474_32 vgnd vpwr scs8hd_decap_12
XFILLER_327_59 vpwr vgnd scs8hd_fill_2
XFILLER_193_55 vgnd vpwr scs8hd_decap_6
XFILLER_598_3 vgnd vpwr scs8hd_decap_12
XFILLER_423_80 vgnd vpwr scs8hd_fill_1
XFILLER_19_80 vgnd vpwr scs8hd_fill_1
XFILLER_212_29 vpwr vgnd scs8hd_fill_2
XFILLER_499_51 vgnd vpwr scs8hd_decap_8
XFILLER_499_62 vgnd vpwr scs8hd_decap_12
XFILLER_368_44 vgnd vpwr scs8hd_decap_4
XPHY_880 vgnd vpwr scs8hd_decap_3
XPHY_891 vgnd vpwr scs8hd_decap_3
XFILLER_237_15 vgnd vpwr scs8hd_decap_12
XPHY_1490 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_384_32 vgnd vpwr scs8hd_decap_12
XFILLER_237_59 vpwr vgnd scs8hd_fill_2
XFILLER_534_68 vgnd vpwr scs8hd_decap_12
XFILLER_333_80 vgnd vpwr scs8hd_fill_1
XFILLER_403_39 vgnd vpwr scs8hd_decap_12
XFILLER_550_56 vgnd vpwr scs8hd_decap_12
X_09_ address[1] enable address[3] _08_/Y _09_/X vgnd vpwr scs8hd_and4_4
XFILLER_15_27 vgnd vpwr scs8hd_decap_12
XFILLER_278_44 vgnd vpwr scs8hd_decap_12
XFILLER_31_15 vgnd vpwr scs8hd_decap_12
XFILLER_31_59 vpwr vgnd scs8hd_fill_2
XFILLER_147_15 vgnd vpwr scs8hd_decap_12
XFILLER_147_59 vpwr vgnd scs8hd_fill_2
XFILLER_294_32 vgnd vpwr scs8hd_decap_12
XFILLER_508_80 vgnd vpwr scs8hd_fill_1
XFILLER_591_74 vgnd vpwr scs8hd_decap_6
XFILLER_444_68 vgnd vpwr scs8hd_decap_12
XFILLER_313_39 vgnd vpwr scs8hd_decap_12
XFILLER_56_56 vgnd vpwr scs8hd_decap_12
XFILLER_243_80 vgnd vpwr scs8hd_fill_1
XFILLER_460_56 vgnd vpwr scs8hd_decap_12
XFILLER_179_3 vgnd vpwr scs8hd_decap_12
XFILLER_72_44 vgnd vpwr scs8hd_decap_12
XFILLER_346_3 vgnd vpwr scs8hd_decap_12
XPHY_143 vgnd vpwr scs8hd_decap_3
XPHY_132 vgnd vpwr scs8hd_decap_3
XPHY_121 vgnd vpwr scs8hd_decap_3
XPHY_110 vgnd vpwr scs8hd_decap_3
XFILLER_188_44 vgnd vpwr scs8hd_decap_12
XPHY_176 vgnd vpwr scs8hd_decap_3
XPHY_165 vgnd vpwr scs8hd_decap_3
XPHY_154 vgnd vpwr scs8hd_decap_3
XPHY_198 vgnd vpwr scs8hd_decap_3
XPHY_187 vgnd vpwr scs8hd_decap_3
XFILLER_513_3 vgnd vpwr scs8hd_decap_12
XFILLER_418_80 vgnd vpwr scs8hd_fill_1
XFILLER_97_74 vgnd vpwr scs8hd_decap_6
XFILLER_354_68 vgnd vpwr scs8hd_decap_12
XFILLER_504_27 vgnd vpwr scs8hd_decap_4
XFILLER_223_39 vgnd vpwr scs8hd_decap_12
XFILLER_153_80 vgnd vpwr scs8hd_fill_1
XFILLER_370_56 vgnd vpwr scs8hd_decap_12
XFILLER_520_15 vgnd vpwr scs8hd_decap_12
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_94_3 vgnd vpwr scs8hd_decap_12
XFILLER_328_80 vgnd vpwr scs8hd_fill_1
XFILLER_264_68 vgnd vpwr scs8hd_decap_12
XFILLER_414_27 vgnd vpwr scs8hd_decap_4
XFILLER_133_39 vgnd vpwr scs8hd_decap_12
XFILLER_280_56 vgnd vpwr scs8hd_decap_12
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
XFILLER_430_15 vgnd vpwr scs8hd_decap_12
XANTENNA__15__D address[2] vgnd vpwr scs8hd_diode_2
XFILLER_238_80 vgnd vpwr scs8hd_fill_1
XFILLER_174_68 vgnd vpwr scs8hd_decap_12
XFILLER_107_62 vgnd vpwr scs8hd_decap_12
XFILLER_107_51 vgnd vpwr scs8hd_decap_8
XFILLER_324_27 vgnd vpwr scs8hd_decap_4
XFILLER_296_3 vgnd vpwr scs8hd_decap_12
XFILLER_190_56 vgnd vpwr scs8hd_decap_12
XFILLER_340_15 vgnd vpwr scs8hd_decap_12
XFILLER_463_3 vgnd vpwr scs8hd_decap_12
XFILLER_199_43 vgnd vpwr scs8hd_decap_12
XFILLER_32_80 vgnd vpwr scs8hd_fill_1
XFILLER_148_80 vgnd vpwr scs8hd_fill_1
XFILLER_515_15 vgnd vpwr scs8hd_decap_12
XFILLER_515_59 vpwr vgnd scs8hd_fill_2
XFILLER_234_27 vgnd vpwr scs8hd_decap_4
XFILLER_250_15 vgnd vpwr scs8hd_decap_12
XFILLER_556_44 vgnd vpwr scs8hd_decap_12
XFILLER_409_27 vgnd vpwr scs8hd_decap_12
XFILLER_425_15 vgnd vpwr scs8hd_decap_12
XFILLER_572_32 vgnd vpwr scs8hd_decap_12
XFILLER_208_61 vgnd vpwr scs8hd_decap_12
XFILLER_425_59 vpwr vgnd scs8hd_fill_2
XFILLER_144_27 vgnd vpwr scs8hd_decap_4
XFILLER_160_15 vgnd vpwr scs8hd_decap_12
XFILLER_521_80 vgnd vpwr scs8hd_fill_1
XFILLER_597_62 vgnd vpwr scs8hd_decap_12
XFILLER_597_51 vgnd vpwr scs8hd_decap_8
XFILLER_319_27 vgnd vpwr scs8hd_decap_12
XFILLER_466_44 vgnd vpwr scs8hd_decap_12
XFILLER_211_3 vgnd vpwr scs8hd_decap_4
XFILLER_309_3 vgnd vpwr scs8hd_decap_12
XFILLER_335_15 vgnd vpwr scs8hd_decap_12
XFILLER_78_32 vgnd vpwr scs8hd_decap_12
XFILLER_335_59 vpwr vgnd scs8hd_fill_2
XFILLER_482_32 vgnd vpwr scs8hd_decap_12
XFILLER_580_3 vgnd vpwr scs8hd_decap_12
XFILLER_501_39 vgnd vpwr scs8hd_decap_12
XFILLER_27_80 vgnd vpwr scs8hd_fill_1
XFILLER_431_80 vgnd vpwr scs8hd_fill_1
XFILLER_229_27 vgnd vpwr scs8hd_decap_12
XFILLER_376_44 vgnd vpwr scs8hd_decap_12
XFILLER_57_3 vgnd vpwr scs8hd_decap_12
XFILLER_245_15 vgnd vpwr scs8hd_decap_12
XFILLER_392_32 vgnd vpwr scs8hd_decap_12
XFILLER_245_59 vpwr vgnd scs8hd_fill_2
XFILLER_542_68 vgnd vpwr scs8hd_decap_12
XFILLER_341_80 vgnd vpwr scs8hd_fill_1
XFILLER_411_39 vgnd vpwr scs8hd_decap_12
XPHY_709 vgnd vpwr scs8hd_decap_3
XPHY_1319 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1308 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_27 vgnd vpwr scs8hd_decap_12
XFILLER_139_27 vgnd vpwr scs8hd_decap_12
XFILLER_286_44 vgnd vpwr scs8hd_decap_12
XFILLER_155_15 vgnd vpwr scs8hd_decap_12
XFILLER_155_59 vpwr vgnd scs8hd_fill_2
XFILLER_516_80 vgnd vpwr scs8hd_fill_1
XFILLER_452_68 vgnd vpwr scs8hd_decap_12
XFILLER_602_27 vgnd vpwr scs8hd_decap_4
XFILLER_48_68 vgnd vpwr scs8hd_decap_12
XFILLER_251_80 vgnd vpwr scs8hd_fill_1
XFILLER_321_39 vgnd vpwr scs8hd_decap_12
XFILLER_64_56 vgnd vpwr scs8hd_decap_12
XFILLER_161_3 vgnd vpwr scs8hd_decap_12
XFILLER_259_3 vgnd vpwr scs8hd_decap_12
XFILLER_80_44 vgnd vpwr scs8hd_decap_12
XFILLER_426_3 vgnd vpwr scs8hd_decap_12
XFILLER_196_44 vgnd vpwr scs8hd_decap_12
XFILLER_426_80 vgnd vpwr scs8hd_fill_1
XFILLER_362_68 vgnd vpwr scs8hd_decap_12
XFILLER_512_27 vgnd vpwr scs8hd_decap_4
XFILLER_161_80 vgnd vpwr scs8hd_fill_1
XFILLER_231_39 vgnd vpwr scs8hd_decap_12
XFILLER_336_80 vgnd vpwr scs8hd_fill_1
XFILLER_272_68 vgnd vpwr scs8hd_decap_12
XFILLER_205_62 vgnd vpwr scs8hd_decap_12
XFILLER_422_27 vgnd vpwr scs8hd_decap_4
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XFILLER_141_39 vgnd vpwr scs8hd_decap_12
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XPHY_506 vgnd vpwr scs8hd_decap_3
XPHY_517 vgnd vpwr scs8hd_decap_3
XPHY_1105 vgnd vpwr scs8hd_decap_3
XPHY_528 vgnd vpwr scs8hd_decap_3
XPHY_539 vgnd vpwr scs8hd_decap_3
XPHY_1138 vgnd vpwr scs8hd_decap_3
XPHY_1127 vgnd vpwr scs8hd_decap_3
XPHY_1116 vgnd vpwr scs8hd_decap_3
XPHY_1149 vgnd vpwr scs8hd_decap_3
XFILLER_246_80 vgnd vpwr scs8hd_fill_1
XFILLER_182_68 vgnd vpwr scs8hd_decap_12
XFILLER_115_62 vgnd vpwr scs8hd_decap_12
XFILLER_115_51 vgnd vpwr scs8hd_decap_8
XFILLER_332_27 vgnd vpwr scs8hd_decap_4
XFILLER_376_3 vgnd vpwr scs8hd_decap_12
XFILLER_543_3 vgnd vpwr scs8hd_decap_12
XPHY_1650 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1661 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1672 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1683 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1694 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_507_27 vgnd vpwr scs8hd_decap_12
XFILLER_40_80 vgnd vpwr scs8hd_fill_1
XFILLER_156_80 vgnd vpwr scs8hd_fill_1
XFILLER_523_15 vgnd vpwr scs8hd_decap_12
XFILLER_523_59 vpwr vgnd scs8hd_fill_2
XFILLER_242_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_74 vgnd vpwr scs8hd_decap_6
XFILLER_548_56 vgnd vpwr scs8hd_decap_12
XFILLER_417_27 vgnd vpwr scs8hd_decap_12
XFILLER_564_44 vgnd vpwr scs8hd_decap_12
XFILLER_433_15 vgnd vpwr scs8hd_decap_12
XFILLER_580_32 vgnd vpwr scs8hd_decap_12
XFILLER_29_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_59 vpwr vgnd scs8hd_fill_2
XFILLER_152_27 vgnd vpwr scs8hd_decap_4
XFILLER_433_59 vpwr vgnd scs8hd_fill_2
XFILLER_589_74 vgnd vpwr scs8hd_decap_6
XPHY_303 vgnd vpwr scs8hd_decap_3
XPHY_314 vgnd vpwr scs8hd_decap_3
XPHY_325 vgnd vpwr scs8hd_decap_3
XPHY_336 vgnd vpwr scs8hd_decap_3
XPHY_347 vgnd vpwr scs8hd_decap_3
XPHY_358 vgnd vpwr scs8hd_decap_3
XPHY_369 vgnd vpwr scs8hd_decap_3
XFILLER_458_56 vgnd vpwr scs8hd_decap_12
XFILLER_124_3 vgnd vpwr scs8hd_decap_12
XFILLER_327_27 vgnd vpwr scs8hd_decap_12
XFILLER_474_44 vgnd vpwr scs8hd_decap_12
XFILLER_493_3 vgnd vpwr scs8hd_decap_12
XFILLER_343_15 vgnd vpwr scs8hd_decap_12
XFILLER_490_32 vgnd vpwr scs8hd_decap_12
XFILLER_86_32 vgnd vpwr scs8hd_decap_12
XFILLER_343_59 vpwr vgnd scs8hd_fill_2
XFILLER_499_74 vgnd vpwr scs8hd_decap_6
XFILLER_35_80 vgnd vpwr scs8hd_fill_1
XPHY_870 vgnd vpwr scs8hd_decap_3
XPHY_881 vgnd vpwr scs8hd_decap_3
XPHY_892 vgnd vpwr scs8hd_decap_3
XFILLER_518_15 vgnd vpwr scs8hd_decap_12
XFILLER_237_27 vgnd vpwr scs8hd_decap_12
XPHY_1480 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1491 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_384_44 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ right_width_0_height_0__pin_10_ logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[5] vgnd vpwr scs8hd_ebufn_1
XFILLER_253_15 vgnd vpwr scs8hd_decap_12
XFILLER_253_59 vpwr vgnd scs8hd_fill_2
XFILLER_550_68 vgnd vpwr scs8hd_decap_12
X_08_ address[2] _08_/Y vgnd vpwr scs8hd_inv_8
XFILLER_202_30 vgnd vpwr scs8hd_fill_1
XFILLER_15_39 vgnd vpwr scs8hd_decap_12
XFILLER_278_56 vgnd vpwr scs8hd_decap_12
XFILLER_428_15 vgnd vpwr scs8hd_decap_12
XFILLER_31_27 vgnd vpwr scs8hd_decap_12
XFILLER_147_27 vgnd vpwr scs8hd_decap_12
XFILLER_294_44 vgnd vpwr scs8hd_decap_12
XFILLER_163_15 vgnd vpwr scs8hd_decap_12
XFILLER_524_80 vgnd vpwr scs8hd_fill_1
XFILLER_163_59 vpwr vgnd scs8hd_fill_2
XFILLER_460_68 vgnd vpwr scs8hd_decap_12
XFILLER_56_68 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ right_width_0_height_0__pin_14_ vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_decap_3
XFILLER_72_56 vgnd vpwr scs8hd_decap_12
XPHY_133 vgnd vpwr scs8hd_decap_3
XPHY_122 vgnd vpwr scs8hd_decap_3
XPHY_111 vgnd vpwr scs8hd_decap_3
XFILLER_241_3 vgnd vpwr scs8hd_decap_12
XPHY_166 vgnd vpwr scs8hd_decap_3
XPHY_155 vgnd vpwr scs8hd_decap_3
XPHY_144 vgnd vpwr scs8hd_decap_3
XFILLER_188_56 vgnd vpwr scs8hd_decap_12
XFILLER_339_3 vgnd vpwr scs8hd_decap_12
XPHY_199 vgnd vpwr scs8hd_decap_3
XPHY_188 vgnd vpwr scs8hd_decap_3
XPHY_177 vgnd vpwr scs8hd_decap_3
XFILLER_338_15 vgnd vpwr scs8hd_decap_12
XFILLER_506_3 vgnd vpwr scs8hd_decap_12
XFILLER_434_80 vgnd vpwr scs8hd_fill_1
XFILLER_370_68 vgnd vpwr scs8hd_decap_12
XFILLER_303_51 vgnd vpwr scs8hd_decap_8
XFILLER_303_62 vgnd vpwr scs8hd_decap_12
XFILLER_520_27 vgnd vpwr scs8hd_decap_4
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_87_3 vgnd vpwr scs8hd_decap_12
XFILLER_248_15 vgnd vpwr scs8hd_decap_12
XFILLER_7_51 vgnd vpwr scs8hd_decap_8
XFILLER_7_62 vgnd vpwr scs8hd_decap_12
XFILLER_344_80 vgnd vpwr scs8hd_fill_1
XFILLER_280_68 vgnd vpwr scs8hd_decap_12
XFILLER_213_51 vgnd vpwr scs8hd_decap_8
XFILLER_213_62 vgnd vpwr scs8hd_decap_12
XFILLER_430_27 vgnd vpwr scs8hd_decap_4
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XFILLER_158_15 vgnd vpwr scs8hd_decap_12
XFILLER_519_80 vgnd vpwr scs8hd_fill_1
XFILLER_107_74 vgnd vpwr scs8hd_decap_6
XFILLER_254_80 vgnd vpwr scs8hd_fill_1
XFILLER_191_3 vgnd vpwr scs8hd_decap_12
XFILLER_190_68 vgnd vpwr scs8hd_decap_12
XFILLER_289_3 vgnd vpwr scs8hd_decap_12
XFILLER_123_62 vgnd vpwr scs8hd_decap_12
XFILLER_123_51 vgnd vpwr scs8hd_decap_8
XFILLER_340_27 vgnd vpwr scs8hd_decap_4
XFILLER_456_3 vgnd vpwr scs8hd_decap_12
XFILLER_199_55 vgnd vpwr scs8hd_decap_6
XFILLER_429_80 vgnd vpwr scs8hd_fill_1
XFILLER_515_27 vgnd vpwr scs8hd_decap_12
XFILLER_164_80 vgnd vpwr scs8hd_fill_1
XFILLER_531_15 vgnd vpwr scs8hd_decap_12
XFILLER_531_59 vpwr vgnd scs8hd_fill_2
XFILLER_250_27 vgnd vpwr scs8hd_decap_4
XFILLER_409_39 vgnd vpwr scs8hd_decap_12
XFILLER_556_56 vgnd vpwr scs8hd_decap_12
XFILLER_339_80 vgnd vpwr scs8hd_fill_1
XFILLER_572_44 vgnd vpwr scs8hd_decap_12
XFILLER_208_73 vgnd vpwr scs8hd_decap_8
XFILLER_425_27 vgnd vpwr scs8hd_decap_12
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XFILLER_441_15 vgnd vpwr scs8hd_decap_12
XFILLER_441_59 vpwr vgnd scs8hd_fill_2
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
XFILLER_160_27 vgnd vpwr scs8hd_decap_4
XFILLER_597_74 vgnd vpwr scs8hd_decap_6
XFILLER_249_80 vgnd vpwr scs8hd_fill_1
XFILLER_319_39 vgnd vpwr scs8hd_decap_12
XFILLER_466_56 vgnd vpwr scs8hd_decap_12
XFILLER_335_27 vgnd vpwr scs8hd_decap_12
XFILLER_482_44 vgnd vpwr scs8hd_decap_12
XFILLER_78_44 vgnd vpwr scs8hd_decap_12
XFILLER_573_3 vgnd vpwr scs8hd_decap_12
XFILLER_351_15 vgnd vpwr scs8hd_decap_12
XFILLER_94_32 vgnd vpwr scs8hd_decap_12
XFILLER_351_59 vpwr vgnd scs8hd_fill_2
XFILLER_43_80 vgnd vpwr scs8hd_fill_1
XFILLER_159_80 vgnd vpwr scs8hd_fill_1
XFILLER_229_39 vgnd vpwr scs8hd_decap_12
XFILLER_376_56 vgnd vpwr scs8hd_decap_12
XFILLER_526_15 vgnd vpwr scs8hd_decap_12
XFILLER_245_27 vgnd vpwr scs8hd_decap_12
XFILLER_392_44 vgnd vpwr scs8hd_decap_12
XFILLER_261_15 vgnd vpwr scs8hd_decap_12
XFILLER_261_59 vpwr vgnd scs8hd_fill_2
XFILLER_210_30 vgnd vpwr scs8hd_fill_1
XPHY_1309 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_39 vgnd vpwr scs8hd_decap_12
XFILLER_139_39 vgnd vpwr scs8hd_decap_12
XFILLER_286_56 vgnd vpwr scs8hd_decap_12
XFILLER_436_15 vgnd vpwr scs8hd_decap_12
XFILLER_155_27 vgnd vpwr scs8hd_decap_12
XFILLER_171_15 vgnd vpwr scs8hd_decap_12
XFILLER_171_59 vpwr vgnd scs8hd_fill_2
XFILLER_532_80 vgnd vpwr scs8hd_fill_1
XFILLER_64_68 vgnd vpwr scs8hd_decap_12
XFILLER_401_51 vgnd vpwr scs8hd_decap_8
XFILLER_154_3 vgnd vpwr scs8hd_decap_12
XFILLER_401_62 vgnd vpwr scs8hd_decap_12
XPHY_1810 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_80_56 vgnd vpwr scs8hd_decap_12
XFILLER_321_3 vgnd vpwr scs8hd_decap_12
XFILLER_196_56 vgnd vpwr scs8hd_decap_12
XFILLER_419_3 vgnd vpwr scs8hd_decap_12
XFILLER_346_15 vgnd vpwr scs8hd_decap_12
XFILLER_38_80 vgnd vpwr scs8hd_fill_1
XFILLER_442_80 vgnd vpwr scs8hd_fill_1
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ right_width_0_height_0__pin_10_ vgnd vpwr scs8hd_diode_2
XFILLER_311_51 vgnd vpwr scs8hd_decap_8
XFILLER_311_62 vgnd vpwr scs8hd_decap_12
XFILLER_256_15 vgnd vpwr scs8hd_decap_12
XFILLER_205_30 vgnd vpwr scs8hd_decap_12
XFILLER_205_74 vgnd vpwr scs8hd_decap_6
XFILLER_352_80 vgnd vpwr scs8hd_fill_1
XFILLER_221_51 vgnd vpwr scs8hd_decap_8
XFILLER_578_32 vgnd vpwr scs8hd_decap_12
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XFILLER_221_62 vgnd vpwr scs8hd_decap_12
XPHY_507 vgnd vpwr scs8hd_decap_3
XPHY_518 vgnd vpwr scs8hd_decap_3
XPHY_529 vgnd vpwr scs8hd_decap_3
XPHY_1139 vgnd vpwr scs8hd_decap_3
XPHY_1128 vgnd vpwr scs8hd_decap_3
XPHY_1117 vgnd vpwr scs8hd_decap_3
XPHY_1106 vgnd vpwr scs8hd_decap_3
XFILLER_50_15 vgnd vpwr scs8hd_decap_12
XFILLER_166_15 vgnd vpwr scs8hd_decap_12
XFILLER_527_80 vgnd vpwr scs8hd_fill_1
XFILLER_115_74 vgnd vpwr scs8hd_decap_6
XFILLER_262_80 vgnd vpwr scs8hd_fill_1
XFILLER_271_3 vgnd vpwr scs8hd_decap_12
XFILLER_369_3 vgnd vpwr scs8hd_decap_12
XFILLER_131_51 vgnd vpwr scs8hd_decap_8
XFILLER_131_62 vgnd vpwr scs8hd_decap_12
XFILLER_488_32 vgnd vpwr scs8hd_decap_12
XFILLER_536_3 vgnd vpwr scs8hd_decap_12
XPHY_1640 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1651 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1662 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1673 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1684 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1695 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_437_80 vgnd vpwr scs8hd_fill_1
XFILLER_507_39 vgnd vpwr scs8hd_decap_12
XFILLER_523_27 vgnd vpwr scs8hd_decap_12
XFILLER_172_80 vgnd vpwr scs8hd_fill_1
XFILLER_1_53 vgnd vpwr scs8hd_decap_8
XFILLER_398_32 vgnd vpwr scs8hd_decap_12
XFILLER_548_68 vgnd vpwr scs8hd_decap_12
XFILLER_564_56 vgnd vpwr scs8hd_decap_12
XFILLER_347_80 vgnd vpwr scs8hd_fill_1
XFILLER_417_39 vgnd vpwr scs8hd_decap_12
XFILLER_580_44 vgnd vpwr scs8hd_decap_12
XFILLER_433_27 vgnd vpwr scs8hd_decap_12
XFILLER_29_27 vgnd vpwr scs8hd_decap_12
XFILLER_45_15 vgnd vpwr scs8hd_decap_12
XFILLER_45_59 vpwr vgnd scs8hd_fill_2
XPHY_304 vgnd vpwr scs8hd_decap_3
XPHY_315 vgnd vpwr scs8hd_decap_3
XPHY_326 vgnd vpwr scs8hd_decap_3
XPHY_337 vgnd vpwr scs8hd_decap_3
XPHY_348 vgnd vpwr scs8hd_decap_3
XPHY_359 vgnd vpwr scs8hd_decap_3
XFILLER_458_68 vgnd vpwr scs8hd_decap_12
XFILLER_117_3 vgnd vpwr scs8hd_decap_12
XFILLER_257_80 vgnd vpwr scs8hd_fill_1
XFILLER_327_39 vgnd vpwr scs8hd_decap_12
XFILLER_474_56 vgnd vpwr scs8hd_decap_12
XFILLER_343_27 vgnd vpwr scs8hd_decap_12
XFILLER_490_44 vgnd vpwr scs8hd_decap_12
XFILLER_86_44 vgnd vpwr scs8hd_decap_12
XFILLER_486_3 vgnd vpwr scs8hd_decap_12
XFILLER_368_57 vgnd vpwr scs8hd_decap_12
XPHY_860 vgnd vpwr scs8hd_decap_3
XPHY_871 vgnd vpwr scs8hd_decap_3
XPHY_882 vgnd vpwr scs8hd_decap_3
XPHY_893 vgnd vpwr scs8hd_decap_3
XFILLER_518_27 vgnd vpwr scs8hd_decap_4
XFILLER_51_80 vgnd vpwr scs8hd_fill_1
XPHY_1470 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1481 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1492 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_167_80 vgnd vpwr scs8hd_fill_1
XFILLER_237_39 vgnd vpwr scs8hd_decap_12
XFILLER_384_56 vgnd vpwr scs8hd_decap_12
XFILLER_534_15 vgnd vpwr scs8hd_decap_12
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XFILLER_253_27 vgnd vpwr scs8hd_decap_12
X_07_ _07_/A address[2] _07_/C enable _07_/X vgnd vpwr scs8hd_and4_4
XFILLER_202_20 vpwr vgnd scs8hd_fill_2
XFILLER_278_68 vgnd vpwr scs8hd_decap_12
XFILLER_428_27 vgnd vpwr scs8hd_decap_4
XFILLER_31_39 vgnd vpwr scs8hd_decap_12
XFILLER_147_39 vgnd vpwr scs8hd_decap_12
XFILLER_294_56 vgnd vpwr scs8hd_decap_12
XFILLER_444_15 vgnd vpwr scs8hd_decap_12
XFILLER_163_27 vgnd vpwr scs8hd_decap_12
XFILLER_193_7 vgnd vpwr scs8hd_decap_12
XFILLER_540_80 vgnd vpwr scs8hd_fill_1
XFILLER_72_68 vgnd vpwr scs8hd_decap_12
XPHY_134 vgnd vpwr scs8hd_decap_3
XPHY_123 vgnd vpwr scs8hd_decap_3
XPHY_112 vgnd vpwr scs8hd_decap_3
XPHY_101 vgnd vpwr scs8hd_decap_3
XPHY_167 vgnd vpwr scs8hd_decap_3
XPHY_156 vgnd vpwr scs8hd_decap_3
XPHY_145 vgnd vpwr scs8hd_decap_3
XFILLER_188_68 vgnd vpwr scs8hd_decap_12
XFILLER_234_3 vgnd vpwr scs8hd_decap_12
XPHY_189 vgnd vpwr scs8hd_decap_3
XPHY_178 vgnd vpwr scs8hd_decap_3
XFILLER_338_27 vgnd vpwr scs8hd_decap_4
XFILLER_401_3 vgnd vpwr scs8hd_decap_12
XFILLER_354_15 vgnd vpwr scs8hd_decap_12
XFILLER_303_74 vgnd vpwr scs8hd_decap_6
XFILLER_450_80 vgnd vpwr scs8hd_fill_1
XFILLER_46_80 vgnd vpwr scs8hd_fill_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_529_15 vgnd vpwr scs8hd_decap_12
XFILLER_529_59 vpwr vgnd scs8hd_fill_2
XFILLER_248_27 vgnd vpwr scs8hd_decap_4
XPHY_690 vgnd vpwr scs8hd_decap_3
XFILLER_7_74 vgnd vpwr scs8hd_decap_6
XFILLER_264_15 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ right_width_0_height_0__pin_6_ vgnd vpwr scs8hd_diode_2
XFILLER_213_74 vgnd vpwr scs8hd_decap_6
XFILLER_360_80 vgnd vpwr scs8hd_fill_1
XFILLER_586_32 vgnd vpwr scs8hd_decap_12
XFILLER_439_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_158_27 vgnd vpwr scs8hd_decap_4
XFILLER_439_59 vpwr vgnd scs8hd_fill_2
XFILLER_206_7 vpwr vgnd scs8hd_fill_2
XFILLER_174_15 vgnd vpwr scs8hd_decap_12
XFILLER_535_80 vgnd vpwr scs8hd_fill_1
XFILLER_184_3 vgnd vpwr scs8hd_decap_12
XFILLER_123_74 vgnd vpwr scs8hd_decap_6
XFILLER_270_80 vgnd vpwr scs8hd_fill_1
XFILLER_351_3 vgnd vpwr scs8hd_decap_12
XFILLER_449_3 vgnd vpwr scs8hd_decap_12
XFILLER_349_15 vgnd vpwr scs8hd_decap_12
XFILLER_496_32 vgnd vpwr scs8hd_decap_12
XFILLER_349_59 vpwr vgnd scs8hd_fill_2
XFILLER_218_19 vgnd vpwr scs8hd_decap_12
XFILLER_445_80 vgnd vpwr scs8hd_fill_1
XFILLER_515_39 vgnd vpwr scs8hd_decap_12
XFILLER_531_27 vgnd vpwr scs8hd_decap_12
XFILLER_259_15 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_259_59 vpwr vgnd scs8hd_fill_2
XFILLER_556_68 vgnd vpwr scs8hd_decap_12
XFILLER_572_56 vgnd vpwr scs8hd_decap_12
XFILLER_355_80 vgnd vpwr scs8hd_fill_1
XFILLER_425_39 vgnd vpwr scs8hd_decap_12
XFILLER_441_27 vgnd vpwr scs8hd_decap_12
XFILLER_37_27 vgnd vpwr scs8hd_decap_12
XFILLER_53_15 vgnd vpwr scs8hd_decap_12
XFILLER_53_59 vpwr vgnd scs8hd_fill_2
XFILLER_169_15 vgnd vpwr scs8hd_decap_12
XFILLER_169_59 vpwr vgnd scs8hd_fill_2
XFILLER_466_68 vgnd vpwr scs8hd_decap_12
XFILLER_265_80 vgnd vpwr scs8hd_fill_1
XFILLER_335_39 vgnd vpwr scs8hd_decap_12
XFILLER_78_56 vgnd vpwr scs8hd_decap_12
XFILLER_482_56 vgnd vpwr scs8hd_decap_12
XFILLER_399_3 vgnd vpwr scs8hd_decap_12
XFILLER_351_27 vgnd vpwr scs8hd_decap_12
XFILLER_566_3 vgnd vpwr scs8hd_decap_12
XFILLER_94_44 vgnd vpwr scs8hd_decap_12
XFILLER_376_68 vgnd vpwr scs8hd_decap_12
XFILLER_526_27 vgnd vpwr scs8hd_decap_4
XFILLER_309_51 vgnd vpwr scs8hd_decap_8
XFILLER_309_62 vgnd vpwr scs8hd_decap_12
XFILLER_175_80 vgnd vpwr scs8hd_fill_1
XFILLER_245_39 vgnd vpwr scs8hd_decap_12
XFILLER_392_56 vgnd vpwr scs8hd_decap_12
XFILLER_542_15 vgnd vpwr scs8hd_decap_12
XFILLER_261_27 vgnd vpwr scs8hd_decap_12
XFILLER_286_68 vgnd vpwr scs8hd_decap_12
XFILLER_219_62 vgnd vpwr scs8hd_decap_12
XFILLER_436_27 vgnd vpwr scs8hd_decap_4
XFILLER_155_39 vgnd vpwr scs8hd_decap_12
XFILLER_48_15 vgnd vpwr scs8hd_decap_12
XFILLER_452_15 vgnd vpwr scs8hd_decap_12
XFILLER_171_27 vgnd vpwr scs8hd_decap_12
XFILLER_104_32 vgnd vpwr scs8hd_decap_12
XFILLER_401_74 vgnd vpwr scs8hd_decap_6
XPHY_1800 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_147_3 vgnd vpwr scs8hd_decap_12
XPHY_1811 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_80_68 vgnd vpwr scs8hd_decap_12
XFILLER_13_51 vgnd vpwr scs8hd_decap_8
XFILLER_129_51 vgnd vpwr scs8hd_decap_8
XFILLER_13_62 vgnd vpwr scs8hd_decap_12
XFILLER_196_68 vgnd vpwr scs8hd_decap_12
XFILLER_314_3 vgnd vpwr scs8hd_decap_12
XFILLER_129_62 vgnd vpwr scs8hd_decap_12
XFILLER_346_27 vgnd vpwr scs8hd_decap_4
XFILLER_362_15 vgnd vpwr scs8hd_decap_12
XFILLER_311_74 vgnd vpwr scs8hd_decap_6
XFILLER_54_80 vgnd vpwr scs8hd_fill_1
XFILLER_537_15 vgnd vpwr scs8hd_decap_12
XFILLER_537_59 vpwr vgnd scs8hd_fill_2
XFILLER_62_3 vgnd vpwr scs8hd_decap_12
XFILLER_256_27 vgnd vpwr scs8hd_decap_4
XFILLER_272_15 vgnd vpwr scs8hd_decap_12
XFILLER_205_42 vgnd vpwr scs8hd_decap_12
XFILLER_578_44 vgnd vpwr scs8hd_decap_12
XFILLER_221_74 vgnd vpwr scs8hd_decap_6
XPHY_508 vgnd vpwr scs8hd_decap_3
XPHY_519 vgnd vpwr scs8hd_decap_3
XPHY_1129 vgnd vpwr scs8hd_decap_3
XPHY_1118 vgnd vpwr scs8hd_decap_3
XPHY_1107 vgnd vpwr scs8hd_decap_3
XFILLER_594_32 vgnd vpwr scs8hd_decap_12
XFILLER_447_15 vgnd vpwr scs8hd_decap_12
XFILLER_50_27 vgnd vpwr scs8hd_decap_4
XFILLER_447_59 vpwr vgnd scs8hd_fill_2
XFILLER_166_27 vgnd vpwr scs8hd_decap_4
XFILLER_182_15 vgnd vpwr scs8hd_decap_12
XFILLER_543_80 vgnd vpwr scs8hd_fill_1
XFILLER_264_3 vgnd vpwr scs8hd_decap_12
XFILLER_131_74 vgnd vpwr scs8hd_decap_6
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ right_width_0_height_0__pin_2_ vgnd vpwr scs8hd_diode_2
XFILLER_488_44 vgnd vpwr scs8hd_decap_12
XFILLER_431_3 vgnd vpwr scs8hd_decap_12
XFILLER_529_3 vgnd vpwr scs8hd_decap_12
XFILLER_357_15 vgnd vpwr scs8hd_decap_12
XPHY_1630 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1641 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1652 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_357_59 vpwr vgnd scs8hd_fill_2
XPHY_1663 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1674 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1685 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1696 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_523_39 vgnd vpwr scs8hd_decap_12
XFILLER_453_80 vgnd vpwr scs8hd_fill_1
XFILLER_49_80 vgnd vpwr scs8hd_fill_1
X_23_ gfpga_pad_GPIO_PAD[4] right_width_0_height_0__pin_9_ vgnd vpwr scs8hd_buf_2
XFILLER_398_44 vgnd vpwr scs8hd_decap_12
XFILLER_267_15 vgnd vpwr scs8hd_decap_12
XFILLER_267_59 vpwr vgnd scs8hd_fill_2
XFILLER_564_68 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _12_/Y vgnd vpwr scs8hd_diode_2
XFILLER_433_39 vgnd vpwr scs8hd_decap_12
XFILLER_580_56 vgnd vpwr scs8hd_decap_12
XFILLER_29_39 vgnd vpwr scs8hd_decap_12
XFILLER_363_80 vgnd vpwr scs8hd_fill_1
XFILLER_45_27 vgnd vpwr scs8hd_decap_12
XFILLER_232_73 vgnd vpwr scs8hd_decap_8
XPHY_305 vgnd vpwr scs8hd_decap_3
XPHY_316 vgnd vpwr scs8hd_decap_3
XFILLER_61_15 vgnd vpwr scs8hd_decap_12
XPHY_327 vgnd vpwr scs8hd_decap_3
XPHY_338 vgnd vpwr scs8hd_decap_3
XPHY_349 vgnd vpwr scs8hd_decap_3
XFILLER_61_59 vpwr vgnd scs8hd_fill_2
XFILLER_177_15 vgnd vpwr scs8hd_decap_12
XFILLER_177_59 vpwr vgnd scs8hd_fill_2
XFILLER_538_80 vgnd vpwr scs8hd_fill_1
XFILLER_407_51 vgnd vpwr scs8hd_decap_8
XFILLER_474_68 vgnd vpwr scs8hd_decap_12
XFILLER_407_62 vgnd vpwr scs8hd_decap_12
XFILLER_343_39 vgnd vpwr scs8hd_decap_12
XFILLER_86_56 vgnd vpwr scs8hd_decap_12
XFILLER_273_80 vgnd vpwr scs8hd_fill_1
XFILLER_490_56 vgnd vpwr scs8hd_decap_12
XFILLER_381_3 vgnd vpwr scs8hd_decap_12
XFILLER_479_3 vgnd vpwr scs8hd_decap_12
XFILLER_368_69 vgnd vpwr scs8hd_decap_12
XPHY_850 vgnd vpwr scs8hd_decap_3
XPHY_861 vgnd vpwr scs8hd_decap_3
XPHY_872 vgnd vpwr scs8hd_decap_3
XPHY_1460 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_883 vgnd vpwr scs8hd_decap_3
XPHY_894 vgnd vpwr scs8hd_decap_3
XPHY_1471 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1482 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1493 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_448_80 vgnd vpwr scs8hd_fill_1
XFILLER_384_68 vgnd vpwr scs8hd_decap_12
XFILLER_534_27 vgnd vpwr scs8hd_decap_4
XFILLER_317_51 vgnd vpwr scs8hd_decap_8
XFILLER_317_62 vgnd vpwr scs8hd_decap_12
XFILLER_183_80 vgnd vpwr scs8hd_fill_1
XFILLER_253_39 vgnd vpwr scs8hd_decap_12
XFILLER_550_15 vgnd vpwr scs8hd_decap_12
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
X_06_ address[1] _07_/C vgnd vpwr scs8hd_inv_8
XFILLER_202_32 vgnd vpwr scs8hd_decap_12
XFILLER_358_80 vgnd vpwr scs8hd_fill_1
XFILLER_294_68 vgnd vpwr scs8hd_decap_12
XFILLER_227_51 vgnd vpwr scs8hd_decap_8
XFILLER_227_62 vgnd vpwr scs8hd_decap_12
XFILLER_444_27 vgnd vpwr scs8hd_decap_4
XFILLER_163_39 vgnd vpwr scs8hd_decap_12
XFILLER_460_15 vgnd vpwr scs8hd_decap_12
XFILLER_56_15 vgnd vpwr scs8hd_decap_12
XFILLER_112_32 vgnd vpwr scs8hd_decap_12
XPHY_124 vgnd vpwr scs8hd_decap_3
XPHY_113 vgnd vpwr scs8hd_decap_3
XPHY_102 vgnd vpwr scs8hd_decap_3
XPHY_157 vgnd vpwr scs8hd_decap_3
XPHY_146 vgnd vpwr scs8hd_decap_3
XPHY_135 vgnd vpwr scs8hd_decap_3
XPHY_179 vgnd vpwr scs8hd_decap_3
XPHY_168 vgnd vpwr scs8hd_decap_3
XFILLER_227_3 vgnd vpwr scs8hd_decap_12
XFILLER_268_80 vgnd vpwr scs8hd_fill_1
XFILLER_21_51 vgnd vpwr scs8hd_decap_8
XFILLER_21_62 vgnd vpwr scs8hd_decap_12
XFILLER_137_51 vgnd vpwr scs8hd_decap_8
XFILLER_137_62 vgnd vpwr scs8hd_decap_12
XFILLER_354_27 vgnd vpwr scs8hd_decap_4
XFILLER_596_3 vgnd vpwr scs8hd_decap_12
XFILLER_370_15 vgnd vpwr scs8hd_decap_12
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_529_27 vgnd vpwr scs8hd_decap_12
XFILLER_62_80 vgnd vpwr scs8hd_fill_1
XPHY_680 vgnd vpwr scs8hd_decap_3
XFILLER_178_80 vgnd vpwr scs8hd_fill_1
XPHY_691 vgnd vpwr scs8hd_decap_3
XFILLER_545_15 vgnd vpwr scs8hd_decap_12
XPHY_1290 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_545_59 vpwr vgnd scs8hd_fill_2
XFILLER_264_27 vgnd vpwr scs8hd_decap_4
XFILLER_280_15 vgnd vpwr scs8hd_decap_12
XFILLER_439_27 vgnd vpwr scs8hd_decap_12
XFILLER_586_44 vgnd vpwr scs8hd_decap_12
XFILLER_455_15 vgnd vpwr scs8hd_decap_12
XFILLER_174_27 vgnd vpwr scs8hd_decap_4
XFILLER_455_59 vpwr vgnd scs8hd_fill_2
XFILLER_190_15 vgnd vpwr scs8hd_decap_4
XFILLER_551_80 vgnd vpwr scs8hd_fill_1
XFILLER_177_3 vgnd vpwr scs8hd_decap_12
XFILLER_344_3 vgnd vpwr scs8hd_decap_12
XFILLER_349_27 vgnd vpwr scs8hd_decap_12
XFILLER_496_44 vgnd vpwr scs8hd_decap_12
XFILLER_511_3 vgnd vpwr scs8hd_decap_12
XFILLER_365_15 vgnd vpwr scs8hd_decap_12
XFILLER_365_59 vpwr vgnd scs8hd_fill_2
XFILLER_531_39 vgnd vpwr scs8hd_decap_12
XFILLER_57_80 vgnd vpwr scs8hd_fill_1
XFILLER_461_80 vgnd vpwr scs8hd_fill_1
XFILLER_259_27 vgnd vpwr scs8hd_decap_12
XFILLER_92_3 vgnd vpwr scs8hd_decap_12
XFILLER_275_15 vgnd vpwr scs8hd_decap_12
XFILLER_275_59 vpwr vgnd scs8hd_fill_2
XFILLER_572_68 vgnd vpwr scs8hd_decap_12
XFILLER_505_51 vgnd vpwr scs8hd_decap_8
XFILLER_505_62 vgnd vpwr scs8hd_decap_12
XFILLER_37_39 vgnd vpwr scs8hd_decap_12
XFILLER_371_80 vgnd vpwr scs8hd_fill_1
XFILLER_441_39 vgnd vpwr scs8hd_decap_12
XFILLER_53_27 vgnd vpwr scs8hd_decap_12
XFILLER_169_27 vgnd vpwr scs8hd_decap_12
XFILLER_185_15 vgnd vpwr scs8hd_decap_3
XFILLER_546_80 vgnd vpwr scs8hd_fill_1
XFILLER_482_68 vgnd vpwr scs8hd_decap_12
XFILLER_78_68 vgnd vpwr scs8hd_decap_12
XFILLER_415_51 vgnd vpwr scs8hd_decap_8
XFILLER_415_62 vgnd vpwr scs8hd_decap_12
XFILLER_294_3 vgnd vpwr scs8hd_decap_12
XFILLER_281_80 vgnd vpwr scs8hd_fill_1
XFILLER_351_39 vgnd vpwr scs8hd_decap_12
XFILLER_559_3 vgnd vpwr scs8hd_decap_12
XFILLER_94_56 vgnd vpwr scs8hd_decap_12
XFILLER_461_3 vgnd vpwr scs8hd_decap_12
XFILLER_300_32 vgnd vpwr scs8hd_decap_12
XFILLER_309_74 vgnd vpwr scs8hd_decap_6
XFILLER_456_80 vgnd vpwr scs8hd_fill_1
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XFILLER_392_68 vgnd vpwr scs8hd_decap_12
XFILLER_542_27 vgnd vpwr scs8hd_decap_4
XFILLER_325_51 vgnd vpwr scs8hd_decap_8
XFILLER_325_62 vgnd vpwr scs8hd_decap_12
XFILLER_191_80 vgnd vpwr scs8hd_fill_1
XFILLER_261_39 vgnd vpwr scs8hd_decap_12
XFILLER_210_32 vgnd vpwr scs8hd_decap_12
XFILLER_219_41 vgnd vpwr scs8hd_decap_12
XFILLER_219_74 vgnd vpwr scs8hd_decap_6
XFILLER_366_80 vgnd vpwr scs8hd_fill_1
XFILLER_235_51 vgnd vpwr scs8hd_decap_8
XFILLER_235_62 vgnd vpwr scs8hd_decap_12
XFILLER_452_27 vgnd vpwr scs8hd_decap_4
XFILLER_48_27 vgnd vpwr scs8hd_decap_4
XFILLER_171_39 vgnd vpwr scs8hd_decap_12
XFILLER_104_44 vgnd vpwr scs8hd_decap_12
XFILLER_64_15 vgnd vpwr scs8hd_decap_12
XFILLER_120_32 vgnd vpwr scs8hd_decap_12
XPHY_1801 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1812 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_196_14 vpwr vgnd scs8hd_fill_2
XFILLER_13_74 vgnd vpwr scs8hd_decap_6
XFILLER_129_74 vgnd vpwr scs8hd_decap_6
XFILLER_276_80 vgnd vpwr scs8hd_fill_1
XFILLER_307_3 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_145_51 vgnd vpwr scs8hd_decap_8
XFILLER_145_62 vgnd vpwr scs8hd_decap_12
XFILLER_362_27 vgnd vpwr scs8hd_decap_4
XFILLER_537_27 vgnd vpwr scs8hd_decap_12
XFILLER_70_80 vgnd vpwr scs8hd_fill_1
XFILLER_186_80 vgnd vpwr scs8hd_fill_1
XFILLER_55_3 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _05_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_553_15 vgnd vpwr scs8hd_decap_12
XFILLER_553_59 vpwr vgnd scs8hd_fill_2
XFILLER_272_27 vgnd vpwr scs8hd_decap_4
XFILLER_205_54 vgnd vpwr scs8hd_decap_6
XFILLER_578_56 vgnd vpwr scs8hd_decap_12
XPHY_509 vgnd vpwr scs8hd_decap_3
XPHY_1119 vgnd vpwr scs8hd_decap_3
XPHY_1108 vgnd vpwr scs8hd_decap_3
XFILLER_447_27 vgnd vpwr scs8hd_decap_12
XFILLER_594_44 vgnd vpwr scs8hd_decap_12
XFILLER_59_15 vgnd vpwr scs8hd_decap_12
XFILLER_463_15 vgnd vpwr scs8hd_decap_12
XFILLER_59_59 vpwr vgnd scs8hd_fill_2
XFILLER_182_27 vgnd vpwr scs8hd_decap_4
XFILLER_463_59 vpwr vgnd scs8hd_fill_2
XFILLER_257_3 vgnd vpwr scs8hd_decap_12
XFILLER_488_56 vgnd vpwr scs8hd_decap_12
XPHY_1620 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1631 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_424_3 vgnd vpwr scs8hd_decap_12
XPHY_1642 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_357_27 vgnd vpwr scs8hd_decap_12
XPHY_1653 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1664 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1675 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1686 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1697 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_373_15 vgnd vpwr scs8hd_decap_12
XFILLER_373_59 vpwr vgnd scs8hd_fill_2
X_22_ gfpga_pad_GPIO_PAD[3] right_width_0_height_0__pin_7_ vgnd vpwr scs8hd_buf_2
XFILLER_65_80 vgnd vpwr scs8hd_fill_1
XFILLER_398_56 vgnd vpwr scs8hd_decap_12
XFILLER_548_15 vgnd vpwr scs8hd_decap_12
XFILLER_267_27 vgnd vpwr scs8hd_decap_12
XFILLER_283_15 vgnd vpwr scs8hd_decap_12
XFILLER_283_59 vpwr vgnd scs8hd_fill_2
XFILLER_580_68 vgnd vpwr scs8hd_decap_12
XFILLER_513_51 vgnd vpwr scs8hd_decap_8
XFILLER_513_62 vgnd vpwr scs8hd_decap_12
XFILLER_45_39 vgnd vpwr scs8hd_decap_12
XPHY_306 vgnd vpwr scs8hd_decap_3
XPHY_317 vgnd vpwr scs8hd_decap_3
XPHY_328 vgnd vpwr scs8hd_decap_3
XPHY_339 vgnd vpwr scs8hd_decap_3
XFILLER_458_15 vgnd vpwr scs8hd_decap_12
XFILLER_61_27 vgnd vpwr scs8hd_decap_12
XFILLER_177_27 vgnd vpwr scs8hd_decap_12
XFILLER_554_80 vgnd vpwr scs8hd_fill_1
XFILLER_407_74 vgnd vpwr scs8hd_decap_6
XFILLER_490_68 vgnd vpwr scs8hd_decap_12
XFILLER_86_68 vgnd vpwr scs8hd_decap_12
XFILLER_423_51 vgnd vpwr scs8hd_decap_8
XFILLER_423_62 vgnd vpwr scs8hd_decap_12
XFILLER_19_51 vgnd vpwr scs8hd_decap_8
XFILLER_19_62 vgnd vpwr scs8hd_decap_12
XFILLER_374_3 vgnd vpwr scs8hd_decap_12
XFILLER_541_3 vgnd vpwr scs8hd_decap_12
XFILLER_368_15 vgnd vpwr scs8hd_decap_12
XFILLER_368_48 vgnd vpwr scs8hd_fill_1
XPHY_840 vgnd vpwr scs8hd_decap_3
XPHY_851 vgnd vpwr scs8hd_decap_3
XPHY_862 vgnd vpwr scs8hd_decap_3
XPHY_1450 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_873 vgnd vpwr scs8hd_decap_3
XPHY_884 vgnd vpwr scs8hd_decap_3
XPHY_895 vgnd vpwr scs8hd_decap_3
XPHY_1461 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1472 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1483 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1494 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_317_74 vgnd vpwr scs8hd_decap_6
XFILLER_464_80 vgnd vpwr scs8hd_fill_1
XFILLER_550_27 vgnd vpwr scs8hd_decap_4
XFILLER_333_51 vgnd vpwr scs8hd_decap_8
XFILLER_333_62 vgnd vpwr scs8hd_decap_12
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
X_05_ _07_/A address[2] address[1] enable _05_/X vgnd vpwr scs8hd_and4_4
XFILLER_202_44 vgnd vpwr scs8hd_decap_12
XFILLER_278_15 vgnd vpwr scs8hd_decap_12
XFILLER_227_74 vgnd vpwr scs8hd_decap_6
XFILLER_374_80 vgnd vpwr scs8hd_fill_1
XFILLER_243_51 vgnd vpwr scs8hd_decap_8
XFILLER_460_27 vgnd vpwr scs8hd_decap_4
XFILLER_56_27 vgnd vpwr scs8hd_decap_4
XFILLER_243_62 vgnd vpwr scs8hd_decap_12
XFILLER_112_44 vgnd vpwr scs8hd_decap_12
XFILLER_72_15 vgnd vpwr scs8hd_decap_12
XPHY_125 vgnd vpwr scs8hd_decap_3
XPHY_114 vgnd vpwr scs8hd_decap_3
XPHY_103 vgnd vpwr scs8hd_decap_3
XFILLER_188_15 vgnd vpwr scs8hd_decap_4
XPHY_158 vgnd vpwr scs8hd_decap_3
XPHY_147 vgnd vpwr scs8hd_decap_3
XPHY_136 vgnd vpwr scs8hd_decap_3
XFILLER_549_80 vgnd vpwr scs8hd_fill_1
XPHY_169 vgnd vpwr scs8hd_decap_3
XFILLER_122_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_74 vgnd vpwr scs8hd_decap_6
XFILLER_137_74 vgnd vpwr scs8hd_decap_6
XFILLER_284_80 vgnd vpwr scs8hd_fill_1
XFILLER_589_3 vgnd vpwr scs8hd_decap_12
XFILLER_491_3 vgnd vpwr scs8hd_decap_12
XFILLER_153_51 vgnd vpwr scs8hd_decap_8
XFILLER_153_62 vgnd vpwr scs8hd_decap_12
XFILLER_370_27 vgnd vpwr scs8hd_decap_4
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_529_39 vgnd vpwr scs8hd_decap_12
XPHY_670 vgnd vpwr scs8hd_decap_3
XFILLER_459_80 vgnd vpwr scs8hd_fill_1
XPHY_681 vgnd vpwr scs8hd_decap_3
XPHY_692 vgnd vpwr scs8hd_decap_3
XPHY_1291 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_545_27 vgnd vpwr scs8hd_decap_12
XFILLER_194_80 vgnd vpwr scs8hd_fill_1
XFILLER_561_15 vgnd vpwr scs8hd_decap_12
XFILLER_561_59 vpwr vgnd scs8hd_fill_2
XFILLER_280_27 vgnd vpwr scs8hd_decap_4
XFILLER_586_56 vgnd vpwr scs8hd_decap_12
XFILLER_369_80 vgnd vpwr scs8hd_fill_1
XFILLER_439_39 vgnd vpwr scs8hd_decap_12
XFILLER_455_27 vgnd vpwr scs8hd_decap_12
XFILLER_471_15 vgnd vpwr scs8hd_decap_12
XFILLER_67_15 vgnd vpwr scs8hd_decap_12
XFILLER_471_59 vpwr vgnd scs8hd_fill_2
XFILLER_67_59 vpwr vgnd scs8hd_fill_2
XFILLER_279_80 vgnd vpwr scs8hd_fill_1
XFILLER_337_3 vgnd vpwr scs8hd_decap_12
XFILLER_349_39 vgnd vpwr scs8hd_decap_12
XFILLER_496_56 vgnd vpwr scs8hd_decap_12
XFILLER_504_3 vgnd vpwr scs8hd_decap_12
XFILLER_365_27 vgnd vpwr scs8hd_decap_12
XFILLER_381_15 vgnd vpwr scs8hd_decap_12
XFILLER_381_59 vpwr vgnd scs8hd_fill_2
XFILLER_73_80 vgnd vpwr scs8hd_fill_1
XFILLER_189_80 vgnd vpwr scs8hd_fill_1
XFILLER_259_39 vgnd vpwr scs8hd_decap_12
XFILLER_556_15 vgnd vpwr scs8hd_decap_12
XFILLER_85_3 vgnd vpwr scs8hd_decap_12
XFILLER_275_27 vgnd vpwr scs8hd_decap_12
XFILLER_208_32 vgnd vpwr scs8hd_decap_3
XFILLER_291_15 vgnd vpwr scs8hd_decap_12
XFILLER_291_59 vpwr vgnd scs8hd_fill_2
XFILLER_505_74 vgnd vpwr scs8hd_decap_6
XFILLER_521_51 vgnd vpwr scs8hd_decap_8
XFILLER_521_62 vgnd vpwr scs8hd_decap_12
XFILLER_53_39 vgnd vpwr scs8hd_decap_12
XFILLER_169_39 vgnd vpwr scs8hd_decap_12
XFILLER_466_15 vgnd vpwr scs8hd_decap_12
XFILLER_211_7 vgnd vpwr scs8hd_fill_1
XFILLER_118_32 vgnd vpwr scs8hd_decap_12
XFILLER_562_80 vgnd vpwr scs8hd_fill_1
XFILLER_415_74 vgnd vpwr scs8hd_decap_6
XFILLER_287_3 vgnd vpwr scs8hd_decap_12
XFILLER_94_68 vgnd vpwr scs8hd_decap_12
XFILLER_431_51 vgnd vpwr scs8hd_decap_8
XFILLER_27_51 vgnd vpwr scs8hd_decap_8
XFILLER_27_62 vgnd vpwr scs8hd_decap_12
XFILLER_431_62 vgnd vpwr scs8hd_decap_12
XFILLER_454_3 vgnd vpwr scs8hd_decap_12
XFILLER_300_44 vgnd vpwr scs8hd_decap_12
XFILLER_376_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XFILLER_68_80 vgnd vpwr scs8hd_fill_1
XFILLER_325_74 vgnd vpwr scs8hd_decap_6
XFILLER_472_80 vgnd vpwr scs8hd_fill_1
XFILLER_341_51 vgnd vpwr scs8hd_decap_8
XFILLER_341_62 vgnd vpwr scs8hd_decap_12
XFILLER_210_22 vpwr vgnd scs8hd_fill_2
XFILLER_210_44 vgnd vpwr scs8hd_decap_12
XFILLER_286_15 vgnd vpwr scs8hd_decap_12
XFILLER_219_53 vgnd vpwr scs8hd_decap_8
XFILLER_235_74 vgnd vpwr scs8hd_decap_6
XFILLER_382_80 vgnd vpwr scs8hd_fill_1
XFILLER_104_56 vgnd vpwr scs8hd_decap_12
XFILLER_64_27 vgnd vpwr scs8hd_decap_4
XFILLER_251_51 vgnd vpwr scs8hd_decap_8
XFILLER_251_62 vgnd vpwr scs8hd_decap_12
XFILLER_120_44 vgnd vpwr scs8hd_decap_12
XPHY_1813 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1802 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_80_15 vgnd vpwr scs8hd_decap_12
XFILLER_557_80 vgnd vpwr scs8hd_fill_1
XFILLER_145_74 vgnd vpwr scs8hd_decap_6
XFILLER_292_80 vgnd vpwr scs8hd_fill_1
XFILLER_571_3 vgnd vpwr scs8hd_decap_12
XFILLER_161_51 vgnd vpwr scs8hd_decap_8
XFILLER_161_62 vgnd vpwr scs8hd_decap_12
XFILLER_537_39 vgnd vpwr scs8hd_decap_12
XFILLER_467_80 vgnd vpwr scs8hd_fill_1
XFILLER_553_27 vgnd vpwr scs8hd_decap_12
XFILLER_48_3 vgnd vpwr scs8hd_decap_12
XFILLER_205_22 vpwr vgnd scs8hd_fill_2
XFILLER_578_68 vgnd vpwr scs8hd_decap_12
XPHY_1109 vgnd vpwr scs8hd_decap_3
XFILLER_594_56 vgnd vpwr scs8hd_decap_12
XFILLER_377_80 vgnd vpwr scs8hd_fill_1
XFILLER_447_39 vgnd vpwr scs8hd_decap_12
XFILLER_463_27 vgnd vpwr scs8hd_decap_12
XFILLER_59_27 vgnd vpwr scs8hd_decap_12
XFILLER_75_15 vgnd vpwr scs8hd_decap_12
XFILLER_75_59 vpwr vgnd scs8hd_fill_2
XFILLER_152_3 vgnd vpwr scs8hd_decap_12
XFILLER_488_68 vgnd vpwr scs8hd_decap_12
XPHY_1610 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1621 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1632 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1643 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_287_80 vgnd vpwr scs8hd_fill_1
XFILLER_357_39 vgnd vpwr scs8hd_decap_12
XFILLER_417_3 vgnd vpwr scs8hd_decap_12
XPHY_1654 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1665 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1676 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1687 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1698 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_373_27 vgnd vpwr scs8hd_decap_12
XFILLER_306_32 vgnd vpwr scs8hd_decap_12
XFILLER_603_63 vgnd vpwr scs8hd_decap_12
X_21_ gfpga_pad_GPIO_PAD[2] right_width_0_height_0__pin_5_ vgnd vpwr scs8hd_buf_2
XFILLER_398_68 vgnd vpwr scs8hd_decap_12
XFILLER_548_27 vgnd vpwr scs8hd_decap_4
XFILLER_81_80 vgnd vpwr scs8hd_fill_1
XFILLER_197_80 vgnd vpwr scs8hd_fill_1
XFILLER_267_39 vgnd vpwr scs8hd_decap_12
XFILLER_564_15 vgnd vpwr scs8hd_decap_12
XFILLER_283_27 vgnd vpwr scs8hd_decap_12
XFILLER_216_32 vgnd vpwr scs8hd_decap_12
XFILLER_513_74 vgnd vpwr scs8hd_decap_6
XPHY_307 vgnd vpwr scs8hd_decap_3
XPHY_318 vgnd vpwr scs8hd_decap_3
XPHY_329 vgnd vpwr scs8hd_decap_3
XFILLER_458_27 vgnd vpwr scs8hd_decap_4
XFILLER_61_39 vgnd vpwr scs8hd_decap_12
XFILLER_177_39 vgnd vpwr scs8hd_decap_12
XFILLER_474_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_126_32 vgnd vpwr scs8hd_decap_12
XFILLER_570_80 vgnd vpwr scs8hd_fill_1
XFILLER_19_74 vgnd vpwr scs8hd_decap_6
XFILLER_423_74 vgnd vpwr scs8hd_decap_6
XFILLER_367_3 vgnd vpwr scs8hd_decap_12
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
XFILLER_534_3 vgnd vpwr scs8hd_decap_12
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
XFILLER_368_27 vgnd vpwr scs8hd_decap_4
XPHY_830 vgnd vpwr scs8hd_decap_3
XPHY_841 vgnd vpwr scs8hd_decap_3
XPHY_852 vgnd vpwr scs8hd_decap_3
XPHY_863 vgnd vpwr scs8hd_decap_3
Xlogical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _13_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_1440 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1451 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_874 vgnd vpwr scs8hd_decap_3
XPHY_885 vgnd vpwr scs8hd_decap_3
XPHY_896 vgnd vpwr scs8hd_decap_3
XPHY_1462 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1473 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1484 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1495 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_384_15 vgnd vpwr scs8hd_decap_12
XFILLER_333_74 vgnd vpwr scs8hd_decap_6
XFILLER_480_80 vgnd vpwr scs8hd_fill_1
XFILLER_76_80 vgnd vpwr scs8hd_fill_1
X_04_ address[3] _07_/A vgnd vpwr scs8hd_buf_1
XFILLER_559_15 vgnd vpwr scs8hd_decap_12
XFILLER_202_56 vgnd vpwr scs8hd_decap_12
XFILLER_559_59 vpwr vgnd scs8hd_fill_2
XFILLER_278_27 vgnd vpwr scs8hd_decap_4
XFILLER_294_15 vgnd vpwr scs8hd_decap_12
XFILLER_243_74 vgnd vpwr scs8hd_decap_6
XFILLER_390_80 vgnd vpwr scs8hd_fill_1
XFILLER_112_56 vgnd vpwr scs8hd_decap_12
XFILLER_469_15 vgnd vpwr scs8hd_decap_12
XFILLER_72_27 vgnd vpwr scs8hd_decap_4
XPHY_115 vgnd vpwr scs8hd_decap_3
XPHY_104 vgnd vpwr scs8hd_decap_3
XFILLER_469_59 vpwr vgnd scs8hd_fill_2
XPHY_148 vgnd vpwr scs8hd_decap_3
XPHY_137 vgnd vpwr scs8hd_decap_3
XPHY_126 vgnd vpwr scs8hd_decap_3
XPHY_159 vgnd vpwr scs8hd_decap_3
XFILLER_565_80 vgnd vpwr scs8hd_fill_1
XFILLER_115_3 vgnd vpwr scs8hd_decap_12
XFILLER_484_3 vgnd vpwr scs8hd_decap_12
XFILLER_153_74 vgnd vpwr scs8hd_decap_6
XFILLER_379_15 vgnd vpwr scs8hd_decap_12
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_379_59 vpwr vgnd scs8hd_fill_2
XPHY_660 vgnd vpwr scs8hd_decap_3
XPHY_671 vgnd vpwr scs8hd_decap_3
XPHY_682 vgnd vpwr scs8hd_decap_3
XPHY_693 vgnd vpwr scs8hd_decap_3
XPHY_1292 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_545_39 vgnd vpwr scs8hd_decap_12
XFILLER_475_80 vgnd vpwr scs8hd_fill_1
XFILLER_561_27 vgnd vpwr scs8hd_decap_12
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
XFILLER_289_15 vgnd vpwr scs8hd_decap_12
XFILLER_289_59 vpwr vgnd scs8hd_fill_2
XFILLER_586_68 vgnd vpwr scs8hd_decap_12
XFILLER_519_51 vgnd vpwr scs8hd_decap_8
XFILLER_519_62 vgnd vpwr scs8hd_decap_12
XFILLER_385_80 vgnd vpwr scs8hd_fill_1
XFILLER_455_39 vgnd vpwr scs8hd_decap_12
XFILLER_471_27 vgnd vpwr scs8hd_decap_12
XFILLER_67_27 vgnd vpwr scs8hd_decap_12
XFILLER_404_32 vgnd vpwr scs8hd_decap_12
XFILLER_83_15 vgnd vpwr scs8hd_decap_12
XFILLER_83_59 vpwr vgnd scs8hd_fill_2
XFILLER_232_3 vgnd vpwr scs8hd_decap_12
XFILLER_429_51 vgnd vpwr scs8hd_decap_8
XFILLER_496_68 vgnd vpwr scs8hd_decap_12
XFILLER_429_62 vgnd vpwr scs8hd_decap_12
XFILLER_295_80 vgnd vpwr scs8hd_fill_1
XFILLER_365_39 vgnd vpwr scs8hd_decap_12
XFILLER_381_27 vgnd vpwr scs8hd_decap_12
XFILLER_314_32 vgnd vpwr scs8hd_decap_12
XFILLER_339_51 vgnd vpwr scs8hd_decap_8
XFILLER_556_27 vgnd vpwr scs8hd_decap_4
XFILLER_78_3 vgnd vpwr scs8hd_decap_12
XPHY_490 vgnd vpwr scs8hd_decap_3
XFILLER_339_62 vgnd vpwr scs8hd_decap_12
XFILLER_275_39 vgnd vpwr scs8hd_decap_12
XFILLER_208_11 vpwr vgnd scs8hd_fill_2
XFILLER_572_15 vgnd vpwr scs8hd_decap_12
XFILLER_291_27 vgnd vpwr scs8hd_decap_12
XFILLER_224_32 vgnd vpwr scs8hd_decap_12
XFILLER_521_74 vgnd vpwr scs8hd_decap_6
XFILLER_249_51 vgnd vpwr scs8hd_decap_8
XFILLER_249_62 vgnd vpwr scs8hd_decap_12
XFILLER_466_27 vgnd vpwr scs8hd_decap_4
XFILLER_118_44 vgnd vpwr scs8hd_decap_12
XFILLER_78_15 vgnd vpwr scs8hd_decap_12
XFILLER_482_15 vgnd vpwr scs8hd_decap_12
XFILLER_134_32 vgnd vpwr scs8hd_decap_12
XFILLER_182_3 vgnd vpwr scs8hd_decap_12
XFILLER_431_74 vgnd vpwr scs8hd_decap_6
XFILLER_27_74 vgnd vpwr scs8hd_decap_6
XFILLER_447_3 vgnd vpwr scs8hd_decap_12
XFILLER_300_56 vgnd vpwr scs8hd_decap_12
XFILLER_43_62 vgnd vpwr scs8hd_decap_12
XFILLER_43_51 vgnd vpwr scs8hd_decap_8
XFILLER_159_51 vgnd vpwr scs8hd_decap_8
XFILLER_159_62 vgnd vpwr scs8hd_decap_12
XFILLER_376_27 vgnd vpwr scs8hd_decap_4
XFILLER_392_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_56 vgnd vpwr scs8hd_decap_12
XFILLER_341_74 vgnd vpwr scs8hd_decap_6
XFILLER_84_80 vgnd vpwr scs8hd_fill_1
XFILLER_210_12 vgnd vpwr scs8hd_fill_1
Xlogical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ right_width_0_height_0__pin_12_ logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[6] vgnd vpwr scs8hd_ebufn_1
XFILLER_567_15 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_210_56 vgnd vpwr scs8hd_decap_12
XFILLER_567_59 vpwr vgnd scs8hd_fill_2
XFILLER_286_27 vgnd vpwr scs8hd_decap_4
XFILLER_104_68 vgnd vpwr scs8hd_decap_12
XFILLER_251_74 vgnd vpwr scs8hd_decap_6
XFILLER_120_56 vgnd vpwr scs8hd_decap_12
XFILLER_477_15 vgnd vpwr scs8hd_decap_12
XPHY_1803 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_80_27 vgnd vpwr scs8hd_decap_4
XFILLER_477_59 vpwr vgnd scs8hd_fill_2
XFILLER_573_80 vgnd vpwr scs8hd_fill_1
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XFILLER_397_3 vgnd vpwr scs8hd_decap_12
XFILLER_564_3 vgnd vpwr scs8hd_decap_12
XFILLER_161_74 vgnd vpwr scs8hd_decap_6
XFILLER_387_15 vgnd vpwr scs8hd_decap_12
XFILLER_387_59 vpwr vgnd scs8hd_fill_2
XFILLER_553_39 vgnd vpwr scs8hd_decap_12
XFILLER_79_80 vgnd vpwr scs8hd_fill_1
XFILLER_483_80 vgnd vpwr scs8hd_fill_1
XFILLER_502_32 vgnd vpwr scs8hd_decap_12
XFILLER_297_15 vgnd vpwr scs8hd_decap_12
XFILLER_297_59 vpwr vgnd scs8hd_fill_2
XFILLER_594_68 vgnd vpwr scs8hd_decap_12
XFILLER_527_62 vgnd vpwr scs8hd_decap_12
XFILLER_527_51 vgnd vpwr scs8hd_decap_8
XFILLER_59_39 vgnd vpwr scs8hd_decap_12
XFILLER_393_80 vgnd vpwr scs8hd_fill_1
XFILLER_463_39 vgnd vpwr scs8hd_decap_12
XFILLER_75_27 vgnd vpwr scs8hd_decap_12
XFILLER_412_32 vgnd vpwr scs8hd_decap_12
XFILLER_91_15 vgnd vpwr scs8hd_decap_12
XFILLER_91_59 vpwr vgnd scs8hd_fill_2
XPHY_1600 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_568_80 vgnd vpwr scs8hd_fill_1
XFILLER_145_3 vgnd vpwr scs8hd_decap_12
XPHY_1611 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1622 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1633 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1644 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1655 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1666 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_312_3 vgnd vpwr scs8hd_decap_12
XPHY_1677 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1688 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1699 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_437_51 vgnd vpwr scs8hd_decap_8
XFILLER_437_62 vgnd vpwr scs8hd_decap_12
XFILLER_373_39 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_306_44 vgnd vpwr scs8hd_decap_12
X_20_ gfpga_pad_GPIO_PAD[1] right_width_0_height_0__pin_3_ vgnd vpwr scs8hd_buf_2
XFILLER_603_75 vgnd vpwr scs8hd_decap_6
XFILLER_322_32 vgnd vpwr scs8hd_decap_12
XFILLER_478_80 vgnd vpwr scs8hd_fill_1
XFILLER_564_27 vgnd vpwr scs8hd_decap_4
XFILLER_60_3 vgnd vpwr scs8hd_decap_12
XFILLER_347_51 vgnd vpwr scs8hd_decap_8
XFILLER_347_62 vgnd vpwr scs8hd_decap_12
XFILLER_283_39 vgnd vpwr scs8hd_decap_12
XFILLER_580_15 vgnd vpwr scs8hd_decap_12
XFILLER_216_44 vgnd vpwr scs8hd_decap_12
XFILLER_232_32 vgnd vpwr scs8hd_decap_12
XPHY_308 vgnd vpwr scs8hd_decap_3
XPHY_319 vgnd vpwr scs8hd_decap_3
XFILLER_388_80 vgnd vpwr scs8hd_fill_1
XFILLER_257_51 vgnd vpwr scs8hd_decap_8
XFILLER_257_62 vgnd vpwr scs8hd_decap_12
XFILLER_474_27 vgnd vpwr scs8hd_decap_4
XFILLER_10_44 vgnd vpwr scs8hd_decap_12
XFILLER_126_44 vgnd vpwr scs8hd_decap_12
XFILLER_490_15 vgnd vpwr scs8hd_decap_12
XFILLER_86_15 vgnd vpwr scs8hd_decap_12
XFILLER_142_32 vgnd vpwr scs8hd_decap_12
XFILLER_262_3 vgnd vpwr scs8hd_decap_12
XFILLER_35_74 vgnd vpwr scs8hd_decap_6
XPHY_820 vgnd vpwr scs8hd_decap_3
XFILLER_527_3 vgnd vpwr scs8hd_decap_12
XFILLER_298_80 vgnd vpwr scs8hd_fill_1
XPHY_831 vgnd vpwr scs8hd_decap_3
XPHY_842 vgnd vpwr scs8hd_decap_3
XPHY_853 vgnd vpwr scs8hd_decap_3
XPHY_1430 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1441 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_864 vgnd vpwr scs8hd_decap_3
XPHY_875 vgnd vpwr scs8hd_decap_3
XPHY_886 vgnd vpwr scs8hd_decap_3
XPHY_897 vgnd vpwr scs8hd_decap_3
XFILLER_51_62 vgnd vpwr scs8hd_decap_12
XFILLER_51_51 vgnd vpwr scs8hd_decap_8
XPHY_1452 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1463 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1474 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1485 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_167_51 vgnd vpwr scs8hd_decap_8
XFILLER_167_62 vgnd vpwr scs8hd_decap_12
XPHY_1496 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_384_27 vgnd vpwr scs8hd_decap_4
XFILLER_202_24 vgnd vpwr scs8hd_decap_6
XFILLER_559_27 vgnd vpwr scs8hd_decap_12
XFILLER_202_68 vgnd vpwr scs8hd_decap_12
XFILLER_92_80 vgnd vpwr scs8hd_fill_1
XFILLER_575_15 vgnd vpwr scs8hd_decap_12
XFILLER_575_59 vpwr vgnd scs8hd_fill_2
XFILLER_294_27 vgnd vpwr scs8hd_decap_4
XFILLER_112_68 vgnd vpwr scs8hd_decap_12
XFILLER_469_27 vgnd vpwr scs8hd_decap_12
XPHY_116 vgnd vpwr scs8hd_decap_3
XPHY_105 vgnd vpwr scs8hd_decap_3
XPHY_149 vgnd vpwr scs8hd_decap_3
XPHY_138 vgnd vpwr scs8hd_decap_3
XPHY_127 vgnd vpwr scs8hd_decap_3
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_485_15 vgnd vpwr scs8hd_decap_12
XFILLER_485_59 vpwr vgnd scs8hd_fill_2
XFILLER_108_3 vgnd vpwr scs8hd_decap_12
XFILLER_581_80 vgnd vpwr scs8hd_fill_1
XFILLER_477_3 vgnd vpwr scs8hd_decap_12
XFILLER_600_32 vgnd vpwr scs8hd_decap_12
XFILLER_379_27 vgnd vpwr scs8hd_decap_12
XPHY_7 vgnd vpwr scs8hd_decap_3
XPHY_650 vgnd vpwr scs8hd_decap_3
XPHY_661 vgnd vpwr scs8hd_decap_3
XPHY_672 vgnd vpwr scs8hd_decap_3
XPHY_683 vgnd vpwr scs8hd_decap_3
XPHY_694 vgnd vpwr scs8hd_decap_3
XFILLER_395_15 vgnd vpwr scs8hd_decap_12
XPHY_1293 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_395_59 vpwr vgnd scs8hd_fill_2
XFILLER_561_39 vgnd vpwr scs8hd_decap_12
XFILLER_491_80 vgnd vpwr scs8hd_fill_1
XFILLER_87_80 vgnd vpwr scs8hd_fill_1
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
XFILLER_289_27 vgnd vpwr scs8hd_decap_12
XFILLER_510_32 vgnd vpwr scs8hd_decap_12
XFILLER_519_74 vgnd vpwr scs8hd_decap_6
XFILLER_535_62 vgnd vpwr scs8hd_decap_12
XFILLER_535_51 vgnd vpwr scs8hd_decap_8
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _05_/X vgnd vpwr scs8hd_diode_2
XFILLER_67_39 vgnd vpwr scs8hd_decap_12
XFILLER_471_39 vgnd vpwr scs8hd_decap_12
XFILLER_190_29 vpwr vgnd scs8hd_fill_2
XFILLER_404_44 vgnd vpwr scs8hd_decap_12
XFILLER_83_27 vgnd vpwr scs8hd_decap_12
XFILLER_420_32 vgnd vpwr scs8hd_decap_12
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
XFILLER_576_80 vgnd vpwr scs8hd_fill_1
XFILLER_225_3 vgnd vpwr scs8hd_decap_8
XFILLER_429_74 vgnd vpwr scs8hd_decap_6
XFILLER_445_51 vgnd vpwr scs8hd_decap_8
XFILLER_445_62 vgnd vpwr scs8hd_decap_12
XFILLER_594_3 vgnd vpwr scs8hd_decap_12
XFILLER_381_39 vgnd vpwr scs8hd_decap_12
XFILLER_314_44 vgnd vpwr scs8hd_decap_12
XFILLER_330_32 vgnd vpwr scs8hd_decap_12
XFILLER_189_60 vgnd vpwr scs8hd_fill_1
XPHY_480 vgnd vpwr scs8hd_decap_3
XPHY_491 vgnd vpwr scs8hd_decap_3
XFILLER_339_74 vgnd vpwr scs8hd_decap_6
XFILLER_486_80 vgnd vpwr scs8hd_fill_1
XPHY_1090 vgnd vpwr scs8hd_decap_3
XFILLER_208_23 vpwr vgnd scs8hd_fill_2
XFILLER_572_27 vgnd vpwr scs8hd_decap_4
XFILLER_355_51 vgnd vpwr scs8hd_decap_8
XFILLER_355_62 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_291_39 vgnd vpwr scs8hd_decap_12
XFILLER_224_44 vgnd vpwr scs8hd_decap_12
XFILLER_240_32 vgnd vpwr scs8hd_decap_12
XFILLER_249_74 vgnd vpwr scs8hd_decap_6
XFILLER_396_80 vgnd vpwr scs8hd_fill_1
XFILLER_118_56 vgnd vpwr scs8hd_decap_12
XFILLER_265_51 vgnd vpwr scs8hd_decap_8
XFILLER_265_62 vgnd vpwr scs8hd_decap_12
XFILLER_482_27 vgnd vpwr scs8hd_decap_4
XFILLER_78_27 vgnd vpwr scs8hd_decap_4
XFILLER_134_44 vgnd vpwr scs8hd_decap_12
XFILLER_94_15 vgnd vpwr scs8hd_decap_12
XFILLER_175_3 vgnd vpwr scs8hd_decap_12
XFILLER_150_32 vgnd vpwr scs8hd_decap_12
XFILLER_342_3 vgnd vpwr scs8hd_decap_12
XFILLER_43_74 vgnd vpwr scs8hd_decap_6
XFILLER_300_68 vgnd vpwr scs8hd_decap_12
XFILLER_159_74 vgnd vpwr scs8hd_decap_6
XFILLER_175_51 vgnd vpwr scs8hd_decap_8
XFILLER_175_62 vgnd vpwr scs8hd_decap_12
XFILLER_392_27 vgnd vpwr scs8hd_decap_4
XFILLER_4_68 vgnd vpwr scs8hd_decap_12
XFILLER_567_27 vgnd vpwr scs8hd_decap_12
XFILLER_90_3 vgnd vpwr scs8hd_decap_12
XFILLER_210_68 vgnd vpwr scs8hd_decap_12
XFILLER_583_15 vgnd vpwr scs8hd_decap_12
XFILLER_583_59 vpwr vgnd scs8hd_fill_2
XPHY_1804 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_120_68 vgnd vpwr scs8hd_decap_12
XFILLER_477_27 vgnd vpwr scs8hd_decap_12
XFILLER_89_15 vgnd vpwr scs8hd_decap_12
XFILLER_493_15 vgnd vpwr scs8hd_decap_12
XFILLER_493_59 vpwr vgnd scs8hd_fill_2
XFILLER_89_59 vpwr vgnd scs8hd_fill_2
XFILLER_292_3 vgnd vpwr scs8hd_decap_12
XFILLER_557_3 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_387_27 vgnd vpwr scs8hd_decap_12
XFILLER_95_80 vgnd vpwr scs8hd_fill_1
XFILLER_502_44 vgnd vpwr scs8hd_decap_12
XFILLER_578_15 vgnd vpwr scs8hd_decap_12
XFILLER_297_27 vgnd vpwr scs8hd_decap_12
XFILLER_527_74 vgnd vpwr scs8hd_decap_6
XFILLER_543_62 vgnd vpwr scs8hd_decap_12
XFILLER_543_51 vgnd vpwr scs8hd_decap_8
XFILLER_75_39 vgnd vpwr scs8hd_decap_12
XFILLER_412_44 vgnd vpwr scs8hd_decap_12
XFILLER_488_15 vgnd vpwr scs8hd_decap_12
XFILLER_91_27 vgnd vpwr scs8hd_decap_12
XFILLER_24_32 vgnd vpwr scs8hd_decap_12
XPHY_1601 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1612 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1623 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1634 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_138_3 vgnd vpwr scs8hd_decap_12
XPHY_1645 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1656 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1667 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1678 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1689 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_584_80 vgnd vpwr scs8hd_fill_1
XFILLER_305_3 vgnd vpwr scs8hd_decap_12
XFILLER_437_74 vgnd vpwr scs8hd_decap_6
XFILLER_306_56 vgnd vpwr scs8hd_decap_12
XFILLER_453_51 vgnd vpwr scs8hd_decap_8
XFILLER_49_62 vgnd vpwr scs8hd_decap_12
XFILLER_49_51 vgnd vpwr scs8hd_decap_8
XFILLER_453_62 vgnd vpwr scs8hd_decap_12
XFILLER_603_32 vgnd vpwr scs8hd_decap_12
XFILLER_322_44 vgnd vpwr scs8hd_decap_12
XFILLER_398_15 vgnd vpwr scs8hd_decap_12
XFILLER_347_74 vgnd vpwr scs8hd_decap_6
XFILLER_53_3 vgnd vpwr scs8hd_decap_12
XFILLER_494_80 vgnd vpwr scs8hd_fill_1
XFILLER_580_27 vgnd vpwr scs8hd_decap_4
XFILLER_216_56 vgnd vpwr scs8hd_decap_12
XFILLER_363_51 vgnd vpwr scs8hd_decap_8
XFILLER_363_62 vgnd vpwr scs8hd_decap_12
XFILLER_232_44 vgnd vpwr scs8hd_decap_12
XFILLER_101_15 vgnd vpwr scs8hd_decap_12
XPHY_309 vgnd vpwr scs8hd_decap_3
XFILLER_101_59 vpwr vgnd scs8hd_fill_2
XFILLER_257_74 vgnd vpwr scs8hd_decap_6
XFILLER_10_56 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_273_51 vgnd vpwr scs8hd_decap_8
XFILLER_126_56 vgnd vpwr scs8hd_decap_12
XFILLER_86_27 vgnd vpwr scs8hd_decap_4
XFILLER_273_62 vgnd vpwr scs8hd_decap_12
XFILLER_490_27 vgnd vpwr scs8hd_decap_4
XFILLER_142_44 vgnd vpwr scs8hd_decap_12
XFILLER_255_3 vgnd vpwr scs8hd_decap_12
XFILLER_579_80 vgnd vpwr scs8hd_fill_1
XPHY_810 vgnd vpwr scs8hd_decap_3
XPHY_821 vgnd vpwr scs8hd_decap_3
XPHY_832 vgnd vpwr scs8hd_decap_3
XPHY_843 vgnd vpwr scs8hd_decap_3
XPHY_854 vgnd vpwr scs8hd_decap_3
XPHY_1420 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1431 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1442 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_422_3 vgnd vpwr scs8hd_decap_12
XPHY_865 vgnd vpwr scs8hd_decap_3
XPHY_876 vgnd vpwr scs8hd_decap_3
XPHY_887 vgnd vpwr scs8hd_decap_3
XPHY_1453 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1464 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1475 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_898 vgnd vpwr scs8hd_decap_3
XFILLER_51_74 vgnd vpwr scs8hd_decap_6
XPHY_1486 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1497 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_167_74 vgnd vpwr scs8hd_decap_6
XFILLER_183_62 vgnd vpwr scs8hd_decap_12
XFILLER_559_39 vgnd vpwr scs8hd_decap_12
XFILLER_489_80 vgnd vpwr scs8hd_fill_1
XFILLER_575_27 vgnd vpwr scs8hd_decap_12
XFILLER_508_32 vgnd vpwr scs8hd_decap_12
XFILLER_591_15 vgnd vpwr scs8hd_decap_12
XFILLER_591_59 vpwr vgnd scs8hd_fill_2
XPHY_106 vgnd vpwr scs8hd_decap_3
XFILLER_399_80 vgnd vpwr scs8hd_fill_1
XFILLER_469_39 vgnd vpwr scs8hd_decap_12
XPHY_139 vgnd vpwr scs8hd_decap_3
XPHY_128 vgnd vpwr scs8hd_decap_3
XPHY_117 vgnd vpwr scs8hd_decap_3
XFILLER_188_29 vpwr vgnd scs8hd_fill_2
XFILLER_485_27 vgnd vpwr scs8hd_decap_12
XFILLER_418_32 vgnd vpwr scs8hd_decap_12
XFILLER_97_15 vgnd vpwr scs8hd_decap_12
XFILLER_97_59 vpwr vgnd scs8hd_fill_2
XFILLER_372_3 vgnd vpwr scs8hd_decap_12
XFILLER_600_44 vgnd vpwr scs8hd_decap_12
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_379_39 vgnd vpwr scs8hd_decap_12
XFILLER_102_80 vgnd vpwr scs8hd_fill_1
XPHY_640 vgnd vpwr scs8hd_decap_3
XPHY_651 vgnd vpwr scs8hd_decap_3
XPHY_662 vgnd vpwr scs8hd_decap_3
XPHY_1250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_673 vgnd vpwr scs8hd_decap_3
XPHY_684 vgnd vpwr scs8hd_decap_3
XPHY_695 vgnd vpwr scs8hd_decap_3
XFILLER_395_27 vgnd vpwr scs8hd_decap_12
XPHY_1283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_328_32 vgnd vpwr scs8hd_decap_12
XPHY_1294 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_3 vgnd vpwr scs8hd_decap_12
XFILLER_289_39 vgnd vpwr scs8hd_decap_12
XFILLER_510_44 vgnd vpwr scs8hd_decap_12
XFILLER_586_15 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_238_32 vgnd vpwr scs8hd_decap_12
XFILLER_535_74 vgnd vpwr scs8hd_decap_6
XFILLER_551_51 vgnd vpwr scs8hd_decap_8
XFILLER_551_62 vgnd vpwr scs8hd_decap_12
XFILLER_404_56 vgnd vpwr scs8hd_decap_12
XFILLER_83_39 vgnd vpwr scs8hd_decap_12
XFILLER_16_44 vgnd vpwr scs8hd_decap_12
XFILLER_420_44 vgnd vpwr scs8hd_decap_12
XFILLER_496_15 vgnd vpwr scs8hd_decap_12
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XFILLER_148_32 vgnd vpwr scs8hd_decap_12
XFILLER_120_3 vgnd vpwr scs8hd_decap_12
XFILLER_592_80 vgnd vpwr scs8hd_fill_1
XFILLER_445_74 vgnd vpwr scs8hd_decap_6
XFILLER_587_3 vgnd vpwr scs8hd_decap_12
XFILLER_57_62 vgnd vpwr scs8hd_decap_12
XFILLER_57_51 vgnd vpwr scs8hd_decap_8
XFILLER_314_56 vgnd vpwr scs8hd_decap_12
XFILLER_461_51 vgnd vpwr scs8hd_decap_8
XFILLER_461_62 vgnd vpwr scs8hd_decap_12
XFILLER_330_44 vgnd vpwr scs8hd_decap_12
XPHY_470 vgnd vpwr scs8hd_decap_3
XPHY_481 vgnd vpwr scs8hd_decap_3
XPHY_492 vgnd vpwr scs8hd_decap_3
XPHY_1091 vgnd vpwr scs8hd_decap_3
XPHY_1080 vgnd vpwr scs8hd_decap_3
XFILLER_98_80 vgnd vpwr scs8hd_fill_1
XFILLER_355_74 vgnd vpwr scs8hd_decap_6
XFILLER_224_56 vgnd vpwr scs8hd_decap_12
XFILLER_371_51 vgnd vpwr scs8hd_decap_8
XFILLER_371_62 vgnd vpwr scs8hd_decap_12
XFILLER_240_44 vgnd vpwr scs8hd_decap_12
XFILLER_118_68 vgnd vpwr scs8hd_decap_12
XFILLER_265_74 vgnd vpwr scs8hd_decap_6
XFILLER_94_27 vgnd vpwr scs8hd_decap_4
XFILLER_134_56 vgnd vpwr scs8hd_decap_12
XFILLER_281_51 vgnd vpwr scs8hd_decap_8
XFILLER_281_62 vgnd vpwr scs8hd_decap_12
XFILLER_150_44 vgnd vpwr scs8hd_decap_12
XFILLER_168_3 vgnd vpwr scs8hd_decap_12
XFILLER_587_80 vgnd vpwr scs8hd_fill_1
XFILLER_335_3 vgnd vpwr scs8hd_decap_12
XFILLER_502_3 vgnd vpwr scs8hd_decap_12
XFILLER_175_74 vgnd vpwr scs8hd_decap_6
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_191_51 vgnd vpwr scs8hd_decap_8
XFILLER_191_62 vgnd vpwr scs8hd_decap_12
XFILLER_567_39 vgnd vpwr scs8hd_decap_12
XFILLER_497_80 vgnd vpwr scs8hd_fill_1
XFILLER_83_3 vgnd vpwr scs8hd_decap_12
XFILLER_583_27 vgnd vpwr scs8hd_decap_12
XFILLER_516_32 vgnd vpwr scs8hd_decap_12
XFILLER_104_15 vgnd vpwr scs8hd_decap_12
XPHY_1805 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_477_39 vgnd vpwr scs8hd_decap_12
XFILLER_196_18 vgnd vpwr scs8hd_decap_12
XFILLER_200_80 vgnd vpwr scs8hd_fill_1
XFILLER_493_27 vgnd vpwr scs8hd_decap_12
XFILLER_89_27 vgnd vpwr scs8hd_decap_12
XFILLER_426_32 vgnd vpwr scs8hd_decap_12
XFILLER_285_3 vgnd vpwr scs8hd_decap_12
XFILLER_452_3 vgnd vpwr scs8hd_decap_12
XFILLER_387_39 vgnd vpwr scs8hd_decap_12
XFILLER_110_80 vgnd vpwr scs8hd_fill_1
XFILLER_336_32 vgnd vpwr scs8hd_decap_12
XFILLER_205_14 vpwr vgnd scs8hd_fill_2
XFILLER_502_56 vgnd vpwr scs8hd_decap_12
XFILLER_578_27 vgnd vpwr scs8hd_decap_4
XFILLER_297_39 vgnd vpwr scs8hd_decap_12
XFILLER_594_15 vgnd vpwr scs8hd_decap_12
XFILLER_246_32 vgnd vpwr scs8hd_decap_12
XFILLER_543_74 vgnd vpwr scs8hd_decap_6
XFILLER_412_56 vgnd vpwr scs8hd_decap_12
XFILLER_488_27 vgnd vpwr scs8hd_decap_4
XFILLER_91_39 vgnd vpwr scs8hd_decap_12
XFILLER_24_44 vgnd vpwr scs8hd_decap_12
XPHY_1602 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1613 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1624 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1635 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1646 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1657 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1668 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1679 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
XFILLER_156_32 vgnd vpwr scs8hd_decap_12
XFILLER_200_3 vpwr vgnd scs8hd_fill_2
XFILLER_306_68 vgnd vpwr scs8hd_decap_12
XFILLER_453_74 vgnd vpwr scs8hd_decap_6
XFILLER_603_44 vgnd vpwr scs8hd_decap_12
XFILLER_49_74 vgnd vpwr scs8hd_decap_6
XFILLER_1_15 vgnd vpwr scs8hd_decap_12
XFILLER_105_80 vgnd vpwr scs8hd_fill_1
XFILLER_65_51 vgnd vpwr scs8hd_decap_8
XFILLER_322_56 vgnd vpwr scs8hd_decap_12
XFILLER_65_62 vgnd vpwr scs8hd_decap_12
XFILLER_398_27 vgnd vpwr scs8hd_decap_4
XFILLER_46_3 vgnd vpwr scs8hd_decap_12
XFILLER_216_68 vgnd vpwr scs8hd_decap_12
XFILLER_363_74 vgnd vpwr scs8hd_decap_6
XFILLER_589_15 vgnd vpwr scs8hd_decap_12
XFILLER_232_56 vgnd vpwr scs8hd_decap_12
XFILLER_589_59 vpwr vgnd scs8hd_fill_2
XFILLER_101_27 vgnd vpwr scs8hd_decap_12
XFILLER_193_19 vgnd vpwr scs8hd_decap_12
XFILLER_10_68 vgnd vpwr scs8hd_decap_12
XFILLER_126_68 vgnd vpwr scs8hd_decap_12
XFILLER_273_74 vgnd vpwr scs8hd_decap_6
XFILLER_142_56 vgnd vpwr scs8hd_decap_12
XFILLER_499_15 vgnd vpwr scs8hd_decap_12
XFILLER_499_59 vpwr vgnd scs8hd_fill_2
XFILLER_150_3 vgnd vpwr scs8hd_decap_12
XPHY_800 vgnd vpwr scs8hd_decap_3
XPHY_811 vgnd vpwr scs8hd_decap_3
XFILLER_248_3 vgnd vpwr scs8hd_decap_12
XPHY_822 vgnd vpwr scs8hd_decap_3
XPHY_833 vgnd vpwr scs8hd_decap_3
XPHY_844 vgnd vpwr scs8hd_decap_3
XPHY_1410 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1421 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1432 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_855 vgnd vpwr scs8hd_decap_3
XPHY_866 vgnd vpwr scs8hd_decap_3
XPHY_877 vgnd vpwr scs8hd_decap_3
XPHY_888 vgnd vpwr scs8hd_decap_3
XFILLER_595_80 vgnd vpwr scs8hd_fill_1
XPHY_1443 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1454 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1465 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1476 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_415_3 vgnd vpwr scs8hd_decap_12
XPHY_899 vgnd vpwr scs8hd_decap_3
XPHY_1487 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1498 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_183_41 vgnd vpwr scs8hd_decap_12
XFILLER_183_74 vgnd vpwr scs8hd_decap_6
XFILLER_575_39 vgnd vpwr scs8hd_decap_12
XFILLER_508_44 vgnd vpwr scs8hd_decap_12
XFILLER_591_27 vgnd vpwr scs8hd_decap_12
XFILLER_524_32 vgnd vpwr scs8hd_decap_12
XFILLER_2_80 vgnd vpwr scs8hd_fill_1
XFILLER_112_15 vgnd vpwr scs8hd_decap_12
XPHY_107 vgnd vpwr scs8hd_decap_3
XFILLER_549_51 vgnd vpwr scs8hd_decap_8
XPHY_129 vgnd vpwr scs8hd_decap_3
XPHY_118 vgnd vpwr scs8hd_decap_3
XFILLER_549_62 vgnd vpwr scs8hd_decap_12
XFILLER_485_39 vgnd vpwr scs8hd_decap_12
XFILLER_418_44 vgnd vpwr scs8hd_decap_12
XFILLER_97_27 vgnd vpwr scs8hd_decap_12
XANTENNA__10__A _07_/C vgnd vpwr scs8hd_diode_2
XFILLER_434_32 vgnd vpwr scs8hd_decap_12
XFILLER_198_3 vgnd vpwr scs8hd_decap_12
XFILLER_365_3 vgnd vpwr scs8hd_decap_12
XFILLER_600_56 vgnd vpwr scs8hd_decap_12
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_532_3 vgnd vpwr scs8hd_decap_12
XFILLER_459_51 vgnd vpwr scs8hd_decap_8
XPHY_630 vgnd vpwr scs8hd_decap_3
XPHY_641 vgnd vpwr scs8hd_decap_3
XPHY_652 vgnd vpwr scs8hd_decap_3
XFILLER_459_62 vgnd vpwr scs8hd_decap_12
XPHY_1240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_663 vgnd vpwr scs8hd_decap_3
XPHY_674 vgnd vpwr scs8hd_decap_3
XPHY_685 vgnd vpwr scs8hd_decap_3
XPHY_696 vgnd vpwr scs8hd_decap_3
XFILLER_395_39 vgnd vpwr scs8hd_decap_12
XPHY_1284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1295 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_328_44 vgnd vpwr scs8hd_decap_12
XFILLER_344_32 vgnd vpwr scs8hd_decap_12
XFILLER_510_56 vgnd vpwr scs8hd_decap_12
XFILLER_586_27 vgnd vpwr scs8hd_decap_4
XFILLER_369_51 vgnd vpwr scs8hd_decap_8
XFILLER_369_62 vgnd vpwr scs8hd_decap_12
XFILLER_238_44 vgnd vpwr scs8hd_decap_12
XFILLER_107_15 vgnd vpwr scs8hd_decap_12
XFILLER_254_32 vgnd vpwr scs8hd_decap_12
XFILLER_107_59 vpwr vgnd scs8hd_fill_2
XFILLER_551_74 vgnd vpwr scs8hd_decap_6
XFILLER_404_68 vgnd vpwr scs8hd_decap_12
XFILLER_203_80 vgnd vpwr scs8hd_fill_1
XFILLER_420_56 vgnd vpwr scs8hd_decap_12
XFILLER_16_56 vgnd vpwr scs8hd_decap_12
XFILLER_279_51 vgnd vpwr scs8hd_decap_8
XFILLER_279_62 vgnd vpwr scs8hd_decap_12
XFILLER_496_27 vgnd vpwr scs8hd_decap_4
XANTENNA__05__A _07_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_148_44 vgnd vpwr scs8hd_decap_12
XFILLER_113_3 vgnd vpwr scs8hd_decap_12
XFILLER_164_32 vgnd vpwr scs8hd_decap_12
XFILLER_482_3 vgnd vpwr scs8hd_decap_12
XFILLER_314_68 vgnd vpwr scs8hd_decap_12
XFILLER_461_74 vgnd vpwr scs8hd_decap_6
XFILLER_57_74 vgnd vpwr scs8hd_decap_6
XFILLER_113_80 vgnd vpwr scs8hd_fill_1
XFILLER_330_56 vgnd vpwr scs8hd_decap_12
XFILLER_73_62 vgnd vpwr scs8hd_decap_12
XFILLER_73_51 vgnd vpwr scs8hd_decap_8
XFILLER_189_40 vgnd vpwr scs8hd_decap_12
XFILLER_189_62 vgnd vpwr scs8hd_decap_12
XPHY_460 vgnd vpwr scs8hd_decap_3
XPHY_471 vgnd vpwr scs8hd_decap_3
XPHY_482 vgnd vpwr scs8hd_decap_3
XPHY_493 vgnd vpwr scs8hd_decap_3
XPHY_1092 vgnd vpwr scs8hd_decap_3
XPHY_1081 vgnd vpwr scs8hd_decap_3
XPHY_1070 vgnd vpwr scs8hd_decap_3
XFILLER_224_68 vgnd vpwr scs8hd_decap_12
XFILLER_371_74 vgnd vpwr scs8hd_decap_6
XFILLER_597_15 vgnd vpwr scs8hd_decap_12
XFILLER_240_56 vgnd vpwr scs8hd_decap_12
XFILLER_597_59 vpwr vgnd scs8hd_fill_2
XFILLER_134_68 vgnd vpwr scs8hd_decap_12
XFILLER_281_74 vgnd vpwr scs8hd_decap_6
XFILLER_150_56 vgnd vpwr scs8hd_decap_12
XFILLER_300_15 vgnd vpwr scs8hd_decap_12
XFILLER_230_3 vgnd vpwr scs8hd_decap_12
XFILLER_328_3 vgnd vpwr scs8hd_decap_12
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XFILLER_108_80 vgnd vpwr scs8hd_fill_1
XFILLER_191_74 vgnd vpwr scs8hd_decap_6
XFILLER_210_26 vgnd vpwr scs8hd_decap_4
XFILLER_76_3 vgnd vpwr scs8hd_decap_12
XPHY_290 vgnd vpwr scs8hd_decap_3
XFILLER_219_13 vpwr vgnd scs8hd_fill_2
XFILLER_583_39 vgnd vpwr scs8hd_decap_12
XFILLER_516_44 vgnd vpwr scs8hd_decap_12
XFILLER_532_32 vgnd vpwr scs8hd_decap_12
XFILLER_104_27 vgnd vpwr scs8hd_decap_4
XFILLER_120_15 vgnd vpwr scs8hd_decap_12
XPHY_1806 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_557_62 vgnd vpwr scs8hd_decap_12
XFILLER_557_51 vgnd vpwr scs8hd_decap_8
XFILLER_89_39 vgnd vpwr scs8hd_decap_12
XFILLER_493_39 vgnd vpwr scs8hd_decap_12
XFILLER_426_44 vgnd vpwr scs8hd_decap_12
XFILLER_442_32 vgnd vpwr scs8hd_decap_12
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_180_3 vgnd vpwr scs8hd_decap_12
XFILLER_278_3 vgnd vpwr scs8hd_decap_12
XFILLER_598_80 vgnd vpwr scs8hd_fill_1
XFILLER_445_3 vgnd vpwr scs8hd_decap_12
XFILLER_467_51 vgnd vpwr scs8hd_decap_8
XFILLER_467_62 vgnd vpwr scs8hd_decap_12
XFILLER_336_44 vgnd vpwr scs8hd_decap_12
XFILLER_205_26 vpwr vgnd scs8hd_fill_2
XFILLER_352_32 vgnd vpwr scs8hd_decap_12
XFILLER_502_68 vgnd vpwr scs8hd_decap_12
XFILLER_301_80 vgnd vpwr scs8hd_fill_1
XFILLER_594_27 vgnd vpwr scs8hd_decap_4
XFILLER_377_51 vgnd vpwr scs8hd_decap_8
XFILLER_377_62 vgnd vpwr scs8hd_decap_12
XFILLER_246_44 vgnd vpwr scs8hd_decap_12
XFILLER_5_80 vgnd vpwr scs8hd_fill_1
XFILLER_115_15 vgnd vpwr scs8hd_decap_12
XFILLER_262_32 vgnd vpwr scs8hd_decap_12
XFILLER_115_59 vpwr vgnd scs8hd_fill_2
XFILLER_412_68 vgnd vpwr scs8hd_decap_12
XFILLER_211_80 vgnd vpwr scs8hd_fill_1
XFILLER_24_56 vgnd vpwr scs8hd_decap_12
XPHY_1603 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1614 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1625 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_287_51 vgnd vpwr scs8hd_decap_8
XFILLER_287_62 vgnd vpwr scs8hd_decap_12
XPHY_1636 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1647 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1658 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__13__A address[1] vgnd vpwr scs8hd_diode_2
XPHY_1669 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XFILLER_156_44 vgnd vpwr scs8hd_decap_12
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XFILLER_172_32 vgnd vpwr scs8hd_decap_12
XFILLER_395_3 vgnd vpwr scs8hd_decap_12
XFILLER_603_56 vgnd vpwr scs8hd_decap_6
XFILLER_562_3 vgnd vpwr scs8hd_decap_12
XFILLER_1_27 vgnd vpwr scs8hd_decap_12
XFILLER_1_49 vpwr vgnd scs8hd_fill_2
XFILLER_322_68 vgnd vpwr scs8hd_decap_12
XFILLER_65_74 vgnd vpwr scs8hd_decap_6
XFILLER_121_80 vgnd vpwr scs8hd_fill_1
XFILLER_81_62 vgnd vpwr scs8hd_decap_12
XFILLER_81_51 vgnd vpwr scs8hd_decap_8
XFILLER_197_51 vgnd vpwr scs8hd_decap_8
XFILLER_197_62 vgnd vpwr scs8hd_decap_12
XFILLER_39_3 vgnd vpwr scs8hd_decap_12
XFILLER_589_27 vgnd vpwr scs8hd_decap_12
XFILLER_232_68 vgnd vpwr scs8hd_fill_1
XFILLER_101_39 vgnd vpwr scs8hd_decap_12
XFILLER_206_80 vgnd vpwr scs8hd_fill_1
XFILLER_499_27 vgnd vpwr scs8hd_decap_12
XFILLER_142_68 vgnd vpwr scs8hd_decap_12
XANTENNA__08__A address[2] vgnd vpwr scs8hd_diode_2
XPHY_801 vgnd vpwr scs8hd_decap_3
XPHY_812 vgnd vpwr scs8hd_decap_3
XPHY_823 vgnd vpwr scs8hd_decap_3
XPHY_834 vgnd vpwr scs8hd_decap_3
XPHY_845 vgnd vpwr scs8hd_decap_3
XFILLER_143_3 vgnd vpwr scs8hd_decap_12
XPHY_1400 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1411 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1422 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1433 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_856 vgnd vpwr scs8hd_decap_3
XPHY_867 vgnd vpwr scs8hd_decap_3
XPHY_878 vgnd vpwr scs8hd_decap_3
XPHY_1444 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1455 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1466 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_889 vgnd vpwr scs8hd_decap_3
XPHY_1477 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1488 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1499 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_310_3 vgnd vpwr scs8hd_decap_12
XFILLER_408_3 vgnd vpwr scs8hd_decap_12
XFILLER_183_53 vgnd vpwr scs8hd_decap_8
XFILLER_116_80 vgnd vpwr scs8hd_fill_1
XFILLER_508_56 vgnd vpwr scs8hd_decap_12
XFILLER_591_39 vgnd vpwr scs8hd_decap_12
XFILLER_524_44 vgnd vpwr scs8hd_decap_12
XFILLER_540_32 vgnd vpwr scs8hd_decap_12
XFILLER_112_27 vgnd vpwr scs8hd_decap_4
XPHY_119 vgnd vpwr scs8hd_decap_3
XPHY_108 vgnd vpwr scs8hd_decap_3
XFILLER_549_74 vgnd vpwr scs8hd_decap_6
XFILLER_565_62 vgnd vpwr scs8hd_decap_12
XFILLER_565_51 vgnd vpwr scs8hd_decap_8
XFILLER_418_56 vgnd vpwr scs8hd_decap_12
XFILLER_97_39 vgnd vpwr scs8hd_decap_12
XANTENNA__10__B enable vgnd vpwr scs8hd_diode_2
XFILLER_434_44 vgnd vpwr scs8hd_decap_12
XFILLER_303_15 vgnd vpwr scs8hd_decap_12
XFILLER_450_32 vgnd vpwr scs8hd_decap_12
XFILLER_46_32 vgnd vpwr scs8hd_decap_12
XFILLER_303_59 vpwr vgnd scs8hd_fill_2
XFILLER_260_3 vgnd vpwr scs8hd_decap_12
XFILLER_358_3 vgnd vpwr scs8hd_decap_12
XFILLER_600_68 vgnd vpwr scs8hd_decap_12
XPHY_620 vgnd vpwr scs8hd_decap_3
XFILLER_525_3 vgnd vpwr scs8hd_decap_12
XPHY_631 vgnd vpwr scs8hd_decap_3
XPHY_642 vgnd vpwr scs8hd_decap_3
XPHY_653 vgnd vpwr scs8hd_decap_3
XFILLER_459_74 vgnd vpwr scs8hd_decap_6
XPHY_1230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_664 vgnd vpwr scs8hd_decap_3
XPHY_675 vgnd vpwr scs8hd_decap_3
XPHY_686 vgnd vpwr scs8hd_decap_3
XPHY_1274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XPHY_697 vgnd vpwr scs8hd_decap_3
XPHY_1296 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_59 vpwr vgnd scs8hd_fill_2
XFILLER_328_56 vgnd vpwr scs8hd_decap_12
XFILLER_475_51 vgnd vpwr scs8hd_decap_8
XFILLER_475_62 vgnd vpwr scs8hd_decap_12
XFILLER_344_44 vgnd vpwr scs8hd_decap_12
XFILLER_213_15 vgnd vpwr scs8hd_decap_12
XFILLER_213_59 vpwr vgnd scs8hd_fill_2
XFILLER_360_32 vgnd vpwr scs8hd_decap_12
XFILLER_510_68 vgnd vpwr scs8hd_decap_12
XFILLER_369_74 vgnd vpwr scs8hd_decap_6
XFILLER_238_56 vgnd vpwr scs8hd_decap_12
XFILLER_385_51 vgnd vpwr scs8hd_decap_8
XFILLER_385_62 vgnd vpwr scs8hd_decap_12
XFILLER_107_27 vgnd vpwr scs8hd_decap_12
XFILLER_254_44 vgnd vpwr scs8hd_decap_12
XFILLER_123_15 vgnd vpwr scs8hd_decap_12
XFILLER_123_59 vpwr vgnd scs8hd_fill_2
XFILLER_270_32 vgnd vpwr scs8hd_decap_12
XFILLER_199_19 vgnd vpwr scs8hd_decap_12
XFILLER_16_68 vgnd vpwr scs8hd_decap_12
XFILLER_420_68 vgnd vpwr scs8hd_decap_12
XFILLER_279_74 vgnd vpwr scs8hd_decap_6
XANTENNA__05__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
XFILLER_148_56 vgnd vpwr scs8hd_decap_12
XFILLER_295_62 vgnd vpwr scs8hd_decap_12
XFILLER_106_3 vgnd vpwr scs8hd_decap_12
XANTENNA__21__A gfpga_pad_GPIO_PAD[2] vgnd vpwr scs8hd_diode_2
XFILLER_164_44 vgnd vpwr scs8hd_decap_12
XFILLER_475_3 vgnd vpwr scs8hd_decap_12
XFILLER_180_32 vgnd vpwr scs8hd_decap_12
XFILLER_73_74 vgnd vpwr scs8hd_decap_6
XFILLER_330_68 vgnd vpwr scs8hd_decap_12
XFILLER_189_52 vgnd vpwr scs8hd_decap_8
XFILLER_189_74 vgnd vpwr scs8hd_decap_6
XPHY_450 vgnd vpwr scs8hd_decap_3
XPHY_461 vgnd vpwr scs8hd_decap_3
XPHY_472 vgnd vpwr scs8hd_decap_3
XPHY_483 vgnd vpwr scs8hd_decap_3
XPHY_494 vgnd vpwr scs8hd_decap_3
XPHY_1082 vgnd vpwr scs8hd_decap_3
XPHY_1071 vgnd vpwr scs8hd_decap_3
XPHY_1060 vgnd vpwr scs8hd_decap_3
XPHY_1093 vgnd vpwr scs8hd_decap_3
XFILLER_208_15 vpwr vgnd scs8hd_fill_2
XFILLER_208_37 vgnd vpwr scs8hd_decap_12
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
XFILLER_304_80 vgnd vpwr scs8hd_fill_1
XFILLER_597_27 vgnd vpwr scs8hd_decap_12
XFILLER_240_68 vgnd vpwr scs8hd_decap_12
XFILLER_118_15 vgnd vpwr scs8hd_decap_12
XFILLER_8_80 vgnd vpwr scs8hd_fill_1
XFILLER_214_80 vgnd vpwr scs8hd_fill_1
XFILLER_150_68 vgnd vpwr scs8hd_decap_12
XANTENNA__16__A gfpga_pad_GPIO_PAD[5] vgnd vpwr scs8hd_diode_2
XFILLER_300_27 vgnd vpwr scs8hd_decap_4
XFILLER_223_3 vgnd vpwr scs8hd_decap_12
XFILLER_592_3 vgnd vpwr scs8hd_decap_12
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XFILLER_124_80 vgnd vpwr scs8hd_fill_1
XPHY_280 vgnd vpwr scs8hd_decap_3
XPHY_291 vgnd vpwr scs8hd_decap_3
XFILLER_69_3 vgnd vpwr scs8hd_decap_12
XFILLER_516_56 vgnd vpwr scs8hd_decap_12
XFILLER_532_44 vgnd vpwr scs8hd_decap_12
XFILLER_401_15 vgnd vpwr scs8hd_decap_12
XFILLER_401_59 vpwr vgnd scs8hd_fill_2
XFILLER_120_27 vgnd vpwr scs8hd_decap_4
XPHY_1807 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_557_74 vgnd vpwr scs8hd_decap_6
XFILLER_573_51 vgnd vpwr scs8hd_decap_8
XFILLER_209_80 vgnd vpwr scs8hd_fill_1
XFILLER_426_56 vgnd vpwr scs8hd_decap_12
XFILLER_573_62 vgnd vpwr scs8hd_decap_12
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XFILLER_442_44 vgnd vpwr scs8hd_decap_12
XFILLER_173_3 vgnd vpwr scs8hd_decap_12
XFILLER_311_15 vgnd vpwr scs8hd_decap_12
XFILLER_54_32 vgnd vpwr scs8hd_decap_12
XFILLER_311_59 vpwr vgnd scs8hd_fill_2
XFILLER_340_3 vgnd vpwr scs8hd_decap_12
XFILLER_438_3 vgnd vpwr scs8hd_decap_12
XFILLER_467_74 vgnd vpwr scs8hd_decap_6
XFILLER_119_80 vgnd vpwr scs8hd_fill_1
XFILLER_483_51 vgnd vpwr scs8hd_decap_8
XFILLER_79_62 vgnd vpwr scs8hd_decap_12
XFILLER_79_51 vgnd vpwr scs8hd_decap_8
XFILLER_336_56 vgnd vpwr scs8hd_decap_12
XFILLER_483_62 vgnd vpwr scs8hd_decap_12
XFILLER_352_44 vgnd vpwr scs8hd_decap_12
XFILLER_221_15 vgnd vpwr scs8hd_decap_12
XFILLER_221_59 vpwr vgnd scs8hd_fill_2
XFILLER_377_74 vgnd vpwr scs8hd_decap_6
XFILLER_393_51 vgnd vpwr scs8hd_decap_8
XFILLER_246_56 vgnd vpwr scs8hd_decap_12
XFILLER_393_62 vgnd vpwr scs8hd_decap_12
XFILLER_115_27 vgnd vpwr scs8hd_decap_12
XFILLER_262_44 vgnd vpwr scs8hd_decap_12
XFILLER_131_15 vgnd vpwr scs8hd_decap_12
XFILLER_131_59 vpwr vgnd scs8hd_fill_2
XPHY_1604 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1615 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_68 vgnd vpwr scs8hd_decap_12
XPHY_1626 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1637 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1648 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__13__B _14_/B vgnd vpwr scs8hd_diode_2
XFILLER_287_74 vgnd vpwr scs8hd_decap_6
XPHY_1659 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XFILLER_156_56 vgnd vpwr scs8hd_decap_12
XFILLER_306_15 vgnd vpwr scs8hd_decap_12
XFILLER_172_44 vgnd vpwr scs8hd_decap_12
XFILLER_290_3 vgnd vpwr scs8hd_decap_12
XFILLER_388_3 vgnd vpwr scs8hd_decap_12
XFILLER_1_39 vgnd vpwr scs8hd_decap_6
XFILLER_555_3 vgnd vpwr scs8hd_decap_12
XFILLER_402_80 vgnd vpwr scs8hd_fill_1
XFILLER_81_74 vgnd vpwr scs8hd_decap_6
XFILLER_197_74 vgnd vpwr scs8hd_decap_6
XFILLER_216_15 vgnd vpwr scs8hd_decap_12
XFILLER_589_39 vgnd vpwr scs8hd_decap_12
XFILLER_312_80 vgnd vpwr scs8hd_fill_1
XFILLER_538_32 vgnd vpwr scs8hd_decap_12
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_126_15 vgnd vpwr scs8hd_decap_12
XFILLER_499_39 vgnd vpwr scs8hd_decap_12
XFILLER_222_80 vgnd vpwr scs8hd_fill_1
XPHY_802 vgnd vpwr scs8hd_decap_3
XPHY_813 vgnd vpwr scs8hd_decap_3
XPHY_824 vgnd vpwr scs8hd_decap_3
XPHY_835 vgnd vpwr scs8hd_decap_3
XPHY_1401 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1412 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1423 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_846 vgnd vpwr scs8hd_decap_3
XPHY_857 vgnd vpwr scs8hd_decap_3
XPHY_868 vgnd vpwr scs8hd_decap_3
XPHY_879 vgnd vpwr scs8hd_decap_3
XFILLER_448_32 vgnd vpwr scs8hd_decap_12
XFILLER_136_3 vgnd vpwr scs8hd_decap_12
XPHY_1434 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1445 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1456 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1467 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1478 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1489 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_303_3 vgnd vpwr scs8hd_decap_12
XFILLER_132_80 vgnd vpwr scs8hd_fill_1
XFILLER_358_32 vgnd vpwr scs8hd_decap_12
XFILLER_508_68 vgnd vpwr scs8hd_decap_12
XFILLER_51_3 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ right_width_0_height_0__pin_14_ logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[7] vgnd vpwr scs8hd_ebufn_1
XFILLER_307_80 vgnd vpwr scs8hd_fill_1
XFILLER_524_56 vgnd vpwr scs8hd_decap_12
XFILLER_540_44 vgnd vpwr scs8hd_decap_12
XPHY_109 vgnd vpwr scs8hd_decap_3
XFILLER_268_32 vgnd vpwr scs8hd_decap_12
XFILLER_565_74 vgnd vpwr scs8hd_decap_6
XFILLER_418_68 vgnd vpwr scs8hd_decap_12
XANTENNA__10__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_581_62 vgnd vpwr scs8hd_decap_12
XFILLER_581_51 vgnd vpwr scs8hd_decap_8
XFILLER_217_80 vgnd vpwr scs8hd_fill_1
XFILLER_434_56 vgnd vpwr scs8hd_decap_12
XFILLER_303_27 vgnd vpwr scs8hd_decap_12
XANTENNA__19__A gfpga_pad_GPIO_PAD[0] vgnd vpwr scs8hd_diode_2
XFILLER_450_44 vgnd vpwr scs8hd_decap_12
XFILLER_46_44 vgnd vpwr scs8hd_decap_12
XFILLER_253_3 vgnd vpwr scs8hd_decap_12
XPHY_610 vgnd vpwr scs8hd_decap_3
XFILLER_62_32 vgnd vpwr scs8hd_decap_12
XPHY_621 vgnd vpwr scs8hd_decap_3
XPHY_632 vgnd vpwr scs8hd_decap_3
XPHY_643 vgnd vpwr scs8hd_decap_3
XPHY_1220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_178_32 vgnd vpwr scs8hd_decap_12
XPHY_654 vgnd vpwr scs8hd_decap_3
XPHY_665 vgnd vpwr scs8hd_decap_3
XPHY_676 vgnd vpwr scs8hd_decap_3
XPHY_687 vgnd vpwr scs8hd_decap_3
XFILLER_420_3 vgnd vpwr scs8hd_decap_12
XFILLER_518_3 vgnd vpwr scs8hd_decap_12
XPHY_1275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_27 vgnd vpwr scs8hd_decap_12
XPHY_698 vgnd vpwr scs8hd_decap_3
XPHY_1297 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1286 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_194_20 vgnd vpwr scs8hd_decap_8
XFILLER_328_68 vgnd vpwr scs8hd_decap_12
XFILLER_475_74 vgnd vpwr scs8hd_decap_6
XFILLER_11_80 vgnd vpwr scs8hd_fill_1
XFILLER_127_80 vgnd vpwr scs8hd_fill_1
XFILLER_87_51 vgnd vpwr scs8hd_decap_8
XFILLER_344_56 vgnd vpwr scs8hd_decap_12
XFILLER_491_51 vgnd vpwr scs8hd_decap_8
XFILLER_491_62 vgnd vpwr scs8hd_decap_12
XFILLER_87_62 vgnd vpwr scs8hd_decap_12
XFILLER_213_27 vgnd vpwr scs8hd_decap_12
XFILLER_360_44 vgnd vpwr scs8hd_decap_12
XFILLER_99_3 vgnd vpwr scs8hd_decap_12
XFILLER_238_68 vgnd vpwr scs8hd_decap_12
XFILLER_385_74 vgnd vpwr scs8hd_decap_6
XFILLER_107_39 vgnd vpwr scs8hd_decap_12
XFILLER_254_56 vgnd vpwr scs8hd_decap_12
XFILLER_404_15 vgnd vpwr scs8hd_decap_12
XFILLER_123_27 vgnd vpwr scs8hd_decap_12
XFILLER_270_44 vgnd vpwr scs8hd_decap_12
XFILLER_500_80 vgnd vpwr scs8hd_fill_1
XANTENNA__05__C address[1] vgnd vpwr scs8hd_diode_2
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XFILLER_148_68 vgnd vpwr scs8hd_decap_12
XFILLER_295_74 vgnd vpwr scs8hd_decap_6
XFILLER_164_56 vgnd vpwr scs8hd_decap_12
XFILLER_314_15 vgnd vpwr scs8hd_decap_12
XFILLER_180_44 vgnd vpwr scs8hd_decap_12
XFILLER_370_3 vgnd vpwr scs8hd_decap_12
XFILLER_180_66 vgnd vpwr scs8hd_decap_12
XFILLER_468_3 vgnd vpwr scs8hd_decap_12
XFILLER_410_80 vgnd vpwr scs8hd_fill_1
XPHY_440 vgnd vpwr scs8hd_decap_3
XPHY_451 vgnd vpwr scs8hd_decap_3
XPHY_462 vgnd vpwr scs8hd_decap_3
XPHY_1050 vgnd vpwr scs8hd_decap_3
XPHY_473 vgnd vpwr scs8hd_decap_3
XPHY_484 vgnd vpwr scs8hd_decap_3
XPHY_495 vgnd vpwr scs8hd_decap_3
XPHY_1083 vgnd vpwr scs8hd_decap_3
XPHY_1072 vgnd vpwr scs8hd_decap_3
XPHY_1061 vgnd vpwr scs8hd_decap_3
XPHY_1094 vgnd vpwr scs8hd_decap_3
XFILLER_208_27 vgnd vpwr scs8hd_decap_4
XFILLER_208_49 vgnd vpwr scs8hd_decap_12
XFILLER_224_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
XFILLER_597_39 vgnd vpwr scs8hd_decap_12
XFILLER_320_80 vgnd vpwr scs8hd_fill_1
XFILLER_546_32 vgnd vpwr scs8hd_decap_12
XFILLER_118_27 vgnd vpwr scs8hd_decap_4
XFILLER_134_15 vgnd vpwr scs8hd_decap_12
XFILLER_309_15 vgnd vpwr scs8hd_decap_12
XFILLER_216_3 vgnd vpwr scs8hd_decap_12
XFILLER_309_59 vpwr vgnd scs8hd_fill_2
XFILLER_456_32 vgnd vpwr scs8hd_decap_12
XFILLER_585_3 vgnd vpwr scs8hd_decap_12
XFILLER_405_80 vgnd vpwr scs8hd_fill_1
XFILLER_140_80 vgnd vpwr scs8hd_fill_1
XPHY_270 vgnd vpwr scs8hd_decap_3
XPHY_281 vgnd vpwr scs8hd_decap_3
XPHY_292 vgnd vpwr scs8hd_decap_3
XFILLER_366_32 vgnd vpwr scs8hd_decap_12
XFILLER_516_68 vgnd vpwr scs8hd_decap_12
XFILLER_532_56 vgnd vpwr scs8hd_decap_12
XFILLER_315_80 vgnd vpwr scs8hd_fill_1
XFILLER_401_27 vgnd vpwr scs8hd_decap_12
XPHY_1808 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
XFILLER_129_15 vgnd vpwr scs8hd_decap_12
XFILLER_13_59 vpwr vgnd scs8hd_fill_2
XFILLER_276_32 vgnd vpwr scs8hd_decap_12
XFILLER_129_59 vpwr vgnd scs8hd_fill_2
XFILLER_573_74 vgnd vpwr scs8hd_decap_6
XFILLER_426_68 vgnd vpwr scs8hd_decap_12
XFILLER_225_80 vgnd vpwr scs8hd_fill_1
XFILLER_442_56 vgnd vpwr scs8hd_decap_12
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
XFILLER_311_27 vgnd vpwr scs8hd_decap_12
XFILLER_54_44 vgnd vpwr scs8hd_decap_12
XFILLER_166_3 vgnd vpwr scs8hd_decap_12
XFILLER_333_3 vgnd vpwr scs8hd_decap_12
XFILLER_70_32 vgnd vpwr scs8hd_decap_12
XFILLER_186_32 vgnd vpwr scs8hd_decap_12
XFILLER_500_3 vgnd vpwr scs8hd_decap_12
XFILLER_336_68 vgnd vpwr scs8hd_decap_12
XFILLER_483_74 vgnd vpwr scs8hd_decap_6
XFILLER_79_74 vgnd vpwr scs8hd_decap_6
XFILLER_135_80 vgnd vpwr scs8hd_fill_1
XFILLER_352_56 vgnd vpwr scs8hd_decap_12
XFILLER_95_62 vgnd vpwr scs8hd_decap_12
XFILLER_95_51 vgnd vpwr scs8hd_decap_8
XFILLER_502_15 vgnd vpwr scs8hd_decap_12
XFILLER_221_27 vgnd vpwr scs8hd_decap_12
XFILLER_81_3 vgnd vpwr scs8hd_decap_12
XFILLER_246_68 vgnd vpwr scs8hd_decap_12
XFILLER_393_74 vgnd vpwr scs8hd_decap_6
XFILLER_115_39 vgnd vpwr scs8hd_decap_12
XFILLER_262_56 vgnd vpwr scs8hd_decap_12
XFILLER_412_15 vgnd vpwr scs8hd_decap_12
XFILLER_131_27 vgnd vpwr scs8hd_decap_12
XPHY_1605 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1616 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1627 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1638 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1649 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__13__C _07_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XFILLER_156_68 vgnd vpwr scs8hd_decap_12
XFILLER_306_27 vgnd vpwr scs8hd_decap_4
XFILLER_172_56 vgnd vpwr scs8hd_decap_12
XFILLER_283_3 vgnd vpwr scs8hd_decap_12
XFILLER_322_15 vgnd vpwr scs8hd_decap_12
XFILLER_450_3 vgnd vpwr scs8hd_decap_12
XFILLER_548_3 vgnd vpwr scs8hd_decap_12
XFILLER_14_80 vgnd vpwr scs8hd_fill_1
XFILLER_216_27 vgnd vpwr scs8hd_decap_4
XFILLER_232_15 vgnd vpwr scs8hd_decap_12
XFILLER_538_44 vgnd vpwr scs8hd_decap_12
XFILLER_407_15 vgnd vpwr scs8hd_decap_12
XFILLER_554_32 vgnd vpwr scs8hd_decap_12
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XFILLER_126_27 vgnd vpwr scs8hd_decap_4
XFILLER_407_59 vpwr vgnd scs8hd_fill_2
XFILLER_142_15 vgnd vpwr scs8hd_decap_12
XFILLER_503_80 vgnd vpwr scs8hd_fill_1
XFILLER_579_51 vgnd vpwr scs8hd_decap_8
XFILLER_579_62 vgnd vpwr scs8hd_decap_12
XPHY_803 vgnd vpwr scs8hd_decap_3
XPHY_814 vgnd vpwr scs8hd_decap_3
XPHY_825 vgnd vpwr scs8hd_decap_3
XPHY_836 vgnd vpwr scs8hd_decap_3
XPHY_1402 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1413 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1424 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_847 vgnd vpwr scs8hd_decap_3
XPHY_858 vgnd vpwr scs8hd_decap_3
XPHY_869 vgnd vpwr scs8hd_decap_3
XPHY_1435 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1446 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1457 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_448_44 vgnd vpwr scs8hd_decap_12
XFILLER_129_3 vgnd vpwr scs8hd_decap_12
XPHY_1468 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1479 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_317_15 vgnd vpwr scs8hd_decap_12
XFILLER_464_32 vgnd vpwr scs8hd_decap_12
XFILLER_317_59 vpwr vgnd scs8hd_fill_2
XFILLER_498_3 vgnd vpwr scs8hd_decap_12
XFILLER_413_80 vgnd vpwr scs8hd_fill_1
XFILLER_489_51 vgnd vpwr scs8hd_decap_8
XFILLER_489_62 vgnd vpwr scs8hd_decap_12
XPHY_90 vgnd vpwr scs8hd_decap_3
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _13_/Y vgnd vpwr scs8hd_diode_2
XFILLER_358_44 vgnd vpwr scs8hd_decap_12
XFILLER_227_15 vgnd vpwr scs8hd_decap_12
XFILLER_374_32 vgnd vpwr scs8hd_decap_12
XFILLER_227_59 vpwr vgnd scs8hd_fill_2
XFILLER_44_3 vgnd vpwr scs8hd_decap_12
XFILLER_524_68 vgnd vpwr scs8hd_decap_12
XFILLER_540_56 vgnd vpwr scs8hd_decap_12
XFILLER_323_80 vgnd vpwr scs8hd_fill_1
XFILLER_399_51 vgnd vpwr scs8hd_decap_8
XFILLER_399_62 vgnd vpwr scs8hd_decap_12
XFILLER_268_44 vgnd vpwr scs8hd_decap_12
XFILLER_21_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_59 vpwr vgnd scs8hd_fill_2
XFILLER_137_15 vgnd vpwr scs8hd_decap_12
XFILLER_284_32 vgnd vpwr scs8hd_decap_12
XFILLER_137_59 vpwr vgnd scs8hd_fill_2
XANTENNA__10__D _08_/Y vgnd vpwr scs8hd_diode_2
XFILLER_581_74 vgnd vpwr scs8hd_decap_6
XFILLER_434_68 vgnd vpwr scs8hd_decap_12
XFILLER_233_80 vgnd vpwr scs8hd_fill_1
XFILLER_303_39 vgnd vpwr scs8hd_decap_12
XFILLER_450_56 vgnd vpwr scs8hd_decap_12
XFILLER_600_15 vgnd vpwr scs8hd_decap_12
XFILLER_46_56 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _07_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_600 vgnd vpwr scs8hd_decap_3
XPHY_611 vgnd vpwr scs8hd_decap_3
XFILLER_62_44 vgnd vpwr scs8hd_decap_12
XFILLER_246_3 vgnd vpwr scs8hd_decap_12
XPHY_622 vgnd vpwr scs8hd_decap_3
XPHY_633 vgnd vpwr scs8hd_decap_3
XPHY_644 vgnd vpwr scs8hd_decap_3
XPHY_1210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_178_44 vgnd vpwr scs8hd_decap_12
XPHY_655 vgnd vpwr scs8hd_decap_3
XPHY_666 vgnd vpwr scs8hd_decap_3
XPHY_677 vgnd vpwr scs8hd_decap_3
XPHY_1265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_688 vgnd vpwr scs8hd_decap_3
XPHY_699 vgnd vpwr scs8hd_decap_3
XFILLER_413_3 vgnd vpwr scs8hd_decap_12
XPHY_1298 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1287 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_39 vgnd vpwr scs8hd_decap_12
XFILLER_194_32 vgnd vpwr scs8hd_decap_12
XFILLER_408_80 vgnd vpwr scs8hd_fill_1
XFILLER_344_68 vgnd vpwr scs8hd_decap_12
XFILLER_491_74 vgnd vpwr scs8hd_decap_6
XFILLER_87_74 vgnd vpwr scs8hd_decap_6
XFILLER_143_80 vgnd vpwr scs8hd_fill_1
XFILLER_213_39 vgnd vpwr scs8hd_decap_12
XFILLER_360_56 vgnd vpwr scs8hd_decap_12
XFILLER_510_15 vgnd vpwr scs8hd_decap_12
XFILLER_318_80 vgnd vpwr scs8hd_fill_1
XFILLER_254_68 vgnd vpwr scs8hd_decap_12
XFILLER_404_27 vgnd vpwr scs8hd_decap_4
XFILLER_123_39 vgnd vpwr scs8hd_decap_12
XFILLER_270_56 vgnd vpwr scs8hd_decap_12
XFILLER_420_15 vgnd vpwr scs8hd_decap_12
XFILLER_16_15 vgnd vpwr scs8hd_decap_12
XANTENNA__05__D enable vgnd vpwr scs8hd_diode_2
XFILLER_218_7 vgnd vpwr scs8hd_decap_12
XFILLER_228_80 vgnd vpwr scs8hd_fill_1
XFILLER_164_68 vgnd vpwr scs8hd_decap_12
XFILLER_314_27 vgnd vpwr scs8hd_decap_4
XFILLER_196_3 vgnd vpwr scs8hd_decap_8
XFILLER_180_56 vgnd vpwr scs8hd_decap_8
XFILLER_180_78 vgnd vpwr scs8hd_decap_3
XFILLER_330_15 vgnd vpwr scs8hd_decap_12
XFILLER_363_3 vgnd vpwr scs8hd_decap_12
XFILLER_530_3 vgnd vpwr scs8hd_decap_12
XPHY_430 vgnd vpwr scs8hd_decap_3
XPHY_441 vgnd vpwr scs8hd_decap_3
XPHY_452 vgnd vpwr scs8hd_decap_3
XPHY_463 vgnd vpwr scs8hd_decap_3
XPHY_474 vgnd vpwr scs8hd_decap_3
XPHY_485 vgnd vpwr scs8hd_decap_3
XPHY_1040 vgnd vpwr scs8hd_decap_3
XPHY_1073 vgnd vpwr scs8hd_decap_3
XPHY_1062 vgnd vpwr scs8hd_decap_3
XPHY_1051 vgnd vpwr scs8hd_decap_3
XPHY_496 vgnd vpwr scs8hd_decap_3
XPHY_1095 vgnd vpwr scs8hd_decap_3
XPHY_1084 vgnd vpwr scs8hd_decap_3
XFILLER_22_80 vgnd vpwr scs8hd_fill_1
XFILLER_138_80 vgnd vpwr scs8hd_fill_1
XFILLER_505_15 vgnd vpwr scs8hd_decap_12
XFILLER_224_27 vgnd vpwr scs8hd_decap_4
XFILLER_505_59 vpwr vgnd scs8hd_fill_2
XFILLER_240_15 vgnd vpwr scs8hd_decap_12
XFILLER_601_80 vgnd vpwr scs8hd_fill_1
XFILLER_546_44 vgnd vpwr scs8hd_decap_12
XFILLER_562_32 vgnd vpwr scs8hd_decap_12
XFILLER_415_15 vgnd vpwr scs8hd_decap_12
XFILLER_415_59 vpwr vgnd scs8hd_fill_2
XFILLER_134_27 vgnd vpwr scs8hd_decap_4
XFILLER_150_15 vgnd vpwr scs8hd_decap_12
XFILLER_511_80 vgnd vpwr scs8hd_fill_1
XFILLER_587_62 vgnd vpwr scs8hd_decap_12
XFILLER_587_51 vgnd vpwr scs8hd_decap_8
XFILLER_309_27 vgnd vpwr scs8hd_decap_12
XFILLER_456_44 vgnd vpwr scs8hd_decap_12
XFILLER_111_3 vgnd vpwr scs8hd_decap_12
XFILLER_209_3 vgnd vpwr scs8hd_decap_4
XFILLER_325_15 vgnd vpwr scs8hd_decap_12
XFILLER_472_32 vgnd vpwr scs8hd_decap_12
XFILLER_68_32 vgnd vpwr scs8hd_decap_12
XFILLER_325_59 vpwr vgnd scs8hd_fill_2
XFILLER_480_3 vgnd vpwr scs8hd_decap_12
XFILLER_578_3 vgnd vpwr scs8hd_decap_12
XFILLER_421_80 vgnd vpwr scs8hd_fill_1
XFILLER_17_80 vgnd vpwr scs8hd_fill_1
XFILLER_497_51 vgnd vpwr scs8hd_decap_8
XFILLER_497_62 vgnd vpwr scs8hd_decap_12
XPHY_260 vgnd vpwr scs8hd_decap_3
XPHY_271 vgnd vpwr scs8hd_decap_3
XPHY_282 vgnd vpwr scs8hd_decap_3
XPHY_293 vgnd vpwr scs8hd_decap_3
XFILLER_366_44 vgnd vpwr scs8hd_decap_12
XFILLER_235_15 vgnd vpwr scs8hd_decap_12
XFILLER_382_32 vgnd vpwr scs8hd_decap_12
XFILLER_235_59 vpwr vgnd scs8hd_fill_2
XFILLER_532_68 vgnd vpwr scs8hd_decap_12
XFILLER_331_80 vgnd vpwr scs8hd_fill_1
XFILLER_401_39 vgnd vpwr scs8hd_decap_12
XPHY_1809 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_13_27 vgnd vpwr scs8hd_decap_12
XFILLER_129_27 vgnd vpwr scs8hd_decap_12
XFILLER_276_44 vgnd vpwr scs8hd_decap_12
XFILLER_145_15 vgnd vpwr scs8hd_decap_12
XFILLER_292_32 vgnd vpwr scs8hd_decap_12
XFILLER_145_59 vpwr vgnd scs8hd_fill_2
XFILLER_506_80 vgnd vpwr scs8hd_fill_1
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_442_68 vgnd vpwr scs8hd_decap_12
XFILLER_241_80 vgnd vpwr scs8hd_fill_1
XFILLER_311_39 vgnd vpwr scs8hd_decap_12
XFILLER_54_56 vgnd vpwr scs8hd_decap_12
XFILLER_159_3 vgnd vpwr scs8hd_decap_12
XFILLER_70_44 vgnd vpwr scs8hd_decap_12
XFILLER_326_3 vgnd vpwr scs8hd_decap_12
XFILLER_186_44 vgnd vpwr scs8hd_decap_12
XFILLER_205_18 vpwr vgnd scs8hd_fill_2
XFILLER_416_80 vgnd vpwr scs8hd_fill_1
XFILLER_95_74 vgnd vpwr scs8hd_decap_6
XFILLER_352_68 vgnd vpwr scs8hd_decap_12
XFILLER_502_27 vgnd vpwr scs8hd_decap_4
XFILLER_221_39 vgnd vpwr scs8hd_decap_12
XFILLER_151_80 vgnd vpwr scs8hd_fill_1
XFILLER_74_3 vgnd vpwr scs8hd_decap_12
XFILLER_326_80 vgnd vpwr scs8hd_fill_1
XFILLER_262_68 vgnd vpwr scs8hd_decap_12
XFILLER_412_27 vgnd vpwr scs8hd_decap_4
XFILLER_131_39 vgnd vpwr scs8hd_decap_12
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
XPHY_1606 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1617 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1628 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1639 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__13__D _08_/Y vgnd vpwr scs8hd_diode_2
XFILLER_200_7 vgnd vpwr scs8hd_decap_3
XFILLER_236_80 vgnd vpwr scs8hd_fill_1
XFILLER_603_15 vgnd vpwr scs8hd_decap_12
XFILLER_105_51 vgnd vpwr scs8hd_decap_8
XFILLER_172_68 vgnd vpwr scs8hd_decap_12
XFILLER_105_62 vgnd vpwr scs8hd_decap_12
XFILLER_322_27 vgnd vpwr scs8hd_decap_4
XFILLER_276_3 vgnd vpwr scs8hd_decap_12
XFILLER_443_3 vgnd vpwr scs8hd_decap_12
XFILLER_30_80 vgnd vpwr scs8hd_fill_1
XFILLER_146_80 vgnd vpwr scs8hd_fill_1
XFILLER_513_15 vgnd vpwr scs8hd_decap_12
XFILLER_513_59 vpwr vgnd scs8hd_fill_2
XFILLER_232_27 vgnd vpwr scs8hd_decap_4
XFILLER_538_56 vgnd vpwr scs8hd_decap_12
XFILLER_554_44 vgnd vpwr scs8hd_decap_12
XFILLER_407_27 vgnd vpwr scs8hd_decap_12
XFILLER_570_32 vgnd vpwr scs8hd_decap_12
XFILLER_423_15 vgnd vpwr scs8hd_decap_12
XFILLER_19_15 vgnd vpwr scs8hd_decap_12
XFILLER_423_59 vpwr vgnd scs8hd_fill_2
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
XFILLER_142_27 vgnd vpwr scs8hd_decap_4
XFILLER_579_74 vgnd vpwr scs8hd_decap_6
XPHY_804 vgnd vpwr scs8hd_decap_3
XPHY_815 vgnd vpwr scs8hd_decap_3
XPHY_826 vgnd vpwr scs8hd_decap_3
XPHY_1403 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1414 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_837 vgnd vpwr scs8hd_decap_3
XPHY_848 vgnd vpwr scs8hd_decap_3
XPHY_859 vgnd vpwr scs8hd_decap_3
XFILLER_595_62 vgnd vpwr scs8hd_decap_12
XFILLER_595_51 vgnd vpwr scs8hd_decap_8
XPHY_1425 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1436 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1447 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1458 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_448_56 vgnd vpwr scs8hd_decap_12
XPHY_1469 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_317_27 vgnd vpwr scs8hd_decap_12
XFILLER_464_44 vgnd vpwr scs8hd_decap_12
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XFILLER_333_15 vgnd vpwr scs8hd_decap_12
XFILLER_393_3 vgnd vpwr scs8hd_decap_12
XFILLER_76_32 vgnd vpwr scs8hd_decap_12
XFILLER_333_59 vpwr vgnd scs8hd_fill_2
XFILLER_480_32 vgnd vpwr scs8hd_decap_12
XFILLER_560_3 vgnd vpwr scs8hd_decap_12
XFILLER_489_74 vgnd vpwr scs8hd_decap_6
XPHY_91 vgnd vpwr scs8hd_decap_3
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_25_80 vgnd vpwr scs8hd_fill_1
XFILLER_358_56 vgnd vpwr scs8hd_decap_12
XFILLER_508_15 vgnd vpwr scs8hd_decap_12
XFILLER_227_27 vgnd vpwr scs8hd_decap_12
XFILLER_374_44 vgnd vpwr scs8hd_decap_12
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
XFILLER_243_15 vgnd vpwr scs8hd_decap_12
XFILLER_243_59 vpwr vgnd scs8hd_fill_2
XFILLER_390_32 vgnd vpwr scs8hd_decap_12
XFILLER_540_68 vgnd vpwr scs8hd_decap_12
XFILLER_399_74 vgnd vpwr scs8hd_decap_6
XFILLER_268_56 vgnd vpwr scs8hd_decap_12
XFILLER_418_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_27 vgnd vpwr scs8hd_decap_12
XFILLER_137_27 vgnd vpwr scs8hd_decap_12
XFILLER_284_44 vgnd vpwr scs8hd_decap_12
XFILLER_153_15 vgnd vpwr scs8hd_decap_12
XFILLER_153_59 vpwr vgnd scs8hd_fill_2
XFILLER_514_80 vgnd vpwr scs8hd_fill_1
XFILLER_46_68 vgnd vpwr scs8hd_decap_12
XFILLER_450_68 vgnd vpwr scs8hd_decap_12
XFILLER_600_27 vgnd vpwr scs8hd_decap_4
XPHY_601 vgnd vpwr scs8hd_decap_3
XPHY_612 vgnd vpwr scs8hd_decap_3
XPHY_623 vgnd vpwr scs8hd_decap_3
XPHY_634 vgnd vpwr scs8hd_decap_3
XPHY_1200 vgnd vpwr scs8hd_decap_3
XFILLER_62_56 vgnd vpwr scs8hd_decap_12
XPHY_1211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_141_3 vgnd vpwr scs8hd_decap_12
XFILLER_239_3 vgnd vpwr scs8hd_decap_12
XPHY_645 vgnd vpwr scs8hd_decap_3
XPHY_656 vgnd vpwr scs8hd_decap_3
XPHY_667 vgnd vpwr scs8hd_decap_3
XPHY_678 vgnd vpwr scs8hd_decap_3
XPHY_1266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_178_56 vgnd vpwr scs8hd_decap_12
XFILLER_328_15 vgnd vpwr scs8hd_decap_12
XPHY_689 vgnd vpwr scs8hd_decap_3
XPHY_1299 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1288 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_406_3 vgnd vpwr scs8hd_decap_12
XFILLER_194_44 vgnd vpwr scs8hd_decap_12
XFILLER_424_80 vgnd vpwr scs8hd_fill_1
XFILLER_360_68 vgnd vpwr scs8hd_decap_12
XFILLER_510_27 vgnd vpwr scs8hd_decap_4
XFILLER_238_15 vgnd vpwr scs8hd_decap_12
XFILLER_334_80 vgnd vpwr scs8hd_fill_1
XFILLER_270_68 vgnd vpwr scs8hd_decap_12
XFILLER_203_62 vgnd vpwr scs8hd_decap_12
XFILLER_420_27 vgnd vpwr scs8hd_decap_4
XFILLER_16_27 vgnd vpwr scs8hd_decap_4
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XFILLER_148_15 vgnd vpwr scs8hd_decap_12
XFILLER_509_80 vgnd vpwr scs8hd_fill_1
XFILLER_244_80 vgnd vpwr scs8hd_fill_1
XFILLER_189_3 vgnd vpwr scs8hd_decap_8
XFILLER_113_62 vgnd vpwr scs8hd_decap_12
XFILLER_113_51 vgnd vpwr scs8hd_decap_8
XFILLER_330_27 vgnd vpwr scs8hd_decap_4
XFILLER_189_11 vpwr vgnd scs8hd_fill_2
XFILLER_356_3 vgnd vpwr scs8hd_decap_12
XFILLER_523_3 vgnd vpwr scs8hd_decap_12
XPHY_420 vgnd vpwr scs8hd_decap_3
XPHY_431 vgnd vpwr scs8hd_decap_3
XPHY_442 vgnd vpwr scs8hd_decap_3
XPHY_453 vgnd vpwr scs8hd_decap_3
XPHY_464 vgnd vpwr scs8hd_decap_3
XPHY_475 vgnd vpwr scs8hd_decap_3
XPHY_486 vgnd vpwr scs8hd_decap_3
XPHY_1030 vgnd vpwr scs8hd_decap_3
XPHY_1041 vgnd vpwr scs8hd_decap_3
XPHY_1074 vgnd vpwr scs8hd_decap_3
XPHY_1063 vgnd vpwr scs8hd_decap_3
XPHY_1052 vgnd vpwr scs8hd_decap_3
XPHY_497 vgnd vpwr scs8hd_decap_3
XPHY_1096 vgnd vpwr scs8hd_decap_3
XPHY_1085 vgnd vpwr scs8hd_decap_3
XFILLER_419_80 vgnd vpwr scs8hd_fill_1
XFILLER_505_27 vgnd vpwr scs8hd_decap_12
XFILLER_154_80 vgnd vpwr scs8hd_fill_1
XFILLER_521_15 vgnd vpwr scs8hd_decap_12
XFILLER_240_27 vgnd vpwr scs8hd_decap_4
XFILLER_521_59 vpwr vgnd scs8hd_fill_2
XFILLER_329_80 vgnd vpwr scs8hd_fill_1
XFILLER_546_56 vgnd vpwr scs8hd_decap_12
XFILLER_415_27 vgnd vpwr scs8hd_decap_12
XFILLER_562_44 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _14_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_431_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_59 vpwr vgnd scs8hd_fill_2
XFILLER_150_27 vgnd vpwr scs8hd_decap_4
XFILLER_431_59 vpwr vgnd scs8hd_fill_2
XFILLER_587_74 vgnd vpwr scs8hd_decap_6
XFILLER_239_80 vgnd vpwr scs8hd_fill_1
XFILLER_309_39 vgnd vpwr scs8hd_decap_12
XFILLER_456_56 vgnd vpwr scs8hd_decap_12
XFILLER_104_3 vgnd vpwr scs8hd_decap_12
XFILLER_325_27 vgnd vpwr scs8hd_decap_12
XFILLER_68_44 vgnd vpwr scs8hd_decap_12
XFILLER_472_44 vgnd vpwr scs8hd_decap_12
XFILLER_341_15 vgnd vpwr scs8hd_decap_12
XFILLER_473_3 vgnd vpwr scs8hd_decap_12
XFILLER_84_32 vgnd vpwr scs8hd_decap_12
XFILLER_341_59 vpwr vgnd scs8hd_fill_2
XPHY_261 vgnd vpwr scs8hd_decap_3
XPHY_250 vgnd vpwr scs8hd_decap_3
XFILLER_497_74 vgnd vpwr scs8hd_decap_6
XPHY_272 vgnd vpwr scs8hd_decap_3
XPHY_283 vgnd vpwr scs8hd_decap_3
XPHY_294 vgnd vpwr scs8hd_decap_3
XFILLER_33_80 vgnd vpwr scs8hd_fill_1
XFILLER_149_80 vgnd vpwr scs8hd_fill_1
XFILLER_219_17 vgnd vpwr scs8hd_decap_12
XFILLER_366_56 vgnd vpwr scs8hd_decap_12
XFILLER_516_15 vgnd vpwr scs8hd_decap_12
XFILLER_235_27 vgnd vpwr scs8hd_decap_12
XFILLER_382_44 vgnd vpwr scs8hd_decap_12
XFILLER_251_15 vgnd vpwr scs8hd_decap_12
XFILLER_251_59 vpwr vgnd scs8hd_fill_2
XFILLER_200_30 vgnd vpwr scs8hd_fill_1
XFILLER_13_39 vgnd vpwr scs8hd_decap_12
XFILLER_129_39 vgnd vpwr scs8hd_decap_12
XFILLER_276_56 vgnd vpwr scs8hd_decap_12
XFILLER_426_15 vgnd vpwr scs8hd_decap_12
XFILLER_145_27 vgnd vpwr scs8hd_decap_12
XFILLER_292_44 vgnd vpwr scs8hd_decap_12
XFILLER_225_60 vgnd vpwr scs8hd_fill_1
XFILLER_161_15 vgnd vpwr scs8hd_decap_12
XFILLER_522_80 vgnd vpwr scs8hd_fill_1
XFILLER_161_59 vpwr vgnd scs8hd_fill_2
XFILLER_54_68 vgnd vpwr scs8hd_decap_12
XFILLER_70_56 vgnd vpwr scs8hd_decap_12
XFILLER_221_3 vgnd vpwr scs8hd_decap_12
XFILLER_186_56 vgnd vpwr scs8hd_decap_12
XFILLER_319_3 vgnd vpwr scs8hd_decap_12
XFILLER_336_15 vgnd vpwr scs8hd_decap_12
XFILLER_590_3 vgnd vpwr scs8hd_decap_12
XFILLER_432_80 vgnd vpwr scs8hd_fill_1
XFILLER_28_80 vgnd vpwr scs8hd_fill_1
XFILLER_301_51 vgnd vpwr scs8hd_decap_8
XFILLER_301_62 vgnd vpwr scs8hd_decap_12
XFILLER_67_3 vgnd vpwr scs8hd_decap_12
XFILLER_246_15 vgnd vpwr scs8hd_decap_12
XFILLER_5_62 vgnd vpwr scs8hd_decap_12
XFILLER_5_51 vgnd vpwr scs8hd_decap_8
XFILLER_342_80 vgnd vpwr scs8hd_fill_1
XFILLER_568_32 vgnd vpwr scs8hd_decap_12
XFILLER_211_51 vpwr vgnd scs8hd_fill_2
XFILLER_211_62 vgnd vpwr scs8hd_decap_12
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XPHY_1607 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1618 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1629 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_156_15 vgnd vpwr scs8hd_decap_12
XFILLER_517_80 vgnd vpwr scs8hd_fill_1
XFILLER_603_27 vgnd vpwr scs8hd_decap_4
XFILLER_105_74 vgnd vpwr scs8hd_decap_6
XFILLER_252_80 vgnd vpwr scs8hd_fill_1
XFILLER_171_3 vgnd vpwr scs8hd_decap_12
XFILLER_269_3 vgnd vpwr scs8hd_decap_12
XFILLER_121_62 vgnd vpwr scs8hd_decap_12
XFILLER_121_51 vgnd vpwr scs8hd_decap_8
XFILLER_478_32 vgnd vpwr scs8hd_decap_12
XFILLER_436_3 vgnd vpwr scs8hd_decap_12
XFILLER_603_3 vgnd vpwr scs8hd_decap_12
XFILLER_427_80 vgnd vpwr scs8hd_fill_1
XFILLER_513_27 vgnd vpwr scs8hd_decap_12
XFILLER_162_80 vgnd vpwr scs8hd_fill_1
XFILLER_388_32 vgnd vpwr scs8hd_decap_12
XFILLER_538_68 vgnd vpwr scs8hd_decap_12
XFILLER_407_39 vgnd vpwr scs8hd_decap_12
XFILLER_554_56 vgnd vpwr scs8hd_decap_12
XFILLER_337_80 vgnd vpwr scs8hd_fill_1
XFILLER_570_44 vgnd vpwr scs8hd_decap_12
XFILLER_19_27 vgnd vpwr scs8hd_decap_12
XFILLER_423_27 vgnd vpwr scs8hd_decap_12
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XFILLER_298_32 vgnd vpwr scs8hd_decap_12
XPHY_805 vgnd vpwr scs8hd_decap_3
XPHY_816 vgnd vpwr scs8hd_decap_3
XPHY_827 vgnd vpwr scs8hd_decap_3
XPHY_1404 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1415 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_838 vgnd vpwr scs8hd_decap_3
XPHY_849 vgnd vpwr scs8hd_decap_3
XPHY_1426 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1437 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1448 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_595_74 vgnd vpwr scs8hd_decap_6
XPHY_1459 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_448_68 vgnd vpwr scs8hd_decap_12
XFILLER_317_39 vgnd vpwr scs8hd_decap_12
XFILLER_247_80 vgnd vpwr scs8hd_fill_1
XFILLER_464_56 vgnd vpwr scs8hd_decap_12
XFILLER_333_27 vgnd vpwr scs8hd_decap_12
XFILLER_386_3 vgnd vpwr scs8hd_decap_12
XFILLER_480_44 vgnd vpwr scs8hd_decap_12
XFILLER_76_44 vgnd vpwr scs8hd_decap_12
XFILLER_553_3 vgnd vpwr scs8hd_decap_12
XFILLER_92_32 vgnd vpwr scs8hd_decap_12
XPHY_92 vgnd vpwr scs8hd_decap_3
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XFILLER_358_68 vgnd vpwr scs8hd_decap_12
XFILLER_508_27 vgnd vpwr scs8hd_decap_4
XFILLER_41_80 vgnd vpwr scs8hd_fill_1
XFILLER_157_80 vgnd vpwr scs8hd_fill_1
XFILLER_227_39 vgnd vpwr scs8hd_decap_12
XFILLER_374_56 vgnd vpwr scs8hd_decap_12
XFILLER_524_15 vgnd vpwr scs8hd_decap_12
XFILLER_243_27 vgnd vpwr scs8hd_decap_12
XFILLER_390_44 vgnd vpwr scs8hd_decap_12
XFILLER_268_68 vgnd vpwr scs8hd_decap_12
XFILLER_418_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_39 vgnd vpwr scs8hd_decap_12
XFILLER_137_39 vgnd vpwr scs8hd_decap_12
XFILLER_284_56 vgnd vpwr scs8hd_decap_12
XFILLER_217_50 vgnd vpwr scs8hd_decap_8
XFILLER_434_15 vgnd vpwr scs8hd_decap_12
XFILLER_153_27 vgnd vpwr scs8hd_decap_12
XFILLER_530_80 vgnd vpwr scs8hd_fill_1
XPHY_602 vgnd vpwr scs8hd_decap_3
XPHY_613 vgnd vpwr scs8hd_decap_3
XPHY_624 vgnd vpwr scs8hd_decap_3
XPHY_635 vgnd vpwr scs8hd_decap_3
XPHY_1201 vgnd vpwr scs8hd_decap_3
XFILLER_62_68 vgnd vpwr scs8hd_decap_12
XPHY_1212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_646 vgnd vpwr scs8hd_decap_3
XPHY_657 vgnd vpwr scs8hd_decap_3
XPHY_668 vgnd vpwr scs8hd_decap_3
XPHY_1256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_134_3 vgnd vpwr scs8hd_decap_12
XFILLER_178_68 vgnd vpwr scs8hd_decap_12
XPHY_679 vgnd vpwr scs8hd_decap_3
XPHY_1289 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_328_27 vgnd vpwr scs8hd_decap_4
XFILLER_194_12 vpwr vgnd scs8hd_fill_2
XFILLER_301_3 vgnd vpwr scs8hd_decap_12
XFILLER_194_56 vgnd vpwr scs8hd_decap_12
XFILLER_344_15 vgnd vpwr scs8hd_decap_12
XFILLER_36_80 vgnd vpwr scs8hd_fill_1
XFILLER_440_80 vgnd vpwr scs8hd_fill_1
XFILLER_519_15 vgnd vpwr scs8hd_decap_12
XFILLER_519_59 vpwr vgnd scs8hd_fill_2
XFILLER_238_27 vgnd vpwr scs8hd_decap_4
XPHY_1790 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_254_15 vgnd vpwr scs8hd_decap_12
XFILLER_203_30 vpwr vgnd scs8hd_fill_2
XFILLER_203_74 vgnd vpwr scs8hd_decap_6
XFILLER_350_80 vgnd vpwr scs8hd_fill_1
XFILLER_429_15 vgnd vpwr scs8hd_decap_12
XFILLER_576_32 vgnd vpwr scs8hd_decap_12
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XFILLER_148_27 vgnd vpwr scs8hd_decap_4
XFILLER_295_11 vgnd vpwr scs8hd_decap_12
XFILLER_429_59 vpwr vgnd scs8hd_fill_2
XFILLER_164_15 vgnd vpwr scs8hd_decap_12
XFILLER_525_80 vgnd vpwr scs8hd_fill_1
XFILLER_113_74 vgnd vpwr scs8hd_decap_6
XFILLER_260_80 vgnd vpwr scs8hd_fill_1
XPHY_410 vgnd vpwr scs8hd_decap_3
XFILLER_251_3 vgnd vpwr scs8hd_decap_12
XFILLER_349_3 vgnd vpwr scs8hd_decap_12
XPHY_421 vgnd vpwr scs8hd_decap_3
XPHY_432 vgnd vpwr scs8hd_decap_3
XPHY_443 vgnd vpwr scs8hd_decap_3
XFILLER_339_15 vgnd vpwr scs8hd_decap_12
XPHY_454 vgnd vpwr scs8hd_decap_3
XPHY_465 vgnd vpwr scs8hd_decap_3
XPHY_476 vgnd vpwr scs8hd_decap_3
XFILLER_486_32 vgnd vpwr scs8hd_decap_12
XPHY_1020 vgnd vpwr scs8hd_decap_3
XFILLER_516_3 vgnd vpwr scs8hd_decap_12
XPHY_1031 vgnd vpwr scs8hd_decap_3
XPHY_1064 vgnd vpwr scs8hd_decap_3
XPHY_1053 vgnd vpwr scs8hd_decap_3
XPHY_487 vgnd vpwr scs8hd_decap_3
XPHY_498 vgnd vpwr scs8hd_decap_3
XFILLER_339_59 vpwr vgnd scs8hd_fill_2
XPHY_1042 vgnd vpwr scs8hd_decap_3
XPHY_1097 vgnd vpwr scs8hd_decap_3
XPHY_1086 vgnd vpwr scs8hd_decap_3
XPHY_1075 vgnd vpwr scs8hd_decap_3
XFILLER_208_19 vpwr vgnd scs8hd_fill_2
XFILLER_435_80 vgnd vpwr scs8hd_fill_1
XFILLER_505_39 vgnd vpwr scs8hd_decap_12
XFILLER_521_27 vgnd vpwr scs8hd_decap_12
XFILLER_170_80 vgnd vpwr scs8hd_fill_1
XFILLER_97_3 vgnd vpwr scs8hd_decap_12
XFILLER_249_15 vgnd vpwr scs8hd_decap_12
XFILLER_396_32 vgnd vpwr scs8hd_decap_12
XFILLER_249_59 vpwr vgnd scs8hd_fill_2
XFILLER_546_68 vgnd vpwr scs8hd_decap_12
XFILLER_562_56 vgnd vpwr scs8hd_decap_12
XFILLER_345_80 vgnd vpwr scs8hd_fill_1
XFILLER_415_39 vgnd vpwr scs8hd_decap_12
XFILLER_27_27 vgnd vpwr scs8hd_decap_12
XFILLER_431_27 vgnd vpwr scs8hd_decap_12
XFILLER_43_15 vgnd vpwr scs8hd_decap_12
XFILLER_43_59 vpwr vgnd scs8hd_fill_2
XFILLER_159_15 vgnd vpwr scs8hd_decap_12
XFILLER_159_59 vpwr vgnd scs8hd_fill_2
XFILLER_456_68 vgnd vpwr scs8hd_decap_12
XFILLER_255_80 vgnd vpwr scs8hd_fill_1
XFILLER_325_39 vgnd vpwr scs8hd_decap_12
XFILLER_472_56 vgnd vpwr scs8hd_decap_12
XFILLER_68_56 vgnd vpwr scs8hd_decap_12
XFILLER_299_3 vgnd vpwr scs8hd_decap_12
XFILLER_341_27 vgnd vpwr scs8hd_decap_12
XFILLER_84_44 vgnd vpwr scs8hd_decap_12
XFILLER_466_3 vgnd vpwr scs8hd_decap_12
XPHY_251 vgnd vpwr scs8hd_decap_3
XPHY_240 vgnd vpwr scs8hd_decap_3
XPHY_262 vgnd vpwr scs8hd_decap_3
XPHY_273 vgnd vpwr scs8hd_decap_3
XPHY_284 vgnd vpwr scs8hd_decap_3
XPHY_295 vgnd vpwr scs8hd_decap_3
XFILLER_219_29 vgnd vpwr scs8hd_decap_12
XFILLER_366_68 vgnd vpwr scs8hd_decap_12
XFILLER_516_27 vgnd vpwr scs8hd_decap_4
XFILLER_235_39 vgnd vpwr scs8hd_decap_12
XFILLER_382_56 vgnd vpwr scs8hd_decap_12
XFILLER_532_15 vgnd vpwr scs8hd_decap_12
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_251_27 vgnd vpwr scs8hd_decap_12
XFILLER_276_68 vgnd vpwr scs8hd_decap_12
XFILLER_209_62 vgnd vpwr scs8hd_decap_12
XFILLER_426_27 vgnd vpwr scs8hd_decap_4
XFILLER_145_39 vgnd vpwr scs8hd_decap_12
XFILLER_292_56 vgnd vpwr scs8hd_decap_12
XFILLER_442_15 vgnd vpwr scs8hd_decap_12
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XFILLER_161_27 vgnd vpwr scs8hd_decap_12
XFILLER_70_68 vgnd vpwr scs8hd_decap_12
XFILLER_186_68 vgnd vpwr scs8hd_decap_12
XFILLER_214_3 vgnd vpwr scs8hd_decap_12
XFILLER_119_62 vgnd vpwr scs8hd_decap_12
XFILLER_119_51 vgnd vpwr scs8hd_decap_8
XFILLER_336_27 vgnd vpwr scs8hd_decap_4
XFILLER_583_3 vgnd vpwr scs8hd_decap_12
XFILLER_352_15 vgnd vpwr scs8hd_decap_12
XFILLER_44_80 vgnd vpwr scs8hd_fill_1
XFILLER_301_74 vgnd vpwr scs8hd_decap_6
XFILLER_527_15 vgnd vpwr scs8hd_decap_12
XFILLER_527_59 vpwr vgnd scs8hd_fill_2
XFILLER_246_27 vgnd vpwr scs8hd_decap_4
XFILLER_5_74 vgnd vpwr scs8hd_decap_6
XFILLER_262_15 vgnd vpwr scs8hd_decap_12
XFILLER_568_44 vgnd vpwr scs8hd_decap_12
XFILLER_211_74 vgnd vpwr scs8hd_decap_6
XPHY_1608 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1619 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_584_32 vgnd vpwr scs8hd_decap_12
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XFILLER_437_15 vgnd vpwr scs8hd_decap_12
XFILLER_156_27 vgnd vpwr scs8hd_decap_4
XFILLER_437_59 vpwr vgnd scs8hd_fill_2
XFILLER_172_15 vgnd vpwr scs8hd_decap_12
XFILLER_533_80 vgnd vpwr scs8hd_fill_1
XFILLER_164_3 vgnd vpwr scs8hd_decap_12
XFILLER_121_74 vgnd vpwr scs8hd_decap_6
XFILLER_478_44 vgnd vpwr scs8hd_decap_12
XFILLER_331_3 vgnd vpwr scs8hd_decap_12
XFILLER_429_3 vgnd vpwr scs8hd_decap_12
XFILLER_347_15 vgnd vpwr scs8hd_decap_12
XFILLER_494_32 vgnd vpwr scs8hd_decap_12
XFILLER_347_59 vpwr vgnd scs8hd_fill_2
XFILLER_443_80 vgnd vpwr scs8hd_fill_1
XFILLER_513_39 vgnd vpwr scs8hd_decap_12
XFILLER_39_80 vgnd vpwr scs8hd_fill_1
XFILLER_388_44 vgnd vpwr scs8hd_decap_12
XFILLER_257_15 vgnd vpwr scs8hd_decap_12
XFILLER_257_59 vpwr vgnd scs8hd_fill_2
XFILLER_554_68 vgnd vpwr scs8hd_decap_12
XFILLER_206_30 vgnd vpwr scs8hd_fill_1
XFILLER_570_56 vgnd vpwr scs8hd_decap_12
XFILLER_353_80 vgnd vpwr scs8hd_fill_1
XFILLER_423_39 vgnd vpwr scs8hd_decap_12
XFILLER_19_39 vgnd vpwr scs8hd_decap_12
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XFILLER_298_44 vgnd vpwr scs8hd_decap_12
XPHY_806 vgnd vpwr scs8hd_decap_3
XPHY_817 vgnd vpwr scs8hd_decap_3
XPHY_1405 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_828 vgnd vpwr scs8hd_decap_3
XPHY_839 vgnd vpwr scs8hd_decap_3
XFILLER_51_15 vgnd vpwr scs8hd_decap_12
XPHY_1416 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1427 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1438 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1449 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_59 vpwr vgnd scs8hd_fill_2
XFILLER_167_15 vgnd vpwr scs8hd_decap_12
XFILLER_528_80 vgnd vpwr scs8hd_fill_1
XFILLER_167_59 vpwr vgnd scs8hd_fill_2
XFILLER_464_68 vgnd vpwr scs8hd_decap_12
XFILLER_263_80 vgnd vpwr scs8hd_fill_1
XFILLER_333_39 vgnd vpwr scs8hd_decap_12
XFILLER_480_56 vgnd vpwr scs8hd_decap_12
XFILLER_76_56 vgnd vpwr scs8hd_decap_12
XFILLER_281_3 vgnd vpwr scs8hd_decap_12
XFILLER_379_3 vgnd vpwr scs8hd_decap_12
XFILLER_546_3 vgnd vpwr scs8hd_decap_12
XFILLER_92_44 vgnd vpwr scs8hd_decap_12
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XPHY_93 vgnd vpwr scs8hd_decap_3
XFILLER_438_80 vgnd vpwr scs8hd_fill_1
XFILLER_374_68 vgnd vpwr scs8hd_decap_12
XFILLER_524_27 vgnd vpwr scs8hd_decap_4
XFILLER_307_51 vgnd vpwr scs8hd_decap_8
XFILLER_307_62 vgnd vpwr scs8hd_decap_12
XFILLER_173_80 vgnd vpwr scs8hd_fill_1
XFILLER_243_39 vgnd vpwr scs8hd_decap_12
XFILLER_390_56 vgnd vpwr scs8hd_decap_12
XFILLER_540_15 vgnd vpwr scs8hd_decap_12
XFILLER_348_80 vgnd vpwr scs8hd_fill_1
XFILLER_284_68 vgnd vpwr scs8hd_decap_12
XFILLER_434_27 vgnd vpwr scs8hd_decap_4
XFILLER_217_62 vgnd vpwr scs8hd_decap_12
XFILLER_153_39 vgnd vpwr scs8hd_decap_12
XFILLER_46_15 vgnd vpwr scs8hd_decap_12
XFILLER_450_15 vgnd vpwr scs8hd_decap_12
XFILLER_102_32 vgnd vpwr scs8hd_decap_12
XPHY_603 vgnd vpwr scs8hd_decap_3
XPHY_614 vgnd vpwr scs8hd_decap_3
XPHY_625 vgnd vpwr scs8hd_decap_3
XPHY_1202 vgnd vpwr scs8hd_decap_3
XPHY_1213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_636 vgnd vpwr scs8hd_decap_3
XPHY_647 vgnd vpwr scs8hd_decap_3
XPHY_658 vgnd vpwr scs8hd_decap_3
XPHY_669 vgnd vpwr scs8hd_decap_3
XPHY_1257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_127_3 vgnd vpwr scs8hd_decap_12
XPHY_1279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_258_80 vgnd vpwr scs8hd_fill_1
XFILLER_11_51 vgnd vpwr scs8hd_decap_8
XFILLER_127_51 vgnd vpwr scs8hd_decap_8
XFILLER_11_62 vgnd vpwr scs8hd_decap_12
XFILLER_194_68 vgnd vpwr scs8hd_decap_12
XFILLER_127_62 vgnd vpwr scs8hd_decap_12
XFILLER_344_27 vgnd vpwr scs8hd_decap_4
XFILLER_496_3 vgnd vpwr scs8hd_decap_12
XFILLER_360_15 vgnd vpwr scs8hd_decap_12
XFILLER_519_27 vgnd vpwr scs8hd_decap_12
XFILLER_52_80 vgnd vpwr scs8hd_fill_1
XPHY_1791 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1780 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_168_80 vgnd vpwr scs8hd_fill_1
XFILLER_535_15 vgnd vpwr scs8hd_decap_12
XFILLER_535_59 vpwr vgnd scs8hd_fill_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_254_27 vgnd vpwr scs8hd_decap_4
XFILLER_270_15 vgnd vpwr scs8hd_decap_12
XFILLER_576_44 vgnd vpwr scs8hd_decap_12
XFILLER_429_27 vgnd vpwr scs8hd_decap_12
XFILLER_295_23 vgnd vpwr scs8hd_decap_12
XFILLER_592_32 vgnd vpwr scs8hd_decap_12
XFILLER_445_15 vgnd vpwr scs8hd_decap_12
XFILLER_445_59 vpwr vgnd scs8hd_fill_2
XFILLER_164_27 vgnd vpwr scs8hd_decap_4
XFILLER_180_15 vgnd vpwr scs8hd_decap_12
XFILLER_541_80 vgnd vpwr scs8hd_fill_1
XPHY_400 vgnd vpwr scs8hd_decap_3
XPHY_411 vgnd vpwr scs8hd_decap_3
XPHY_422 vgnd vpwr scs8hd_decap_3
XPHY_433 vgnd vpwr scs8hd_decap_3
XPHY_444 vgnd vpwr scs8hd_decap_3
XFILLER_244_3 vgnd vpwr scs8hd_decap_12
XPHY_455 vgnd vpwr scs8hd_decap_3
XPHY_466 vgnd vpwr scs8hd_decap_3
XPHY_477 vgnd vpwr scs8hd_decap_3
XFILLER_339_27 vgnd vpwr scs8hd_decap_12
XFILLER_486_44 vgnd vpwr scs8hd_decap_12
XPHY_1010 vgnd vpwr scs8hd_decap_3
XPHY_1021 vgnd vpwr scs8hd_decap_3
XPHY_1032 vgnd vpwr scs8hd_decap_3
XPHY_1065 vgnd vpwr scs8hd_decap_3
XPHY_1054 vgnd vpwr scs8hd_decap_3
XPHY_1043 vgnd vpwr scs8hd_decap_3
XPHY_488 vgnd vpwr scs8hd_decap_3
XPHY_499 vgnd vpwr scs8hd_decap_3
XFILLER_411_3 vgnd vpwr scs8hd_decap_12
XPHY_1098 vgnd vpwr scs8hd_decap_3
XPHY_1087 vgnd vpwr scs8hd_decap_3
XPHY_1076 vgnd vpwr scs8hd_decap_3
XFILLER_509_3 vgnd vpwr scs8hd_decap_12
XFILLER_355_15 vgnd vpwr scs8hd_decap_12
XFILLER_98_32 vgnd vpwr scs8hd_decap_12
XFILLER_355_59 vpwr vgnd scs8hd_fill_2
XFILLER_451_80 vgnd vpwr scs8hd_fill_1
XFILLER_521_39 vgnd vpwr scs8hd_decap_12
XFILLER_47_80 vgnd vpwr scs8hd_fill_1
Xlogical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ right_width_0_height_0__pin_0_ logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[0] vgnd vpwr scs8hd_ebufn_1
XFILLER_249_27 vgnd vpwr scs8hd_decap_12
XFILLER_396_44 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _07_/X vgnd vpwr scs8hd_diode_2
XFILLER_265_15 vgnd vpwr scs8hd_decap_12
XFILLER_265_59 vpwr vgnd scs8hd_fill_2
XFILLER_562_68 vgnd vpwr scs8hd_decap_12
XFILLER_431_39 vgnd vpwr scs8hd_decap_12
XFILLER_27_39 vgnd vpwr scs8hd_decap_12
XFILLER_361_80 vgnd vpwr scs8hd_fill_1
XFILLER_43_27 vgnd vpwr scs8hd_decap_12
XFILLER_230_73 vgnd vpwr scs8hd_decap_8
XFILLER_159_27 vgnd vpwr scs8hd_decap_12
XFILLER_175_15 vgnd vpwr scs8hd_decap_12
XFILLER_175_59 vpwr vgnd scs8hd_fill_2
XFILLER_536_80 vgnd vpwr scs8hd_fill_1
XFILLER_68_68 vgnd vpwr scs8hd_decap_12
XFILLER_405_51 vgnd vpwr scs8hd_decap_8
XFILLER_472_68 vgnd vpwr scs8hd_decap_12
XFILLER_405_62 vgnd vpwr scs8hd_decap_12
XFILLER_341_39 vgnd vpwr scs8hd_decap_12
XFILLER_84_56 vgnd vpwr scs8hd_decap_12
XFILLER_271_80 vgnd vpwr scs8hd_fill_1
XFILLER_361_3 vgnd vpwr scs8hd_decap_12
XFILLER_459_3 vgnd vpwr scs8hd_decap_12
XPHY_252 vgnd vpwr scs8hd_decap_3
XPHY_241 vgnd vpwr scs8hd_decap_3
XPHY_230 vgnd vpwr scs8hd_decap_3
XPHY_263 vgnd vpwr scs8hd_decap_3
XPHY_274 vgnd vpwr scs8hd_decap_3
XPHY_285 vgnd vpwr scs8hd_decap_3
XPHY_296 vgnd vpwr scs8hd_decap_3
XFILLER_446_80 vgnd vpwr scs8hd_fill_1
XFILLER_315_51 vgnd vpwr scs8hd_decap_8
XFILLER_382_68 vgnd vpwr scs8hd_decap_12
XFILLER_532_27 vgnd vpwr scs8hd_decap_4
XFILLER_315_62 vgnd vpwr scs8hd_decap_12
XFILLER_251_39 vgnd vpwr scs8hd_decap_12
XFILLER_181_80 vgnd vpwr scs8hd_fill_1
XFILLER_200_32 vgnd vpwr scs8hd_decap_12
XFILLER_209_74 vgnd vpwr scs8hd_decap_6
XFILLER_356_80 vgnd vpwr scs8hd_fill_1
XFILLER_292_68 vgnd vpwr scs8hd_decap_12
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
XFILLER_225_62 vgnd vpwr scs8hd_decap_12
XFILLER_442_27 vgnd vpwr scs8hd_decap_4
XFILLER_161_39 vgnd vpwr scs8hd_decap_12
XFILLER_54_15 vgnd vpwr scs8hd_decap_12
XFILLER_110_32 vgnd vpwr scs8hd_decap_12
XFILLER_119_74 vgnd vpwr scs8hd_decap_6
XFILLER_266_80 vgnd vpwr scs8hd_fill_1
XFILLER_135_51 vgnd vpwr scs8hd_decap_8
XFILLER_135_62 vgnd vpwr scs8hd_decap_12
XFILLER_352_27 vgnd vpwr scs8hd_decap_4
XFILLER_576_3 vgnd vpwr scs8hd_decap_12
XFILLER_527_27 vgnd vpwr scs8hd_decap_12
XFILLER_60_80 vgnd vpwr scs8hd_fill_1
XFILLER_176_80 vgnd vpwr scs8hd_fill_1
XFILLER_543_15 vgnd vpwr scs8hd_decap_12
XFILLER_543_59 vpwr vgnd scs8hd_fill_2
XFILLER_262_27 vgnd vpwr scs8hd_decap_4
XFILLER_568_56 vgnd vpwr scs8hd_decap_12
XPHY_1609 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_584_44 vgnd vpwr scs8hd_decap_12
XFILLER_437_27 vgnd vpwr scs8hd_decap_12
XFILLER_453_15 vgnd vpwr scs8hd_decap_12
XFILLER_49_15 vgnd vpwr scs8hd_decap_12
XFILLER_453_59 vpwr vgnd scs8hd_fill_2
XFILLER_49_59 vpwr vgnd scs8hd_fill_2
XFILLER_172_27 vgnd vpwr scs8hd_decap_4
XFILLER_157_3 vgnd vpwr scs8hd_decap_12
XFILLER_478_56 vgnd vpwr scs8hd_decap_12
XFILLER_324_3 vgnd vpwr scs8hd_decap_12
XFILLER_347_27 vgnd vpwr scs8hd_decap_12
XFILLER_494_44 vgnd vpwr scs8hd_decap_12
XFILLER_363_15 vgnd vpwr scs8hd_decap_12
XFILLER_363_59 vpwr vgnd scs8hd_fill_2
XFILLER_55_80 vgnd vpwr scs8hd_fill_1
XFILLER_388_56 vgnd vpwr scs8hd_decap_12
XFILLER_538_15 vgnd vpwr scs8hd_decap_12
XFILLER_257_27 vgnd vpwr scs8hd_decap_12
XFILLER_72_3 vgnd vpwr scs8hd_decap_12
XFILLER_273_15 vgnd vpwr scs8hd_decap_12
XFILLER_273_59 vpwr vgnd scs8hd_fill_2
XFILLER_570_68 vgnd vpwr scs8hd_decap_12
XFILLER_503_51 vgnd vpwr scs8hd_decap_8
XFILLER_503_62 vgnd vpwr scs8hd_decap_12
XFILLER_35_39 vgnd vpwr scs8hd_decap_12
XPHY_807 vgnd vpwr scs8hd_decap_3
XPHY_818 vgnd vpwr scs8hd_decap_3
XPHY_1406 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_298_56 vgnd vpwr scs8hd_decap_12
XPHY_829 vgnd vpwr scs8hd_decap_3
XFILLER_51_27 vgnd vpwr scs8hd_decap_12
XPHY_1417 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1428 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1439 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_448_15 vgnd vpwr scs8hd_decap_12
XFILLER_167_27 vgnd vpwr scs8hd_decap_12
XFILLER_183_15 vgnd vpwr scs8hd_decap_12
XFILLER_183_37 vpwr vgnd scs8hd_fill_2
XFILLER_544_80 vgnd vpwr scs8hd_fill_1
XFILLER_480_68 vgnd vpwr scs8hd_decap_12
XFILLER_76_68 vgnd vpwr scs8hd_decap_12
XFILLER_413_51 vgnd vpwr scs8hd_decap_8
XFILLER_413_62 vgnd vpwr scs8hd_decap_12
XFILLER_274_3 vgnd vpwr scs8hd_decap_12
XFILLER_539_3 vgnd vpwr scs8hd_decap_12
XFILLER_92_56 vgnd vpwr scs8hd_decap_12
XFILLER_441_3 vgnd vpwr scs8hd_decap_12
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_decap_3
XFILLER_358_15 vgnd vpwr scs8hd_decap_12
XFILLER_307_74 vgnd vpwr scs8hd_decap_6
XFILLER_454_80 vgnd vpwr scs8hd_fill_1
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_390_68 vgnd vpwr scs8hd_decap_12
XFILLER_540_27 vgnd vpwr scs8hd_decap_4
XFILLER_323_51 vgnd vpwr scs8hd_decap_8
XFILLER_323_62 vgnd vpwr scs8hd_decap_12
XFILLER_268_15 vgnd vpwr scs8hd_decap_12
XFILLER_217_74 vgnd vpwr scs8hd_decap_6
XFILLER_364_80 vgnd vpwr scs8hd_fill_1
XFILLER_233_51 vgnd vpwr scs8hd_decap_8
XFILLER_233_62 vgnd vpwr scs8hd_decap_12
XFILLER_450_27 vgnd vpwr scs8hd_decap_4
XFILLER_46_27 vgnd vpwr scs8hd_decap_4
XFILLER_102_44 vgnd vpwr scs8hd_decap_12
XFILLER_62_15 vgnd vpwr scs8hd_decap_12
XPHY_604 vgnd vpwr scs8hd_decap_3
XPHY_615 vgnd vpwr scs8hd_decap_3
XPHY_626 vgnd vpwr scs8hd_decap_3
XPHY_1203 vgnd vpwr scs8hd_decap_3
XPHY_1214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_178_15 vgnd vpwr scs8hd_decap_12
XPHY_637 vgnd vpwr scs8hd_decap_3
XPHY_648 vgnd vpwr scs8hd_decap_3
XPHY_659 vgnd vpwr scs8hd_decap_3
XFILLER_539_80 vgnd vpwr scs8hd_fill_1
XPHY_1247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_74 vgnd vpwr scs8hd_decap_6
XFILLER_127_74 vgnd vpwr scs8hd_decap_6
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_274_80 vgnd vpwr scs8hd_fill_1
XFILLER_391_3 vgnd vpwr scs8hd_decap_12
XFILLER_489_3 vgnd vpwr scs8hd_decap_12
XFILLER_143_51 vgnd vpwr scs8hd_decap_8
XFILLER_143_62 vgnd vpwr scs8hd_decap_12
XFILLER_360_27 vgnd vpwr scs8hd_decap_4
XFILLER_449_80 vgnd vpwr scs8hd_fill_1
XFILLER_519_39 vgnd vpwr scs8hd_decap_12
XPHY_1770 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1792 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1781 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_535_27 vgnd vpwr scs8hd_decap_12
XFILLER_551_15 vgnd vpwr scs8hd_decap_12
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_551_59 vpwr vgnd scs8hd_fill_2
XFILLER_270_27 vgnd vpwr scs8hd_decap_4
XFILLER_359_80 vgnd vpwr scs8hd_fill_1
XFILLER_429_39 vgnd vpwr scs8hd_decap_12
XFILLER_576_56 vgnd vpwr scs8hd_decap_12
XFILLER_295_35 vgnd vpwr scs8hd_decap_12
XFILLER_445_27 vgnd vpwr scs8hd_decap_12
XFILLER_592_44 vgnd vpwr scs8hd_decap_12
XFILLER_57_15 vgnd vpwr scs8hd_decap_12
XFILLER_461_15 vgnd vpwr scs8hd_decap_12
XFILLER_57_59 vpwr vgnd scs8hd_fill_2
XFILLER_180_27 vgnd vpwr scs8hd_decap_4
XFILLER_461_59 vpwr vgnd scs8hd_fill_2
XPHY_401 vgnd vpwr scs8hd_decap_3
XPHY_412 vgnd vpwr scs8hd_decap_3
XPHY_423 vgnd vpwr scs8hd_decap_3
XPHY_434 vgnd vpwr scs8hd_decap_3
XPHY_445 vgnd vpwr scs8hd_decap_3
XPHY_456 vgnd vpwr scs8hd_decap_3
XPHY_467 vgnd vpwr scs8hd_decap_3
XFILLER_237_3 vgnd vpwr scs8hd_decap_12
XFILLER_339_39 vgnd vpwr scs8hd_decap_12
XPHY_1000 vgnd vpwr scs8hd_decap_3
XPHY_1011 vgnd vpwr scs8hd_decap_3
XPHY_1022 vgnd vpwr scs8hd_decap_3
XPHY_1055 vgnd vpwr scs8hd_decap_3
XPHY_1044 vgnd vpwr scs8hd_decap_3
XPHY_478 vgnd vpwr scs8hd_decap_3
XPHY_489 vgnd vpwr scs8hd_decap_3
XFILLER_269_80 vgnd vpwr scs8hd_fill_1
XFILLER_486_56 vgnd vpwr scs8hd_decap_12
XPHY_1033 vgnd vpwr scs8hd_decap_3
XPHY_1099 vgnd vpwr scs8hd_decap_3
XPHY_1088 vgnd vpwr scs8hd_decap_3
XPHY_1077 vgnd vpwr scs8hd_decap_3
XPHY_1066 vgnd vpwr scs8hd_decap_3
XFILLER_355_27 vgnd vpwr scs8hd_decap_12
XFILLER_404_3 vgnd vpwr scs8hd_decap_12
XFILLER_98_44 vgnd vpwr scs8hd_decap_12
XFILLER_371_15 vgnd vpwr scs8hd_decap_12
XFILLER_371_59 vpwr vgnd scs8hd_fill_2
XFILLER_601_62 vgnd vpwr scs8hd_decap_12
XFILLER_601_51 vgnd vpwr scs8hd_decap_8
XFILLER_63_80 vgnd vpwr scs8hd_fill_1
XFILLER_249_39 vgnd vpwr scs8hd_decap_12
XFILLER_179_80 vgnd vpwr scs8hd_fill_1
XFILLER_396_56 vgnd vpwr scs8hd_decap_12
XPHY_990 vgnd vpwr scs8hd_decap_3
XFILLER_546_15 vgnd vpwr scs8hd_decap_12
XFILLER_265_27 vgnd vpwr scs8hd_decap_12
XFILLER_281_15 vgnd vpwr scs8hd_decap_12
XFILLER_281_59 vpwr vgnd scs8hd_fill_2
XFILLER_511_51 vgnd vpwr scs8hd_decap_8
XFILLER_511_62 vgnd vpwr scs8hd_decap_12
XFILLER_43_39 vgnd vpwr scs8hd_decap_12
XFILLER_159_39 vgnd vpwr scs8hd_decap_12
XFILLER_456_15 vgnd vpwr scs8hd_decap_12
XFILLER_175_27 vgnd vpwr scs8hd_decap_12
XFILLER_209_7 vgnd vpwr scs8hd_fill_1
XFILLER_108_32 vgnd vpwr scs8hd_decap_12
XFILLER_191_15 vgnd vpwr scs8hd_decap_12
XFILLER_552_80 vgnd vpwr scs8hd_fill_1
XFILLER_191_59 vpwr vgnd scs8hd_fill_2
XFILLER_405_74 vgnd vpwr scs8hd_decap_6
XFILLER_187_3 vgnd vpwr scs8hd_decap_12
XFILLER_84_68 vgnd vpwr scs8hd_decap_12
XFILLER_421_51 vgnd vpwr scs8hd_decap_8
XFILLER_421_62 vgnd vpwr scs8hd_decap_12
XFILLER_17_51 vgnd vpwr scs8hd_decap_8
XFILLER_17_62 vgnd vpwr scs8hd_decap_12
XFILLER_354_3 vgnd vpwr scs8hd_decap_12
XPHY_242 vgnd vpwr scs8hd_decap_3
XPHY_231 vgnd vpwr scs8hd_decap_3
XPHY_220 vgnd vpwr scs8hd_decap_3
XFILLER_521_3 vgnd vpwr scs8hd_decap_12
XPHY_264 vgnd vpwr scs8hd_decap_3
XPHY_253 vgnd vpwr scs8hd_decap_3
XPHY_275 vgnd vpwr scs8hd_decap_3
XPHY_286 vgnd vpwr scs8hd_decap_3
XPHY_297 vgnd vpwr scs8hd_decap_3
XFILLER_366_15 vgnd vpwr scs8hd_decap_12
XFILLER_165_71 vgnd vpwr scs8hd_decap_8
XFILLER_315_74 vgnd vpwr scs8hd_decap_6
XFILLER_462_80 vgnd vpwr scs8hd_fill_1
XFILLER_58_80 vgnd vpwr scs8hd_fill_1
XFILLER_331_51 vgnd vpwr scs8hd_decap_8
XFILLER_331_62 vgnd vpwr scs8hd_decap_12
XFILLER_200_44 vgnd vpwr scs8hd_decap_12
XFILLER_276_15 vgnd vpwr scs8hd_decap_12
XFILLER_209_31 vpwr vgnd scs8hd_fill_2
XFILLER_225_74 vgnd vpwr scs8hd_decap_6
XFILLER_372_80 vgnd vpwr scs8hd_fill_1
XFILLER_241_51 vgnd vpwr scs8hd_decap_8
XFILLER_241_62 vgnd vpwr scs8hd_decap_12
XFILLER_598_32 vgnd vpwr scs8hd_decap_12
XFILLER_54_27 vgnd vpwr scs8hd_decap_4
XFILLER_110_44 vgnd vpwr scs8hd_decap_12
XFILLER_70_15 vgnd vpwr scs8hd_decap_12
XFILLER_186_15 vgnd vpwr scs8hd_decap_12
XFILLER_547_80 vgnd vpwr scs8hd_fill_1
XFILLER_102_3 vgnd vpwr scs8hd_decap_12
XFILLER_135_74 vgnd vpwr scs8hd_decap_6
XFILLER_282_80 vgnd vpwr scs8hd_fill_1
XFILLER_569_3 vgnd vpwr scs8hd_decap_12
XFILLER_471_3 vgnd vpwr scs8hd_decap_12
XFILLER_151_51 vgnd vpwr scs8hd_decap_8
XFILLER_151_62 vgnd vpwr scs8hd_decap_12
XFILLER_527_39 vgnd vpwr scs8hd_decap_12
XFILLER_457_80 vgnd vpwr scs8hd_fill_1
XFILLER_543_27 vgnd vpwr scs8hd_decap_12
XFILLER_192_80 vgnd vpwr scs8hd_fill_1
XFILLER_568_68 vgnd vpwr scs8hd_decap_12
XFILLER_584_56 vgnd vpwr scs8hd_decap_12
XFILLER_367_80 vgnd vpwr scs8hd_fill_1
XFILLER_437_39 vgnd vpwr scs8hd_decap_12
XFILLER_49_27 vgnd vpwr scs8hd_decap_12
XFILLER_453_27 vgnd vpwr scs8hd_decap_12
XFILLER_65_15 vgnd vpwr scs8hd_decap_12
XFILLER_65_59 vpwr vgnd scs8hd_fill_2
XFILLER_478_68 vgnd vpwr scs8hd_decap_12
XFILLER_277_80 vgnd vpwr scs8hd_fill_1
XFILLER_317_3 vgnd vpwr scs8hd_decap_12
XFILLER_347_39 vgnd vpwr scs8hd_decap_12
XFILLER_494_56 vgnd vpwr scs8hd_decap_12
XFILLER_363_27 vgnd vpwr scs8hd_decap_12
XFILLER_388_68 vgnd vpwr scs8hd_decap_12
XFILLER_538_27 vgnd vpwr scs8hd_decap_4
XFILLER_71_80 vgnd vpwr scs8hd_fill_1
XFILLER_187_80 vgnd vpwr scs8hd_fill_1
XFILLER_257_39 vgnd vpwr scs8hd_decap_12
XFILLER_554_15 vgnd vpwr scs8hd_decap_12
XFILLER_65_3 vgnd vpwr scs8hd_decap_12
XFILLER_273_27 vgnd vpwr scs8hd_decap_12
XFILLER_206_32 vgnd vpwr scs8hd_decap_12
XFILLER_503_74 vgnd vpwr scs8hd_decap_6
XPHY_808 vgnd vpwr scs8hd_decap_3
XFILLER_298_68 vgnd vpwr scs8hd_decap_12
XPHY_819 vgnd vpwr scs8hd_decap_3
XPHY_1407 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1418 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1429 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_448_27 vgnd vpwr scs8hd_decap_4
XFILLER_51_39 vgnd vpwr scs8hd_decap_12
XFILLER_167_39 vgnd vpwr scs8hd_decap_12
XFILLER_464_15 vgnd vpwr scs8hd_decap_12
XFILLER_183_27 vgnd vpwr scs8hd_decap_8
XFILLER_116_32 vgnd vpwr scs8hd_decap_12
XFILLER_413_74 vgnd vpwr scs8hd_decap_6
XFILLER_560_80 vgnd vpwr scs8hd_fill_1
XFILLER_267_3 vgnd vpwr scs8hd_decap_12
XFILLER_92_68 vgnd vpwr scs8hd_decap_12
XPHY_40 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XFILLER_25_51 vgnd vpwr scs8hd_decap_8
XFILLER_25_62 vgnd vpwr scs8hd_decap_12
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_434_3 vgnd vpwr scs8hd_decap_12
XPHY_95 vgnd vpwr scs8hd_decap_3
XPHY_84 vgnd vpwr scs8hd_decap_3
XFILLER_358_27 vgnd vpwr scs8hd_decap_4
XFILLER_601_3 vgnd vpwr scs8hd_decap_12
XFILLER_374_15 vgnd vpwr scs8hd_decap_12
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XFILLER_66_80 vgnd vpwr scs8hd_fill_1
XFILLER_323_74 vgnd vpwr scs8hd_decap_6
XFILLER_470_80 vgnd vpwr scs8hd_fill_1
XFILLER_549_15 vgnd vpwr scs8hd_decap_12
XFILLER_549_59 vpwr vgnd scs8hd_fill_2
XFILLER_268_27 vgnd vpwr scs8hd_decap_4
XFILLER_284_15 vgnd vpwr scs8hd_decap_12
XFILLER_233_74 vgnd vpwr scs8hd_decap_6
XFILLER_380_80 vgnd vpwr scs8hd_fill_1
XFILLER_459_15 vgnd vpwr scs8hd_decap_12
XFILLER_102_56 vgnd vpwr scs8hd_decap_12
XFILLER_62_27 vgnd vpwr scs8hd_decap_4
XPHY_605 vgnd vpwr scs8hd_decap_3
XPHY_616 vgnd vpwr scs8hd_decap_3
XPHY_1204 vgnd vpwr scs8hd_decap_3
XFILLER_178_27 vgnd vpwr scs8hd_decap_4
XPHY_627 vgnd vpwr scs8hd_decap_3
XPHY_638 vgnd vpwr scs8hd_decap_3
XPHY_649 vgnd vpwr scs8hd_decap_3
XFILLER_459_59 vpwr vgnd scs8hd_fill_2
XPHY_1248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_555_80 vgnd vpwr scs8hd_fill_1
XFILLER_384_3 vgnd vpwr scs8hd_decap_12
XFILLER_143_74 vgnd vpwr scs8hd_decap_6
XFILLER_290_80 vgnd vpwr scs8hd_fill_1
XFILLER_551_3 vgnd vpwr scs8hd_decap_12
XFILLER_369_15 vgnd vpwr scs8hd_decap_12
XFILLER_369_59 vpwr vgnd scs8hd_fill_2
XPHY_1760 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1793 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1782 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1771 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_535_39 vgnd vpwr scs8hd_decap_12
XFILLER_465_80 vgnd vpwr scs8hd_fill_1
XFILLER_184_70 vgnd vpwr scs8hd_decap_8
XFILLER_551_27 vgnd vpwr scs8hd_decap_12
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
XFILLER_203_22 vpwr vgnd scs8hd_fill_2
XFILLER_279_15 vgnd vpwr scs8hd_decap_12
XFILLER_279_59 vpwr vgnd scs8hd_fill_2
XFILLER_576_68 vgnd vpwr scs8hd_decap_12
XFILLER_295_47 vgnd vpwr scs8hd_decap_12
XFILLER_509_51 vgnd vpwr scs8hd_decap_8
XFILLER_509_62 vgnd vpwr scs8hd_decap_12
XFILLER_592_56 vgnd vpwr scs8hd_decap_12
XFILLER_375_80 vgnd vpwr scs8hd_fill_1
XFILLER_445_39 vgnd vpwr scs8hd_decap_12
XFILLER_461_27 vgnd vpwr scs8hd_decap_12
XFILLER_57_27 vgnd vpwr scs8hd_decap_12
XFILLER_73_15 vgnd vpwr scs8hd_decap_12
XFILLER_73_59 vpwr vgnd scs8hd_fill_2
XFILLER_189_15 vpwr vgnd scs8hd_fill_2
XPHY_402 vgnd vpwr scs8hd_decap_3
XPHY_413 vgnd vpwr scs8hd_decap_3
XPHY_424 vgnd vpwr scs8hd_decap_3
XPHY_435 vgnd vpwr scs8hd_decap_3
XPHY_446 vgnd vpwr scs8hd_decap_3
XPHY_457 vgnd vpwr scs8hd_decap_3
XPHY_468 vgnd vpwr scs8hd_decap_3
XPHY_1001 vgnd vpwr scs8hd_decap_3
XPHY_1012 vgnd vpwr scs8hd_decap_3
XPHY_1023 vgnd vpwr scs8hd_decap_3
XPHY_1056 vgnd vpwr scs8hd_decap_3
XPHY_1045 vgnd vpwr scs8hd_decap_3
XFILLER_132_3 vgnd vpwr scs8hd_decap_12
XPHY_479 vgnd vpwr scs8hd_decap_3
XFILLER_486_68 vgnd vpwr scs8hd_decap_12
XPHY_1034 vgnd vpwr scs8hd_decap_3
XPHY_1089 vgnd vpwr scs8hd_decap_3
XPHY_1078 vgnd vpwr scs8hd_decap_3
XPHY_1067 vgnd vpwr scs8hd_decap_3
XFILLER_419_51 vgnd vpwr scs8hd_decap_8
XFILLER_419_62 vgnd vpwr scs8hd_decap_12
XFILLER_285_80 vgnd vpwr scs8hd_fill_1
XFILLER_355_39 vgnd vpwr scs8hd_decap_12
XFILLER_98_56 vgnd vpwr scs8hd_decap_12
XFILLER_599_3 vgnd vpwr scs8hd_decap_12
XFILLER_371_27 vgnd vpwr scs8hd_decap_12
XFILLER_304_32 vgnd vpwr scs8hd_decap_12
XFILLER_601_74 vgnd vpwr scs8hd_decap_6
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
XFILLER_396_68 vgnd vpwr scs8hd_decap_12
XPHY_980 vgnd vpwr scs8hd_decap_3
XFILLER_546_27 vgnd vpwr scs8hd_decap_4
XFILLER_329_51 vgnd vpwr scs8hd_decap_8
XFILLER_329_62 vgnd vpwr scs8hd_decap_12
XPHY_991 vgnd vpwr scs8hd_decap_3
XPHY_1590 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_195_80 vgnd vpwr scs8hd_fill_1
XFILLER_265_39 vgnd vpwr scs8hd_decap_12
XFILLER_562_15 vgnd vpwr scs8hd_decap_12
XFILLER_281_27 vgnd vpwr scs8hd_decap_12
XFILLER_214_32 vgnd vpwr scs8hd_decap_12
X_19_ gfpga_pad_GPIO_PAD[0] right_width_0_height_0__pin_1_ vgnd vpwr scs8hd_buf_2
XFILLER_511_74 vgnd vpwr scs8hd_decap_6
XFILLER_239_51 vgnd vpwr scs8hd_decap_8
XFILLER_239_62 vgnd vpwr scs8hd_decap_12
XFILLER_456_27 vgnd vpwr scs8hd_decap_4
XFILLER_175_39 vgnd vpwr scs8hd_decap_12
XFILLER_108_44 vgnd vpwr scs8hd_decap_12
XFILLER_472_15 vgnd vpwr scs8hd_decap_12
XFILLER_68_15 vgnd vpwr scs8hd_decap_12
XFILLER_191_27 vgnd vpwr scs8hd_decap_12
XFILLER_124_32 vgnd vpwr scs8hd_decap_12
XFILLER_17_74 vgnd vpwr scs8hd_decap_6
XFILLER_421_74 vgnd vpwr scs8hd_decap_6
XPHY_210 vgnd vpwr scs8hd_decap_3
XFILLER_347_3 vgnd vpwr scs8hd_decap_12
XPHY_243 vgnd vpwr scs8hd_decap_3
XPHY_232 vgnd vpwr scs8hd_decap_3
XPHY_221 vgnd vpwr scs8hd_decap_3
XPHY_254 vgnd vpwr scs8hd_decap_3
XFILLER_33_51 vgnd vpwr scs8hd_decap_8
XPHY_265 vgnd vpwr scs8hd_decap_3
XPHY_276 vgnd vpwr scs8hd_decap_3
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XPHY_287 vgnd vpwr scs8hd_decap_3
XPHY_298 vgnd vpwr scs8hd_decap_3
XFILLER_149_51 vgnd vpwr scs8hd_decap_8
XFILLER_149_62 vgnd vpwr scs8hd_decap_12
XFILLER_366_27 vgnd vpwr scs8hd_decap_4
XFILLER_514_3 vgnd vpwr scs8hd_decap_12
XFILLER_382_15 vgnd vpwr scs8hd_decap_12
XFILLER_331_74 vgnd vpwr scs8hd_decap_6
XFILLER_74_80 vgnd vpwr scs8hd_fill_1
XFILLER_95_3 vgnd vpwr scs8hd_decap_12
XFILLER_200_12 vgnd vpwr scs8hd_decap_12
XFILLER_557_15 vgnd vpwr scs8hd_decap_12
XFILLER_200_56 vgnd vpwr scs8hd_decap_12
XFILLER_557_59 vpwr vgnd scs8hd_fill_2
XFILLER_276_27 vgnd vpwr scs8hd_decap_4
XFILLER_292_15 vgnd vpwr scs8hd_decap_12
XFILLER_225_20 vgnd vpwr scs8hd_decap_12
XFILLER_598_44 vgnd vpwr scs8hd_decap_12
XFILLER_241_74 vgnd vpwr scs8hd_decap_6
XFILLER_110_56 vgnd vpwr scs8hd_decap_12
XFILLER_467_15 vgnd vpwr scs8hd_decap_12
XFILLER_70_27 vgnd vpwr scs8hd_decap_4
XFILLER_467_59 vpwr vgnd scs8hd_fill_2
XFILLER_186_27 vgnd vpwr scs8hd_decap_4
XFILLER_563_80 vgnd vpwr scs8hd_fill_1
XFILLER_297_3 vgnd vpwr scs8hd_decap_12
XFILLER_464_3 vgnd vpwr scs8hd_decap_12
XFILLER_151_74 vgnd vpwr scs8hd_decap_6
XFILLER_377_15 vgnd vpwr scs8hd_decap_12
XFILLER_377_59 vpwr vgnd scs8hd_fill_2
XFILLER_543_39 vgnd vpwr scs8hd_decap_12
XFILLER_473_80 vgnd vpwr scs8hd_fill_1
XFILLER_69_80 vgnd vpwr scs8hd_fill_1
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XFILLER_211_55 vgnd vpwr scs8hd_decap_6
XFILLER_287_15 vgnd vpwr scs8hd_decap_12
XFILLER_287_59 vpwr vgnd scs8hd_fill_2
XFILLER_584_68 vgnd vpwr scs8hd_decap_12
XFILLER_517_51 vgnd vpwr scs8hd_decap_8
XFILLER_517_62 vgnd vpwr scs8hd_decap_12
XFILLER_383_80 vgnd vpwr scs8hd_fill_1
XFILLER_453_39 vgnd vpwr scs8hd_decap_12
XFILLER_49_39 vgnd vpwr scs8hd_decap_12
XFILLER_65_27 vgnd vpwr scs8hd_decap_12
XFILLER_402_32 vgnd vpwr scs8hd_decap_12
XFILLER_81_15 vgnd vpwr scs8hd_decap_12
XFILLER_81_59 vpwr vgnd scs8hd_fill_2
XFILLER_197_15 vgnd vpwr scs8hd_decap_12
XFILLER_558_80 vgnd vpwr scs8hd_fill_1
XFILLER_197_59 vpwr vgnd scs8hd_fill_2
XFILLER_212_3 vgnd vpwr scs8hd_decap_6
XFILLER_494_68 vgnd vpwr scs8hd_decap_12
XFILLER_427_51 vgnd vpwr scs8hd_decap_8
XFILLER_427_62 vgnd vpwr scs8hd_decap_12
XFILLER_293_80 vgnd vpwr scs8hd_fill_1
XFILLER_363_39 vgnd vpwr scs8hd_decap_12
XFILLER_581_3 vgnd vpwr scs8hd_decap_12
XFILLER_312_32 vgnd vpwr scs8hd_decap_12
XFILLER_468_80 vgnd vpwr scs8hd_fill_1
XFILLER_337_51 vgnd vpwr scs8hd_decap_8
XFILLER_554_27 vgnd vpwr scs8hd_decap_4
XFILLER_58_3 vgnd vpwr scs8hd_decap_12
XFILLER_337_62 vgnd vpwr scs8hd_decap_12
XFILLER_273_39 vgnd vpwr scs8hd_decap_12
XFILLER_206_11 vpwr vgnd scs8hd_fill_2
XFILLER_206_22 vpwr vgnd scs8hd_fill_2
XFILLER_570_15 vgnd vpwr scs8hd_decap_12
XFILLER_206_44 vgnd vpwr scs8hd_decap_12
XFILLER_222_32 vgnd vpwr scs8hd_decap_12
XPHY_809 vgnd vpwr scs8hd_decap_3
XPHY_1408 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1419 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_378_80 vgnd vpwr scs8hd_fill_1
XFILLER_247_51 vgnd vpwr scs8hd_decap_8
XFILLER_247_62 vgnd vpwr scs8hd_decap_12
XFILLER_464_27 vgnd vpwr scs8hd_decap_4
XFILLER_116_44 vgnd vpwr scs8hd_decap_12
XFILLER_76_15 vgnd vpwr scs8hd_decap_12
XFILLER_480_15 vgnd vpwr scs8hd_decap_12
XFILLER_132_32 vgnd vpwr scs8hd_decap_12
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_162_3 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_25_74 vgnd vpwr scs8hd_decap_6
XFILLER_288_80 vgnd vpwr scs8hd_fill_1
XFILLER_427_3 vgnd vpwr scs8hd_decap_12
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
XFILLER_157_51 vgnd vpwr scs8hd_decap_8
XFILLER_157_62 vgnd vpwr scs8hd_decap_12
XFILLER_374_27 vgnd vpwr scs8hd_decap_4
XFILLER_390_15 vgnd vpwr scs8hd_decap_12
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XFILLER_549_27 vgnd vpwr scs8hd_decap_12
XFILLER_82_80 vgnd vpwr scs8hd_fill_1
XFILLER_198_80 vgnd vpwr scs8hd_fill_1
XFILLER_565_15 vgnd vpwr scs8hd_decap_12
XFILLER_565_59 vpwr vgnd scs8hd_fill_2
XFILLER_284_27 vgnd vpwr scs8hd_decap_4
XFILLER_102_68 vgnd vpwr scs8hd_decap_12
XPHY_606 vgnd vpwr scs8hd_decap_3
XPHY_617 vgnd vpwr scs8hd_decap_3
XFILLER_459_27 vgnd vpwr scs8hd_decap_12
XPHY_1205 vgnd vpwr scs8hd_decap_3
XPHY_628 vgnd vpwr scs8hd_decap_3
XPHY_639 vgnd vpwr scs8hd_decap_3
XPHY_1216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_475_15 vgnd vpwr scs8hd_decap_12
XFILLER_475_59 vpwr vgnd scs8hd_fill_2
XFILLER_194_16 vpwr vgnd scs8hd_fill_2
XFILLER_571_80 vgnd vpwr scs8hd_fill_1
XFILLER_377_3 vgnd vpwr scs8hd_decap_12
XFILLER_544_3 vgnd vpwr scs8hd_decap_12
XFILLER_369_27 vgnd vpwr scs8hd_decap_12
XPHY_1761 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1750 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_385_15 vgnd vpwr scs8hd_decap_12
XPHY_1794 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1783 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1772 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_385_59 vpwr vgnd scs8hd_fill_2
XFILLER_551_39 vgnd vpwr scs8hd_decap_12
XFILLER_77_80 vgnd vpwr scs8hd_fill_1
XFILLER_481_80 vgnd vpwr scs8hd_fill_1
XFILLER_203_34 vgnd vpwr scs8hd_decap_12
XFILLER_279_27 vgnd vpwr scs8hd_decap_12
XFILLER_500_32 vgnd vpwr scs8hd_decap_12
XFILLER_295_59 vpwr vgnd scs8hd_fill_2
XFILLER_509_74 vgnd vpwr scs8hd_decap_6
XFILLER_592_68 vgnd vpwr scs8hd_decap_12
XFILLER_525_51 vgnd vpwr scs8hd_decap_8
XFILLER_525_62 vgnd vpwr scs8hd_decap_12
XFILLER_461_39 vgnd vpwr scs8hd_decap_12
XFILLER_57_39 vgnd vpwr scs8hd_decap_12
XFILLER_391_80 vgnd vpwr scs8hd_fill_1
XFILLER_73_27 vgnd vpwr scs8hd_decap_12
XFILLER_410_32 vgnd vpwr scs8hd_decap_12
XPHY_403 vgnd vpwr scs8hd_decap_3
XPHY_414 vgnd vpwr scs8hd_decap_3
XPHY_425 vgnd vpwr scs8hd_decap_3
XPHY_436 vgnd vpwr scs8hd_decap_3
XPHY_447 vgnd vpwr scs8hd_decap_3
XPHY_458 vgnd vpwr scs8hd_decap_3
XPHY_1002 vgnd vpwr scs8hd_decap_3
XPHY_1013 vgnd vpwr scs8hd_decap_3
XPHY_1046 vgnd vpwr scs8hd_decap_3
XPHY_469 vgnd vpwr scs8hd_decap_3
XPHY_1024 vgnd vpwr scs8hd_decap_3
XPHY_1035 vgnd vpwr scs8hd_decap_3
XPHY_1079 vgnd vpwr scs8hd_decap_3
XPHY_1068 vgnd vpwr scs8hd_decap_3
XPHY_1057 vgnd vpwr scs8hd_decap_3
XFILLER_566_80 vgnd vpwr scs8hd_fill_1
XFILLER_125_3 vgnd vpwr scs8hd_decap_12
XFILLER_419_74 vgnd vpwr scs8hd_decap_6
XFILLER_98_68 vgnd vpwr scs8hd_decap_12
XFILLER_435_51 vgnd vpwr scs8hd_decap_8
XFILLER_435_62 vgnd vpwr scs8hd_decap_12
XFILLER_494_3 vgnd vpwr scs8hd_decap_12
XFILLER_371_39 vgnd vpwr scs8hd_decap_12
XFILLER_304_44 vgnd vpwr scs8hd_decap_12
XFILLER_320_32 vgnd vpwr scs8hd_decap_12
XPHY_970 vgnd vpwr scs8hd_decap_3
XPHY_981 vgnd vpwr scs8hd_decap_3
XFILLER_8_44 vgnd vpwr scs8hd_decap_12
XPHY_992 vgnd vpwr scs8hd_decap_3
XFILLER_329_74 vgnd vpwr scs8hd_decap_6
XPHY_1580 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1591 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_476_80 vgnd vpwr scs8hd_fill_1
XFILLER_562_27 vgnd vpwr scs8hd_decap_4
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XFILLER_345_51 vgnd vpwr scs8hd_decap_8
XFILLER_345_62 vgnd vpwr scs8hd_decap_12
XFILLER_281_39 vgnd vpwr scs8hd_decap_12
XFILLER_214_44 vgnd vpwr scs8hd_decap_12
X_18_ gfpga_pad_GPIO_PAD[7] right_width_0_height_0__pin_15_ vgnd vpwr scs8hd_buf_2
XFILLER_230_32 vgnd vpwr scs8hd_decap_12
XFILLER_239_74 vgnd vpwr scs8hd_decap_6
XFILLER_386_80 vgnd vpwr scs8hd_fill_1
XFILLER_108_56 vgnd vpwr scs8hd_decap_12
XFILLER_255_51 vgnd vpwr scs8hd_decap_8
XFILLER_255_62 vgnd vpwr scs8hd_decap_12
XFILLER_472_27 vgnd vpwr scs8hd_decap_4
XFILLER_68_27 vgnd vpwr scs8hd_decap_4
XFILLER_191_39 vgnd vpwr scs8hd_decap_12
XFILLER_124_44 vgnd vpwr scs8hd_decap_12
XFILLER_84_15 vgnd vpwr scs8hd_decap_12
XFILLER_140_32 vgnd vpwr scs8hd_decap_12
XPHY_200 vgnd vpwr scs8hd_decap_3
XPHY_233 vgnd vpwr scs8hd_decap_3
XPHY_222 vgnd vpwr scs8hd_decap_3
XPHY_211 vgnd vpwr scs8hd_decap_3
XFILLER_242_3 vgnd vpwr scs8hd_decap_12
XPHY_266 vgnd vpwr scs8hd_decap_3
XPHY_255 vgnd vpwr scs8hd_decap_3
XPHY_244 vgnd vpwr scs8hd_decap_3
XPHY_277 vgnd vpwr scs8hd_decap_3
XFILLER_33_74 vgnd vpwr scs8hd_decap_6
XPHY_288 vgnd vpwr scs8hd_decap_3
XPHY_299 vgnd vpwr scs8hd_decap_3
XFILLER_149_74 vgnd vpwr scs8hd_decap_6
XFILLER_296_80 vgnd vpwr scs8hd_fill_1
XFILLER_507_3 vgnd vpwr scs8hd_decap_12
XFILLER_165_51 vgnd vpwr scs8hd_decap_8
XFILLER_165_62 vgnd vpwr scs8hd_decap_6
XFILLER_382_27 vgnd vpwr scs8hd_decap_4
XFILLER_181_72 vgnd vpwr scs8hd_decap_8
XFILLER_200_24 vgnd vpwr scs8hd_decap_6
XFILLER_557_27 vgnd vpwr scs8hd_decap_12
XFILLER_200_68 vgnd vpwr scs8hd_decap_12
XFILLER_90_80 vgnd vpwr scs8hd_fill_1
XFILLER_88_3 vgnd vpwr scs8hd_decap_12
XFILLER_573_15 vgnd vpwr scs8hd_decap_12
XFILLER_573_59 vpwr vgnd scs8hd_fill_2
XFILLER_292_27 vgnd vpwr scs8hd_decap_4
XFILLER_225_32 vgnd vpwr scs8hd_decap_12
XFILLER_598_56 vgnd vpwr scs8hd_decap_12
XFILLER_110_68 vgnd vpwr scs8hd_decap_12
XFILLER_467_27 vgnd vpwr scs8hd_decap_12
XFILLER_483_15 vgnd vpwr scs8hd_decap_12
XFILLER_79_15 vgnd vpwr scs8hd_decap_12
XFILLER_79_59 vpwr vgnd scs8hd_fill_2
XFILLER_483_59 vpwr vgnd scs8hd_fill_2
XFILLER_192_3 vgnd vpwr scs8hd_decap_12
XFILLER_457_3 vgnd vpwr scs8hd_decap_12
XFILLER_377_27 vgnd vpwr scs8hd_decap_12
XFILLER_393_15 vgnd vpwr scs8hd_decap_12
XFILLER_393_59 vpwr vgnd scs8hd_fill_2
XFILLER_85_80 vgnd vpwr scs8hd_fill_1
XFILLER_211_23 vpwr vgnd scs8hd_fill_2
XFILLER_568_15 vgnd vpwr scs8hd_decap_12
XFILLER_287_27 vgnd vpwr scs8hd_decap_12
XFILLER_517_74 vgnd vpwr scs8hd_decap_6
XFILLER_533_62 vgnd vpwr scs8hd_decap_12
XFILLER_533_51 vgnd vpwr scs8hd_decap_8
XFILLER_65_39 vgnd vpwr scs8hd_decap_12
XFILLER_402_44 vgnd vpwr scs8hd_decap_12
XFILLER_81_27 vgnd vpwr scs8hd_decap_12
XFILLER_478_15 vgnd vpwr scs8hd_decap_12
XFILLER_197_27 vgnd vpwr scs8hd_decap_12
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
XFILLER_574_80 vgnd vpwr scs8hd_fill_1
XFILLER_427_74 vgnd vpwr scs8hd_decap_6
XFILLER_39_51 vgnd vpwr scs8hd_decap_8
XFILLER_443_51 vgnd vpwr scs8hd_decap_8
XFILLER_443_62 vgnd vpwr scs8hd_decap_12
XFILLER_574_3 vgnd vpwr scs8hd_decap_12
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XFILLER_312_44 vgnd vpwr scs8hd_decap_12
XFILLER_388_15 vgnd vpwr scs8hd_decap_12
XFILLER_337_74 vgnd vpwr scs8hd_decap_6
XFILLER_484_80 vgnd vpwr scs8hd_fill_1
XFILLER_570_27 vgnd vpwr scs8hd_decap_4
XFILLER_206_56 vgnd vpwr scs8hd_decap_12
XFILLER_353_51 vgnd vpwr scs8hd_decap_8
XFILLER_353_62 vgnd vpwr scs8hd_decap_12
XFILLER_222_44 vgnd vpwr scs8hd_decap_12
XFILLER_298_15 vgnd vpwr scs8hd_decap_12
XPHY_1409 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_247_74 vgnd vpwr scs8hd_decap_6
XFILLER_394_80 vgnd vpwr scs8hd_fill_1
XFILLER_116_56 vgnd vpwr scs8hd_decap_12
XFILLER_263_51 vgnd vpwr scs8hd_decap_8
XFILLER_263_62 vgnd vpwr scs8hd_decap_12
XFILLER_480_27 vgnd vpwr scs8hd_decap_4
XFILLER_76_27 vgnd vpwr scs8hd_decap_4
XFILLER_132_44 vgnd vpwr scs8hd_decap_12
XFILLER_92_15 vgnd vpwr scs8hd_decap_12
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_569_80 vgnd vpwr scs8hd_fill_1
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_64 vgnd vpwr scs8hd_decap_3
XFILLER_155_3 vgnd vpwr scs8hd_decap_12
XPHY_97 vgnd vpwr scs8hd_decap_3
XPHY_86 vgnd vpwr scs8hd_decap_3
XPHY_75 vgnd vpwr scs8hd_decap_3
XFILLER_322_3 vgnd vpwr scs8hd_decap_12
XFILLER_41_74 vgnd vpwr scs8hd_decap_6
XFILLER_157_74 vgnd vpwr scs8hd_decap_6
XFILLER_173_51 vgnd vpwr scs8hd_decap_8
XFILLER_173_62 vgnd vpwr scs8hd_decap_12
XFILLER_390_27 vgnd vpwr scs8hd_decap_4
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XFILLER_549_39 vgnd vpwr scs8hd_decap_12
XFILLER_479_80 vgnd vpwr scs8hd_fill_1
XFILLER_565_27 vgnd vpwr scs8hd_decap_12
XFILLER_70_3 vgnd vpwr scs8hd_decap_12
XFILLER_217_22 vpwr vgnd scs8hd_fill_2
XFILLER_581_15 vgnd vpwr scs8hd_decap_12
XFILLER_581_59 vpwr vgnd scs8hd_fill_2
XPHY_607 vgnd vpwr scs8hd_decap_3
XFILLER_459_39 vgnd vpwr scs8hd_decap_12
XPHY_618 vgnd vpwr scs8hd_decap_3
XPHY_629 vgnd vpwr scs8hd_decap_3
XFILLER_389_80 vgnd vpwr scs8hd_fill_1
XPHY_1206 vgnd vpwr scs8hd_decap_3
XPHY_1217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_475_27 vgnd vpwr scs8hd_decap_12
XFILLER_194_28 vgnd vpwr scs8hd_decap_3
XFILLER_408_32 vgnd vpwr scs8hd_decap_12
XFILLER_87_15 vgnd vpwr scs8hd_decap_12
XFILLER_491_15 vgnd vpwr scs8hd_decap_12
XFILLER_87_59 vpwr vgnd scs8hd_fill_2
XFILLER_491_59 vpwr vgnd scs8hd_fill_2
XFILLER_272_3 vgnd vpwr scs8hd_decap_12
XFILLER_537_3 vgnd vpwr scs8hd_decap_12
XFILLER_369_39 vgnd vpwr scs8hd_decap_12
XFILLER_299_80 vgnd vpwr scs8hd_fill_1
XPHY_1751 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1740 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1795 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1784 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1773 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1762 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_385_27 vgnd vpwr scs8hd_decap_12
XFILLER_318_32 vgnd vpwr scs8hd_decap_12
XFILLER_203_46 vgnd vpwr scs8hd_decap_12
XFILLER_93_80 vgnd vpwr scs8hd_fill_1
XFILLER_500_44 vgnd vpwr scs8hd_decap_12
XFILLER_279_39 vgnd vpwr scs8hd_decap_12
XFILLER_576_15 vgnd vpwr scs8hd_decap_12
XFILLER_228_32 vgnd vpwr scs8hd_decap_12
XFILLER_525_74 vgnd vpwr scs8hd_decap_6
XFILLER_541_62 vgnd vpwr scs8hd_decap_12
XFILLER_541_51 vgnd vpwr scs8hd_decap_8
XFILLER_73_39 vgnd vpwr scs8hd_decap_12
XFILLER_189_28 vgnd vpwr scs8hd_decap_12
XFILLER_410_44 vgnd vpwr scs8hd_decap_12
XPHY_404 vgnd vpwr scs8hd_decap_3
XPHY_415 vgnd vpwr scs8hd_decap_3
XPHY_426 vgnd vpwr scs8hd_decap_3
XPHY_437 vgnd vpwr scs8hd_decap_3
XPHY_448 vgnd vpwr scs8hd_decap_3
XPHY_459 vgnd vpwr scs8hd_decap_3
XFILLER_486_15 vgnd vpwr scs8hd_decap_12
XPHY_1003 vgnd vpwr scs8hd_decap_3
XPHY_1014 vgnd vpwr scs8hd_decap_3
XPHY_1047 vgnd vpwr scs8hd_decap_3
XPHY_1025 vgnd vpwr scs8hd_decap_3
XPHY_1036 vgnd vpwr scs8hd_decap_3
XPHY_1069 vgnd vpwr scs8hd_decap_3
XPHY_1058 vgnd vpwr scs8hd_decap_3
XFILLER_22_32 vgnd vpwr scs8hd_decap_12
XFILLER_138_32 vgnd vpwr scs8hd_decap_12
XFILLER_118_3 vgnd vpwr scs8hd_decap_12
XFILLER_582_80 vgnd vpwr scs8hd_fill_1
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XFILLER_435_74 vgnd vpwr scs8hd_decap_6
XFILLER_487_3 vgnd vpwr scs8hd_decap_12
XFILLER_304_56 vgnd vpwr scs8hd_decap_12
XFILLER_451_51 vgnd vpwr scs8hd_decap_8
XFILLER_451_62 vgnd vpwr scs8hd_decap_12
XFILLER_47_62 vgnd vpwr scs8hd_decap_12
XFILLER_47_51 vgnd vpwr scs8hd_decap_8
XFILLER_320_44 vgnd vpwr scs8hd_decap_12
XFILLER_396_15 vgnd vpwr scs8hd_decap_12
XPHY_960 vgnd vpwr scs8hd_decap_3
XPHY_971 vgnd vpwr scs8hd_decap_3
XFILLER_8_56 vgnd vpwr scs8hd_decap_12
XPHY_982 vgnd vpwr scs8hd_decap_3
XPHY_993 vgnd vpwr scs8hd_decap_3
XPHY_1570 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1581 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1592 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_345_74 vgnd vpwr scs8hd_decap_6
XFILLER_492_80 vgnd vpwr scs8hd_fill_1
XFILLER_88_80 vgnd vpwr scs8hd_fill_1
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
XFILLER_214_56 vgnd vpwr scs8hd_decap_12
XFILLER_361_51 vgnd vpwr scs8hd_decap_8
XFILLER_361_62 vgnd vpwr scs8hd_decap_12
X_17_ gfpga_pad_GPIO_PAD[6] right_width_0_height_0__pin_13_ vgnd vpwr scs8hd_buf_2
XFILLER_230_44 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_108_68 vgnd vpwr scs8hd_decap_12
XFILLER_255_74 vgnd vpwr scs8hd_decap_6
XFILLER_124_56 vgnd vpwr scs8hd_decap_12
XFILLER_271_51 vgnd vpwr scs8hd_decap_8
XFILLER_84_27 vgnd vpwr scs8hd_decap_4
XFILLER_271_62 vgnd vpwr scs8hd_decap_12
XPHY_201 vgnd vpwr scs8hd_decap_3
XFILLER_140_44 vgnd vpwr scs8hd_decap_12
XPHY_234 vgnd vpwr scs8hd_decap_3
XPHY_223 vgnd vpwr scs8hd_decap_3
XPHY_212 vgnd vpwr scs8hd_decap_3
XPHY_256 vgnd vpwr scs8hd_decap_3
XPHY_245 vgnd vpwr scs8hd_decap_3
XPHY_267 vgnd vpwr scs8hd_decap_3
XFILLER_235_3 vgnd vpwr scs8hd_decap_12
XFILLER_577_80 vgnd vpwr scs8hd_fill_1
XPHY_278 vgnd vpwr scs8hd_decap_3
XPHY_289 vgnd vpwr scs8hd_decap_3
XFILLER_402_3 vgnd vpwr scs8hd_decap_12
XFILLER_181_51 vgnd vpwr scs8hd_decap_8
XFILLER_181_62 vpwr vgnd scs8hd_fill_2
XFILLER_557_39 vgnd vpwr scs8hd_decap_12
XPHY_790 vgnd vpwr scs8hd_decap_3
XFILLER_487_80 vgnd vpwr scs8hd_fill_1
XFILLER_573_27 vgnd vpwr scs8hd_decap_12
XFILLER_506_32 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _09_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_225_11 vgnd vpwr scs8hd_decap_3
XFILLER_225_44 vgnd vpwr scs8hd_decap_12
XFILLER_598_68 vgnd vpwr scs8hd_decap_12
XFILLER_397_80 vgnd vpwr scs8hd_fill_1
XFILLER_467_39 vgnd vpwr scs8hd_decap_12
XFILLER_79_27 vgnd vpwr scs8hd_decap_12
XFILLER_483_27 vgnd vpwr scs8hd_decap_12
XFILLER_416_32 vgnd vpwr scs8hd_decap_12
XFILLER_95_15 vgnd vpwr scs8hd_decap_12
XFILLER_95_59 vpwr vgnd scs8hd_fill_2
XFILLER_185_3 vgnd vpwr scs8hd_decap_12
XFILLER_352_3 vgnd vpwr scs8hd_decap_12
XFILLER_377_39 vgnd vpwr scs8hd_decap_12
XFILLER_100_80 vgnd vpwr scs8hd_fill_1
XFILLER_393_27 vgnd vpwr scs8hd_decap_12
XFILLER_326_32 vgnd vpwr scs8hd_decap_12
XFILLER_568_27 vgnd vpwr scs8hd_decap_4
XFILLER_211_46 vgnd vpwr scs8hd_decap_3
XFILLER_287_39 vgnd vpwr scs8hd_decap_12
XFILLER_584_15 vgnd vpwr scs8hd_decap_12
XFILLER_236_32 vgnd vpwr scs8hd_decap_12
XFILLER_533_74 vgnd vpwr scs8hd_decap_6
XFILLER_402_56 vgnd vpwr scs8hd_decap_12
XFILLER_478_27 vgnd vpwr scs8hd_decap_4
XFILLER_81_39 vgnd vpwr scs8hd_decap_12
XFILLER_14_44 vgnd vpwr scs8hd_decap_12
XFILLER_197_39 vgnd vpwr scs8hd_decap_12
XFILLER_494_15 vgnd vpwr scs8hd_decap_12
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XFILLER_146_32 vgnd vpwr scs8hd_decap_12
XFILLER_100_3 vgnd vpwr scs8hd_decap_12
XFILLER_590_80 vgnd vpwr scs8hd_fill_1
XFILLER_39_74 vgnd vpwr scs8hd_decap_6
XFILLER_443_74 vgnd vpwr scs8hd_decap_6
XFILLER_567_3 vgnd vpwr scs8hd_decap_12
XFILLER_55_62 vgnd vpwr scs8hd_decap_12
XFILLER_55_51 vgnd vpwr scs8hd_decap_8
XFILLER_312_56 vgnd vpwr scs8hd_decap_12
XFILLER_388_27 vgnd vpwr scs8hd_decap_4
Xlogical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ right_width_0_height_0__pin_2_ logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[1] vgnd vpwr scs8hd_ebufn_1
XFILLER_96_80 vgnd vpwr scs8hd_fill_1
XFILLER_206_68 vgnd vpwr scs8hd_decap_12
XFILLER_353_74 vgnd vpwr scs8hd_decap_6
XFILLER_579_15 vgnd vpwr scs8hd_decap_12
XFILLER_222_56 vgnd vpwr scs8hd_decap_12
XFILLER_579_59 vpwr vgnd scs8hd_fill_2
XFILLER_298_27 vgnd vpwr scs8hd_decap_4
XFILLER_116_68 vgnd vpwr scs8hd_decap_12
XFILLER_263_74 vgnd vpwr scs8hd_decap_6
XFILLER_92_27 vgnd vpwr scs8hd_decap_4
XFILLER_132_56 vgnd vpwr scs8hd_decap_12
XFILLER_489_15 vgnd vpwr scs8hd_decap_12
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XFILLER_489_59 vpwr vgnd scs8hd_fill_2
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_decap_3
XPHY_76 vgnd vpwr scs8hd_decap_3
XFILLER_148_3 vgnd vpwr scs8hd_decap_12
XFILLER_585_80 vgnd vpwr scs8hd_fill_1
XFILLER_315_3 vgnd vpwr scs8hd_decap_12
XFILLER_173_74 vgnd vpwr scs8hd_decap_6
XFILLER_399_15 vgnd vpwr scs8hd_decap_12
XFILLER_399_59 vpwr vgnd scs8hd_fill_2
XFILLER_565_39 vgnd vpwr scs8hd_decap_12
XFILLER_495_80 vgnd vpwr scs8hd_fill_1
XFILLER_63_3 vgnd vpwr scs8hd_decap_12
XFILLER_581_27 vgnd vpwr scs8hd_decap_12
XFILLER_514_32 vgnd vpwr scs8hd_decap_12
XFILLER_102_15 vgnd vpwr scs8hd_decap_12
XPHY_608 vgnd vpwr scs8hd_decap_3
XPHY_619 vgnd vpwr scs8hd_decap_3
XPHY_1207 vgnd vpwr scs8hd_decap_3
XFILLER_539_62 vgnd vpwr scs8hd_decap_12
XFILLER_539_51 vgnd vpwr scs8hd_decap_8
XPHY_1218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_475_39 vgnd vpwr scs8hd_decap_12
XFILLER_408_44 vgnd vpwr scs8hd_decap_12
XFILLER_491_27 vgnd vpwr scs8hd_decap_12
XFILLER_87_27 vgnd vpwr scs8hd_decap_12
XFILLER_424_32 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _14_/Y vgnd vpwr scs8hd_diode_2
XFILLER_265_3 vgnd vpwr scs8hd_decap_12
XFILLER_432_3 vgnd vpwr scs8hd_decap_12
XFILLER_449_51 vgnd vpwr scs8hd_decap_8
XFILLER_449_62 vgnd vpwr scs8hd_decap_12
XPHY_1752 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1741 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1730 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1785 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1774 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1763 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_385_39 vgnd vpwr scs8hd_decap_12
XPHY_1796 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_318_44 vgnd vpwr scs8hd_decap_12
XFILLER_334_32 vgnd vpwr scs8hd_decap_12
XFILLER_203_14 vpwr vgnd scs8hd_fill_2
XFILLER_203_58 vgnd vpwr scs8hd_decap_3
XFILLER_500_56 vgnd vpwr scs8hd_decap_12
XFILLER_576_27 vgnd vpwr scs8hd_decap_4
XFILLER_359_51 vgnd vpwr scs8hd_decap_8
XFILLER_359_62 vgnd vpwr scs8hd_decap_12
XFILLER_592_15 vgnd vpwr scs8hd_decap_12
XFILLER_228_44 vgnd vpwr scs8hd_decap_12
XFILLER_244_32 vgnd vpwr scs8hd_decap_12
XFILLER_541_74 vgnd vpwr scs8hd_decap_6
XPHY_405 vgnd vpwr scs8hd_decap_3
XPHY_416 vgnd vpwr scs8hd_decap_3
XFILLER_410_56 vgnd vpwr scs8hd_decap_12
XPHY_427 vgnd vpwr scs8hd_decap_3
XPHY_438 vgnd vpwr scs8hd_decap_3
XPHY_449 vgnd vpwr scs8hd_decap_3
XFILLER_269_51 vgnd vpwr scs8hd_decap_8
XFILLER_486_27 vgnd vpwr scs8hd_decap_4
XPHY_1004 vgnd vpwr scs8hd_decap_3
XFILLER_269_62 vgnd vpwr scs8hd_decap_12
XPHY_1015 vgnd vpwr scs8hd_decap_3
XPHY_1026 vgnd vpwr scs8hd_decap_3
XPHY_1037 vgnd vpwr scs8hd_decap_3
XPHY_1059 vgnd vpwr scs8hd_decap_3
XPHY_1048 vgnd vpwr scs8hd_decap_3
XFILLER_22_44 vgnd vpwr scs8hd_decap_12
XFILLER_98_15 vgnd vpwr scs8hd_decap_12
XFILLER_138_44 vgnd vpwr scs8hd_decap_12
XFILLER_154_32 vgnd vpwr scs8hd_decap_12
XFILLER_382_3 vgnd vpwr scs8hd_decap_12
XFILLER_304_68 vgnd vpwr scs8hd_decap_12
XFILLER_451_74 vgnd vpwr scs8hd_decap_6
XFILLER_47_74 vgnd vpwr scs8hd_decap_6
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ right_width_0_height_0__pin_12_ vgnd vpwr scs8hd_diode_2
XFILLER_103_80 vgnd vpwr scs8hd_fill_1
XFILLER_63_51 vgnd vpwr scs8hd_decap_8
XFILLER_320_56 vgnd vpwr scs8hd_decap_12
XFILLER_63_62 vgnd vpwr scs8hd_decap_12
XFILLER_179_51 vgnd vpwr scs8hd_decap_8
XFILLER_396_27 vgnd vpwr scs8hd_decap_4
XFILLER_179_62 vgnd vpwr scs8hd_decap_12
XPHY_950 vgnd vpwr scs8hd_decap_3
XPHY_961 vgnd vpwr scs8hd_decap_3
XPHY_972 vgnd vpwr scs8hd_decap_3
XPHY_1560 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_983 vgnd vpwr scs8hd_decap_3
XPHY_994 vgnd vpwr scs8hd_decap_3
XFILLER_8_68 vgnd vpwr scs8hd_decap_12
XPHY_1571 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1582 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1593 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XFILLER_214_68 vgnd vpwr scs8hd_decap_12
XFILLER_361_74 vgnd vpwr scs8hd_decap_6
X_16_ gfpga_pad_GPIO_PAD[5] right_width_0_height_0__pin_11_ vgnd vpwr scs8hd_buf_2
XFILLER_587_15 vgnd vpwr scs8hd_decap_12
XFILLER_230_56 vgnd vpwr scs8hd_decap_12
XFILLER_587_59 vpwr vgnd scs8hd_fill_2
XFILLER_124_68 vgnd vpwr scs8hd_decap_12
XFILLER_271_74 vgnd vpwr scs8hd_decap_6
XFILLER_140_56 vgnd vpwr scs8hd_decap_12
XFILLER_497_15 vgnd vpwr scs8hd_decap_12
XPHY_224 vgnd vpwr scs8hd_decap_3
XPHY_213 vgnd vpwr scs8hd_decap_3
XPHY_202 vgnd vpwr scs8hd_decap_3
XFILLER_497_59 vpwr vgnd scs8hd_fill_2
XPHY_257 vgnd vpwr scs8hd_decap_3
XPHY_246 vgnd vpwr scs8hd_decap_3
XPHY_235 vgnd vpwr scs8hd_decap_3
XPHY_268 vgnd vpwr scs8hd_decap_3
XFILLER_130_3 vgnd vpwr scs8hd_decap_12
XPHY_279 vgnd vpwr scs8hd_decap_3
XFILLER_228_3 vgnd vpwr scs8hd_decap_12
XFILLER_593_80 vgnd vpwr scs8hd_fill_1
XFILLER_597_3 vgnd vpwr scs8hd_decap_12
XPHY_780 vgnd vpwr scs8hd_decap_3
XPHY_791 vgnd vpwr scs8hd_decap_3
XPHY_1390 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_573_39 vgnd vpwr scs8hd_decap_12
XFILLER_209_46 vgnd vpwr scs8hd_decap_12
XFILLER_99_80 vgnd vpwr scs8hd_fill_1
XFILLER_506_44 vgnd vpwr scs8hd_decap_12
XFILLER_225_56 vgnd vpwr scs8hd_decap_4
XFILLER_522_32 vgnd vpwr scs8hd_decap_12
XFILLER_110_15 vgnd vpwr scs8hd_decap_12
XFILLER_547_51 vgnd vpwr scs8hd_decap_8
XFILLER_547_62 vgnd vpwr scs8hd_decap_12
XFILLER_483_39 vgnd vpwr scs8hd_decap_12
XFILLER_79_39 vgnd vpwr scs8hd_decap_12
XFILLER_416_44 vgnd vpwr scs8hd_decap_12
XFILLER_95_27 vgnd vpwr scs8hd_decap_12
XFILLER_28_32 vgnd vpwr scs8hd_decap_12
XFILLER_432_32 vgnd vpwr scs8hd_decap_12
XFILLER_178_3 vgnd vpwr scs8hd_decap_12
XFILLER_345_3 vgnd vpwr scs8hd_decap_12
XFILLER_588_80 vgnd vpwr scs8hd_fill_1
XFILLER_457_51 vgnd vpwr scs8hd_decap_8
XFILLER_512_3 vgnd vpwr scs8hd_decap_12
XFILLER_457_62 vgnd vpwr scs8hd_decap_12
XFILLER_393_39 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_326_44 vgnd vpwr scs8hd_decap_12
XFILLER_342_32 vgnd vpwr scs8hd_decap_12
XFILLER_498_80 vgnd vpwr scs8hd_fill_1
XFILLER_93_3 vgnd vpwr scs8hd_decap_12
XFILLER_367_51 vpwr vgnd scs8hd_fill_2
XFILLER_584_27 vgnd vpwr scs8hd_decap_4
XFILLER_367_62 vgnd vpwr scs8hd_decap_12
XFILLER_236_44 vgnd vpwr scs8hd_decap_12
XFILLER_105_15 vgnd vpwr scs8hd_decap_12
XFILLER_252_32 vgnd vpwr scs8hd_decap_12
XFILLER_105_59 vpwr vgnd scs8hd_fill_2
XFILLER_402_68 vgnd vpwr scs8hd_decap_12
XFILLER_201_80 vgnd vpwr scs8hd_fill_1
XFILLER_14_56 vgnd vpwr scs8hd_decap_12
XFILLER_277_51 vgnd vpwr scs8hd_decap_8
XFILLER_277_62 vgnd vpwr scs8hd_decap_12
XFILLER_494_27 vgnd vpwr scs8hd_decap_4
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XFILLER_146_44 vgnd vpwr scs8hd_decap_12
XFILLER_162_32 vgnd vpwr scs8hd_decap_12
XFILLER_462_3 vgnd vpwr scs8hd_decap_12
XFILLER_312_68 vgnd vpwr scs8hd_decap_12
XFILLER_55_74 vgnd vpwr scs8hd_decap_6
XFILLER_111_80 vgnd vpwr scs8hd_fill_1
XFILLER_71_62 vgnd vpwr scs8hd_decap_12
XFILLER_71_51 vgnd vpwr scs8hd_decap_8
XFILLER_187_51 vgnd vpwr scs8hd_decap_8
XFILLER_187_62 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _15_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_579_27 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ right_width_0_height_0__pin_8_ vgnd vpwr scs8hd_diode_2
XFILLER_222_68 vgnd vpwr scs8hd_decap_12
XFILLER_595_15 vgnd vpwr scs8hd_decap_12
XFILLER_595_59 vpwr vgnd scs8hd_fill_2
XFILLER_132_68 vgnd vpwr scs8hd_decap_12
XFILLER_489_27 vgnd vpwr scs8hd_decap_12
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_decap_3
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_decap_3
XFILLER_210_3 vgnd vpwr scs8hd_decap_3
XFILLER_308_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_106_80 vgnd vpwr scs8hd_fill_1
XFILLER_399_27 vgnd vpwr scs8hd_decap_12
XFILLER_56_3 vgnd vpwr scs8hd_decap_12
XFILLER_581_39 vgnd vpwr scs8hd_decap_12
XFILLER_514_44 vgnd vpwr scs8hd_decap_12
XFILLER_530_32 vgnd vpwr scs8hd_decap_12
XFILLER_102_27 vgnd vpwr scs8hd_decap_4
XPHY_609 vgnd vpwr scs8hd_decap_3
XPHY_1208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_539_74 vgnd vpwr scs8hd_decap_6
XFILLER_555_62 vgnd vpwr scs8hd_decap_12
XFILLER_555_51 vgnd vpwr scs8hd_decap_8
XFILLER_408_56 vgnd vpwr scs8hd_decap_12
XFILLER_87_39 vgnd vpwr scs8hd_decap_12
XFILLER_491_39 vgnd vpwr scs8hd_decap_12
XFILLER_424_44 vgnd vpwr scs8hd_decap_12
XFILLER_440_32 vgnd vpwr scs8hd_decap_12
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XFILLER_160_3 vgnd vpwr scs8hd_decap_12
XFILLER_258_3 vgnd vpwr scs8hd_decap_12
XFILLER_596_80 vgnd vpwr scs8hd_fill_1
XPHY_1742 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1731 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_425_3 vgnd vpwr scs8hd_decap_12
XFILLER_449_74 vgnd vpwr scs8hd_decap_6
XPHY_1720 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1786 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1775 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1764 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1753 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1797 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_318_56 vgnd vpwr scs8hd_decap_12
XFILLER_465_51 vgnd vpwr scs8hd_decap_8
XFILLER_465_62 vgnd vpwr scs8hd_decap_12
XFILLER_184_30 vgnd vpwr scs8hd_fill_1
XFILLER_334_44 vgnd vpwr scs8hd_decap_12
XFILLER_203_26 vpwr vgnd scs8hd_fill_2
XFILLER_350_32 vgnd vpwr scs8hd_decap_12
XFILLER_500_68 vgnd vpwr scs8hd_decap_12
XFILLER_359_74 vgnd vpwr scs8hd_decap_6
XFILLER_592_27 vgnd vpwr scs8hd_decap_4
XFILLER_228_56 vgnd vpwr scs8hd_decap_12
XFILLER_375_51 vgnd vpwr scs8hd_decap_8
XFILLER_375_62 vgnd vpwr scs8hd_decap_12
XFILLER_244_44 vgnd vpwr scs8hd_decap_12
XFILLER_3_80 vgnd vpwr scs8hd_fill_1
XFILLER_113_15 vgnd vpwr scs8hd_decap_12
XFILLER_260_32 vgnd vpwr scs8hd_decap_12
XFILLER_113_59 vpwr vgnd scs8hd_fill_2
XPHY_406 vgnd vpwr scs8hd_decap_3
XPHY_417 vgnd vpwr scs8hd_decap_3
XFILLER_410_68 vgnd vpwr scs8hd_decap_12
XPHY_428 vgnd vpwr scs8hd_decap_3
XPHY_439 vgnd vpwr scs8hd_decap_3
XPHY_1005 vgnd vpwr scs8hd_decap_3
XFILLER_269_74 vgnd vpwr scs8hd_decap_6
XPHY_1016 vgnd vpwr scs8hd_decap_3
XPHY_1027 vgnd vpwr scs8hd_decap_3
XPHY_1038 vgnd vpwr scs8hd_decap_3
XPHY_1049 vgnd vpwr scs8hd_decap_3
XFILLER_22_56 vgnd vpwr scs8hd_decap_12
XFILLER_138_56 vgnd vpwr scs8hd_decap_12
XFILLER_285_51 vgnd vpwr scs8hd_decap_8
XFILLER_285_62 vgnd vpwr scs8hd_decap_12
XFILLER_98_27 vgnd vpwr scs8hd_decap_4
XANTENNA__11__A enable vgnd vpwr scs8hd_diode_2
XFILLER_154_44 vgnd vpwr scs8hd_decap_12
XFILLER_170_32 vgnd vpwr scs8hd_decap_12
XFILLER_375_3 vgnd vpwr scs8hd_decap_12
XFILLER_542_3 vgnd vpwr scs8hd_decap_12
XFILLER_320_68 vgnd vpwr scs8hd_decap_12
XFILLER_63_74 vgnd vpwr scs8hd_decap_6
XFILLER_179_74 vgnd vpwr scs8hd_decap_6
XPHY_940 vgnd vpwr scs8hd_decap_3
XPHY_951 vgnd vpwr scs8hd_decap_3
XPHY_962 vgnd vpwr scs8hd_decap_3
XPHY_1550 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_973 vgnd vpwr scs8hd_decap_3
XPHY_984 vgnd vpwr scs8hd_decap_3
XPHY_995 vgnd vpwr scs8hd_decap_3
XPHY_1561 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1572 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1583 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1594 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_195_62 vgnd vpwr scs8hd_decap_12
XFILLER_19_3 vgnd vpwr scs8hd_decap_12
X_15_ address[1] _14_/B _07_/A address[2] _15_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_587_27 vgnd vpwr scs8hd_decap_12
XFILLER_230_68 vgnd vpwr scs8hd_fill_1
XFILLER_108_15 vgnd vpwr scs8hd_decap_12
XFILLER_204_80 vgnd vpwr scs8hd_fill_1
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ right_width_0_height_0__pin_4_ vgnd vpwr scs8hd_diode_2
XFILLER_497_27 vgnd vpwr scs8hd_decap_12
XPHY_225 vgnd vpwr scs8hd_decap_3
XPHY_214 vgnd vpwr scs8hd_decap_3
XPHY_203 vgnd vpwr scs8hd_decap_3
XFILLER_140_68 vgnd vpwr scs8hd_decap_12
XPHY_258 vgnd vpwr scs8hd_decap_3
XPHY_247 vgnd vpwr scs8hd_decap_3
XPHY_236 vgnd vpwr scs8hd_decap_3
XANTENNA__06__A address[1] vgnd vpwr scs8hd_diode_2
XPHY_269 vgnd vpwr scs8hd_decap_3
XFILLER_123_3 vgnd vpwr scs8hd_decap_12
XFILLER_492_3 vgnd vpwr scs8hd_decap_12
XFILLER_114_80 vgnd vpwr scs8hd_fill_1
XPHY_770 vgnd vpwr scs8hd_decap_3
XPHY_781 vgnd vpwr scs8hd_decap_3
XPHY_792 vgnd vpwr scs8hd_decap_3
XPHY_1380 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1391 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_209_58 vgnd vpwr scs8hd_decap_3
XFILLER_506_56 vgnd vpwr scs8hd_decap_12
XFILLER_522_44 vgnd vpwr scs8hd_decap_12
XFILLER_598_15 vgnd vpwr scs8hd_decap_12
XFILLER_110_27 vgnd vpwr scs8hd_decap_4
XFILLER_547_74 vgnd vpwr scs8hd_decap_6
XFILLER_563_62 vgnd vpwr scs8hd_decap_12
XFILLER_563_51 vgnd vpwr scs8hd_decap_8
XFILLER_416_56 vgnd vpwr scs8hd_decap_12
XFILLER_95_39 vgnd vpwr scs8hd_decap_12
XFILLER_432_44 vgnd vpwr scs8hd_decap_12
XFILLER_28_44 vgnd vpwr scs8hd_decap_12
XFILLER_301_15 vgnd vpwr scs8hd_decap_12
XFILLER_44_32 vgnd vpwr scs8hd_decap_12
XFILLER_301_59 vpwr vgnd scs8hd_fill_2
XFILLER_240_3 vgnd vpwr scs8hd_decap_12
XFILLER_338_3 vgnd vpwr scs8hd_decap_12
XFILLER_457_74 vgnd vpwr scs8hd_decap_6
XFILLER_505_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_109_80 vgnd vpwr scs8hd_fill_1
XFILLER_5_59 vpwr vgnd scs8hd_fill_2
XFILLER_326_56 vgnd vpwr scs8hd_decap_12
XFILLER_473_51 vgnd vpwr scs8hd_decap_8
XFILLER_473_62 vgnd vpwr scs8hd_decap_12
XFILLER_69_62 vgnd vpwr scs8hd_decap_12
XFILLER_69_51 vgnd vpwr scs8hd_decap_8
XFILLER_342_44 vgnd vpwr scs8hd_decap_12
XFILLER_86_3 vgnd vpwr scs8hd_decap_12
XFILLER_367_74 vgnd vpwr scs8hd_decap_6
XFILLER_236_56 vgnd vpwr scs8hd_decap_12
XFILLER_383_51 vgnd vpwr scs8hd_decap_8
XFILLER_383_62 vgnd vpwr scs8hd_decap_12
XFILLER_105_27 vgnd vpwr scs8hd_decap_12
XFILLER_252_44 vgnd vpwr scs8hd_decap_12
XFILLER_121_15 vgnd vpwr scs8hd_decap_12
XFILLER_121_59 vpwr vgnd scs8hd_fill_2
XFILLER_14_68 vgnd vpwr scs8hd_decap_12
XFILLER_277_74 vgnd vpwr scs8hd_decap_6
XFILLER_30_56 vgnd vpwr scs8hd_decap_12
XFILLER_146_56 vgnd vpwr scs8hd_decap_12
XFILLER_293_51 vgnd vpwr scs8hd_decap_8
XFILLER_293_62 vgnd vpwr scs8hd_decap_12
XFILLER_162_44 vgnd vpwr scs8hd_decap_12
XFILLER_190_3 vgnd vpwr scs8hd_decap_12
XFILLER_288_3 vgnd vpwr scs8hd_decap_12
XFILLER_455_3 vgnd vpwr scs8hd_decap_12
XFILLER_599_80 vgnd vpwr scs8hd_fill_1
XFILLER_71_74 vgnd vpwr scs8hd_decap_6
XFILLER_187_74 vgnd vpwr scs8hd_decap_6
XFILLER_206_26 vgnd vpwr scs8hd_decap_4
XFILLER_579_39 vgnd vpwr scs8hd_decap_12
XFILLER_302_80 vgnd vpwr scs8hd_fill_1
XFILLER_595_27 vgnd vpwr scs8hd_decap_12
XFILLER_528_32 vgnd vpwr scs8hd_decap_12
XFILLER_116_15 vgnd vpwr scs8hd_decap_12
XFILLER_6_80 vgnd vpwr scs8hd_fill_1
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_489_39 vgnd vpwr scs8hd_decap_12
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_decap_3
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XANTENNA__14__A _07_/C vgnd vpwr scs8hd_diode_2
XFILLER_438_32 vgnd vpwr scs8hd_decap_12
XFILLER_572_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_399_39 vgnd vpwr scs8hd_decap_12
XFILLER_122_80 vgnd vpwr scs8hd_fill_1
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ right_width_0_height_0__pin_0_ vgnd vpwr scs8hd_diode_2
XFILLER_348_32 vgnd vpwr scs8hd_decap_12
XFILLER_217_58 vgnd vpwr scs8hd_decap_3
XFILLER_49_3 vgnd vpwr scs8hd_decap_12
XFILLER_514_56 vgnd vpwr scs8hd_decap_12
XFILLER_530_44 vgnd vpwr scs8hd_decap_12
XPHY_1209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_258_32 vgnd vpwr scs8hd_decap_12
XFILLER_555_74 vgnd vpwr scs8hd_decap_6
XFILLER_408_68 vgnd vpwr scs8hd_decap_12
XFILLER_571_62 vgnd vpwr scs8hd_decap_12
XFILLER_571_51 vgnd vpwr scs8hd_decap_8
XFILLER_207_80 vgnd vpwr scs8hd_fill_1
XFILLER_424_56 vgnd vpwr scs8hd_decap_12
XANTENNA__09__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
XFILLER_440_44 vgnd vpwr scs8hd_decap_12
XFILLER_153_3 vgnd vpwr scs8hd_decap_12
XFILLER_52_32 vgnd vpwr scs8hd_decap_12
XPHY_1743 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1732 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_168_32 vgnd vpwr scs8hd_decap_12
XFILLER_320_3 vgnd vpwr scs8hd_decap_12
XPHY_1710 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1721 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1776 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1765 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1754 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_418_3 vgnd vpwr scs8hd_decap_12
XPHY_1798 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1787 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_318_68 vgnd vpwr scs8hd_decap_12
XFILLER_465_74 vgnd vpwr scs8hd_decap_6
XFILLER_117_80 vgnd vpwr scs8hd_fill_1
XFILLER_334_56 vgnd vpwr scs8hd_decap_12
XFILLER_481_51 vgnd vpwr scs8hd_decap_8
XFILLER_77_62 vgnd vpwr scs8hd_decap_12
XFILLER_77_51 vgnd vpwr scs8hd_decap_8
XFILLER_481_62 vgnd vpwr scs8hd_decap_12
XFILLER_350_44 vgnd vpwr scs8hd_decap_12
XFILLER_228_68 vgnd vpwr scs8hd_decap_12
XFILLER_375_74 vgnd vpwr scs8hd_decap_6
XFILLER_391_51 vgnd vpwr scs8hd_decap_8
XFILLER_244_56 vgnd vpwr scs8hd_decap_12
XFILLER_391_62 vgnd vpwr scs8hd_decap_12
XFILLER_113_27 vgnd vpwr scs8hd_decap_12
XFILLER_260_44 vgnd vpwr scs8hd_decap_12
XPHY_407 vgnd vpwr scs8hd_decap_3
XPHY_418 vgnd vpwr scs8hd_decap_3
XPHY_429 vgnd vpwr scs8hd_decap_3
XPHY_1006 vgnd vpwr scs8hd_decap_3
XPHY_1017 vgnd vpwr scs8hd_decap_3
XPHY_1028 vgnd vpwr scs8hd_decap_3
XPHY_1039 vgnd vpwr scs8hd_decap_3
XFILLER_22_68 vgnd vpwr scs8hd_decap_12
XFILLER_138_68 vgnd vpwr scs8hd_decap_12
XFILLER_285_74 vgnd vpwr scs8hd_decap_6
XFILLER_154_56 vgnd vpwr scs8hd_decap_12
XFILLER_304_15 vgnd vpwr scs8hd_decap_12
XFILLER_170_44 vgnd vpwr scs8hd_decap_12
XFILLER_270_3 vgnd vpwr scs8hd_decap_12
XFILLER_368_3 vgnd vpwr scs8hd_decap_12
XFILLER_535_3 vgnd vpwr scs8hd_decap_12
XPHY_930 vgnd vpwr scs8hd_decap_3
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
XFILLER_400_80 vgnd vpwr scs8hd_fill_1
XPHY_941 vgnd vpwr scs8hd_decap_3
XPHY_952 vgnd vpwr scs8hd_decap_3
XPHY_963 vgnd vpwr scs8hd_decap_3
XPHY_1540 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1551 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_974 vgnd vpwr scs8hd_decap_3
XPHY_985 vgnd vpwr scs8hd_decap_3
XPHY_996 vgnd vpwr scs8hd_decap_3
XPHY_1562 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1573 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1584 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1595 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_195_74 vgnd vpwr scs8hd_decap_6
XFILLER_214_15 vgnd vpwr scs8hd_decap_12
X_14_ _07_/C _14_/B _07_/A address[2] _14_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_587_39 vgnd vpwr scs8hd_decap_12
XFILLER_310_80 vgnd vpwr scs8hd_fill_1
XFILLER_536_32 vgnd vpwr scs8hd_decap_12
XFILLER_108_27 vgnd vpwr scs8hd_decap_4
XFILLER_124_15 vgnd vpwr scs8hd_decap_12
XPHY_215 vgnd vpwr scs8hd_decap_3
XPHY_204 vgnd vpwr scs8hd_decap_3
XFILLER_497_39 vgnd vpwr scs8hd_decap_12
XPHY_259 vgnd vpwr scs8hd_decap_3
XPHY_248 vgnd vpwr scs8hd_decap_3
XPHY_237 vgnd vpwr scs8hd_decap_3
XPHY_226 vgnd vpwr scs8hd_decap_3
XFILLER_220_80 vgnd vpwr scs8hd_fill_1
XANTENNA__22__A gfpga_pad_GPIO_PAD[3] vgnd vpwr scs8hd_diode_2
XFILLER_446_32 vgnd vpwr scs8hd_decap_12
XFILLER_116_3 vgnd vpwr scs8hd_decap_12
XFILLER_485_3 vgnd vpwr scs8hd_decap_12
XFILLER_130_80 vgnd vpwr scs8hd_fill_1
XPHY_760 vgnd vpwr scs8hd_decap_3
XPHY_771 vgnd vpwr scs8hd_decap_3
XPHY_782 vgnd vpwr scs8hd_decap_3
XPHY_793 vgnd vpwr scs8hd_decap_3
XPHY_1370 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1381 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1392 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_356_32 vgnd vpwr scs8hd_decap_12
XFILLER_506_68 vgnd vpwr scs8hd_decap_12
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XFILLER_305_80 vgnd vpwr scs8hd_fill_1
XFILLER_522_56 vgnd vpwr scs8hd_decap_12
XFILLER_598_27 vgnd vpwr scs8hd_decap_4
XFILLER_0_71 vgnd vpwr scs8hd_decap_8
XFILLER_9_80 vgnd vpwr scs8hd_fill_1
XFILLER_119_15 vgnd vpwr scs8hd_decap_12
XFILLER_266_32 vgnd vpwr scs8hd_decap_12
XFILLER_119_59 vpwr vgnd scs8hd_fill_2
XFILLER_563_74 vgnd vpwr scs8hd_decap_6
XFILLER_416_68 vgnd vpwr scs8hd_decap_12
XFILLER_215_80 vgnd vpwr scs8hd_fill_1
XFILLER_28_56 vgnd vpwr scs8hd_decap_12
XFILLER_432_56 vgnd vpwr scs8hd_decap_12
XANTENNA__17__A gfpga_pad_GPIO_PAD[6] vgnd vpwr scs8hd_diode_2
XFILLER_301_27 vgnd vpwr scs8hd_decap_12
XFILLER_44_44 vgnd vpwr scs8hd_decap_12
XFILLER_233_3 vgnd vpwr scs8hd_decap_12
XFILLER_60_32 vgnd vpwr scs8hd_decap_12
XFILLER_176_32 vgnd vpwr scs8hd_decap_12
XFILLER_400_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XFILLER_69_74 vgnd vpwr scs8hd_decap_6
XFILLER_326_68 vgnd vpwr scs8hd_decap_12
XFILLER_473_74 vgnd vpwr scs8hd_decap_6
XFILLER_125_80 vgnd vpwr scs8hd_fill_1
XFILLER_85_62 vgnd vpwr scs8hd_decap_12
XFILLER_85_51 vgnd vpwr scs8hd_decap_8
XFILLER_342_56 vgnd vpwr scs8hd_decap_12
XFILLER_211_38 vgnd vpwr scs8hd_decap_8
XFILLER_79_3 vgnd vpwr scs8hd_decap_12
XPHY_590 vgnd vpwr scs8hd_decap_3
XFILLER_236_68 vgnd vpwr scs8hd_decap_12
XFILLER_383_74 vgnd vpwr scs8hd_decap_6
XFILLER_105_39 vgnd vpwr scs8hd_decap_12
XFILLER_252_56 vgnd vpwr scs8hd_decap_12
XFILLER_402_15 vgnd vpwr scs8hd_decap_12
XFILLER_121_27 vgnd vpwr scs8hd_decap_12
XFILLER_30_68 vgnd vpwr scs8hd_decap_12
XFILLER_146_68 vgnd vpwr scs8hd_decap_12
XFILLER_293_74 vgnd vpwr scs8hd_decap_6
XFILLER_162_56 vgnd vpwr scs8hd_decap_12
XFILLER_183_3 vgnd vpwr scs8hd_decap_12
XFILLER_312_15 vgnd vpwr scs8hd_decap_12
XFILLER_350_3 vgnd vpwr scs8hd_decap_12
XFILLER_448_3 vgnd vpwr scs8hd_decap_12
XFILLER_222_15 vgnd vpwr scs8hd_decap_12
XFILLER_595_39 vgnd vpwr scs8hd_decap_12
XFILLER_528_44 vgnd vpwr scs8hd_decap_12
XFILLER_544_32 vgnd vpwr scs8hd_decap_12
XFILLER_116_27 vgnd vpwr scs8hd_decap_4
XFILLER_132_15 vgnd vpwr scs8hd_decap_12
XPHY_13 vgnd vpwr scs8hd_decap_3
XFILLER_569_62 vgnd vpwr scs8hd_decap_12
XFILLER_569_51 vgnd vpwr scs8hd_decap_8
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XANTENNA__14__B _14_/B vgnd vpwr scs8hd_diode_2
XFILLER_438_44 vgnd vpwr scs8hd_decap_12
XFILLER_307_15 vgnd vpwr scs8hd_decap_12
XFILLER_307_59 vpwr vgnd scs8hd_fill_2
XFILLER_454_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XFILLER_398_3 vgnd vpwr scs8hd_decap_12
XFILLER_565_3 vgnd vpwr scs8hd_decap_12
XFILLER_403_80 vgnd vpwr scs8hd_fill_1
XFILLER_479_51 vgnd vpwr scs8hd_decap_8
XFILLER_479_62 vgnd vpwr scs8hd_decap_12
XFILLER_348_44 vgnd vpwr scs8hd_decap_12
XFILLER_217_26 vpwr vgnd scs8hd_fill_2
XFILLER_364_32 vgnd vpwr scs8hd_decap_12
XFILLER_514_68 vgnd vpwr scs8hd_decap_12
XFILLER_530_56 vgnd vpwr scs8hd_decap_12
XFILLER_313_80 vgnd vpwr scs8hd_fill_1
XFILLER_389_51 vgnd vpwr scs8hd_decap_8
XFILLER_389_62 vgnd vpwr scs8hd_decap_12
XFILLER_258_44 vgnd vpwr scs8hd_decap_12
XFILLER_11_15 vgnd vpwr scs8hd_decap_12
XFILLER_127_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_59 vpwr vgnd scs8hd_fill_2
XFILLER_274_32 vgnd vpwr scs8hd_decap_12
XFILLER_127_59 vpwr vgnd scs8hd_fill_2
XFILLER_571_74 vgnd vpwr scs8hd_decap_6
XFILLER_424_68 vgnd vpwr scs8hd_decap_12
XANTENNA__09__B enable vgnd vpwr scs8hd_diode_2
XFILLER_223_80 vgnd vpwr scs8hd_fill_1
XFILLER_440_56 vgnd vpwr scs8hd_decap_12
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XFILLER_299_51 vgnd vpwr scs8hd_decap_8
XFILLER_299_62 vgnd vpwr scs8hd_decap_12
XPHY_1700 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1733 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_52_44 vgnd vpwr scs8hd_decap_12
XFILLER_146_3 vgnd vpwr scs8hd_decap_12
XPHY_1711 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1722 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1766 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1755 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1744 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_168_44 vgnd vpwr scs8hd_decap_12
XPHY_1799 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1788 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1777 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_313_3 vgnd vpwr scs8hd_decap_12
XFILLER_184_32 vgnd vpwr scs8hd_decap_3
XFILLER_334_68 vgnd vpwr scs8hd_decap_12
XFILLER_481_74 vgnd vpwr scs8hd_decap_6
XFILLER_77_74 vgnd vpwr scs8hd_decap_6
XFILLER_93_51 vgnd vpwr scs8hd_decap_8
XFILLER_133_80 vgnd vpwr scs8hd_fill_1
XFILLER_350_56 vgnd vpwr scs8hd_decap_12
XFILLER_93_62 vgnd vpwr scs8hd_decap_12
XFILLER_500_15 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_3 vgnd vpwr scs8hd_decap_12
XFILLER_308_80 vgnd vpwr scs8hd_fill_1
XFILLER_244_68 vgnd vpwr scs8hd_decap_12
XFILLER_391_74 vgnd vpwr scs8hd_decap_6
XFILLER_113_39 vgnd vpwr scs8hd_decap_12
XFILLER_260_56 vgnd vpwr scs8hd_decap_12
XFILLER_410_15 vgnd vpwr scs8hd_decap_12
XPHY_408 vgnd vpwr scs8hd_decap_3
XPHY_419 vgnd vpwr scs8hd_decap_3
XPHY_1007 vgnd vpwr scs8hd_decap_3
XPHY_1018 vgnd vpwr scs8hd_decap_3
XPHY_1029 vgnd vpwr scs8hd_decap_3
XFILLER_218_80 vgnd vpwr scs8hd_fill_1
XFILLER_154_68 vgnd vpwr scs8hd_decap_12
XFILLER_304_27 vgnd vpwr scs8hd_decap_4
XFILLER_170_56 vgnd vpwr scs8hd_decap_12
XFILLER_263_3 vgnd vpwr scs8hd_decap_12
XFILLER_320_15 vgnd vpwr scs8hd_decap_12
XFILLER_430_3 vgnd vpwr scs8hd_decap_12
XPHY_920 vgnd vpwr scs8hd_decap_3
XFILLER_528_3 vgnd vpwr scs8hd_decap_12
XPHY_931 vgnd vpwr scs8hd_decap_3
XPHY_942 vgnd vpwr scs8hd_decap_3
XPHY_953 vgnd vpwr scs8hd_decap_3
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
XPHY_1530 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1541 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_964 vgnd vpwr scs8hd_decap_3
XPHY_975 vgnd vpwr scs8hd_decap_3
XPHY_986 vgnd vpwr scs8hd_decap_3
XPHY_997 vgnd vpwr scs8hd_decap_3
XPHY_1552 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1563 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1574 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1585 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_195_31 vgnd vpwr scs8hd_decap_12
XPHY_1596 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_80 vgnd vpwr scs8hd_fill_1
XFILLER_128_80 vgnd vpwr scs8hd_fill_1
XFILLER_214_27 vgnd vpwr scs8hd_decap_4
X_13_ address[1] _14_/B _07_/A _08_/Y _13_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_230_15 vgnd vpwr scs8hd_decap_12
XFILLER_536_44 vgnd vpwr scs8hd_decap_12
XFILLER_405_15 vgnd vpwr scs8hd_decap_12
XFILLER_552_32 vgnd vpwr scs8hd_decap_12
XFILLER_124_27 vgnd vpwr scs8hd_decap_4
XFILLER_405_59 vpwr vgnd scs8hd_fill_2
XFILLER_140_15 vgnd vpwr scs8hd_decap_12
XPHY_216 vgnd vpwr scs8hd_decap_3
XPHY_205 vgnd vpwr scs8hd_decap_3
XFILLER_501_80 vgnd vpwr scs8hd_fill_1
XPHY_249 vgnd vpwr scs8hd_decap_3
XPHY_238 vgnd vpwr scs8hd_decap_3
XPHY_227 vgnd vpwr scs8hd_decap_3
XFILLER_577_62 vgnd vpwr scs8hd_decap_12
XFILLER_446_44 vgnd vpwr scs8hd_decap_12
XFILLER_109_3 vgnd vpwr scs8hd_decap_12
XFILLER_315_15 vgnd vpwr scs8hd_decap_12
XFILLER_462_32 vgnd vpwr scs8hd_decap_12
XFILLER_58_32 vgnd vpwr scs8hd_decap_12
XFILLER_315_59 vpwr vgnd scs8hd_fill_2
XFILLER_380_3 vgnd vpwr scs8hd_decap_12
XFILLER_478_3 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _09_/X vgnd vpwr scs8hd_diode_2
XFILLER_411_80 vgnd vpwr scs8hd_fill_1
XFILLER_487_51 vgnd vpwr scs8hd_decap_8
XPHY_750 vgnd vpwr scs8hd_decap_3
XPHY_761 vgnd vpwr scs8hd_decap_3
XPHY_772 vgnd vpwr scs8hd_decap_3
XFILLER_487_62 vgnd vpwr scs8hd_decap_12
XPHY_1360 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_783 vgnd vpwr scs8hd_decap_3
XPHY_794 vgnd vpwr scs8hd_decap_3
XPHY_1371 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1382 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1393 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_209_27 vpwr vgnd scs8hd_fill_2
XFILLER_356_44 vgnd vpwr scs8hd_decap_12
XFILLER_372_32 vgnd vpwr scs8hd_decap_12
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
XFILLER_522_68 vgnd vpwr scs8hd_decap_12
XFILLER_321_80 vgnd vpwr scs8hd_fill_1
XFILLER_397_51 vgnd vpwr scs8hd_decap_8
XFILLER_397_62 vgnd vpwr scs8hd_decap_12
XFILLER_119_27 vgnd vpwr scs8hd_decap_12
XFILLER_266_44 vgnd vpwr scs8hd_decap_12
XFILLER_135_15 vgnd vpwr scs8hd_decap_12
XFILLER_282_32 vgnd vpwr scs8hd_decap_12
XFILLER_135_59 vpwr vgnd scs8hd_fill_2
XFILLER_432_68 vgnd vpwr scs8hd_decap_12
XFILLER_28_68 vgnd vpwr scs8hd_decap_12
XFILLER_301_39 vgnd vpwr scs8hd_decap_12
XFILLER_44_56 vgnd vpwr scs8hd_decap_12
XFILLER_60_44 vgnd vpwr scs8hd_decap_12
XFILLER_226_3 vgnd vpwr scs8hd_decap_8
XFILLER_176_44 vgnd vpwr scs8hd_decap_12
XFILLER_5_39 vgnd vpwr scs8hd_decap_12
XFILLER_595_3 vgnd vpwr scs8hd_decap_12
XFILLER_192_32 vgnd vpwr scs8hd_decap_12
XFILLER_406_80 vgnd vpwr scs8hd_fill_1
XFILLER_342_68 vgnd vpwr scs8hd_decap_12
XFILLER_85_74 vgnd vpwr scs8hd_decap_6
XFILLER_141_80 vgnd vpwr scs8hd_fill_1
XPHY_580 vgnd vpwr scs8hd_decap_3
XPHY_591 vgnd vpwr scs8hd_decap_3
XPHY_1190 vgnd vpwr scs8hd_decap_3
XFILLER_316_80 vgnd vpwr scs8hd_fill_1
XFILLER_252_68 vgnd vpwr scs8hd_decap_12
XFILLER_402_27 vgnd vpwr scs8hd_decap_4
XFILLER_121_39 vgnd vpwr scs8hd_decap_12
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
XFILLER_212_9 vgnd vpwr scs8hd_fill_1
XFILLER_226_80 vgnd vpwr scs8hd_fill_1
XFILLER_162_68 vgnd vpwr scs8hd_decap_12
XFILLER_312_27 vgnd vpwr scs8hd_decap_4
XFILLER_176_3 vgnd vpwr scs8hd_decap_12
XFILLER_343_3 vgnd vpwr scs8hd_decap_12
XFILLER_510_3 vgnd vpwr scs8hd_decap_12
XFILLER_20_80 vgnd vpwr scs8hd_fill_1
XFILLER_136_80 vgnd vpwr scs8hd_fill_1
XFILLER_503_15 vgnd vpwr scs8hd_decap_12
XFILLER_222_27 vgnd vpwr scs8hd_decap_4
XFILLER_503_59 vpwr vgnd scs8hd_fill_2
XFILLER_91_3 vgnd vpwr scs8hd_decap_12
XFILLER_528_56 vgnd vpwr scs8hd_decap_12
XFILLER_544_44 vgnd vpwr scs8hd_decap_12
XFILLER_560_32 vgnd vpwr scs8hd_decap_12
XFILLER_413_15 vgnd vpwr scs8hd_decap_12
XFILLER_132_27 vgnd vpwr scs8hd_decap_4
XFILLER_413_59 vpwr vgnd scs8hd_fill_2
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XFILLER_569_74 vgnd vpwr scs8hd_decap_6
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XANTENNA__14__C _07_/A vgnd vpwr scs8hd_diode_2
XFILLER_585_62 vgnd vpwr scs8hd_decap_12
XFILLER_585_51 vgnd vpwr scs8hd_decap_8
XFILLER_438_56 vgnd vpwr scs8hd_decap_12
XFILLER_307_27 vgnd vpwr scs8hd_decap_12
XFILLER_454_44 vgnd vpwr scs8hd_decap_12
XFILLER_293_3 vgnd vpwr scs8hd_decap_12
XFILLER_323_15 vgnd vpwr scs8hd_decap_12
XFILLER_470_32 vgnd vpwr scs8hd_decap_12
XFILLER_66_32 vgnd vpwr scs8hd_decap_12
XFILLER_323_59 vpwr vgnd scs8hd_fill_2
XFILLER_558_3 vgnd vpwr scs8hd_decap_12
XFILLER_460_3 vgnd vpwr scs8hd_decap_12
XFILLER_479_74 vgnd vpwr scs8hd_decap_6
XFILLER_15_80 vgnd vpwr scs8hd_fill_1
XFILLER_348_56 vgnd vpwr scs8hd_decap_12
XFILLER_495_51 vgnd vpwr scs8hd_decap_8
XFILLER_495_62 vgnd vpwr scs8hd_decap_12
XFILLER_217_38 vgnd vpwr scs8hd_decap_12
XFILLER_364_44 vgnd vpwr scs8hd_decap_12
XFILLER_233_15 vgnd vpwr scs8hd_decap_12
XFILLER_380_32 vgnd vpwr scs8hd_decap_12
XFILLER_233_59 vpwr vgnd scs8hd_fill_2
XFILLER_530_68 vgnd vpwr scs8hd_decap_12
XFILLER_389_74 vgnd vpwr scs8hd_decap_6
XFILLER_258_56 vgnd vpwr scs8hd_decap_12
XFILLER_408_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_27 vgnd vpwr scs8hd_decap_12
XFILLER_127_27 vgnd vpwr scs8hd_decap_12
XFILLER_274_44 vgnd vpwr scs8hd_decap_12
XFILLER_143_15 vgnd vpwr scs8hd_decap_12
XFILLER_290_32 vgnd vpwr scs8hd_decap_12
XFILLER_143_59 vpwr vgnd scs8hd_fill_2
XFILLER_504_80 vgnd vpwr scs8hd_fill_1
XANTENNA__09__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_440_68 vgnd vpwr scs8hd_decap_12
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
XFILLER_299_74 vgnd vpwr scs8hd_decap_6
XPHY_1734 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_52_56 vgnd vpwr scs8hd_decap_12
XPHY_1701 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1712 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1723 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1767 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1756 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1745 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_139_3 vgnd vpwr scs8hd_decap_12
XFILLER_168_56 vgnd vpwr scs8hd_decap_12
XPHY_1789 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1778 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_318_15 vgnd vpwr scs8hd_decap_12
XFILLER_306_3 vgnd vpwr scs8hd_decap_12
XFILLER_184_22 vgnd vpwr scs8hd_decap_8
XFILLER_203_18 vpwr vgnd scs8hd_fill_2
XFILLER_414_80 vgnd vpwr scs8hd_fill_1
XFILLER_93_74 vgnd vpwr scs8hd_decap_6
XFILLER_350_68 vgnd vpwr scs8hd_decap_12
XFILLER_500_27 vgnd vpwr scs8hd_decap_4
XFILLER_228_15 vgnd vpwr scs8hd_decap_12
XFILLER_54_3 vgnd vpwr scs8hd_decap_12
XFILLER_324_80 vgnd vpwr scs8hd_fill_1
XFILLER_260_68 vgnd vpwr scs8hd_decap_12
XFILLER_410_27 vgnd vpwr scs8hd_decap_4
XPHY_409 vgnd vpwr scs8hd_decap_3
XPHY_1008 vgnd vpwr scs8hd_decap_3
XPHY_1019 vgnd vpwr scs8hd_decap_3
XFILLER_22_15 vgnd vpwr scs8hd_decap_12
XFILLER_138_15 vgnd vpwr scs8hd_decap_12
XFILLER_234_80 vgnd vpwr scs8hd_fill_1
XFILLER_601_15 vgnd vpwr scs8hd_decap_12
XFILLER_601_59 vpwr vgnd scs8hd_fill_2
XFILLER_103_51 vgnd vpwr scs8hd_decap_8
XFILLER_170_68 vgnd vpwr scs8hd_decap_12
XFILLER_103_62 vgnd vpwr scs8hd_decap_12
XFILLER_256_3 vgnd vpwr scs8hd_decap_12
XFILLER_320_27 vgnd vpwr scs8hd_decap_4
XPHY_910 vgnd vpwr scs8hd_decap_3
XPHY_921 vgnd vpwr scs8hd_decap_3
XPHY_932 vgnd vpwr scs8hd_decap_3
XPHY_943 vgnd vpwr scs8hd_decap_3
XPHY_954 vgnd vpwr scs8hd_decap_3
XPHY_1520 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1531 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1542 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_423_3 vgnd vpwr scs8hd_decap_12
XPHY_965 vgnd vpwr scs8hd_decap_3
XPHY_976 vgnd vpwr scs8hd_decap_3
XPHY_987 vgnd vpwr scs8hd_decap_3
XPHY_1553 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1564 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1575 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_998 vgnd vpwr scs8hd_decap_3
XFILLER_195_43 vgnd vpwr scs8hd_decap_12
XPHY_1586 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1597 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_409_80 vgnd vpwr scs8hd_fill_1
XFILLER_144_80 vgnd vpwr scs8hd_fill_1
X_12_ _07_/C _14_/B _07_/A _08_/Y _12_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_511_15 vgnd vpwr scs8hd_decap_12
XFILLER_511_59 vpwr vgnd scs8hd_fill_2
XFILLER_230_27 vgnd vpwr scs8hd_decap_4
Xlogical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ right_width_0_height_0__pin_4_ logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[2] vgnd vpwr scs8hd_ebufn_1
XFILLER_536_56 vgnd vpwr scs8hd_decap_12
XFILLER_319_80 vgnd vpwr scs8hd_fill_1
XFILLER_552_44 vgnd vpwr scs8hd_decap_12
XFILLER_405_27 vgnd vpwr scs8hd_decap_12
XFILLER_421_15 vgnd vpwr scs8hd_decap_12
XFILLER_17_15 vgnd vpwr scs8hd_decap_12
XFILLER_421_59 vpwr vgnd scs8hd_fill_2
XFILLER_17_59 vpwr vgnd scs8hd_fill_2
XFILLER_140_27 vgnd vpwr scs8hd_decap_4
XPHY_206 vgnd vpwr scs8hd_decap_3
XPHY_239 vgnd vpwr scs8hd_decap_3
XPHY_228 vgnd vpwr scs8hd_decap_3
XPHY_217 vgnd vpwr scs8hd_decap_3
XFILLER_577_74 vgnd vpwr scs8hd_decap_6
XFILLER_593_62 vgnd vpwr scs8hd_decap_12
XFILLER_593_51 vgnd vpwr scs8hd_decap_8
XFILLER_446_56 vgnd vpwr scs8hd_decap_12
XFILLER_165_68 vgnd vpwr scs8hd_fill_1
XFILLER_165_79 vpwr vgnd scs8hd_fill_2
XFILLER_315_27 vgnd vpwr scs8hd_decap_12
XFILLER_462_44 vgnd vpwr scs8hd_decap_12
XFILLER_58_44 vgnd vpwr scs8hd_decap_12
XFILLER_331_15 vgnd vpwr scs8hd_decap_12
XFILLER_373_3 vgnd vpwr scs8hd_decap_12
XFILLER_74_32 vgnd vpwr scs8hd_decap_12
XFILLER_331_59 vpwr vgnd scs8hd_fill_2
XFILLER_540_3 vgnd vpwr scs8hd_decap_12
XPHY_740 vgnd vpwr scs8hd_decap_3
XPHY_751 vgnd vpwr scs8hd_decap_3
XPHY_762 vgnd vpwr scs8hd_decap_3
XFILLER_487_74 vgnd vpwr scs8hd_decap_6
XPHY_1350 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_773 vgnd vpwr scs8hd_decap_3
XPHY_784 vgnd vpwr scs8hd_decap_3
XPHY_795 vgnd vpwr scs8hd_decap_3
XFILLER_23_80 vgnd vpwr scs8hd_fill_1
XPHY_1361 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1372 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1383 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_139_80 vgnd vpwr scs8hd_fill_1
XPHY_1394 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_356_56 vgnd vpwr scs8hd_decap_12
XFILLER_99_62 vgnd vpwr scs8hd_decap_12
XFILLER_99_51 vgnd vpwr scs8hd_decap_8
XFILLER_506_15 vgnd vpwr scs8hd_decap_12
XFILLER_225_16 vpwr vgnd scs8hd_fill_2
XFILLER_372_44 vgnd vpwr scs8hd_decap_12
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
XFILLER_241_15 vgnd vpwr scs8hd_decap_12
XFILLER_241_59 vpwr vgnd scs8hd_fill_2
XFILLER_602_80 vgnd vpwr scs8hd_fill_1
XFILLER_397_74 vgnd vpwr scs8hd_decap_6
XFILLER_119_39 vgnd vpwr scs8hd_decap_12
XFILLER_266_56 vgnd vpwr scs8hd_decap_12
XFILLER_416_15 vgnd vpwr scs8hd_decap_12
XFILLER_135_27 vgnd vpwr scs8hd_decap_12
XFILLER_282_44 vgnd vpwr scs8hd_decap_12
XFILLER_151_15 vgnd vpwr scs8hd_decap_12
XFILLER_151_59 vpwr vgnd scs8hd_fill_2
XFILLER_512_80 vgnd vpwr scs8hd_fill_1
XFILLER_44_68 vgnd vpwr scs8hd_decap_12
XFILLER_121_3 vgnd vpwr scs8hd_decap_12
XFILLER_60_56 vgnd vpwr scs8hd_decap_12
XFILLER_176_56 vgnd vpwr scs8hd_decap_12
XFILLER_219_3 vgnd vpwr scs8hd_decap_8
XFILLER_326_15 vgnd vpwr scs8hd_decap_12
XFILLER_588_3 vgnd vpwr scs8hd_decap_12
XFILLER_192_44 vgnd vpwr scs8hd_decap_12
XFILLER_490_3 vgnd vpwr scs8hd_decap_12
XFILLER_18_80 vgnd vpwr scs8hd_fill_1
XFILLER_422_80 vgnd vpwr scs8hd_fill_1
XPHY_570 vgnd vpwr scs8hd_decap_3
XPHY_581 vgnd vpwr scs8hd_decap_3
XPHY_592 vgnd vpwr scs8hd_decap_3
XFILLER_367_55 vgnd vpwr scs8hd_decap_6
XPHY_1191 vgnd vpwr scs8hd_decap_3
XPHY_1180 vgnd vpwr scs8hd_decap_3
XFILLER_236_15 vgnd vpwr scs8hd_decap_12
XFILLER_332_80 vgnd vpwr scs8hd_fill_1
XFILLER_558_32 vgnd vpwr scs8hd_decap_12
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XFILLER_201_62 vgnd vpwr scs8hd_decap_12
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
XFILLER_146_15 vgnd vpwr scs8hd_decap_12
XFILLER_507_80 vgnd vpwr scs8hd_fill_1
XFILLER_295_7 vpwr vgnd scs8hd_fill_2
XFILLER_242_80 vgnd vpwr scs8hd_fill_1
XFILLER_169_3 vgnd vpwr scs8hd_decap_12
XFILLER_111_62 vgnd vpwr scs8hd_decap_12
XFILLER_111_51 vgnd vpwr scs8hd_decap_8
XFILLER_468_32 vgnd vpwr scs8hd_decap_12
XFILLER_336_3 vgnd vpwr scs8hd_decap_12
XFILLER_503_3 vgnd vpwr scs8hd_decap_12
XFILLER_417_80 vgnd vpwr scs8hd_fill_1
XFILLER_503_27 vgnd vpwr scs8hd_decap_12
XFILLER_152_80 vgnd vpwr scs8hd_fill_1
XFILLER_378_32 vgnd vpwr scs8hd_decap_12
XFILLER_84_3 vgnd vpwr scs8hd_decap_12
XFILLER_528_68 vgnd vpwr scs8hd_decap_12
XFILLER_544_56 vgnd vpwr scs8hd_decap_12
XFILLER_327_80 vgnd vpwr scs8hd_fill_1
XFILLER_413_27 vgnd vpwr scs8hd_decap_12
XFILLER_560_44 vgnd vpwr scs8hd_decap_12
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XFILLER_25_15 vgnd vpwr scs8hd_decap_12
XPHY_48 vgnd vpwr scs8hd_decap_3
XFILLER_25_59 vpwr vgnd scs8hd_fill_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_288_32 vgnd vpwr scs8hd_decap_12
XANTENNA__14__D address[2] vgnd vpwr scs8hd_diode_2
XFILLER_585_74 vgnd vpwr scs8hd_decap_6
XFILLER_438_68 vgnd vpwr scs8hd_decap_12
XFILLER_237_80 vgnd vpwr scs8hd_fill_1
XFILLER_307_39 vgnd vpwr scs8hd_decap_12
XFILLER_454_56 vgnd vpwr scs8hd_decap_12
XFILLER_323_27 vgnd vpwr scs8hd_decap_12
XFILLER_66_44 vgnd vpwr scs8hd_decap_12
XFILLER_286_3 vgnd vpwr scs8hd_decap_12
XFILLER_470_44 vgnd vpwr scs8hd_decap_12
XFILLER_453_3 vgnd vpwr scs8hd_decap_12
XFILLER_82_32 vgnd vpwr scs8hd_decap_12
XFILLER_198_32 vgnd vpwr scs8hd_decap_12
XFILLER_348_68 vgnd vpwr scs8hd_decap_12
XFILLER_495_74 vgnd vpwr scs8hd_decap_6
XFILLER_31_80 vgnd vpwr scs8hd_fill_1
XFILLER_147_80 vgnd vpwr scs8hd_fill_1
XFILLER_364_56 vgnd vpwr scs8hd_decap_12
XFILLER_514_15 vgnd vpwr scs8hd_decap_12
XFILLER_233_27 vgnd vpwr scs8hd_decap_12
XFILLER_380_44 vgnd vpwr scs8hd_decap_12
XFILLER_258_68 vgnd vpwr scs8hd_decap_12
XFILLER_408_27 vgnd vpwr scs8hd_decap_4
XFILLER_11_39 vgnd vpwr scs8hd_decap_12
XFILLER_127_39 vgnd vpwr scs8hd_decap_12
XFILLER_274_56 vgnd vpwr scs8hd_decap_12
XFILLER_424_15 vgnd vpwr scs8hd_decap_12
XFILLER_143_27 vgnd vpwr scs8hd_decap_12
XFILLER_290_44 vgnd vpwr scs8hd_decap_12
XANTENNA__09__D _08_/Y vgnd vpwr scs8hd_diode_2
XFILLER_520_80 vgnd vpwr scs8hd_fill_1
XPHY_1702 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1713 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1724 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1757 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1746 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1735 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_52_68 vgnd vpwr scs8hd_decap_12
XPHY_1779 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1768 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_168_68 vgnd vpwr scs8hd_decap_12
XFILLER_318_27 vgnd vpwr scs8hd_decap_4
XFILLER_201_3 vpwr vgnd scs8hd_fill_2
XFILLER_184_78 vgnd vpwr scs8hd_decap_3
XFILLER_334_15 vgnd vpwr scs8hd_decap_12
XFILLER_570_3 vgnd vpwr scs8hd_decap_12
XFILLER_430_80 vgnd vpwr scs8hd_fill_1
XFILLER_26_80 vgnd vpwr scs8hd_fill_1
XFILLER_509_15 vgnd vpwr scs8hd_decap_12
XFILLER_509_59 vpwr vgnd scs8hd_fill_2
XFILLER_228_27 vgnd vpwr scs8hd_decap_4
XFILLER_47_3 vgnd vpwr scs8hd_decap_12
XFILLER_244_15 vgnd vpwr scs8hd_decap_12
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
XFILLER_3_51 vgnd vpwr scs8hd_decap_8
XFILLER_340_80 vgnd vpwr scs8hd_fill_1
XPHY_1009 vgnd vpwr scs8hd_decap_3
XFILLER_566_32 vgnd vpwr scs8hd_decap_12
XFILLER_419_15 vgnd vpwr scs8hd_decap_12
XFILLER_22_27 vgnd vpwr scs8hd_decap_4
XFILLER_419_59 vpwr vgnd scs8hd_fill_2
XFILLER_138_27 vgnd vpwr scs8hd_decap_4
XFILLER_154_15 vgnd vpwr scs8hd_decap_12
XFILLER_515_80 vgnd vpwr scs8hd_fill_1
XFILLER_601_27 vgnd vpwr scs8hd_decap_12
XFILLER_103_74 vgnd vpwr scs8hd_decap_6
XFILLER_250_80 vgnd vpwr scs8hd_fill_1
XFILLER_151_3 vgnd vpwr scs8hd_decap_12
XPHY_900 vgnd vpwr scs8hd_decap_3
XPHY_911 vgnd vpwr scs8hd_decap_3
XFILLER_249_3 vgnd vpwr scs8hd_decap_12
XPHY_922 vgnd vpwr scs8hd_decap_3
XPHY_933 vgnd vpwr scs8hd_decap_3
XPHY_944 vgnd vpwr scs8hd_decap_3
XPHY_1510 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1521 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1532 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_329_15 vgnd vpwr scs8hd_decap_12
XFILLER_476_32 vgnd vpwr scs8hd_decap_12
XPHY_955 vgnd vpwr scs8hd_decap_3
XPHY_966 vgnd vpwr scs8hd_decap_3
XPHY_977 vgnd vpwr scs8hd_decap_3
XPHY_988 vgnd vpwr scs8hd_decap_3
XFILLER_329_59 vpwr vgnd scs8hd_fill_2
XPHY_1543 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1554 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1565 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1576 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_416_3 vgnd vpwr scs8hd_decap_12
XPHY_999 vgnd vpwr scs8hd_decap_3
XFILLER_195_55 vgnd vpwr scs8hd_decap_6
XPHY_1587 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1598 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_425_80 vgnd vpwr scs8hd_fill_1
X_11_ enable _14_/B vgnd vpwr scs8hd_inv_8
XFILLER_511_27 vgnd vpwr scs8hd_decap_12
XFILLER_160_80 vgnd vpwr scs8hd_fill_1
XFILLER_239_15 vgnd vpwr scs8hd_decap_12
XFILLER_239_59 vpwr vgnd scs8hd_fill_2
XFILLER_386_32 vgnd vpwr scs8hd_decap_12
XFILLER_536_68 vgnd vpwr scs8hd_decap_12
XFILLER_405_39 vgnd vpwr scs8hd_decap_12
XFILLER_552_56 vgnd vpwr scs8hd_decap_12
XFILLER_335_80 vgnd vpwr scs8hd_fill_1
XFILLER_421_27 vgnd vpwr scs8hd_decap_12
XFILLER_17_27 vgnd vpwr scs8hd_decap_12
XPHY_207 vgnd vpwr scs8hd_decap_3
XPHY_229 vgnd vpwr scs8hd_decap_3
XPHY_218 vgnd vpwr scs8hd_decap_3
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XFILLER_33_59 vpwr vgnd scs8hd_fill_2
XFILLER_149_15 vgnd vpwr scs8hd_decap_12
XFILLER_149_59 vpwr vgnd scs8hd_fill_2
XFILLER_296_32 vgnd vpwr scs8hd_decap_12
XFILLER_593_74 vgnd vpwr scs8hd_decap_6
XFILLER_446_68 vgnd vpwr scs8hd_decap_12
XFILLER_315_39 vgnd vpwr scs8hd_decap_12
XFILLER_58_56 vgnd vpwr scs8hd_decap_12
XFILLER_245_80 vgnd vpwr scs8hd_fill_1
XFILLER_462_56 vgnd vpwr scs8hd_decap_12
XFILLER_199_3 vpwr vgnd scs8hd_fill_2
XFILLER_331_27 vgnd vpwr scs8hd_decap_12
XFILLER_366_3 vgnd vpwr scs8hd_decap_12
XFILLER_74_44 vgnd vpwr scs8hd_decap_12
XFILLER_533_3 vgnd vpwr scs8hd_decap_12
XFILLER_90_32 vgnd vpwr scs8hd_decap_12
XPHY_730 vgnd vpwr scs8hd_decap_3
XPHY_741 vgnd vpwr scs8hd_decap_3
XPHY_752 vgnd vpwr scs8hd_decap_3
XPHY_763 vgnd vpwr scs8hd_decap_3
XPHY_1340 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1351 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_774 vgnd vpwr scs8hd_decap_3
XPHY_785 vgnd vpwr scs8hd_decap_3
XPHY_796 vgnd vpwr scs8hd_decap_3
XPHY_1362 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1373 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1384 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1395 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_99_74 vgnd vpwr scs8hd_decap_6
XFILLER_356_68 vgnd vpwr scs8hd_decap_12
XFILLER_506_27 vgnd vpwr scs8hd_decap_4
XFILLER_155_80 vgnd vpwr scs8hd_fill_1
XFILLER_372_56 vgnd vpwr scs8hd_decap_12
XFILLER_522_15 vgnd vpwr scs8hd_decap_12
XFILLER_241_27 vgnd vpwr scs8hd_decap_12
XFILLER_266_68 vgnd vpwr scs8hd_decap_12
XFILLER_416_27 vgnd vpwr scs8hd_decap_4
XFILLER_135_39 vgnd vpwr scs8hd_decap_12
XFILLER_282_56 vgnd vpwr scs8hd_decap_12
XFILLER_432_15 vgnd vpwr scs8hd_decap_12
XFILLER_28_15 vgnd vpwr scs8hd_decap_12
XFILLER_151_27 vgnd vpwr scs8hd_decap_12
XFILLER_231_71 vgnd vpwr scs8hd_decap_8
XFILLER_60_68 vgnd vpwr scs8hd_decap_12
XFILLER_114_3 vgnd vpwr scs8hd_decap_12
XFILLER_176_68 vgnd vpwr scs8hd_decap_12
XFILLER_109_62 vgnd vpwr scs8hd_decap_12
XFILLER_109_51 vgnd vpwr scs8hd_decap_8
XFILLER_326_27 vgnd vpwr scs8hd_decap_4
XFILLER_192_56 vgnd vpwr scs8hd_decap_12
XFILLER_342_15 vgnd vpwr scs8hd_decap_12
XFILLER_483_3 vgnd vpwr scs8hd_decap_12
XFILLER_211_19 vpwr vgnd scs8hd_fill_2
XFILLER_34_80 vgnd vpwr scs8hd_fill_1
XPHY_560 vgnd vpwr scs8hd_decap_3
XPHY_571 vgnd vpwr scs8hd_decap_3
XPHY_582 vgnd vpwr scs8hd_decap_3
XPHY_593 vgnd vpwr scs8hd_decap_3
XPHY_1192 vgnd vpwr scs8hd_decap_3
XPHY_1181 vgnd vpwr scs8hd_decap_3
XPHY_1170 vgnd vpwr scs8hd_decap_3
XFILLER_517_15 vgnd vpwr scs8hd_decap_12
XFILLER_517_59 vpwr vgnd scs8hd_fill_2
XFILLER_236_27 vgnd vpwr scs8hd_decap_4
XFILLER_252_15 vgnd vpwr scs8hd_decap_12
XFILLER_558_44 vgnd vpwr scs8hd_decap_12
XFILLER_201_74 vgnd vpwr scs8hd_decap_6
XFILLER_427_15 vgnd vpwr scs8hd_decap_12
XFILLER_574_32 vgnd vpwr scs8hd_decap_12
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
XFILLER_427_59 vpwr vgnd scs8hd_fill_2
XFILLER_146_27 vgnd vpwr scs8hd_decap_4
XFILLER_162_15 vgnd vpwr scs8hd_decap_12
XFILLER_523_80 vgnd vpwr scs8hd_fill_1
XFILLER_599_51 vgnd vpwr scs8hd_decap_8
XFILLER_599_62 vgnd vpwr scs8hd_decap_12
XFILLER_111_74 vgnd vpwr scs8hd_decap_6
XFILLER_468_44 vgnd vpwr scs8hd_decap_12
XFILLER_231_3 vgnd vpwr scs8hd_decap_12
XFILLER_329_3 vgnd vpwr scs8hd_decap_12
XFILLER_337_15 vgnd vpwr scs8hd_decap_12
XFILLER_484_32 vgnd vpwr scs8hd_decap_12
XFILLER_337_59 vpwr vgnd scs8hd_fill_2
XFILLER_29_80 vgnd vpwr scs8hd_fill_1
XFILLER_433_80 vgnd vpwr scs8hd_fill_1
XFILLER_503_39 vgnd vpwr scs8hd_decap_12
XFILLER_378_44 vgnd vpwr scs8hd_decap_12
XFILLER_77_3 vgnd vpwr scs8hd_decap_12
XPHY_390 vgnd vpwr scs8hd_decap_3
XFILLER_247_15 vgnd vpwr scs8hd_decap_12
XFILLER_394_32 vgnd vpwr scs8hd_decap_12
XFILLER_247_59 vpwr vgnd scs8hd_fill_2
XFILLER_544_68 vgnd vpwr scs8hd_decap_12
XFILLER_560_56 vgnd vpwr scs8hd_decap_12
XFILLER_343_80 vgnd vpwr scs8hd_fill_1
XFILLER_413_39 vgnd vpwr scs8hd_decap_12
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_25_27 vgnd vpwr scs8hd_decap_12
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_288_44 vgnd vpwr scs8hd_decap_12
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XFILLER_157_15 vgnd vpwr scs8hd_decap_12
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_210_8 vpwr vgnd scs8hd_fill_2
XFILLER_157_59 vpwr vgnd scs8hd_fill_2
XFILLER_518_80 vgnd vpwr scs8hd_fill_1
XFILLER_454_68 vgnd vpwr scs8hd_decap_12
XFILLER_253_80 vgnd vpwr scs8hd_fill_1
XFILLER_323_39 vgnd vpwr scs8hd_decap_12
XFILLER_470_56 vgnd vpwr scs8hd_decap_12
XFILLER_66_56 vgnd vpwr scs8hd_decap_12
XFILLER_181_3 vgnd vpwr scs8hd_decap_12
XFILLER_279_3 vgnd vpwr scs8hd_decap_12
XFILLER_82_44 vgnd vpwr scs8hd_decap_12
XFILLER_446_3 vgnd vpwr scs8hd_decap_12
XFILLER_198_44 vgnd vpwr scs8hd_decap_12
XFILLER_428_80 vgnd vpwr scs8hd_fill_1
XFILLER_364_68 vgnd vpwr scs8hd_decap_12
XFILLER_514_27 vgnd vpwr scs8hd_decap_4
XFILLER_163_80 vgnd vpwr scs8hd_fill_1
XFILLER_233_39 vgnd vpwr scs8hd_decap_12
XFILLER_380_56 vgnd vpwr scs8hd_decap_12
XFILLER_530_15 vgnd vpwr scs8hd_decap_12
XFILLER_338_80 vgnd vpwr scs8hd_fill_1
XFILLER_274_68 vgnd vpwr scs8hd_decap_12
XFILLER_207_62 vgnd vpwr scs8hd_decap_12
XFILLER_424_27 vgnd vpwr scs8hd_decap_4
XFILLER_143_39 vgnd vpwr scs8hd_decap_12
XFILLER_290_56 vgnd vpwr scs8hd_decap_12
XFILLER_440_15 vgnd vpwr scs8hd_decap_12
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XPHY_1703 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1714 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1725 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1758 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1747 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1736 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1769 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_248_80 vgnd vpwr scs8hd_fill_1
XFILLER_184_46 vgnd vpwr scs8hd_decap_12
XFILLER_117_62 vgnd vpwr scs8hd_decap_12
XFILLER_117_51 vgnd vpwr scs8hd_decap_8
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XFILLER_334_27 vgnd vpwr scs8hd_decap_4
XFILLER_396_3 vgnd vpwr scs8hd_decap_12
XFILLER_563_3 vgnd vpwr scs8hd_decap_12
XFILLER_350_15 vgnd vpwr scs8hd_decap_12
XFILLER_509_27 vgnd vpwr scs8hd_decap_12
XFILLER_42_80 vgnd vpwr scs8hd_fill_1
XFILLER_158_80 vgnd vpwr scs8hd_fill_1
XFILLER_525_15 vgnd vpwr scs8hd_decap_12
XFILLER_525_59 vpwr vgnd scs8hd_fill_2
XFILLER_244_27 vgnd vpwr scs8hd_decap_4
XFILLER_3_74 vgnd vpwr scs8hd_decap_6
XFILLER_260_15 vgnd vpwr scs8hd_decap_12
XFILLER_419_27 vgnd vpwr scs8hd_decap_12
XFILLER_566_44 vgnd vpwr scs8hd_decap_12
XFILLER_582_32 vgnd vpwr scs8hd_decap_12
XFILLER_435_15 vgnd vpwr scs8hd_decap_12
XFILLER_154_27 vgnd vpwr scs8hd_decap_4
XFILLER_435_59 vpwr vgnd scs8hd_fill_2
XFILLER_170_15 vgnd vpwr scs8hd_decap_12
XFILLER_601_39 vgnd vpwr scs8hd_decap_12
XFILLER_531_80 vgnd vpwr scs8hd_fill_1
XPHY_901 vgnd vpwr scs8hd_decap_3
XPHY_912 vgnd vpwr scs8hd_decap_3
XPHY_1500 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_923 vgnd vpwr scs8hd_decap_3
XPHY_934 vgnd vpwr scs8hd_decap_3
XPHY_945 vgnd vpwr scs8hd_decap_3
XFILLER_144_3 vgnd vpwr scs8hd_decap_12
XPHY_1511 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1522 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1533 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_329_27 vgnd vpwr scs8hd_decap_12
XPHY_956 vgnd vpwr scs8hd_decap_3
XPHY_967 vgnd vpwr scs8hd_decap_3
XPHY_978 vgnd vpwr scs8hd_decap_3
XPHY_1544 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1555 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1566 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_476_44 vgnd vpwr scs8hd_decap_12
XPHY_989 vgnd vpwr scs8hd_decap_3
XFILLER_311_3 vgnd vpwr scs8hd_decap_12
XPHY_1577 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1588 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1599 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_409_3 vgnd vpwr scs8hd_decap_12
XFILLER_345_15 vgnd vpwr scs8hd_decap_12
XFILLER_492_32 vgnd vpwr scs8hd_decap_12
XFILLER_88_32 vgnd vpwr scs8hd_decap_12
XFILLER_345_59 vpwr vgnd scs8hd_fill_2
X_10_ _07_/C enable address[3] _08_/Y _10_/X vgnd vpwr scs8hd_and4_4
XFILLER_441_80 vgnd vpwr scs8hd_fill_1
XFILLER_511_39 vgnd vpwr scs8hd_decap_12
XFILLER_37_80 vgnd vpwr scs8hd_fill_1
XFILLER_239_27 vgnd vpwr scs8hd_decap_12
XFILLER_386_44 vgnd vpwr scs8hd_decap_12
XFILLER_255_15 vgnd vpwr scs8hd_decap_12
XFILLER_255_59 vpwr vgnd scs8hd_fill_2
XFILLER_552_68 vgnd vpwr scs8hd_decap_12
XFILLER_204_30 vgnd vpwr scs8hd_fill_1
XFILLER_351_80 vgnd vpwr scs8hd_fill_1
XFILLER_421_39 vgnd vpwr scs8hd_decap_12
XFILLER_17_39 vgnd vpwr scs8hd_decap_12
XPHY_219 vgnd vpwr scs8hd_decap_3
XPHY_208 vgnd vpwr scs8hd_decap_3
XFILLER_577_43 vgnd vpwr scs8hd_decap_12
XFILLER_33_27 vgnd vpwr scs8hd_decap_12
XFILLER_149_27 vgnd vpwr scs8hd_decap_12
XFILLER_296_44 vgnd vpwr scs8hd_decap_12
XFILLER_229_71 vgnd vpwr scs8hd_decap_8
XFILLER_165_15 vgnd vpwr scs8hd_decap_12
XFILLER_526_80 vgnd vpwr scs8hd_fill_1
XFILLER_165_59 vpwr vgnd scs8hd_fill_2
XFILLER_462_68 vgnd vpwr scs8hd_decap_12
XFILLER_58_68 vgnd vpwr scs8hd_decap_12
XFILLER_261_80 vgnd vpwr scs8hd_fill_1
XFILLER_331_39 vgnd vpwr scs8hd_decap_12
XFILLER_74_56 vgnd vpwr scs8hd_decap_12
XFILLER_261_3 vgnd vpwr scs8hd_decap_12
XFILLER_359_3 vgnd vpwr scs8hd_decap_12
XPHY_720 vgnd vpwr scs8hd_decap_3
XFILLER_526_3 vgnd vpwr scs8hd_decap_12
XFILLER_90_44 vgnd vpwr scs8hd_decap_12
XPHY_731 vgnd vpwr scs8hd_decap_3
XPHY_742 vgnd vpwr scs8hd_decap_3
XPHY_753 vgnd vpwr scs8hd_decap_3
XPHY_1341 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1330 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_764 vgnd vpwr scs8hd_decap_3
XPHY_775 vgnd vpwr scs8hd_decap_3
XPHY_786 vgnd vpwr scs8hd_decap_3
XPHY_1352 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1363 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1374 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_797 vgnd vpwr scs8hd_decap_3
XPHY_1385 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1396 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_436_80 vgnd vpwr scs8hd_fill_1
XFILLER_372_68 vgnd vpwr scs8hd_decap_12
XFILLER_522_27 vgnd vpwr scs8hd_decap_4
XFILLER_305_51 vgnd vpwr scs8hd_decap_8
XFILLER_305_62 vgnd vpwr scs8hd_decap_12
XFILLER_171_80 vgnd vpwr scs8hd_fill_1
XFILLER_241_39 vgnd vpwr scs8hd_decap_12
XFILLER_9_51 vgnd vpwr scs8hd_decap_8
XFILLER_9_62 vgnd vpwr scs8hd_decap_12
XFILLER_346_80 vgnd vpwr scs8hd_fill_1
XFILLER_282_68 vgnd vpwr scs8hd_decap_12
XFILLER_215_51 vgnd vpwr scs8hd_decap_8
XFILLER_215_62 vgnd vpwr scs8hd_decap_12
XFILLER_432_27 vgnd vpwr scs8hd_decap_4
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XFILLER_151_39 vgnd vpwr scs8hd_decap_12
XFILLER_44_15 vgnd vpwr scs8hd_decap_12
XFILLER_100_32 vgnd vpwr scs8hd_decap_12
XFILLER_109_74 vgnd vpwr scs8hd_decap_6
XFILLER_107_3 vgnd vpwr scs8hd_decap_12
XFILLER_256_80 vgnd vpwr scs8hd_fill_1
XFILLER_192_68 vgnd vpwr scs8hd_decap_12
XFILLER_125_51 vgnd vpwr scs8hd_decap_8
XFILLER_342_27 vgnd vpwr scs8hd_decap_4
XFILLER_125_62 vgnd vpwr scs8hd_decap_12
XFILLER_476_3 vgnd vpwr scs8hd_decap_12
XPHY_550 vgnd vpwr scs8hd_decap_3
XPHY_561 vgnd vpwr scs8hd_decap_3
XPHY_572 vgnd vpwr scs8hd_decap_3
XPHY_583 vgnd vpwr scs8hd_decap_3
XPHY_594 vgnd vpwr scs8hd_decap_3
XPHY_1193 vgnd vpwr scs8hd_decap_3
XPHY_1182 vgnd vpwr scs8hd_decap_3
XPHY_1171 vgnd vpwr scs8hd_decap_3
XPHY_1160 vgnd vpwr scs8hd_decap_3
XFILLER_517_27 vgnd vpwr scs8hd_decap_12
XFILLER_50_80 vgnd vpwr scs8hd_fill_1
XFILLER_533_15 vgnd vpwr scs8hd_decap_12
XFILLER_533_59 vpwr vgnd scs8hd_fill_2
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
XFILLER_252_27 vgnd vpwr scs8hd_decap_4
XFILLER_558_56 vgnd vpwr scs8hd_decap_12
XFILLER_574_44 vgnd vpwr scs8hd_decap_12
XFILLER_427_27 vgnd vpwr scs8hd_decap_12
XFILLER_590_32 vgnd vpwr scs8hd_decap_12
XFILLER_39_15 vgnd vpwr scs8hd_decap_12
XFILLER_443_15 vgnd vpwr scs8hd_decap_12
XFILLER_443_59 vpwr vgnd scs8hd_fill_2
XFILLER_39_59 vpwr vgnd scs8hd_fill_2
XFILLER_162_27 vgnd vpwr scs8hd_decap_4
XFILLER_599_74 vgnd vpwr scs8hd_decap_6
XFILLER_468_56 vgnd vpwr scs8hd_decap_12
XFILLER_224_3 vgnd vpwr scs8hd_decap_12
XFILLER_337_27 vgnd vpwr scs8hd_decap_12
XFILLER_484_44 vgnd vpwr scs8hd_decap_12
XFILLER_593_3 vgnd vpwr scs8hd_decap_12
XFILLER_353_15 vgnd vpwr scs8hd_decap_12
XFILLER_96_32 vgnd vpwr scs8hd_decap_12
XFILLER_353_59 vpwr vgnd scs8hd_fill_2
XFILLER_45_80 vgnd vpwr scs8hd_fill_1
XFILLER_378_56 vgnd vpwr scs8hd_decap_12
XFILLER_528_15 vgnd vpwr scs8hd_decap_12
XPHY_380 vgnd vpwr scs8hd_decap_3
XPHY_391 vgnd vpwr scs8hd_decap_3
XFILLER_247_27 vgnd vpwr scs8hd_decap_12
XFILLER_394_44 vgnd vpwr scs8hd_decap_12
XFILLER_263_15 vgnd vpwr scs8hd_decap_12
XFILLER_263_59 vpwr vgnd scs8hd_fill_2
XFILLER_560_68 vgnd vpwr scs8hd_decap_12
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_25_39 vgnd vpwr scs8hd_decap_12
XFILLER_288_56 vgnd vpwr scs8hd_decap_12
XFILLER_438_15 vgnd vpwr scs8hd_decap_12
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XFILLER_157_27 vgnd vpwr scs8hd_decap_12
XFILLER_173_15 vgnd vpwr scs8hd_decap_12
XFILLER_173_59 vpwr vgnd scs8hd_fill_2
XFILLER_534_80 vgnd vpwr scs8hd_fill_1
XFILLER_66_68 vgnd vpwr scs8hd_decap_12
XFILLER_403_51 vgnd vpwr scs8hd_decap_8
XFILLER_470_68 vgnd vpwr scs8hd_decap_12
XFILLER_174_3 vgnd vpwr scs8hd_decap_12
XFILLER_403_62 vgnd vpwr scs8hd_decap_12
XFILLER_82_56 vgnd vpwr scs8hd_decap_12
XFILLER_198_56 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _10_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_341_3 vgnd vpwr scs8hd_decap_12
XFILLER_439_3 vgnd vpwr scs8hd_decap_12
XFILLER_348_15 vgnd vpwr scs8hd_decap_12
XFILLER_444_80 vgnd vpwr scs8hd_fill_1
XFILLER_313_51 vgnd vpwr scs8hd_decap_8
XFILLER_380_68 vgnd vpwr scs8hd_decap_12
XFILLER_530_27 vgnd vpwr scs8hd_decap_4
XFILLER_313_62 vgnd vpwr scs8hd_decap_12
XFILLER_258_15 vgnd vpwr scs8hd_decap_12
XFILLER_207_74 vgnd vpwr scs8hd_decap_6
XFILLER_354_80 vgnd vpwr scs8hd_fill_1
XFILLER_223_51 vgnd vpwr scs8hd_decap_8
XFILLER_290_68 vgnd vpwr scs8hd_decap_12
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XFILLER_223_62 vgnd vpwr scs8hd_decap_12
XFILLER_440_27 vgnd vpwr scs8hd_decap_4
XFILLER_52_15 vgnd vpwr scs8hd_decap_12
XFILLER_168_15 vgnd vpwr scs8hd_decap_12
XPHY_1704 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1715 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1748 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1737 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1726 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1759 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_529_80 vgnd vpwr scs8hd_fill_1
XFILLER_184_58 vgnd vpwr scs8hd_decap_12
XFILLER_117_74 vgnd vpwr scs8hd_decap_6
XFILLER_264_80 vgnd vpwr scs8hd_fill_1
XFILLER_291_3 vgnd vpwr scs8hd_decap_12
XFILLER_389_3 vgnd vpwr scs8hd_decap_12
XFILLER_133_51 vgnd vpwr scs8hd_decap_8
XFILLER_133_62 vgnd vpwr scs8hd_decap_12
XFILLER_350_27 vgnd vpwr scs8hd_decap_4
XFILLER_556_3 vgnd vpwr scs8hd_decap_12
XFILLER_439_80 vgnd vpwr scs8hd_fill_1
XFILLER_509_39 vgnd vpwr scs8hd_decap_12
XFILLER_525_27 vgnd vpwr scs8hd_decap_12
XFILLER_174_80 vgnd vpwr scs8hd_fill_1
XFILLER_541_15 vgnd vpwr scs8hd_decap_12
XFILLER_541_59 vpwr vgnd scs8hd_fill_2
XFILLER_260_27 vgnd vpwr scs8hd_decap_4
XFILLER_566_56 vgnd vpwr scs8hd_decap_12
XFILLER_349_80 vgnd vpwr scs8hd_fill_1
XFILLER_419_39 vgnd vpwr scs8hd_decap_12
XFILLER_582_44 vgnd vpwr scs8hd_decap_12
XFILLER_435_27 vgnd vpwr scs8hd_decap_12
XFILLER_451_15 vgnd vpwr scs8hd_decap_12
XFILLER_47_15 vgnd vpwr scs8hd_decap_12
XFILLER_451_59 vpwr vgnd scs8hd_fill_2
XFILLER_47_59 vpwr vgnd scs8hd_fill_2
XFILLER_170_27 vgnd vpwr scs8hd_decap_4
XPHY_902 vgnd vpwr scs8hd_decap_3
XPHY_913 vgnd vpwr scs8hd_decap_3
XPHY_924 vgnd vpwr scs8hd_decap_3
XPHY_935 vgnd vpwr scs8hd_decap_3
XPHY_1501 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1512 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1523 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_946 vgnd vpwr scs8hd_decap_3
XPHY_957 vgnd vpwr scs8hd_decap_3
XPHY_968 vgnd vpwr scs8hd_decap_3
XPHY_979 vgnd vpwr scs8hd_decap_3
XFILLER_137_3 vgnd vpwr scs8hd_decap_12
XFILLER_259_80 vgnd vpwr scs8hd_fill_1
XPHY_1534 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_329_39 vgnd vpwr scs8hd_decap_12
XPHY_1545 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1556 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1567 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_476_56 vgnd vpwr scs8hd_decap_12
XPHY_1578 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1589 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_304_3 vgnd vpwr scs8hd_decap_12
XFILLER_345_27 vgnd vpwr scs8hd_decap_12
XFILLER_492_44 vgnd vpwr scs8hd_decap_12
XFILLER_88_44 vgnd vpwr scs8hd_decap_12
XFILLER_361_15 vgnd vpwr scs8hd_decap_12
XFILLER_361_59 vpwr vgnd scs8hd_fill_2
XFILLER_53_80 vgnd vpwr scs8hd_fill_1
XFILLER_169_80 vgnd vpwr scs8hd_fill_1
XFILLER_239_39 vgnd vpwr scs8hd_decap_12
XFILLER_386_56 vgnd vpwr scs8hd_decap_12
XFILLER_536_15 vgnd vpwr scs8hd_decap_12
XFILLER_52_3 vgnd vpwr scs8hd_decap_12
XFILLER_255_27 vgnd vpwr scs8hd_decap_12
XFILLER_271_15 vgnd vpwr scs8hd_decap_12
XFILLER_204_20 vpwr vgnd scs8hd_fill_2
XFILLER_271_59 vpwr vgnd scs8hd_fill_2
XFILLER_220_30 vgnd vpwr scs8hd_fill_1
XFILLER_501_51 vgnd vpwr scs8hd_decap_8
XFILLER_501_62 vgnd vpwr scs8hd_decap_12
XPHY_209 vgnd vpwr scs8hd_decap_3
XFILLER_577_55 vgnd vpwr scs8hd_decap_6
XFILLER_33_39 vgnd vpwr scs8hd_decap_12
XFILLER_149_39 vgnd vpwr scs8hd_decap_12
XFILLER_296_56 vgnd vpwr scs8hd_decap_12
XFILLER_446_15 vgnd vpwr scs8hd_decap_12
XFILLER_165_27 vgnd vpwr scs8hd_decap_12
XFILLER_181_15 vgnd vpwr scs8hd_decap_12
XFILLER_542_80 vgnd vpwr scs8hd_fill_1
XFILLER_74_68 vgnd vpwr scs8hd_decap_12
XFILLER_411_51 vgnd vpwr scs8hd_decap_8
XFILLER_411_62 vgnd vpwr scs8hd_decap_12
XFILLER_254_3 vgnd vpwr scs8hd_decap_12
XPHY_710 vgnd vpwr scs8hd_decap_3
XPHY_721 vgnd vpwr scs8hd_decap_3
XPHY_732 vgnd vpwr scs8hd_decap_3
XPHY_743 vgnd vpwr scs8hd_decap_3
XPHY_754 vgnd vpwr scs8hd_decap_3
XPHY_1331 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1320 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_90_56 vgnd vpwr scs8hd_decap_12
XPHY_1342 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_765 vgnd vpwr scs8hd_decap_3
XPHY_776 vgnd vpwr scs8hd_decap_3
XPHY_787 vgnd vpwr scs8hd_decap_3
XFILLER_421_3 vgnd vpwr scs8hd_decap_12
XFILLER_519_3 vgnd vpwr scs8hd_decap_12
XPHY_1353 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1364 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1375 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_798 vgnd vpwr scs8hd_decap_3
XPHY_1386 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1397 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_356_15 vgnd vpwr scs8hd_decap_12
XFILLER_305_74 vgnd vpwr scs8hd_decap_6
XFILLER_452_80 vgnd vpwr scs8hd_fill_1
XFILLER_48_80 vgnd vpwr scs8hd_fill_1
XFILLER_0_32 vgnd vpwr scs8hd_decap_4
XFILLER_321_51 vgnd vpwr scs8hd_decap_8
XFILLER_321_62 vgnd vpwr scs8hd_decap_12
XFILLER_9_74 vgnd vpwr scs8hd_decap_6
XFILLER_266_15 vgnd vpwr scs8hd_decap_12
XFILLER_215_74 vgnd vpwr scs8hd_decap_6
XFILLER_362_80 vgnd vpwr scs8hd_fill_1
XFILLER_588_32 vgnd vpwr scs8hd_decap_12
XFILLER_231_51 vgnd vpwr scs8hd_decap_8
XFILLER_231_62 vgnd vpwr scs8hd_decap_6
XFILLER_44_27 vgnd vpwr scs8hd_decap_4
XFILLER_100_44 vgnd vpwr scs8hd_decap_12
XFILLER_60_15 vgnd vpwr scs8hd_decap_12
XFILLER_176_15 vgnd vpwr scs8hd_decap_12
XFILLER_537_80 vgnd vpwr scs8hd_fill_1
XFILLER_125_74 vgnd vpwr scs8hd_decap_6
XFILLER_272_80 vgnd vpwr scs8hd_fill_1
XFILLER_371_3 vgnd vpwr scs8hd_decap_12
XFILLER_469_3 vgnd vpwr scs8hd_decap_12
XFILLER_141_51 vgnd vpwr scs8hd_decap_8
XFILLER_141_62 vgnd vpwr scs8hd_decap_12
XFILLER_498_32 vgnd vpwr scs8hd_decap_12
XPHY_540 vgnd vpwr scs8hd_decap_3
XPHY_551 vgnd vpwr scs8hd_decap_3
XPHY_562 vgnd vpwr scs8hd_decap_3
XPHY_1150 vgnd vpwr scs8hd_decap_3
XPHY_573 vgnd vpwr scs8hd_decap_3
XPHY_584 vgnd vpwr scs8hd_decap_3
XPHY_595 vgnd vpwr scs8hd_decap_3
XFILLER_367_47 vpwr vgnd scs8hd_fill_2
XPHY_1183 vgnd vpwr scs8hd_decap_3
XPHY_1172 vgnd vpwr scs8hd_decap_3
XPHY_1161 vgnd vpwr scs8hd_decap_3
XPHY_1194 vgnd vpwr scs8hd_decap_3
XFILLER_447_80 vgnd vpwr scs8hd_fill_1
XFILLER_517_39 vgnd vpwr scs8hd_decap_12
XFILLER_533_27 vgnd vpwr scs8hd_decap_12
XFILLER_182_80 vgnd vpwr scs8hd_fill_1
XFILLER_15_3 vgnd vpwr scs8hd_decap_12
XFILLER_558_68 vgnd vpwr scs8hd_decap_12
XFILLER_357_80 vgnd vpwr scs8hd_fill_1
XFILLER_427_39 vgnd vpwr scs8hd_decap_12
XFILLER_574_56 vgnd vpwr scs8hd_decap_12
XFILLER_443_27 vgnd vpwr scs8hd_decap_12
XFILLER_590_44 vgnd vpwr scs8hd_decap_12
XFILLER_39_27 vgnd vpwr scs8hd_decap_12
XFILLER_55_15 vgnd vpwr scs8hd_decap_12
XFILLER_55_59 vpwr vgnd scs8hd_fill_2
XFILLER_468_68 vgnd vpwr scs8hd_decap_12
XFILLER_217_3 vpwr vgnd scs8hd_fill_2
XFILLER_267_80 vgnd vpwr scs8hd_fill_1
XFILLER_337_39 vgnd vpwr scs8hd_decap_12
XFILLER_484_56 vgnd vpwr scs8hd_decap_12
XFILLER_353_27 vgnd vpwr scs8hd_decap_12
XFILLER_586_3 vgnd vpwr scs8hd_decap_12
XFILLER_96_44 vgnd vpwr scs8hd_decap_12
XPHY_370 vgnd vpwr scs8hd_decap_3
XFILLER_378_68 vgnd vpwr scs8hd_decap_12
XFILLER_528_27 vgnd vpwr scs8hd_decap_4
XPHY_381 vgnd vpwr scs8hd_decap_3
XPHY_392 vgnd vpwr scs8hd_decap_3
XFILLER_61_80 vgnd vpwr scs8hd_fill_1
XFILLER_247_39 vgnd vpwr scs8hd_decap_12
XFILLER_177_80 vgnd vpwr scs8hd_fill_1
XFILLER_394_56 vgnd vpwr scs8hd_decap_12
XFILLER_544_15 vgnd vpwr scs8hd_decap_12
XFILLER_263_27 vgnd vpwr scs8hd_decap_12
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_288_68 vgnd vpwr scs8hd_decap_12
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_438_27 vgnd vpwr scs8hd_decap_4
XFILLER_157_39 vgnd vpwr scs8hd_decap_12
XFILLER_454_15 vgnd vpwr scs8hd_decap_12
XFILLER_173_27 vgnd vpwr scs8hd_decap_12
XFILLER_106_32 vgnd vpwr scs8hd_decap_12
XFILLER_550_80 vgnd vpwr scs8hd_fill_1
XFILLER_403_74 vgnd vpwr scs8hd_decap_6
XFILLER_167_3 vgnd vpwr scs8hd_decap_12
XFILLER_82_68 vgnd vpwr scs8hd_decap_12
XFILLER_15_51 vgnd vpwr scs8hd_decap_8
XFILLER_15_62 vgnd vpwr scs8hd_decap_12
XFILLER_198_68 vgnd vpwr scs8hd_decap_12
XFILLER_334_3 vgnd vpwr scs8hd_decap_12
XFILLER_348_27 vgnd vpwr scs8hd_decap_4
XFILLER_501_3 vgnd vpwr scs8hd_decap_12
XFILLER_364_15 vgnd vpwr scs8hd_decap_12
XFILLER_313_74 vgnd vpwr scs8hd_decap_6
XFILLER_460_80 vgnd vpwr scs8hd_fill_1
XFILLER_56_80 vgnd vpwr scs8hd_fill_1
XFILLER_539_15 vgnd vpwr scs8hd_decap_12
XFILLER_539_59 vpwr vgnd scs8hd_fill_2
XFILLER_82_3 vgnd vpwr scs8hd_decap_12
XFILLER_258_27 vgnd vpwr scs8hd_decap_4
XFILLER_274_15 vgnd vpwr scs8hd_decap_12
XFILLER_207_31 vpwr vgnd scs8hd_fill_2
XFILLER_223_74 vgnd vpwr scs8hd_decap_6
XFILLER_370_80 vgnd vpwr scs8hd_fill_1
XFILLER_596_32 vgnd vpwr scs8hd_decap_12
XFILLER_449_15 vgnd vpwr scs8hd_decap_12
XFILLER_52_27 vgnd vpwr scs8hd_decap_4
XFILLER_449_59 vpwr vgnd scs8hd_fill_2
XPHY_1705 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1716 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1749 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1738 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_168_27 vgnd vpwr scs8hd_decap_4
XPHY_1727 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_184_15 vgnd vpwr scs8hd_decap_4
XFILLER_545_80 vgnd vpwr scs8hd_fill_1
XFILLER_284_3 vgnd vpwr scs8hd_decap_12
XFILLER_133_74 vgnd vpwr scs8hd_decap_6
XFILLER_280_80 vgnd vpwr scs8hd_fill_1
XFILLER_451_3 vgnd vpwr scs8hd_decap_12
XFILLER_549_3 vgnd vpwr scs8hd_decap_12
XFILLER_359_15 vgnd vpwr scs8hd_decap_12
XFILLER_359_59 vpwr vgnd scs8hd_fill_2
XFILLER_525_39 vgnd vpwr scs8hd_decap_12
XFILLER_455_80 vgnd vpwr scs8hd_fill_1
XFILLER_541_27 vgnd vpwr scs8hd_decap_12
XFILLER_190_80 vgnd vpwr scs8hd_fill_1
XFILLER_269_15 vgnd vpwr scs8hd_decap_12
XFILLER_269_59 vpwr vgnd scs8hd_fill_2
XFILLER_566_68 vgnd vpwr scs8hd_decap_12
XFILLER_435_39 vgnd vpwr scs8hd_decap_12
XFILLER_582_56 vgnd vpwr scs8hd_decap_12
XFILLER_365_80 vgnd vpwr scs8hd_fill_1
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _15_/Y vgnd vpwr scs8hd_diode_2
XFILLER_47_27 vgnd vpwr scs8hd_decap_12
XFILLER_451_27 vgnd vpwr scs8hd_decap_12
XFILLER_63_15 vgnd vpwr scs8hd_decap_12
XFILLER_179_15 vgnd vpwr scs8hd_decap_12
XPHY_903 vgnd vpwr scs8hd_decap_3
XFILLER_63_59 vpwr vgnd scs8hd_fill_2
XPHY_914 vgnd vpwr scs8hd_decap_3
XPHY_925 vgnd vpwr scs8hd_decap_3
XPHY_936 vgnd vpwr scs8hd_decap_3
XFILLER_179_59 vpwr vgnd scs8hd_fill_2
XPHY_1502 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1513 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1524 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_947 vgnd vpwr scs8hd_decap_3
XPHY_958 vgnd vpwr scs8hd_decap_3
XPHY_969 vgnd vpwr scs8hd_decap_3
XPHY_1535 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1546 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1557 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1568 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1579 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_476_68 vgnd vpwr scs8hd_decap_12
XFILLER_409_51 vgnd vpwr scs8hd_decap_8
XFILLER_409_62 vgnd vpwr scs8hd_decap_12
XFILLER_275_80 vgnd vpwr scs8hd_fill_1
XFILLER_345_39 vgnd vpwr scs8hd_decap_12
XFILLER_492_56 vgnd vpwr scs8hd_decap_12
XFILLER_88_56 vgnd vpwr scs8hd_decap_12
XFILLER_499_3 vgnd vpwr scs8hd_decap_12
XFILLER_361_27 vgnd vpwr scs8hd_decap_12
XFILLER_386_68 vgnd vpwr scs8hd_decap_12
XFILLER_536_27 vgnd vpwr scs8hd_decap_4
XFILLER_319_51 vgnd vpwr scs8hd_decap_8
XFILLER_319_62 vgnd vpwr scs8hd_decap_12
XFILLER_185_80 vgnd vpwr scs8hd_fill_1
XFILLER_255_39 vgnd vpwr scs8hd_decap_12
XFILLER_552_15 vgnd vpwr scs8hd_decap_12
XFILLER_45_3 vgnd vpwr scs8hd_decap_12
XFILLER_271_27 vgnd vpwr scs8hd_decap_12
XFILLER_204_32 vgnd vpwr scs8hd_decap_12
XFILLER_501_74 vgnd vpwr scs8hd_decap_6
XFILLER_296_68 vgnd vpwr scs8hd_decap_12
XFILLER_229_51 vgnd vpwr scs8hd_decap_8
XFILLER_229_62 vgnd vpwr scs8hd_decap_6
XFILLER_446_27 vgnd vpwr scs8hd_decap_4
XFILLER_165_39 vgnd vpwr scs8hd_decap_12
XFILLER_462_15 vgnd vpwr scs8hd_decap_12
XFILLER_58_15 vgnd vpwr scs8hd_decap_12
XFILLER_181_27 vgnd vpwr scs8hd_decap_12
XFILLER_114_32 vgnd vpwr scs8hd_decap_12
XFILLER_411_74 vgnd vpwr scs8hd_decap_6
XPHY_700 vgnd vpwr scs8hd_decap_3
XPHY_711 vgnd vpwr scs8hd_decap_3
XFILLER_247_3 vgnd vpwr scs8hd_decap_12
XPHY_722 vgnd vpwr scs8hd_decap_3
XPHY_733 vgnd vpwr scs8hd_decap_3
XPHY_744 vgnd vpwr scs8hd_decap_3
XPHY_1332 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1321 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1310 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_90_68 vgnd vpwr scs8hd_decap_12
XPHY_755 vgnd vpwr scs8hd_decap_3
XPHY_766 vgnd vpwr scs8hd_decap_3
XPHY_777 vgnd vpwr scs8hd_decap_3
XFILLER_23_51 vgnd vpwr scs8hd_decap_8
XFILLER_23_62 vgnd vpwr scs8hd_decap_12
XPHY_1343 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1354 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1365 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_788 vgnd vpwr scs8hd_decap_3
XPHY_799 vgnd vpwr scs8hd_decap_3
XFILLER_414_3 vgnd vpwr scs8hd_decap_12
XFILLER_139_51 vgnd vpwr scs8hd_decap_8
XFILLER_139_62 vgnd vpwr scs8hd_decap_12
XPHY_1376 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1387 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1398 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_356_27 vgnd vpwr scs8hd_decap_4
XFILLER_372_15 vgnd vpwr scs8hd_decap_12
XFILLER_321_74 vgnd vpwr scs8hd_decap_6
XFILLER_64_80 vgnd vpwr scs8hd_fill_1
XFILLER_547_15 vgnd vpwr scs8hd_decap_12
XFILLER_547_59 vpwr vgnd scs8hd_fill_2
XFILLER_266_27 vgnd vpwr scs8hd_decap_4
XFILLER_282_15 vgnd vpwr scs8hd_decap_12
XFILLER_588_44 vgnd vpwr scs8hd_decap_12
XFILLER_457_15 vgnd vpwr scs8hd_decap_12
XFILLER_100_56 vgnd vpwr scs8hd_decap_12
XFILLER_60_27 vgnd vpwr scs8hd_decap_4
XFILLER_176_27 vgnd vpwr scs8hd_decap_4
XFILLER_457_59 vpwr vgnd scs8hd_fill_2
XFILLER_192_15 vgnd vpwr scs8hd_decap_12
XFILLER_553_80 vgnd vpwr scs8hd_fill_1
XFILLER_197_3 vgnd vpwr scs8hd_decap_12
XFILLER_364_3 vgnd vpwr scs8hd_decap_12
XFILLER_141_74 vgnd vpwr scs8hd_decap_6
XFILLER_498_44 vgnd vpwr scs8hd_decap_12
XFILLER_531_3 vgnd vpwr scs8hd_decap_12
XPHY_530 vgnd vpwr scs8hd_decap_3
XPHY_541 vgnd vpwr scs8hd_decap_3
XPHY_552 vgnd vpwr scs8hd_decap_3
XFILLER_367_15 vgnd vpwr scs8hd_decap_12
XPHY_1140 vgnd vpwr scs8hd_decap_3
XPHY_563 vgnd vpwr scs8hd_decap_3
XPHY_574 vgnd vpwr scs8hd_decap_3
XPHY_585 vgnd vpwr scs8hd_decap_3
XPHY_596 vgnd vpwr scs8hd_decap_3
XPHY_1184 vgnd vpwr scs8hd_decap_3
XPHY_1173 vgnd vpwr scs8hd_decap_3
XPHY_1162 vgnd vpwr scs8hd_decap_3
XPHY_1151 vgnd vpwr scs8hd_decap_3
XPHY_1195 vgnd vpwr scs8hd_decap_3
XFILLER_533_39 vgnd vpwr scs8hd_decap_12
XFILLER_59_80 vgnd vpwr scs8hd_fill_1
XFILLER_463_80 vgnd vpwr scs8hd_fill_1
XFILLER_277_15 vgnd vpwr scs8hd_decap_12
XFILLER_277_59 vpwr vgnd scs8hd_fill_2
XFILLER_574_68 vgnd vpwr scs8hd_decap_12
XFILLER_507_51 vgnd vpwr scs8hd_decap_8
XFILLER_507_62 vgnd vpwr scs8hd_decap_12
XFILLER_226_30 vgnd vpwr scs8hd_fill_1
XFILLER_590_56 vgnd vpwr scs8hd_decap_12
XFILLER_39_39 vgnd vpwr scs8hd_decap_12
XFILLER_373_80 vgnd vpwr scs8hd_fill_1
XFILLER_443_39 vgnd vpwr scs8hd_decap_12
XFILLER_55_27 vgnd vpwr scs8hd_decap_12
XFILLER_71_15 vgnd vpwr scs8hd_decap_12
XFILLER_71_59 vpwr vgnd scs8hd_fill_2
XFILLER_187_15 vgnd vpwr scs8hd_decap_12
XFILLER_548_80 vgnd vpwr scs8hd_fill_1
XFILLER_187_59 vpwr vgnd scs8hd_fill_2
XFILLER_112_3 vgnd vpwr scs8hd_decap_12
XFILLER_484_68 vgnd vpwr scs8hd_decap_12
XFILLER_417_51 vgnd vpwr scs8hd_decap_8
XFILLER_417_62 vgnd vpwr scs8hd_decap_12
XFILLER_283_80 vgnd vpwr scs8hd_fill_1
XFILLER_353_39 vgnd vpwr scs8hd_decap_12
XFILLER_96_56 vgnd vpwr scs8hd_decap_12
XFILLER_481_3 vgnd vpwr scs8hd_decap_12
XFILLER_579_3 vgnd vpwr scs8hd_decap_12
XFILLER_302_32 vgnd vpwr scs8hd_decap_12
XPHY_360 vgnd vpwr scs8hd_decap_3
XPHY_371 vgnd vpwr scs8hd_decap_3
XPHY_382 vgnd vpwr scs8hd_decap_3
XPHY_393 vgnd vpwr scs8hd_decap_3
XFILLER_458_80 vgnd vpwr scs8hd_fill_1
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XFILLER_394_68 vgnd vpwr scs8hd_decap_12
XFILLER_544_27 vgnd vpwr scs8hd_decap_4
XFILLER_327_51 vgnd vpwr scs8hd_decap_8
XFILLER_327_62 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ right_width_0_height_0__pin_6_ logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[3] vgnd vpwr scs8hd_ebufn_1
XFILLER_193_80 vgnd vpwr scs8hd_fill_1
XFILLER_263_39 vgnd vpwr scs8hd_decap_12
XFILLER_560_15 vgnd vpwr scs8hd_decap_12
XFILLER_212_32 vgnd vpwr scs8hd_decap_12
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_237_51 vgnd vpwr scs8hd_decap_8
XFILLER_237_62 vgnd vpwr scs8hd_decap_12
XFILLER_454_27 vgnd vpwr scs8hd_decap_4
XFILLER_173_39 vgnd vpwr scs8hd_decap_12
XFILLER_106_44 vgnd vpwr scs8hd_decap_12
XFILLER_470_15 vgnd vpwr scs8hd_decap_12
XFILLER_66_15 vgnd vpwr scs8hd_decap_12
XFILLER_122_32 vgnd vpwr scs8hd_decap_12
XFILLER_15_74 vgnd vpwr scs8hd_decap_6
XFILLER_278_80 vgnd vpwr scs8hd_fill_1
XFILLER_327_3 vgnd vpwr scs8hd_decap_12
XFILLER_31_51 vgnd vpwr scs8hd_decap_8
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XFILLER_147_51 vgnd vpwr scs8hd_decap_8
XFILLER_147_62 vgnd vpwr scs8hd_decap_12
XFILLER_364_27 vgnd vpwr scs8hd_decap_4
XFILLER_380_15 vgnd vpwr scs8hd_decap_12
XFILLER_539_27 vgnd vpwr scs8hd_decap_12
XFILLER_72_80 vgnd vpwr scs8hd_fill_1
XFILLER_188_80 vgnd vpwr scs8hd_fill_1
XPHY_190 vgnd vpwr scs8hd_decap_3
XFILLER_75_3 vgnd vpwr scs8hd_decap_12
XFILLER_555_15 vgnd vpwr scs8hd_decap_12
XFILLER_555_59 vpwr vgnd scs8hd_fill_2
XFILLER_274_27 vgnd vpwr scs8hd_decap_4
XFILLER_290_15 vgnd vpwr scs8hd_decap_12
XFILLER_596_44 vgnd vpwr scs8hd_decap_12
XFILLER_449_27 vgnd vpwr scs8hd_decap_12
XPHY_1706 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1739 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1717 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1728 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_465_15 vgnd vpwr scs8hd_decap_12
XFILLER_465_59 vpwr vgnd scs8hd_fill_2
XFILLER_201_7 vgnd vpwr scs8hd_decap_3
XFILLER_561_80 vgnd vpwr scs8hd_fill_1
XFILLER_277_3 vgnd vpwr scs8hd_decap_12
XFILLER_444_3 vgnd vpwr scs8hd_decap_12
XFILLER_359_27 vgnd vpwr scs8hd_decap_12
XFILLER_375_15 vgnd vpwr scs8hd_decap_12
XFILLER_375_59 vpwr vgnd scs8hd_fill_2
XFILLER_541_39 vgnd vpwr scs8hd_decap_12
XFILLER_471_80 vgnd vpwr scs8hd_fill_1
XFILLER_67_80 vgnd vpwr scs8hd_fill_1
XFILLER_269_27 vgnd vpwr scs8hd_decap_12
XFILLER_285_15 vgnd vpwr scs8hd_decap_12
XFILLER_285_59 vpwr vgnd scs8hd_fill_2
XFILLER_582_68 vgnd vpwr scs8hd_decap_12
XFILLER_515_51 vgnd vpwr scs8hd_decap_8
XFILLER_515_62 vgnd vpwr scs8hd_decap_12
XFILLER_381_80 vgnd vpwr scs8hd_fill_1
XFILLER_451_39 vgnd vpwr scs8hd_decap_12
XFILLER_47_39 vgnd vpwr scs8hd_decap_12
XFILLER_63_27 vgnd vpwr scs8hd_decap_12
XFILLER_179_27 vgnd vpwr scs8hd_decap_12
XFILLER_400_32 vgnd vpwr scs8hd_decap_12
XPHY_904 vgnd vpwr scs8hd_decap_3
XPHY_915 vgnd vpwr scs8hd_decap_3
XPHY_926 vgnd vpwr scs8hd_decap_3
XPHY_1503 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1514 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_937 vgnd vpwr scs8hd_decap_3
XPHY_948 vgnd vpwr scs8hd_decap_3
XPHY_959 vgnd vpwr scs8hd_decap_3
XPHY_1525 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1536 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1547 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1558 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1569 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_556_80 vgnd vpwr scs8hd_fill_1
XFILLER_409_74 vgnd vpwr scs8hd_decap_6
XFILLER_492_68 vgnd vpwr scs8hd_decap_12
XFILLER_88_68 vgnd vpwr scs8hd_decap_12
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XFILLER_425_51 vgnd vpwr scs8hd_decap_8
XFILLER_425_62 vgnd vpwr scs8hd_decap_12
XFILLER_394_3 vgnd vpwr scs8hd_decap_12
XFILLER_291_80 vgnd vpwr scs8hd_fill_1
XFILLER_361_39 vgnd vpwr scs8hd_decap_12
XFILLER_561_3 vgnd vpwr scs8hd_decap_12
XFILLER_310_32 vgnd vpwr scs8hd_decap_12
XFILLER_319_74 vgnd vpwr scs8hd_decap_6
XFILLER_466_80 vgnd vpwr scs8hd_fill_1
XFILLER_552_27 vgnd vpwr scs8hd_decap_4
XFILLER_335_51 vgnd vpwr scs8hd_decap_8
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XFILLER_335_62 vgnd vpwr scs8hd_decap_12
XFILLER_271_39 vgnd vpwr scs8hd_decap_12
XFILLER_204_44 vgnd vpwr scs8hd_decap_12
XFILLER_220_32 vgnd vpwr scs8hd_decap_12
XFILLER_376_80 vgnd vpwr scs8hd_fill_1
XFILLER_245_51 vgnd vpwr scs8hd_decap_8
XFILLER_58_27 vgnd vpwr scs8hd_decap_4
XFILLER_245_62 vgnd vpwr scs8hd_decap_12
XFILLER_462_27 vgnd vpwr scs8hd_decap_4
XFILLER_181_39 vgnd vpwr scs8hd_decap_12
XFILLER_199_7 vgnd vpwr scs8hd_decap_12
XFILLER_114_44 vgnd vpwr scs8hd_decap_12
XFILLER_74_15 vgnd vpwr scs8hd_decap_12
XFILLER_130_32 vgnd vpwr scs8hd_decap_12
XPHY_701 vgnd vpwr scs8hd_decap_3
XPHY_712 vgnd vpwr scs8hd_decap_3
XPHY_723 vgnd vpwr scs8hd_decap_3
XPHY_734 vgnd vpwr scs8hd_decap_3
XPHY_745 vgnd vpwr scs8hd_decap_3
XPHY_1333 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1322 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1311 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1300 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_142_3 vgnd vpwr scs8hd_decap_12
XPHY_756 vgnd vpwr scs8hd_decap_3
XPHY_767 vgnd vpwr scs8hd_decap_3
XPHY_778 vgnd vpwr scs8hd_decap_3
XPHY_1344 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1355 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1366 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_789 vgnd vpwr scs8hd_decap_3
XFILLER_23_74 vgnd vpwr scs8hd_decap_6
XPHY_1377 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1388 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1399 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_407_3 vgnd vpwr scs8hd_decap_12
XFILLER_139_74 vgnd vpwr scs8hd_decap_6
XFILLER_286_80 vgnd vpwr scs8hd_fill_1
XFILLER_155_51 vgnd vpwr scs8hd_decap_8
XFILLER_155_62 vgnd vpwr scs8hd_decap_12
XFILLER_372_27 vgnd vpwr scs8hd_decap_4
XFILLER_0_67 vpwr vgnd scs8hd_fill_2
XFILLER_547_27 vgnd vpwr scs8hd_decap_12
XFILLER_80_80 vgnd vpwr scs8hd_fill_1
XFILLER_196_80 vgnd vpwr scs8hd_fill_1
XFILLER_563_15 vgnd vpwr scs8hd_decap_12
XFILLER_563_59 vpwr vgnd scs8hd_fill_2
XFILLER_282_27 vgnd vpwr scs8hd_decap_4
XFILLER_588_56 vgnd vpwr scs8hd_decap_12
XFILLER_100_68 vgnd vpwr scs8hd_decap_12
XFILLER_457_27 vgnd vpwr scs8hd_decap_12
XFILLER_473_15 vgnd vpwr scs8hd_decap_12
XFILLER_69_15 vgnd vpwr scs8hd_decap_12
XFILLER_473_59 vpwr vgnd scs8hd_fill_2
XFILLER_69_59 vpwr vgnd scs8hd_fill_2
XFILLER_192_27 vgnd vpwr scs8hd_decap_4
XFILLER_357_3 vgnd vpwr scs8hd_decap_12
XFILLER_498_56 vgnd vpwr scs8hd_decap_12
XFILLER_524_3 vgnd vpwr scs8hd_decap_12
XPHY_520 vgnd vpwr scs8hd_decap_3
XPHY_531 vgnd vpwr scs8hd_decap_3
XPHY_542 vgnd vpwr scs8hd_decap_3
XPHY_553 vgnd vpwr scs8hd_decap_3
XPHY_1141 vgnd vpwr scs8hd_decap_3
XPHY_1130 vgnd vpwr scs8hd_decap_3
XPHY_564 vgnd vpwr scs8hd_decap_3
XPHY_575 vgnd vpwr scs8hd_decap_3
XPHY_586 vgnd vpwr scs8hd_decap_3
XFILLER_367_27 vgnd vpwr scs8hd_decap_12
XPHY_1174 vgnd vpwr scs8hd_decap_3
XPHY_1163 vgnd vpwr scs8hd_decap_3
XPHY_1152 vgnd vpwr scs8hd_decap_3
XPHY_597 vgnd vpwr scs8hd_decap_3
XPHY_1196 vgnd vpwr scs8hd_decap_3
XPHY_1185 vgnd vpwr scs8hd_decap_3
XFILLER_383_15 vgnd vpwr scs8hd_decap_12
XFILLER_383_59 vpwr vgnd scs8hd_fill_2
XFILLER_75_80 vgnd vpwr scs8hd_fill_1
XFILLER_201_23 vgnd vpwr scs8hd_decap_12
XFILLER_558_15 vgnd vpwr scs8hd_decap_12
XFILLER_277_27 vgnd vpwr scs8hd_decap_12
XFILLER_293_15 vgnd vpwr scs8hd_decap_12
XFILLER_293_59 vpwr vgnd scs8hd_fill_2
XFILLER_507_74 vgnd vpwr scs8hd_decap_6
XFILLER_590_68 vgnd vpwr scs8hd_decap_12
XFILLER_523_51 vgnd vpwr scs8hd_decap_8
XFILLER_523_62 vgnd vpwr scs8hd_decap_12
XFILLER_55_39 vgnd vpwr scs8hd_decap_12
XFILLER_468_15 vgnd vpwr scs8hd_decap_12
XFILLER_71_27 vgnd vpwr scs8hd_decap_12
XFILLER_187_27 vgnd vpwr scs8hd_decap_12
XFILLER_105_3 vgnd vpwr scs8hd_decap_12
XFILLER_564_80 vgnd vpwr scs8hd_fill_1
XFILLER_417_74 vgnd vpwr scs8hd_decap_6
XFILLER_96_68 vgnd vpwr scs8hd_decap_12
XFILLER_433_51 vgnd vpwr scs8hd_decap_8
XFILLER_29_51 vgnd vpwr scs8hd_decap_8
XFILLER_29_62 vgnd vpwr scs8hd_decap_12
XFILLER_433_62 vgnd vpwr scs8hd_decap_12
XFILLER_474_3 vgnd vpwr scs8hd_decap_12
XFILLER_302_44 vgnd vpwr scs8hd_decap_12
XFILLER_378_15 vgnd vpwr scs8hd_decap_12
XPHY_350 vgnd vpwr scs8hd_decap_3
XPHY_361 vgnd vpwr scs8hd_decap_3
XPHY_372 vgnd vpwr scs8hd_decap_3
XPHY_383 vgnd vpwr scs8hd_decap_3
XPHY_394 vgnd vpwr scs8hd_decap_3
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XFILLER_327_74 vgnd vpwr scs8hd_decap_6
XFILLER_474_80 vgnd vpwr scs8hd_fill_1
XFILLER_560_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_343_51 vgnd vpwr scs8hd_decap_8
XFILLER_343_62 vgnd vpwr scs8hd_decap_12
XFILLER_212_44 vgnd vpwr scs8hd_decap_4
XFILLER_288_15 vgnd vpwr scs8hd_decap_12
XFILLER_237_74 vgnd vpwr scs8hd_decap_6
XFILLER_384_80 vgnd vpwr scs8hd_fill_1
XFILLER_106_56 vgnd vpwr scs8hd_decap_12
XFILLER_66_27 vgnd vpwr scs8hd_decap_4
XFILLER_253_51 vgnd vpwr scs8hd_decap_8
XFILLER_253_62 vgnd vpwr scs8hd_decap_12
XFILLER_470_27 vgnd vpwr scs8hd_decap_4
XFILLER_122_44 vgnd vpwr scs8hd_decap_12
XFILLER_82_15 vgnd vpwr scs8hd_decap_12
XFILLER_198_15 vgnd vpwr scs8hd_decap_12
XFILLER_559_80 vgnd vpwr scs8hd_fill_1
XFILLER_222_3 vgnd vpwr scs8hd_decap_12
XFILLER_31_74 vgnd vpwr scs8hd_decap_6
XFILLER_147_74 vgnd vpwr scs8hd_decap_6
XFILLER_294_80 vgnd vpwr scs8hd_fill_1
XFILLER_591_3 vgnd vpwr scs8hd_decap_12
XFILLER_163_51 vgnd vpwr scs8hd_decap_8
XFILLER_163_62 vgnd vpwr scs8hd_decap_12
XFILLER_380_27 vgnd vpwr scs8hd_decap_4
XFILLER_539_39 vgnd vpwr scs8hd_decap_12
XFILLER_469_80 vgnd vpwr scs8hd_fill_1
XPHY_191 vgnd vpwr scs8hd_decap_3
XPHY_180 vgnd vpwr scs8hd_decap_3
XFILLER_555_27 vgnd vpwr scs8hd_decap_12
XFILLER_68_3 vgnd vpwr scs8hd_decap_12
XFILLER_207_11 vpwr vgnd scs8hd_fill_2
XFILLER_571_15 vgnd vpwr scs8hd_decap_12
XFILLER_571_59 vpwr vgnd scs8hd_fill_2
XFILLER_290_27 vgnd vpwr scs8hd_decap_4
.ends

