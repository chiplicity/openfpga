magic
tech sky130A
magscale 1 2
timestamp 1606929606
<< locali >>
rect 10977 13787 11011 13957
rect 9505 13345 9597 13379
rect 9505 13243 9539 13345
rect 5181 9367 5215 9469
rect 949 1275 983 8789
rect 4905 3383 4939 3689
rect 6745 1479 6779 1853
rect 7113 1683 7147 1785
rect 11069 1479 11103 1785
rect 11713 1411 11747 1853
rect 14473 1411 14507 2057
<< viali >>
rect 11897 17289 11931 17323
rect 12817 17221 12851 17255
rect 5089 17153 5123 17187
rect 6101 17153 6135 17187
rect 6285 17153 6319 17187
rect 7757 17153 7791 17187
rect 8953 17153 8987 17187
rect 10425 17153 10459 17187
rect 14565 17153 14599 17187
rect 1869 17085 1903 17119
rect 2789 17085 2823 17119
rect 7573 17085 7607 17119
rect 10977 17085 11011 17119
rect 11713 17085 11747 17119
rect 12633 17085 12667 17119
rect 2145 17017 2179 17051
rect 3065 17017 3099 17051
rect 4905 17017 4939 17051
rect 7665 17017 7699 17051
rect 10241 17017 10275 17051
rect 13553 17017 13587 17051
rect 13645 17017 13679 17051
rect 4445 16949 4479 16983
rect 4813 16949 4847 16983
rect 5641 16949 5675 16983
rect 6009 16949 6043 16983
rect 7205 16949 7239 16983
rect 8401 16949 8435 16983
rect 8769 16949 8803 16983
rect 8861 16949 8895 16983
rect 9781 16949 9815 16983
rect 10149 16949 10183 16983
rect 11161 16949 11195 16983
rect 3433 16745 3467 16779
rect 6377 16745 6411 16779
rect 9689 16745 9723 16779
rect 10057 16745 10091 16779
rect 13277 16745 13311 16779
rect 14013 16745 14047 16779
rect 8585 16677 8619 16711
rect 1593 16609 1627 16643
rect 1869 16609 1903 16643
rect 2513 16609 2547 16643
rect 2789 16609 2823 16643
rect 3617 16609 3651 16643
rect 4620 16609 4654 16643
rect 6193 16609 6227 16643
rect 7297 16609 7331 16643
rect 8493 16609 8527 16643
rect 10149 16609 10183 16643
rect 10885 16609 10919 16643
rect 11621 16609 11655 16643
rect 12357 16609 12391 16643
rect 13093 16609 13127 16643
rect 13829 16609 13863 16643
rect 14565 16609 14599 16643
rect 4353 16541 4387 16575
rect 7389 16541 7423 16575
rect 7481 16541 7515 16575
rect 8677 16541 8711 16575
rect 10333 16541 10367 16575
rect 5733 16473 5767 16507
rect 11805 16473 11839 16507
rect 12541 16473 12575 16507
rect 6929 16405 6963 16439
rect 8125 16405 8159 16439
rect 11069 16405 11103 16439
rect 1593 16201 1627 16235
rect 3157 16201 3191 16235
rect 6929 16201 6963 16235
rect 13829 16201 13863 16235
rect 5549 16133 5583 16167
rect 8309 16133 8343 16167
rect 11805 16133 11839 16167
rect 13277 16133 13311 16167
rect 2513 16065 2547 16099
rect 3801 16065 3835 16099
rect 4813 16065 4847 16099
rect 4905 16065 4939 16099
rect 6193 16065 6227 16099
rect 7481 16065 7515 16099
rect 9781 16065 9815 16099
rect 11069 16065 11103 16099
rect 12449 16065 12483 16099
rect 14933 16065 14967 16099
rect 1409 15997 1443 16031
rect 2237 15997 2271 16031
rect 6009 15997 6043 16031
rect 8125 15997 8159 16031
rect 9045 15997 9079 16031
rect 9597 15997 9631 16031
rect 11621 15997 11655 16031
rect 12817 15997 12851 16031
rect 13645 15997 13679 16031
rect 14657 15997 14691 16031
rect 5917 15929 5951 15963
rect 7389 15929 7423 15963
rect 10793 15929 10827 15963
rect 13185 15929 13219 15963
rect 3525 15861 3559 15895
rect 3617 15861 3651 15895
rect 4353 15861 4387 15895
rect 4721 15861 4755 15895
rect 7297 15861 7331 15895
rect 8861 15861 8895 15895
rect 9229 15861 9263 15895
rect 9689 15861 9723 15895
rect 10425 15861 10459 15895
rect 10885 15861 10919 15895
rect 2789 15657 2823 15691
rect 3157 15657 3191 15691
rect 5733 15657 5767 15691
rect 7757 15657 7791 15691
rect 8125 15657 8159 15691
rect 9689 15657 9723 15691
rect 10885 15657 10919 15691
rect 11345 15657 11379 15691
rect 12449 15657 12483 15691
rect 13461 15657 13495 15691
rect 6929 15589 6963 15623
rect 1869 15521 1903 15555
rect 3249 15521 3283 15555
rect 4537 15521 4571 15555
rect 5825 15521 5859 15555
rect 10057 15521 10091 15555
rect 10149 15521 10183 15555
rect 11253 15521 11287 15555
rect 13277 15521 13311 15555
rect 14013 15521 14047 15555
rect 2145 15453 2179 15487
rect 3341 15453 3375 15487
rect 4629 15453 4663 15487
rect 4721 15453 4755 15487
rect 5917 15453 5951 15487
rect 7021 15453 7055 15487
rect 7205 15453 7239 15487
rect 8217 15453 8251 15487
rect 8309 15453 8343 15487
rect 8953 15453 8987 15487
rect 10241 15453 10275 15487
rect 11529 15453 11563 15487
rect 12541 15453 12575 15487
rect 12725 15453 12759 15487
rect 14197 15385 14231 15419
rect 4169 15317 4203 15351
rect 5365 15317 5399 15351
rect 6561 15317 6595 15351
rect 12081 15317 12115 15351
rect 5549 15113 5583 15147
rect 8677 15045 8711 15079
rect 12449 15045 12483 15079
rect 14565 15045 14599 15079
rect 2421 14977 2455 15011
rect 2605 14977 2639 15011
rect 3709 14977 3743 15011
rect 4905 14977 4939 15011
rect 9229 14977 9263 15011
rect 11713 14977 11747 15011
rect 13001 14977 13035 15011
rect 5733 14909 5767 14943
rect 6377 14909 6411 14943
rect 6837 14909 6871 14943
rect 10057 14909 10091 14943
rect 13645 14909 13679 14943
rect 14381 14909 14415 14943
rect 3617 14841 3651 14875
rect 4721 14841 4755 14875
rect 7104 14841 7138 14875
rect 9137 14841 9171 14875
rect 11529 14841 11563 14875
rect 12909 14841 12943 14875
rect 1961 14773 1995 14807
rect 2329 14773 2363 14807
rect 3157 14773 3191 14807
rect 3525 14773 3559 14807
rect 4353 14773 4387 14807
rect 4813 14773 4847 14807
rect 6193 14773 6227 14807
rect 8217 14773 8251 14807
rect 9045 14773 9079 14807
rect 9873 14773 9907 14807
rect 11069 14773 11103 14807
rect 11437 14773 11471 14807
rect 12817 14773 12851 14807
rect 13829 14773 13863 14807
rect 1593 14569 1627 14603
rect 4169 14569 4203 14603
rect 10885 14569 10919 14603
rect 12541 14569 12575 14603
rect 14657 14569 14691 14603
rect 2053 14501 2087 14535
rect 4537 14501 4571 14535
rect 5641 14501 5675 14535
rect 11253 14501 11287 14535
rect 13737 14501 13771 14535
rect 1961 14433 1995 14467
rect 3157 14433 3191 14467
rect 5365 14433 5399 14467
rect 6469 14433 6503 14467
rect 7104 14433 7138 14467
rect 9505 14433 9539 14467
rect 10276 14433 10310 14467
rect 10379 14433 10413 14467
rect 11345 14433 11379 14467
rect 12449 14433 12483 14467
rect 13185 14433 13219 14467
rect 13645 14433 13679 14467
rect 14473 14433 14507 14467
rect 2237 14365 2271 14399
rect 3249 14365 3283 14399
rect 3433 14365 3467 14399
rect 4629 14365 4663 14399
rect 4721 14365 4755 14399
rect 6837 14365 6871 14399
rect 8677 14365 8711 14399
rect 11437 14365 11471 14399
rect 12633 14365 12667 14399
rect 13921 14365 13955 14399
rect 2789 14229 2823 14263
rect 6285 14229 6319 14263
rect 8217 14229 8251 14263
rect 9321 14229 9355 14263
rect 12081 14229 12115 14263
rect 13277 14229 13311 14263
rect 3709 14025 3743 14059
rect 7297 14025 7331 14059
rect 11069 14025 11103 14059
rect 12449 14025 12483 14059
rect 2513 13957 2547 13991
rect 10977 13957 11011 13991
rect 3157 13889 3191 13923
rect 4261 13889 4295 13923
rect 7757 13889 7791 13923
rect 7849 13889 7883 13923
rect 1593 13821 1627 13855
rect 2881 13821 2915 13855
rect 4905 13821 4939 13855
rect 9137 13821 9171 13855
rect 11621 13889 11655 13923
rect 13093 13889 13127 13923
rect 13829 13889 13863 13923
rect 14105 13889 14139 13923
rect 1869 13753 1903 13787
rect 4169 13753 4203 13787
rect 5150 13753 5184 13787
rect 8493 13753 8527 13787
rect 9404 13753 9438 13787
rect 10977 13753 11011 13787
rect 13921 13753 13955 13787
rect 2973 13685 3007 13719
rect 4077 13685 4111 13719
rect 6285 13685 6319 13719
rect 7665 13685 7699 13719
rect 10517 13685 10551 13719
rect 11437 13685 11471 13719
rect 11529 13685 11563 13719
rect 12817 13685 12851 13719
rect 12909 13685 12943 13719
rect 2789 13481 2823 13515
rect 7205 13481 7239 13515
rect 7665 13481 7699 13515
rect 8125 13481 8159 13515
rect 3249 13413 3283 13447
rect 13093 13413 13127 13447
rect 14289 13413 14323 13447
rect 1961 13345 1995 13379
rect 3157 13345 3191 13379
rect 4077 13345 4111 13379
rect 6092 13345 6126 13379
rect 8033 13345 8067 13379
rect 8861 13345 8895 13379
rect 9597 13345 9631 13379
rect 9945 13345 9979 13379
rect 11897 13345 11931 13379
rect 14381 13345 14415 13379
rect 2053 13277 2087 13311
rect 2237 13277 2271 13311
rect 3433 13277 3467 13311
rect 4261 13277 4295 13311
rect 5181 13277 5215 13311
rect 5825 13277 5859 13311
rect 8309 13277 8343 13311
rect 9696 13277 9730 13311
rect 11989 13277 12023 13311
rect 12081 13277 12115 13311
rect 13185 13277 13219 13311
rect 13277 13277 13311 13311
rect 14473 13277 14507 13311
rect 1593 13209 1627 13243
rect 9505 13209 9539 13243
rect 11529 13209 11563 13243
rect 11069 13141 11103 13175
rect 12725 13141 12759 13175
rect 13921 13141 13955 13175
rect 1869 12937 1903 12971
rect 4445 12937 4479 12971
rect 6285 12937 6319 12971
rect 8769 12937 8803 12971
rect 10609 12937 10643 12971
rect 13645 12937 13679 12971
rect 15025 12937 15059 12971
rect 11805 12869 11839 12903
rect 2513 12801 2547 12835
rect 6929 12801 6963 12835
rect 9321 12801 9355 12835
rect 11253 12801 11287 12835
rect 13001 12801 13035 12835
rect 14197 12801 14231 12835
rect 3065 12733 3099 12767
rect 4905 12733 4939 12767
rect 5161 12733 5195 12767
rect 7196 12733 7230 12767
rect 11069 12733 11103 12767
rect 11989 12733 12023 12767
rect 14841 12733 14875 12767
rect 2237 12665 2271 12699
rect 3332 12665 3366 12699
rect 9229 12665 9263 12699
rect 14105 12665 14139 12699
rect 2329 12597 2363 12631
rect 8309 12597 8343 12631
rect 9137 12597 9171 12631
rect 9965 12597 9999 12631
rect 10977 12597 11011 12631
rect 12449 12597 12483 12631
rect 12817 12597 12851 12631
rect 12909 12597 12943 12631
rect 14013 12597 14047 12631
rect 1685 12393 1719 12427
rect 5181 12393 5215 12427
rect 5917 12393 5951 12427
rect 6285 12393 6319 12427
rect 9689 12393 9723 12427
rect 10057 12393 10091 12427
rect 10885 12393 10919 12427
rect 11253 12393 11287 12427
rect 12541 12393 12575 12427
rect 13645 12393 13679 12427
rect 14657 12393 14691 12427
rect 2053 12325 2087 12359
rect 5089 12325 5123 12359
rect 6377 12325 6411 12359
rect 7481 12325 7515 12359
rect 10149 12325 10183 12359
rect 2605 12257 2639 12291
rect 3341 12257 3375 12291
rect 7573 12257 7607 12291
rect 11345 12257 11379 12291
rect 12449 12257 12483 12291
rect 13737 12257 13771 12291
rect 14473 12257 14507 12291
rect 2145 12189 2179 12223
rect 2329 12189 2363 12223
rect 4077 12189 4111 12223
rect 4445 12189 4479 12223
rect 5365 12189 5399 12223
rect 6561 12189 6595 12223
rect 7665 12189 7699 12223
rect 8309 12189 8343 12223
rect 8953 12189 8987 12223
rect 10241 12189 10275 12223
rect 11437 12189 11471 12223
rect 12633 12189 12667 12223
rect 13829 12189 13863 12223
rect 7113 12121 7147 12155
rect 12081 12121 12115 12155
rect 4721 12053 4755 12087
rect 13277 12053 13311 12087
rect 6285 11849 6319 11883
rect 8217 11849 8251 11883
rect 10057 11849 10091 11883
rect 10517 11781 10551 11815
rect 12449 11781 12483 11815
rect 2513 11713 2547 11747
rect 3065 11713 3099 11747
rect 4905 11713 4939 11747
rect 6837 11713 6871 11747
rect 11069 11713 11103 11747
rect 13001 11713 13035 11747
rect 14197 11713 14231 11747
rect 2329 11645 2363 11679
rect 3332 11645 3366 11679
rect 7093 11645 7127 11679
rect 8677 11645 8711 11679
rect 8933 11645 8967 11679
rect 12909 11645 12943 11679
rect 14013 11645 14047 11679
rect 14841 11645 14875 11679
rect 5150 11577 5184 11611
rect 10885 11577 10919 11611
rect 1869 11509 1903 11543
rect 2237 11509 2271 11543
rect 4445 11509 4479 11543
rect 10977 11509 11011 11543
rect 11713 11509 11747 11543
rect 12817 11509 12851 11543
rect 13645 11509 13679 11543
rect 14105 11509 14139 11543
rect 15025 11509 15059 11543
rect 5457 11305 5491 11339
rect 6101 11305 6135 11339
rect 7757 11305 7791 11339
rect 8217 11305 8251 11339
rect 8861 11305 8895 11339
rect 11529 11305 11563 11339
rect 12725 11305 12759 11339
rect 13093 11305 13127 11339
rect 13921 11305 13955 11339
rect 14381 11305 14415 11339
rect 1869 11237 1903 11271
rect 6622 11237 6656 11271
rect 11897 11237 11931 11271
rect 11989 11237 12023 11271
rect 1593 11169 1627 11203
rect 2145 11169 2179 11203
rect 2412 11169 2446 11203
rect 4333 11169 4367 11203
rect 6285 11169 6319 11203
rect 9956 11169 9990 11203
rect 13185 11169 13219 11203
rect 14289 11169 14323 11203
rect 4077 11101 4111 11135
rect 6377 11101 6411 11135
rect 9689 11101 9723 11135
rect 12081 11101 12115 11135
rect 13277 11101 13311 11135
rect 14473 11101 14507 11135
rect 3525 11033 3559 11067
rect 11069 10965 11103 10999
rect 1593 10761 1627 10795
rect 1869 10761 1903 10795
rect 4445 10761 4479 10795
rect 6285 10761 6319 10795
rect 8217 10693 8251 10727
rect 10057 10693 10091 10727
rect 11897 10693 11931 10727
rect 15025 10693 15059 10727
rect 2513 10625 2547 10659
rect 3065 10625 3099 10659
rect 4905 10625 4939 10659
rect 6837 10625 6871 10659
rect 8677 10625 8711 10659
rect 13001 10625 13035 10659
rect 14197 10625 14231 10659
rect 1409 10557 1443 10591
rect 2237 10557 2271 10591
rect 10517 10557 10551 10591
rect 14013 10557 14047 10591
rect 14841 10557 14875 10591
rect 3332 10489 3366 10523
rect 5172 10489 5206 10523
rect 7104 10489 7138 10523
rect 8922 10489 8956 10523
rect 10784 10489 10818 10523
rect 12817 10489 12851 10523
rect 14105 10489 14139 10523
rect 2329 10421 2363 10455
rect 12449 10421 12483 10455
rect 12909 10421 12943 10455
rect 13645 10421 13679 10455
rect 1593 10217 1627 10251
rect 5457 10217 5491 10251
rect 11069 10217 11103 10251
rect 11529 10217 11563 10251
rect 11897 10217 11931 10251
rect 13185 10217 13219 10251
rect 13921 10217 13955 10251
rect 2412 10149 2446 10183
rect 6184 10149 6218 10183
rect 8024 10149 8058 10183
rect 14289 10149 14323 10183
rect 1409 10081 1443 10115
rect 2145 10081 2179 10115
rect 4344 10081 4378 10115
rect 9945 10081 9979 10115
rect 11989 10081 12023 10115
rect 13093 10081 13127 10115
rect 4077 10013 4111 10047
rect 5917 10013 5951 10047
rect 7757 10013 7791 10047
rect 9689 10013 9723 10047
rect 12173 10013 12207 10047
rect 13277 10013 13311 10047
rect 14381 10013 14415 10047
rect 14473 10013 14507 10047
rect 7297 9945 7331 9979
rect 9137 9945 9171 9979
rect 12725 9945 12759 9979
rect 3525 9877 3559 9911
rect 1869 9673 1903 9707
rect 12449 9673 12483 9707
rect 4445 9605 4479 9639
rect 10425 9605 10459 9639
rect 13645 9605 13679 9639
rect 2513 9537 2547 9571
rect 3065 9537 3099 9571
rect 5273 9537 5307 9571
rect 13001 9537 13035 9571
rect 14197 9537 14231 9571
rect 2329 9469 2363 9503
rect 5089 9469 5123 9503
rect 5181 9469 5215 9503
rect 9045 9469 9079 9503
rect 10517 9469 10551 9503
rect 12817 9469 12851 9503
rect 14013 9469 14047 9503
rect 14841 9469 14875 9503
rect 2237 9401 2271 9435
rect 3332 9401 3366 9435
rect 5540 9401 5574 9435
rect 7205 9401 7239 9435
rect 8769 9401 8803 9435
rect 9312 9401 9346 9435
rect 10784 9401 10818 9435
rect 12909 9401 12943 9435
rect 4905 9333 4939 9367
rect 5181 9333 5215 9367
rect 6653 9333 6687 9367
rect 11897 9333 11931 9367
rect 14105 9333 14139 9367
rect 15025 9333 15059 9367
rect 13369 9129 13403 9163
rect 6000 9061 6034 9095
rect 9934 9061 9968 9095
rect 1409 8993 1443 9027
rect 2412 8993 2446 9027
rect 4528 8993 4562 9027
rect 5733 8993 5767 9027
rect 7829 8993 7863 9027
rect 9689 8993 9723 9027
rect 11796 8993 11830 9027
rect 13737 8993 13771 9027
rect 2145 8925 2179 8959
rect 4261 8925 4295 8959
rect 7573 8925 7607 8959
rect 11529 8925 11563 8959
rect 13829 8925 13863 8959
rect 14013 8925 14047 8959
rect 14565 8925 14599 8959
rect 5641 8857 5675 8891
rect 11069 8857 11103 8891
rect 949 8789 983 8823
rect 1593 8789 1627 8823
rect 3525 8789 3559 8823
rect 7113 8789 7147 8823
rect 8953 8789 8987 8823
rect 12909 8789 12943 8823
rect 2237 8585 2271 8619
rect 4445 8585 4479 8619
rect 11897 8585 11931 8619
rect 12449 8585 12483 8619
rect 6285 8517 6319 8551
rect 13645 8517 13679 8551
rect 2053 8449 2087 8483
rect 2881 8449 2915 8483
rect 3065 8449 3099 8483
rect 4905 8449 4939 8483
rect 13001 8449 13035 8483
rect 14197 8449 14231 8483
rect 2697 8381 2731 8415
rect 3332 8381 3366 8415
rect 6837 8381 6871 8415
rect 8677 8381 8711 8415
rect 10517 8381 10551 8415
rect 14105 8381 14139 8415
rect 14841 8381 14875 8415
rect 1777 8313 1811 8347
rect 1869 8313 1903 8347
rect 5172 8313 5206 8347
rect 7082 8313 7116 8347
rect 8922 8313 8956 8347
rect 10762 8313 10796 8347
rect 12909 8313 12943 8347
rect 1409 8245 1443 8279
rect 2605 8245 2639 8279
rect 8217 8245 8251 8279
rect 10057 8245 10091 8279
rect 12817 8245 12851 8279
rect 14013 8245 14047 8279
rect 15025 8245 15059 8279
rect 3525 8041 3559 8075
rect 4905 8041 4939 8075
rect 11529 8041 11563 8075
rect 11989 8041 12023 8075
rect 12725 8041 12759 8075
rect 13921 8041 13955 8075
rect 9934 7973 9968 8007
rect 11897 7973 11931 8007
rect 13093 7973 13127 8007
rect 1409 7905 1443 7939
rect 2145 7905 2179 7939
rect 2412 7905 2446 7939
rect 5713 7905 5747 7939
rect 7553 7905 7587 7939
rect 9321 7905 9355 7939
rect 14289 7905 14323 7939
rect 4997 7837 5031 7871
rect 5181 7837 5215 7871
rect 5457 7837 5491 7871
rect 7297 7837 7331 7871
rect 9689 7837 9723 7871
rect 12081 7837 12115 7871
rect 13185 7837 13219 7871
rect 13277 7837 13311 7871
rect 14381 7837 14415 7871
rect 14473 7837 14507 7871
rect 1593 7701 1627 7735
rect 4537 7701 4571 7735
rect 6837 7701 6871 7735
rect 8677 7701 8711 7735
rect 9137 7701 9171 7735
rect 11069 7701 11103 7735
rect 4445 7497 4479 7531
rect 10517 7497 10551 7531
rect 12449 7497 12483 7531
rect 13645 7497 13679 7531
rect 1869 7429 1903 7463
rect 6285 7429 6319 7463
rect 8217 7429 8251 7463
rect 2513 7361 2547 7395
rect 11069 7361 11103 7395
rect 11713 7361 11747 7395
rect 13001 7361 13035 7395
rect 14105 7361 14139 7395
rect 14289 7361 14323 7395
rect 3065 7293 3099 7327
rect 4905 7293 4939 7327
rect 6837 7293 6871 7327
rect 8677 7293 8711 7327
rect 10885 7293 10919 7327
rect 10977 7293 11011 7327
rect 12817 7293 12851 7327
rect 14013 7293 14047 7327
rect 14841 7293 14875 7327
rect 2237 7225 2271 7259
rect 3332 7225 3366 7259
rect 5172 7225 5206 7259
rect 7082 7225 7116 7259
rect 8922 7225 8956 7259
rect 2329 7157 2363 7191
rect 10057 7157 10091 7191
rect 12909 7157 12943 7191
rect 15025 7157 15059 7191
rect 8953 6953 8987 6987
rect 10057 6953 10091 6987
rect 12449 6953 12483 6987
rect 13277 6953 13311 6987
rect 1869 6885 1903 6919
rect 4905 6885 4939 6919
rect 11253 6885 11287 6919
rect 1593 6817 1627 6851
rect 2412 6817 2446 6851
rect 5733 6817 5767 6851
rect 6000 6817 6034 6851
rect 7573 6817 7607 6851
rect 7840 6817 7874 6851
rect 11345 6817 11379 6851
rect 13645 6817 13679 6851
rect 13737 6817 13771 6851
rect 14473 6817 14507 6851
rect 2145 6749 2179 6783
rect 4997 6749 5031 6783
rect 5181 6749 5215 6783
rect 10149 6749 10183 6783
rect 10333 6749 10367 6783
rect 11437 6749 11471 6783
rect 12541 6749 12575 6783
rect 12633 6749 12667 6783
rect 13829 6749 13863 6783
rect 3525 6681 3559 6715
rect 4537 6613 4571 6647
rect 7113 6613 7147 6647
rect 9689 6613 9723 6647
rect 10885 6613 10919 6647
rect 12081 6613 12115 6647
rect 14657 6613 14691 6647
rect 6285 6409 6319 6443
rect 10517 6409 10551 6443
rect 12449 6409 12483 6443
rect 10057 6341 10091 6375
rect 2513 6273 2547 6307
rect 11069 6273 11103 6307
rect 13001 6273 13035 6307
rect 14197 6273 14231 6307
rect 1409 6205 1443 6239
rect 3065 6205 3099 6239
rect 4905 6205 4939 6239
rect 6837 6205 6871 6239
rect 8677 6205 8711 6239
rect 10977 6205 11011 6239
rect 14105 6205 14139 6239
rect 14841 6205 14875 6239
rect 3332 6137 3366 6171
rect 5172 6137 5206 6171
rect 7082 6137 7116 6171
rect 8944 6137 8978 6171
rect 10885 6137 10919 6171
rect 12817 6137 12851 6171
rect 13277 6137 13311 6171
rect 14013 6137 14047 6171
rect 1593 6069 1627 6103
rect 1869 6069 1903 6103
rect 2237 6069 2271 6103
rect 2329 6069 2363 6103
rect 4445 6069 4479 6103
rect 8217 6069 8251 6103
rect 11713 6069 11747 6103
rect 12909 6069 12943 6103
rect 13645 6069 13679 6103
rect 15025 6069 15059 6103
rect 1593 5865 1627 5899
rect 2053 5865 2087 5899
rect 4905 5865 4939 5899
rect 7113 5865 7147 5899
rect 11253 5865 11287 5899
rect 12081 5865 12115 5899
rect 13645 5865 13679 5899
rect 1961 5797 1995 5831
rect 6000 5797 6034 5831
rect 10057 5797 10091 5831
rect 11345 5797 11379 5831
rect 12449 5797 12483 5831
rect 13737 5797 13771 5831
rect 3157 5729 3191 5763
rect 3249 5729 3283 5763
rect 7665 5729 7699 5763
rect 7932 5729 7966 5763
rect 14473 5729 14507 5763
rect 2237 5661 2271 5695
rect 3433 5661 3467 5695
rect 4997 5661 5031 5695
rect 5181 5661 5215 5695
rect 5733 5661 5767 5695
rect 10149 5661 10183 5695
rect 10333 5661 10367 5695
rect 11529 5661 11563 5695
rect 12541 5661 12575 5695
rect 12633 5661 12667 5695
rect 13829 5661 13863 5695
rect 9689 5593 9723 5627
rect 10885 5593 10919 5627
rect 2789 5525 2823 5559
rect 4537 5525 4571 5559
rect 9045 5525 9079 5559
rect 13277 5525 13311 5559
rect 14657 5525 14691 5559
rect 1409 5321 1443 5355
rect 6285 5321 6319 5355
rect 9229 5321 9263 5355
rect 10425 5253 10459 5287
rect 13645 5253 13679 5287
rect 1869 5185 1903 5219
rect 2053 5185 2087 5219
rect 2973 5185 3007 5219
rect 3157 5185 3191 5219
rect 4261 5185 4295 5219
rect 9873 5185 9907 5219
rect 10977 5185 11011 5219
rect 12909 5185 12943 5219
rect 13001 5185 13035 5219
rect 14197 5185 14231 5219
rect 1777 5117 1811 5151
rect 2881 5117 2915 5151
rect 4905 5117 4939 5151
rect 5172 5117 5206 5151
rect 7389 5117 7423 5151
rect 10793 5117 10827 5151
rect 11621 5117 11655 5151
rect 14013 5117 14047 5151
rect 14841 5117 14875 5151
rect 4077 5049 4111 5083
rect 7656 5049 7690 5083
rect 10885 5049 10919 5083
rect 12817 5049 12851 5083
rect 2513 4981 2547 5015
rect 3709 4981 3743 5015
rect 4169 4981 4203 5015
rect 8769 4981 8803 5015
rect 9597 4981 9631 5015
rect 9689 4981 9723 5015
rect 11805 4981 11839 5015
rect 12449 4981 12483 5015
rect 14105 4981 14139 5015
rect 15025 4981 15059 5015
rect 2789 4777 2823 4811
rect 4537 4777 4571 4811
rect 5273 4777 5307 4811
rect 8309 4777 8343 4811
rect 8769 4777 8803 4811
rect 9689 4777 9723 4811
rect 10057 4777 10091 4811
rect 13277 4777 13311 4811
rect 13737 4777 13771 4811
rect 14657 4777 14691 4811
rect 1676 4709 1710 4743
rect 4445 4709 4479 4743
rect 6714 4709 6748 4743
rect 13645 4709 13679 4743
rect 3249 4641 3283 4675
rect 5641 4641 5675 4675
rect 6469 4641 6503 4675
rect 8677 4641 8711 4675
rect 10149 4641 10183 4675
rect 11253 4641 11287 4675
rect 11345 4641 11379 4675
rect 12449 4641 12483 4675
rect 14473 4641 14507 4675
rect 3341 4573 3375 4607
rect 3525 4573 3559 4607
rect 4721 4573 4755 4607
rect 5733 4573 5767 4607
rect 5825 4573 5859 4607
rect 8861 4573 8895 4607
rect 10241 4573 10275 4607
rect 11529 4573 11563 4607
rect 12541 4573 12575 4607
rect 12725 4573 12759 4607
rect 13829 4573 13863 4607
rect 2881 4505 2915 4539
rect 4077 4437 4111 4471
rect 7849 4437 7883 4471
rect 10885 4437 10919 4471
rect 12081 4437 12115 4471
rect 5549 4233 5583 4267
rect 6837 4233 6871 4267
rect 8033 4233 8067 4267
rect 8861 4233 8895 4267
rect 11253 4233 11287 4267
rect 3985 4165 4019 4199
rect 2237 4097 2271 4131
rect 4629 4097 4663 4131
rect 6009 4097 6043 4131
rect 6101 4097 6135 4131
rect 7389 4097 7423 4131
rect 8585 4097 8619 4131
rect 9413 4097 9447 4131
rect 10977 4097 11011 4131
rect 11805 4097 11839 4131
rect 13001 4097 13035 4131
rect 14197 4097 14231 4131
rect 2605 4029 2639 4063
rect 4905 4029 4939 4063
rect 7297 4029 7331 4063
rect 9229 4029 9263 4063
rect 9321 4029 9355 4063
rect 10241 4029 10275 4063
rect 10885 4029 10919 4063
rect 11621 4029 11655 4063
rect 14841 4029 14875 4063
rect 1961 3961 1995 3995
rect 2850 3961 2884 3995
rect 5181 3961 5215 3995
rect 8401 3961 8435 3995
rect 10793 3961 10827 3995
rect 11713 3961 11747 3995
rect 12817 3961 12851 3995
rect 14013 3961 14047 3995
rect 14105 3961 14139 3995
rect 1593 3893 1627 3927
rect 2053 3893 2087 3927
rect 4077 3893 4111 3927
rect 4445 3893 4479 3927
rect 4537 3893 4571 3927
rect 5917 3893 5951 3927
rect 7205 3893 7239 3927
rect 8493 3893 8527 3927
rect 10057 3893 10091 3927
rect 10425 3893 10459 3927
rect 12449 3893 12483 3927
rect 12909 3893 12943 3927
rect 13645 3893 13679 3927
rect 15025 3893 15059 3927
rect 2789 3689 2823 3723
rect 2881 3689 2915 3723
rect 3341 3689 3375 3723
rect 4077 3689 4111 3723
rect 4905 3689 4939 3723
rect 5825 3689 5859 3723
rect 7113 3689 7147 3723
rect 7481 3689 7515 3723
rect 8309 3689 8343 3723
rect 8769 3689 8803 3723
rect 9689 3689 9723 3723
rect 13277 3689 13311 3723
rect 13645 3689 13679 3723
rect 14657 3689 14691 3723
rect 1676 3621 1710 3655
rect 4445 3621 4479 3655
rect 3249 3553 3283 3587
rect 1409 3485 1443 3519
rect 3525 3485 3559 3519
rect 4537 3485 4571 3519
rect 4721 3485 4755 3519
rect 6193 3621 6227 3655
rect 7021 3621 7055 3655
rect 7941 3621 7975 3655
rect 10149 3621 10183 3655
rect 12449 3621 12483 3655
rect 5365 3553 5399 3587
rect 6285 3553 6319 3587
rect 7849 3553 7883 3587
rect 8677 3553 8711 3587
rect 10057 3553 10091 3587
rect 11253 3553 11287 3587
rect 11345 3553 11379 3587
rect 11713 3553 11747 3587
rect 12541 3553 12575 3587
rect 13737 3553 13771 3587
rect 14473 3553 14507 3587
rect 5457 3485 5491 3519
rect 5641 3485 5675 3519
rect 6469 3485 6503 3519
rect 7297 3485 7331 3519
rect 8125 3485 8159 3519
rect 8861 3485 8895 3519
rect 10333 3485 10367 3519
rect 11437 3485 11471 3519
rect 12633 3485 12667 3519
rect 13829 3485 13863 3519
rect 6653 3417 6687 3451
rect 10885 3417 10919 3451
rect 4905 3349 4939 3383
rect 4997 3349 5031 3383
rect 11897 3349 11931 3383
rect 12081 3349 12115 3383
rect 4261 3145 4295 3179
rect 6837 3145 6871 3179
rect 7665 3145 7699 3179
rect 9229 3145 9263 3179
rect 11253 3145 11287 3179
rect 15301 3145 15335 3179
rect 2789 3077 2823 3111
rect 1409 3009 1443 3043
rect 4997 3009 5031 3043
rect 5825 3009 5859 3043
rect 6193 3009 6227 3043
rect 7389 3009 7423 3043
rect 8217 3009 8251 3043
rect 9781 3009 9815 3043
rect 10977 3009 11011 3043
rect 11805 3009 11839 3043
rect 12909 3009 12943 3043
rect 13093 3009 13127 3043
rect 13829 3009 13863 3043
rect 3148 2941 3182 2975
rect 5998 2941 6032 2975
rect 8585 2941 8619 2975
rect 9689 2941 9723 2975
rect 10885 2941 10919 2975
rect 11621 2941 11655 2975
rect 13645 2941 13679 2975
rect 14565 2941 14599 2975
rect 15485 2941 15519 2975
rect 1676 2873 1710 2907
rect 4721 2873 4755 2907
rect 7205 2873 7239 2907
rect 7297 2873 7331 2907
rect 8125 2873 8159 2907
rect 8861 2873 8895 2907
rect 10793 2873 10827 2907
rect 11713 2873 11747 2907
rect 12817 2873 12851 2907
rect 4353 2805 4387 2839
rect 4813 2805 4847 2839
rect 5181 2805 5215 2839
rect 5549 2805 5583 2839
rect 5641 2805 5675 2839
rect 8033 2805 8067 2839
rect 9597 2805 9631 2839
rect 10425 2805 10459 2839
rect 12449 2805 12483 2839
rect 14749 2805 14783 2839
rect 2053 2601 2087 2635
rect 2881 2601 2915 2635
rect 3249 2601 3283 2635
rect 5549 2601 5583 2635
rect 6009 2601 6043 2635
rect 8677 2601 8711 2635
rect 10977 2601 11011 2635
rect 11437 2601 11471 2635
rect 7389 2533 7423 2567
rect 11345 2533 11379 2567
rect 14749 2533 14783 2567
rect 1961 2465 1995 2499
rect 4344 2465 4378 2499
rect 5917 2465 5951 2499
rect 7297 2465 7331 2499
rect 8585 2465 8619 2499
rect 9597 2465 9631 2499
rect 10149 2465 10183 2499
rect 11805 2465 11839 2499
rect 12633 2465 12667 2499
rect 13553 2465 13587 2499
rect 14473 2465 14507 2499
rect 2237 2397 2271 2431
rect 2789 2397 2823 2431
rect 3341 2397 3375 2431
rect 3433 2397 3467 2431
rect 3709 2397 3743 2431
rect 6193 2397 6227 2431
rect 7481 2397 7515 2431
rect 8769 2397 8803 2431
rect 10241 2397 10275 2431
rect 10425 2397 10459 2431
rect 11529 2397 11563 2431
rect 12817 2397 12851 2431
rect 13737 2397 13771 2431
rect 1593 2329 1627 2363
rect 8217 2329 8251 2363
rect 3617 2261 3651 2295
rect 5457 2261 5491 2295
rect 6929 2261 6963 2295
rect 9413 2261 9447 2295
rect 9781 2261 9815 2295
rect 11989 2261 12023 2295
rect 14473 2057 14507 2091
rect 6745 1853 6779 1887
rect 11713 1853 11747 1887
rect 7113 1785 7147 1819
rect 7113 1649 7147 1683
rect 11069 1785 11103 1819
rect 6745 1445 6779 1479
rect 11069 1445 11103 1479
rect 11713 1377 11747 1411
rect 14473 1377 14507 1411
rect 949 1241 983 1275
<< metal1 >>
rect 12250 18776 12256 18828
rect 12308 18816 12314 18828
rect 13906 18816 13912 18828
rect 12308 18788 13912 18816
rect 12308 18776 12314 18788
rect 13906 18776 13912 18788
rect 13964 18776 13970 18828
rect 10594 18232 10600 18284
rect 10652 18272 10658 18284
rect 11054 18272 11060 18284
rect 10652 18244 11060 18272
rect 10652 18232 10658 18244
rect 11054 18232 11060 18244
rect 11112 18232 11118 18284
rect 8294 18164 8300 18216
rect 8352 18204 8358 18216
rect 9582 18204 9588 18216
rect 8352 18176 9588 18204
rect 8352 18164 8358 18176
rect 9582 18164 9588 18176
rect 9640 18164 9646 18216
rect 10502 18164 10508 18216
rect 10560 18204 10566 18216
rect 15102 18204 15108 18216
rect 10560 18176 15108 18204
rect 10560 18164 10566 18176
rect 15102 18164 15108 18176
rect 15160 18164 15166 18216
rect 3418 18096 3424 18148
rect 3476 18136 3482 18148
rect 8846 18136 8852 18148
rect 3476 18108 8852 18136
rect 3476 18096 3482 18108
rect 8846 18096 8852 18108
rect 8904 18096 8910 18148
rect 10686 18096 10692 18148
rect 10744 18136 10750 18148
rect 11422 18136 11428 18148
rect 10744 18108 11428 18136
rect 10744 18096 10750 18108
rect 11422 18096 11428 18108
rect 11480 18096 11486 18148
rect 7466 18028 7472 18080
rect 7524 18068 7530 18080
rect 11146 18068 11152 18080
rect 7524 18040 11152 18068
rect 7524 18028 7530 18040
rect 11146 18028 11152 18040
rect 11204 18028 11210 18080
rect 3510 17960 3516 18012
rect 3568 18000 3574 18012
rect 12802 18000 12808 18012
rect 3568 17972 12808 18000
rect 3568 17960 3574 17972
rect 12802 17960 12808 17972
rect 12860 17960 12866 18012
rect 6086 17892 6092 17944
rect 6144 17932 6150 17944
rect 8938 17932 8944 17944
rect 6144 17904 8944 17932
rect 6144 17892 6150 17904
rect 8938 17892 8944 17904
rect 8996 17892 9002 17944
rect 7098 17824 7104 17876
rect 7156 17864 7162 17876
rect 9674 17864 9680 17876
rect 7156 17836 9680 17864
rect 7156 17824 7162 17836
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 7926 17756 7932 17808
rect 7984 17796 7990 17808
rect 10226 17796 10232 17808
rect 7984 17768 10232 17796
rect 7984 17756 7990 17768
rect 10226 17756 10232 17768
rect 10284 17756 10290 17808
rect 11698 17756 11704 17808
rect 11756 17796 11762 17808
rect 12342 17796 12348 17808
rect 11756 17768 12348 17796
rect 11756 17756 11762 17768
rect 12342 17756 12348 17768
rect 12400 17756 12406 17808
rect 1762 17688 1768 17740
rect 1820 17728 1826 17740
rect 12526 17728 12532 17740
rect 1820 17700 12532 17728
rect 1820 17688 1826 17700
rect 12526 17688 12532 17700
rect 12584 17688 12590 17740
rect 7006 17620 7012 17672
rect 7064 17660 7070 17672
rect 13998 17660 14004 17672
rect 7064 17632 14004 17660
rect 7064 17620 7070 17632
rect 13998 17620 14004 17632
rect 14056 17620 14062 17672
rect 566 17552 572 17604
rect 624 17592 630 17604
rect 11974 17592 11980 17604
rect 624 17564 11980 17592
rect 624 17552 630 17564
rect 11974 17552 11980 17564
rect 12032 17552 12038 17604
rect 13538 17552 13544 17604
rect 13596 17592 13602 17604
rect 14182 17592 14188 17604
rect 13596 17564 14188 17592
rect 13596 17552 13602 17564
rect 14182 17552 14188 17564
rect 14240 17552 14246 17604
rect 4982 17484 4988 17536
rect 5040 17524 5046 17536
rect 6270 17524 6276 17536
rect 5040 17496 6276 17524
rect 5040 17484 5046 17496
rect 6270 17484 6276 17496
rect 6328 17484 6334 17536
rect 6362 17484 6368 17536
rect 6420 17524 6426 17536
rect 10134 17524 10140 17536
rect 6420 17496 10140 17524
rect 6420 17484 6426 17496
rect 10134 17484 10140 17496
rect 10192 17484 10198 17536
rect 1104 17434 15824 17456
rect 1104 17382 3447 17434
rect 3499 17382 3511 17434
rect 3563 17382 3575 17434
rect 3627 17382 3639 17434
rect 3691 17382 8378 17434
rect 8430 17382 8442 17434
rect 8494 17382 8506 17434
rect 8558 17382 8570 17434
rect 8622 17382 13308 17434
rect 13360 17382 13372 17434
rect 13424 17382 13436 17434
rect 13488 17382 13500 17434
rect 13552 17382 15824 17434
rect 1104 17360 15824 17382
rect 4246 17280 4252 17332
rect 4304 17320 4310 17332
rect 11885 17323 11943 17329
rect 11885 17320 11897 17323
rect 4304 17292 11897 17320
rect 4304 17280 4310 17292
rect 11885 17289 11897 17292
rect 11931 17289 11943 17323
rect 11885 17283 11943 17289
rect 7834 17212 7840 17264
rect 7892 17252 7898 17264
rect 12805 17255 12863 17261
rect 12805 17252 12817 17255
rect 7892 17224 12817 17252
rect 7892 17212 7898 17224
rect 12805 17221 12817 17224
rect 12851 17221 12863 17255
rect 12805 17215 12863 17221
rect 5077 17187 5135 17193
rect 5077 17153 5089 17187
rect 5123 17184 5135 17187
rect 5166 17184 5172 17196
rect 5123 17156 5172 17184
rect 5123 17153 5135 17156
rect 5077 17147 5135 17153
rect 5166 17144 5172 17156
rect 5224 17144 5230 17196
rect 5258 17144 5264 17196
rect 5316 17184 5322 17196
rect 6086 17184 6092 17196
rect 5316 17156 6092 17184
rect 5316 17144 5322 17156
rect 6086 17144 6092 17156
rect 6144 17144 6150 17196
rect 6273 17187 6331 17193
rect 6273 17153 6285 17187
rect 6319 17184 6331 17187
rect 6319 17156 6592 17184
rect 6319 17153 6331 17156
rect 6273 17147 6331 17153
rect 1857 17119 1915 17125
rect 1857 17085 1869 17119
rect 1903 17085 1915 17119
rect 1857 17079 1915 17085
rect 2777 17119 2835 17125
rect 2777 17085 2789 17119
rect 2823 17116 2835 17119
rect 5350 17116 5356 17128
rect 2823 17088 5356 17116
rect 2823 17085 2835 17088
rect 2777 17079 2835 17085
rect 1872 16980 1900 17079
rect 5350 17076 5356 17088
rect 5408 17076 5414 17128
rect 6564 17116 6592 17156
rect 6638 17144 6644 17196
rect 6696 17184 6702 17196
rect 7374 17184 7380 17196
rect 6696 17156 7380 17184
rect 6696 17144 6702 17156
rect 7374 17144 7380 17156
rect 7432 17144 7438 17196
rect 7650 17144 7656 17196
rect 7708 17184 7714 17196
rect 7745 17187 7803 17193
rect 7745 17184 7757 17187
rect 7708 17156 7757 17184
rect 7708 17144 7714 17156
rect 7745 17153 7757 17156
rect 7791 17153 7803 17187
rect 7745 17147 7803 17153
rect 8018 17144 8024 17196
rect 8076 17184 8082 17196
rect 8941 17187 8999 17193
rect 8941 17184 8953 17187
rect 8076 17156 8953 17184
rect 8076 17144 8082 17156
rect 8941 17153 8953 17156
rect 8987 17153 8999 17187
rect 10410 17184 10416 17196
rect 10371 17156 10416 17184
rect 8941 17147 8999 17153
rect 10410 17144 10416 17156
rect 10468 17144 10474 17196
rect 12158 17184 12164 17196
rect 10980 17156 12164 17184
rect 7190 17116 7196 17128
rect 6564 17088 7196 17116
rect 7190 17076 7196 17088
rect 7248 17076 7254 17128
rect 7561 17119 7619 17125
rect 7561 17085 7573 17119
rect 7607 17116 7619 17119
rect 10318 17116 10324 17128
rect 7607 17088 10324 17116
rect 7607 17085 7619 17088
rect 7561 17079 7619 17085
rect 10318 17076 10324 17088
rect 10376 17076 10382 17128
rect 10980 17125 11008 17156
rect 12158 17144 12164 17156
rect 12216 17144 12222 17196
rect 13630 17184 13636 17196
rect 12636 17156 13636 17184
rect 10965 17119 11023 17125
rect 10965 17085 10977 17119
rect 11011 17085 11023 17119
rect 10965 17079 11023 17085
rect 11701 17119 11759 17125
rect 11701 17085 11713 17119
rect 11747 17116 11759 17119
rect 11790 17116 11796 17128
rect 11747 17088 11796 17116
rect 11747 17085 11759 17088
rect 11701 17079 11759 17085
rect 11790 17076 11796 17088
rect 11848 17076 11854 17128
rect 12636 17125 12664 17156
rect 13630 17144 13636 17156
rect 13688 17144 13694 17196
rect 14550 17184 14556 17196
rect 14511 17156 14556 17184
rect 14550 17144 14556 17156
rect 14608 17144 14614 17196
rect 12621 17119 12679 17125
rect 12621 17085 12633 17119
rect 12667 17085 12679 17119
rect 12621 17079 12679 17085
rect 2130 17048 2136 17060
rect 2091 17020 2136 17048
rect 2130 17008 2136 17020
rect 2188 17008 2194 17060
rect 3050 17048 3056 17060
rect 3011 17020 3056 17048
rect 3050 17008 3056 17020
rect 3108 17008 3114 17060
rect 4522 17008 4528 17060
rect 4580 17048 4586 17060
rect 4893 17051 4951 17057
rect 4893 17048 4905 17051
rect 4580 17020 4905 17048
rect 4580 17008 4586 17020
rect 4893 17017 4905 17020
rect 4939 17017 4951 17051
rect 4893 17011 4951 17017
rect 4982 17008 4988 17060
rect 5040 17048 5046 17060
rect 7653 17051 7711 17057
rect 5040 17020 6040 17048
rect 5040 17008 5046 17020
rect 4433 16983 4491 16989
rect 4433 16980 4445 16983
rect 1872 16952 4445 16980
rect 4433 16949 4445 16952
rect 4479 16949 4491 16983
rect 4798 16980 4804 16992
rect 4759 16952 4804 16980
rect 4433 16943 4491 16949
rect 4798 16940 4804 16952
rect 4856 16940 4862 16992
rect 5074 16940 5080 16992
rect 5132 16980 5138 16992
rect 6012 16989 6040 17020
rect 7653 17017 7665 17051
rect 7699 17048 7711 17051
rect 8478 17048 8484 17060
rect 7699 17020 8484 17048
rect 7699 17017 7711 17020
rect 7653 17011 7711 17017
rect 8478 17008 8484 17020
rect 8536 17008 8542 17060
rect 8662 17008 8668 17060
rect 8720 17008 8726 17060
rect 10229 17051 10287 17057
rect 10229 17017 10241 17051
rect 10275 17048 10287 17051
rect 12250 17048 12256 17060
rect 10275 17020 12256 17048
rect 10275 17017 10287 17020
rect 10229 17011 10287 17017
rect 12250 17008 12256 17020
rect 12308 17008 12314 17060
rect 12802 17008 12808 17060
rect 12860 17048 12866 17060
rect 13541 17051 13599 17057
rect 13541 17048 13553 17051
rect 12860 17020 13553 17048
rect 12860 17008 12866 17020
rect 13541 17017 13553 17020
rect 13587 17017 13599 17051
rect 13541 17011 13599 17017
rect 13633 17051 13691 17057
rect 13633 17017 13645 17051
rect 13679 17048 13691 17051
rect 13722 17048 13728 17060
rect 13679 17020 13728 17048
rect 13679 17017 13691 17020
rect 13633 17011 13691 17017
rect 13722 17008 13728 17020
rect 13780 17008 13786 17060
rect 5629 16983 5687 16989
rect 5629 16980 5641 16983
rect 5132 16952 5641 16980
rect 5132 16940 5138 16952
rect 5629 16949 5641 16952
rect 5675 16949 5687 16983
rect 5629 16943 5687 16949
rect 5997 16983 6055 16989
rect 5997 16949 6009 16983
rect 6043 16980 6055 16983
rect 6730 16980 6736 16992
rect 6043 16952 6736 16980
rect 6043 16949 6055 16952
rect 5997 16943 6055 16949
rect 6730 16940 6736 16952
rect 6788 16940 6794 16992
rect 7193 16983 7251 16989
rect 7193 16949 7205 16983
rect 7239 16980 7251 16983
rect 7466 16980 7472 16992
rect 7239 16952 7472 16980
rect 7239 16949 7251 16952
rect 7193 16943 7251 16949
rect 7466 16940 7472 16952
rect 7524 16940 7530 16992
rect 7742 16940 7748 16992
rect 7800 16980 7806 16992
rect 8389 16983 8447 16989
rect 8389 16980 8401 16983
rect 7800 16952 8401 16980
rect 7800 16940 7806 16952
rect 8389 16949 8401 16952
rect 8435 16949 8447 16983
rect 8680 16980 8708 17008
rect 8757 16983 8815 16989
rect 8757 16980 8769 16983
rect 8680 16952 8769 16980
rect 8389 16943 8447 16949
rect 8757 16949 8769 16952
rect 8803 16949 8815 16983
rect 8757 16943 8815 16949
rect 8849 16983 8907 16989
rect 8849 16949 8861 16983
rect 8895 16980 8907 16983
rect 8938 16980 8944 16992
rect 8895 16952 8944 16980
rect 8895 16949 8907 16952
rect 8849 16943 8907 16949
rect 8938 16940 8944 16952
rect 8996 16940 9002 16992
rect 9766 16980 9772 16992
rect 9727 16952 9772 16980
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 10137 16983 10195 16989
rect 10137 16949 10149 16983
rect 10183 16980 10195 16983
rect 10686 16980 10692 16992
rect 10183 16952 10692 16980
rect 10183 16949 10195 16952
rect 10137 16943 10195 16949
rect 10686 16940 10692 16952
rect 10744 16940 10750 16992
rect 11146 16980 11152 16992
rect 11107 16952 11152 16980
rect 11146 16940 11152 16952
rect 11204 16940 11210 16992
rect 1104 16890 15824 16912
rect 1104 16838 5912 16890
rect 5964 16838 5976 16890
rect 6028 16838 6040 16890
rect 6092 16838 6104 16890
rect 6156 16838 10843 16890
rect 10895 16838 10907 16890
rect 10959 16838 10971 16890
rect 11023 16838 11035 16890
rect 11087 16838 15824 16890
rect 1104 16816 15824 16838
rect 3326 16736 3332 16788
rect 3384 16776 3390 16788
rect 3421 16779 3479 16785
rect 3421 16776 3433 16779
rect 3384 16748 3433 16776
rect 3384 16736 3390 16748
rect 3421 16745 3433 16748
rect 3467 16745 3479 16779
rect 5626 16776 5632 16788
rect 3421 16739 3479 16745
rect 3620 16748 5632 16776
rect 1578 16640 1584 16652
rect 1539 16612 1584 16640
rect 1578 16600 1584 16612
rect 1636 16600 1642 16652
rect 1854 16640 1860 16652
rect 1815 16612 1860 16640
rect 1854 16600 1860 16612
rect 1912 16600 1918 16652
rect 2406 16600 2412 16652
rect 2464 16640 2470 16652
rect 2501 16643 2559 16649
rect 2501 16640 2513 16643
rect 2464 16612 2513 16640
rect 2464 16600 2470 16612
rect 2501 16609 2513 16612
rect 2547 16609 2559 16643
rect 2501 16603 2559 16609
rect 2777 16643 2835 16649
rect 2777 16609 2789 16643
rect 2823 16640 2835 16643
rect 2958 16640 2964 16652
rect 2823 16612 2964 16640
rect 2823 16609 2835 16612
rect 2777 16603 2835 16609
rect 2958 16600 2964 16612
rect 3016 16600 3022 16652
rect 3620 16649 3648 16748
rect 5626 16736 5632 16748
rect 5684 16736 5690 16788
rect 6270 16736 6276 16788
rect 6328 16776 6334 16788
rect 6365 16779 6423 16785
rect 6365 16776 6377 16779
rect 6328 16748 6377 16776
rect 6328 16736 6334 16748
rect 6365 16745 6377 16748
rect 6411 16745 6423 16779
rect 6365 16739 6423 16745
rect 6730 16736 6736 16788
rect 6788 16776 6794 16788
rect 7098 16776 7104 16788
rect 6788 16748 7104 16776
rect 6788 16736 6794 16748
rect 7098 16736 7104 16748
rect 7156 16736 7162 16788
rect 9674 16776 9680 16788
rect 9635 16748 9680 16776
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 10045 16779 10103 16785
rect 10045 16745 10057 16779
rect 10091 16776 10103 16779
rect 10134 16776 10140 16788
rect 10091 16748 10140 16776
rect 10091 16745 10103 16748
rect 10045 16739 10103 16745
rect 10134 16736 10140 16748
rect 10192 16736 10198 16788
rect 10226 16736 10232 16788
rect 10284 16776 10290 16788
rect 13265 16779 13323 16785
rect 13265 16776 13277 16779
rect 10284 16748 13277 16776
rect 10284 16736 10290 16748
rect 13265 16745 13277 16748
rect 13311 16745 13323 16779
rect 13998 16776 14004 16788
rect 13959 16748 14004 16776
rect 13265 16739 13323 16745
rect 13998 16736 14004 16748
rect 14056 16736 14062 16788
rect 7926 16708 7932 16720
rect 4264 16680 7932 16708
rect 3605 16643 3663 16649
rect 3605 16609 3617 16643
rect 3651 16609 3663 16643
rect 3605 16603 3663 16609
rect 2222 16532 2228 16584
rect 2280 16572 2286 16584
rect 4264 16572 4292 16680
rect 7926 16668 7932 16680
rect 7984 16668 7990 16720
rect 8294 16668 8300 16720
rect 8352 16708 8358 16720
rect 8573 16711 8631 16717
rect 8573 16708 8585 16711
rect 8352 16680 8585 16708
rect 8352 16668 8358 16680
rect 8573 16677 8585 16680
rect 8619 16677 8631 16711
rect 8573 16671 8631 16677
rect 11054 16668 11060 16720
rect 11112 16708 11118 16720
rect 12894 16708 12900 16720
rect 11112 16680 12900 16708
rect 11112 16668 11118 16680
rect 12894 16668 12900 16680
rect 12952 16668 12958 16720
rect 4608 16643 4666 16649
rect 4608 16609 4620 16643
rect 4654 16640 4666 16643
rect 4890 16640 4896 16652
rect 4654 16612 4896 16640
rect 4654 16609 4666 16612
rect 4608 16603 4666 16609
rect 4890 16600 4896 16612
rect 4948 16640 4954 16652
rect 6181 16643 6239 16649
rect 4948 16612 6132 16640
rect 4948 16600 4954 16612
rect 2280 16544 4292 16572
rect 2280 16532 2286 16544
rect 4338 16532 4344 16584
rect 4396 16572 4402 16584
rect 4396 16544 4441 16572
rect 4396 16532 4402 16544
rect 1394 16464 1400 16516
rect 1452 16504 1458 16516
rect 4246 16504 4252 16516
rect 1452 16476 4252 16504
rect 1452 16464 1458 16476
rect 4246 16464 4252 16476
rect 4304 16464 4310 16516
rect 5718 16504 5724 16516
rect 5679 16476 5724 16504
rect 5718 16464 5724 16476
rect 5776 16464 5782 16516
rect 6104 16504 6132 16612
rect 6181 16609 6193 16643
rect 6227 16640 6239 16643
rect 6362 16640 6368 16652
rect 6227 16612 6368 16640
rect 6227 16609 6239 16612
rect 6181 16603 6239 16609
rect 6362 16600 6368 16612
rect 6420 16600 6426 16652
rect 7282 16640 7288 16652
rect 7243 16612 7288 16640
rect 7282 16600 7288 16612
rect 7340 16600 7346 16652
rect 8110 16640 8116 16652
rect 7392 16612 8116 16640
rect 7392 16581 7420 16612
rect 8110 16600 8116 16612
rect 8168 16600 8174 16652
rect 8202 16600 8208 16652
rect 8260 16640 8266 16652
rect 8481 16643 8539 16649
rect 8481 16640 8493 16643
rect 8260 16612 8493 16640
rect 8260 16600 8266 16612
rect 8481 16609 8493 16612
rect 8527 16609 8539 16643
rect 8481 16603 8539 16609
rect 9858 16600 9864 16652
rect 9916 16640 9922 16652
rect 10137 16643 10195 16649
rect 10137 16640 10149 16643
rect 9916 16612 10149 16640
rect 9916 16600 9922 16612
rect 10137 16609 10149 16612
rect 10183 16609 10195 16643
rect 10137 16603 10195 16609
rect 10778 16600 10784 16652
rect 10836 16640 10842 16652
rect 10873 16643 10931 16649
rect 10873 16640 10885 16643
rect 10836 16612 10885 16640
rect 10836 16600 10842 16612
rect 10873 16609 10885 16612
rect 10919 16609 10931 16643
rect 10873 16603 10931 16609
rect 11146 16600 11152 16652
rect 11204 16640 11210 16652
rect 11609 16643 11667 16649
rect 11609 16640 11621 16643
rect 11204 16612 11621 16640
rect 11204 16600 11210 16612
rect 11609 16609 11621 16612
rect 11655 16609 11667 16643
rect 12342 16640 12348 16652
rect 12303 16612 12348 16640
rect 11609 16603 11667 16609
rect 12342 16600 12348 16612
rect 12400 16600 12406 16652
rect 13078 16640 13084 16652
rect 13039 16612 13084 16640
rect 13078 16600 13084 16612
rect 13136 16600 13142 16652
rect 13817 16643 13875 16649
rect 13817 16609 13829 16643
rect 13863 16640 13875 16643
rect 13906 16640 13912 16652
rect 13863 16612 13912 16640
rect 13863 16609 13875 16612
rect 13817 16603 13875 16609
rect 13906 16600 13912 16612
rect 13964 16600 13970 16652
rect 14274 16600 14280 16652
rect 14332 16640 14338 16652
rect 14553 16643 14611 16649
rect 14553 16640 14565 16643
rect 14332 16612 14565 16640
rect 14332 16600 14338 16612
rect 14553 16609 14565 16612
rect 14599 16609 14611 16643
rect 14553 16603 14611 16609
rect 7377 16575 7435 16581
rect 7377 16541 7389 16575
rect 7423 16541 7435 16575
rect 7377 16535 7435 16541
rect 7469 16575 7527 16581
rect 7469 16541 7481 16575
rect 7515 16541 7527 16575
rect 7469 16535 7527 16541
rect 7484 16504 7512 16535
rect 7926 16532 7932 16584
rect 7984 16572 7990 16584
rect 8665 16575 8723 16581
rect 8665 16572 8677 16575
rect 7984 16544 8677 16572
rect 7984 16532 7990 16544
rect 8665 16541 8677 16544
rect 8711 16541 8723 16575
rect 8665 16535 8723 16541
rect 9306 16532 9312 16584
rect 9364 16572 9370 16584
rect 10226 16572 10232 16584
rect 9364 16544 10232 16572
rect 9364 16532 9370 16544
rect 10226 16532 10232 16544
rect 10284 16532 10290 16584
rect 10321 16575 10379 16581
rect 10321 16541 10333 16575
rect 10367 16572 10379 16575
rect 10410 16572 10416 16584
rect 10367 16544 10416 16572
rect 10367 16541 10379 16544
rect 10321 16535 10379 16541
rect 10410 16532 10416 16544
rect 10468 16532 10474 16584
rect 12802 16572 12808 16584
rect 10612 16544 10815 16572
rect 6104 16476 8248 16504
rect 2222 16396 2228 16448
rect 2280 16436 2286 16448
rect 6730 16436 6736 16448
rect 2280 16408 6736 16436
rect 2280 16396 2286 16408
rect 6730 16396 6736 16408
rect 6788 16396 6794 16448
rect 6914 16436 6920 16448
rect 6875 16408 6920 16436
rect 6914 16396 6920 16408
rect 6972 16396 6978 16448
rect 7006 16396 7012 16448
rect 7064 16436 7070 16448
rect 8113 16439 8171 16445
rect 8113 16436 8125 16439
rect 7064 16408 8125 16436
rect 7064 16396 7070 16408
rect 8113 16405 8125 16408
rect 8159 16405 8171 16439
rect 8220 16436 8248 16476
rect 8846 16464 8852 16516
rect 8904 16504 8910 16516
rect 10612 16504 10640 16544
rect 8904 16476 10640 16504
rect 10787 16504 10815 16544
rect 11532 16544 12808 16572
rect 11532 16504 11560 16544
rect 12802 16532 12808 16544
rect 12860 16532 12866 16584
rect 10787 16476 11560 16504
rect 11793 16507 11851 16513
rect 8904 16464 8910 16476
rect 11793 16473 11805 16507
rect 11839 16504 11851 16507
rect 11974 16504 11980 16516
rect 11839 16476 11980 16504
rect 11839 16473 11851 16476
rect 11793 16467 11851 16473
rect 11974 16464 11980 16476
rect 12032 16464 12038 16516
rect 12526 16504 12532 16516
rect 12487 16476 12532 16504
rect 12526 16464 12532 16476
rect 12584 16464 12590 16516
rect 10410 16436 10416 16448
rect 8220 16408 10416 16436
rect 8113 16399 8171 16405
rect 10410 16396 10416 16408
rect 10468 16396 10474 16448
rect 10870 16396 10876 16448
rect 10928 16436 10934 16448
rect 11057 16439 11115 16445
rect 11057 16436 11069 16439
rect 10928 16408 11069 16436
rect 10928 16396 10934 16408
rect 11057 16405 11069 16408
rect 11103 16405 11115 16439
rect 11057 16399 11115 16405
rect 1104 16346 15824 16368
rect 1104 16294 3447 16346
rect 3499 16294 3511 16346
rect 3563 16294 3575 16346
rect 3627 16294 3639 16346
rect 3691 16294 8378 16346
rect 8430 16294 8442 16346
rect 8494 16294 8506 16346
rect 8558 16294 8570 16346
rect 8622 16294 13308 16346
rect 13360 16294 13372 16346
rect 13424 16294 13436 16346
rect 13488 16294 13500 16346
rect 13552 16294 15824 16346
rect 1104 16272 15824 16294
rect 1581 16235 1639 16241
rect 1581 16201 1593 16235
rect 1627 16232 1639 16235
rect 2866 16232 2872 16244
rect 1627 16204 2872 16232
rect 1627 16201 1639 16204
rect 1581 16195 1639 16201
rect 2866 16192 2872 16204
rect 2924 16192 2930 16244
rect 3145 16235 3203 16241
rect 3145 16201 3157 16235
rect 3191 16232 3203 16235
rect 3191 16204 4568 16232
rect 3191 16201 3203 16204
rect 3145 16195 3203 16201
rect 198 16124 204 16176
rect 256 16164 262 16176
rect 4062 16164 4068 16176
rect 256 16136 4068 16164
rect 256 16124 262 16136
rect 4062 16124 4068 16136
rect 4120 16124 4126 16176
rect 4540 16164 4568 16204
rect 4614 16192 4620 16244
rect 4672 16232 4678 16244
rect 6917 16235 6975 16241
rect 4672 16204 6500 16232
rect 4672 16192 4678 16204
rect 4706 16164 4712 16176
rect 4540 16136 4712 16164
rect 4706 16124 4712 16136
rect 4764 16124 4770 16176
rect 4982 16164 4988 16176
rect 4816 16136 4988 16164
rect 2501 16099 2559 16105
rect 2501 16065 2513 16099
rect 2547 16096 2559 16099
rect 2774 16096 2780 16108
rect 2547 16068 2780 16096
rect 2547 16065 2559 16068
rect 2501 16059 2559 16065
rect 2774 16056 2780 16068
rect 2832 16056 2838 16108
rect 3789 16099 3847 16105
rect 3789 16065 3801 16099
rect 3835 16096 3847 16099
rect 3970 16096 3976 16108
rect 3835 16068 3976 16096
rect 3835 16065 3847 16068
rect 3789 16059 3847 16065
rect 3970 16056 3976 16068
rect 4028 16056 4034 16108
rect 4154 16056 4160 16108
rect 4212 16096 4218 16108
rect 4816 16105 4844 16136
rect 4982 16124 4988 16136
rect 5040 16124 5046 16176
rect 5537 16167 5595 16173
rect 5537 16133 5549 16167
rect 5583 16133 5595 16167
rect 6472 16164 6500 16204
rect 6917 16201 6929 16235
rect 6963 16232 6975 16235
rect 6963 16204 8432 16232
rect 6963 16201 6975 16204
rect 6917 16195 6975 16201
rect 8297 16167 8355 16173
rect 8297 16164 8309 16167
rect 6472 16136 8309 16164
rect 5537 16127 5595 16133
rect 8297 16133 8309 16136
rect 8343 16133 8355 16167
rect 8297 16127 8355 16133
rect 4801 16099 4859 16105
rect 4801 16096 4813 16099
rect 4212 16068 4813 16096
rect 4212 16056 4218 16068
rect 4801 16065 4813 16068
rect 4847 16065 4859 16099
rect 4801 16059 4859 16065
rect 4890 16056 4896 16108
rect 4948 16096 4954 16108
rect 4948 16068 4993 16096
rect 4948 16056 4954 16068
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 15997 1455 16031
rect 1397 15991 1455 15997
rect 1412 15960 1440 15991
rect 1670 15988 1676 16040
rect 1728 16028 1734 16040
rect 2225 16031 2283 16037
rect 1728 16000 2176 16028
rect 1728 15988 1734 16000
rect 2148 15960 2176 16000
rect 2225 15997 2237 16031
rect 2271 16028 2283 16031
rect 5552 16028 5580 16127
rect 6181 16099 6239 16105
rect 6181 16065 6193 16099
rect 6227 16096 6239 16099
rect 6730 16096 6736 16108
rect 6227 16068 6736 16096
rect 6227 16065 6239 16068
rect 6181 16059 6239 16065
rect 6730 16056 6736 16068
rect 6788 16056 6794 16108
rect 7098 16056 7104 16108
rect 7156 16096 7162 16108
rect 7469 16099 7527 16105
rect 7469 16096 7481 16099
rect 7156 16068 7481 16096
rect 7156 16056 7162 16068
rect 7469 16065 7481 16068
rect 7515 16096 7527 16099
rect 8404 16096 8432 16204
rect 9582 16192 9588 16244
rect 9640 16232 9646 16244
rect 11238 16232 11244 16244
rect 9640 16204 11244 16232
rect 9640 16192 9646 16204
rect 11238 16192 11244 16204
rect 11296 16192 11302 16244
rect 11330 16192 11336 16244
rect 11388 16232 11394 16244
rect 13817 16235 13875 16241
rect 13817 16232 13829 16235
rect 11388 16204 13829 16232
rect 11388 16192 11394 16204
rect 13817 16201 13829 16204
rect 13863 16201 13875 16235
rect 13817 16195 13875 16201
rect 9674 16124 9680 16176
rect 9732 16164 9738 16176
rect 11793 16167 11851 16173
rect 11793 16164 11805 16167
rect 9732 16136 11805 16164
rect 9732 16124 9738 16136
rect 11793 16133 11805 16136
rect 11839 16133 11851 16167
rect 13265 16167 13323 16173
rect 13265 16164 13277 16167
rect 11793 16127 11851 16133
rect 12452 16136 13277 16164
rect 8846 16096 8852 16108
rect 7515 16068 8340 16096
rect 8404 16068 8852 16096
rect 7515 16065 7527 16068
rect 7469 16059 7527 16065
rect 2271 16000 5580 16028
rect 5997 16031 6055 16037
rect 2271 15997 2283 16000
rect 2225 15991 2283 15997
rect 5997 15997 6009 16031
rect 6043 16028 6055 16031
rect 7742 16028 7748 16040
rect 6043 16000 7748 16028
rect 6043 15997 6055 16000
rect 5997 15991 6055 15997
rect 7742 15988 7748 16000
rect 7800 15988 7806 16040
rect 7834 15988 7840 16040
rect 7892 16028 7898 16040
rect 8113 16031 8171 16037
rect 8113 16028 8125 16031
rect 7892 16000 8125 16028
rect 7892 15988 7898 16000
rect 8113 15997 8125 16000
rect 8159 15997 8171 16031
rect 8312 16028 8340 16068
rect 8846 16056 8852 16068
rect 8904 16056 8910 16108
rect 9306 16056 9312 16108
rect 9364 16096 9370 16108
rect 9769 16099 9827 16105
rect 9769 16096 9781 16099
rect 9364 16068 9781 16096
rect 9364 16056 9370 16068
rect 9769 16065 9781 16068
rect 9815 16065 9827 16099
rect 9769 16059 9827 16065
rect 9950 16056 9956 16108
rect 10008 16096 10014 16108
rect 10318 16096 10324 16108
rect 10008 16068 10324 16096
rect 10008 16056 10014 16068
rect 10318 16056 10324 16068
rect 10376 16056 10382 16108
rect 10410 16056 10416 16108
rect 10468 16096 10474 16108
rect 11057 16099 11115 16105
rect 11057 16096 11069 16099
rect 10468 16068 11069 16096
rect 10468 16056 10474 16068
rect 11057 16065 11069 16068
rect 11103 16096 11115 16099
rect 11103 16068 12020 16096
rect 11103 16065 11115 16068
rect 11057 16059 11115 16065
rect 8938 16028 8944 16040
rect 8312 16000 8944 16028
rect 8113 15991 8171 15997
rect 8938 15988 8944 16000
rect 8996 15988 9002 16040
rect 9033 16031 9091 16037
rect 9033 15997 9045 16031
rect 9079 16028 9091 16031
rect 9490 16028 9496 16040
rect 9079 16000 9496 16028
rect 9079 15997 9091 16000
rect 9033 15991 9091 15997
rect 9490 15988 9496 16000
rect 9548 15988 9554 16040
rect 9585 16031 9643 16037
rect 9585 15997 9597 16031
rect 9631 16028 9643 16031
rect 11609 16031 11667 16037
rect 9631 16000 11560 16028
rect 9631 15997 9643 16000
rect 9585 15991 9643 15997
rect 5442 15960 5448 15972
rect 1412 15932 2084 15960
rect 2148 15932 5448 15960
rect 2056 15892 2084 15932
rect 5442 15920 5448 15932
rect 5500 15920 5506 15972
rect 5905 15963 5963 15969
rect 5905 15929 5917 15963
rect 5951 15960 5963 15963
rect 7190 15960 7196 15972
rect 5951 15932 7196 15960
rect 5951 15929 5963 15932
rect 5905 15923 5963 15929
rect 7190 15920 7196 15932
rect 7248 15920 7254 15972
rect 7377 15963 7435 15969
rect 7377 15929 7389 15963
rect 7423 15960 7435 15963
rect 8662 15960 8668 15972
rect 7423 15932 8668 15960
rect 7423 15929 7435 15932
rect 7377 15923 7435 15929
rect 8662 15920 8668 15932
rect 8720 15920 8726 15972
rect 8772 15932 9812 15960
rect 3142 15892 3148 15904
rect 2056 15864 3148 15892
rect 3142 15852 3148 15864
rect 3200 15852 3206 15904
rect 3510 15892 3516 15904
rect 3471 15864 3516 15892
rect 3510 15852 3516 15864
rect 3568 15852 3574 15904
rect 3605 15895 3663 15901
rect 3605 15861 3617 15895
rect 3651 15892 3663 15895
rect 3878 15892 3884 15904
rect 3651 15864 3884 15892
rect 3651 15861 3663 15864
rect 3605 15855 3663 15861
rect 3878 15852 3884 15864
rect 3936 15852 3942 15904
rect 4338 15892 4344 15904
rect 4299 15864 4344 15892
rect 4338 15852 4344 15864
rect 4396 15852 4402 15904
rect 4709 15895 4767 15901
rect 4709 15861 4721 15895
rect 4755 15892 4767 15895
rect 6270 15892 6276 15904
rect 4755 15864 6276 15892
rect 4755 15861 4767 15864
rect 4709 15855 4767 15861
rect 6270 15852 6276 15864
rect 6328 15852 6334 15904
rect 7285 15895 7343 15901
rect 7285 15861 7297 15895
rect 7331 15892 7343 15895
rect 8772 15892 8800 15932
rect 7331 15864 8800 15892
rect 8849 15895 8907 15901
rect 7331 15861 7343 15864
rect 7285 15855 7343 15861
rect 8849 15861 8861 15895
rect 8895 15892 8907 15895
rect 9030 15892 9036 15904
rect 8895 15864 9036 15892
rect 8895 15861 8907 15864
rect 8849 15855 8907 15861
rect 9030 15852 9036 15864
rect 9088 15852 9094 15904
rect 9214 15892 9220 15904
rect 9175 15864 9220 15892
rect 9214 15852 9220 15864
rect 9272 15852 9278 15904
rect 9582 15852 9588 15904
rect 9640 15892 9646 15904
rect 9677 15895 9735 15901
rect 9677 15892 9689 15895
rect 9640 15864 9689 15892
rect 9640 15852 9646 15864
rect 9677 15861 9689 15864
rect 9723 15861 9735 15895
rect 9784 15892 9812 15932
rect 10042 15920 10048 15972
rect 10100 15960 10106 15972
rect 10778 15960 10784 15972
rect 10100 15932 10784 15960
rect 10100 15920 10106 15932
rect 10778 15920 10784 15932
rect 10836 15920 10842 15972
rect 11054 15960 11060 15972
rect 10888 15932 11060 15960
rect 10226 15892 10232 15904
rect 9784 15864 10232 15892
rect 9677 15855 9735 15861
rect 10226 15852 10232 15864
rect 10284 15852 10290 15904
rect 10410 15892 10416 15904
rect 10371 15864 10416 15892
rect 10410 15852 10416 15864
rect 10468 15852 10474 15904
rect 10686 15852 10692 15904
rect 10744 15892 10750 15904
rect 10888 15901 10916 15932
rect 11054 15920 11060 15932
rect 11112 15920 11118 15972
rect 10873 15895 10931 15901
rect 10873 15892 10885 15895
rect 10744 15864 10885 15892
rect 10744 15852 10750 15864
rect 10873 15861 10885 15864
rect 10919 15861 10931 15895
rect 11532 15892 11560 16000
rect 11609 15997 11621 16031
rect 11655 16028 11667 16031
rect 11882 16028 11888 16040
rect 11655 16000 11888 16028
rect 11655 15997 11667 16000
rect 11609 15991 11667 15997
rect 11882 15988 11888 16000
rect 11940 15988 11946 16040
rect 11992 16028 12020 16068
rect 12066 16056 12072 16108
rect 12124 16096 12130 16108
rect 12452 16105 12480 16136
rect 13265 16133 13277 16136
rect 13311 16133 13323 16167
rect 13265 16127 13323 16133
rect 12437 16099 12495 16105
rect 12437 16096 12449 16099
rect 12124 16068 12449 16096
rect 12124 16056 12130 16068
rect 12437 16065 12449 16068
rect 12483 16065 12495 16099
rect 12437 16059 12495 16065
rect 14921 16099 14979 16105
rect 14921 16065 14933 16099
rect 14967 16096 14979 16099
rect 16758 16096 16764 16108
rect 14967 16068 16764 16096
rect 14967 16065 14979 16068
rect 14921 16059 14979 16065
rect 16758 16056 16764 16068
rect 16816 16056 16822 16108
rect 12526 16028 12532 16040
rect 11992 16000 12532 16028
rect 12526 15988 12532 16000
rect 12584 15988 12590 16040
rect 12805 16031 12863 16037
rect 12805 15997 12817 16031
rect 12851 16028 12863 16031
rect 12894 16028 12900 16040
rect 12851 16000 12900 16028
rect 12851 15997 12863 16000
rect 12805 15991 12863 15997
rect 12894 15988 12900 16000
rect 12952 15988 12958 16040
rect 12986 15988 12992 16040
rect 13044 16028 13050 16040
rect 13633 16031 13691 16037
rect 13633 16028 13645 16031
rect 13044 16000 13645 16028
rect 13044 15988 13050 16000
rect 13633 15997 13645 16000
rect 13679 15997 13691 16031
rect 13633 15991 13691 15997
rect 14550 15988 14556 16040
rect 14608 16028 14614 16040
rect 14645 16031 14703 16037
rect 14645 16028 14657 16031
rect 14608 16000 14657 16028
rect 14608 15988 14614 16000
rect 14645 15997 14657 16000
rect 14691 15997 14703 16031
rect 14645 15991 14703 15997
rect 11974 15920 11980 15972
rect 12032 15960 12038 15972
rect 13173 15963 13231 15969
rect 13173 15960 13185 15963
rect 12032 15932 13185 15960
rect 12032 15920 12038 15932
rect 13173 15929 13185 15932
rect 13219 15960 13231 15963
rect 13722 15960 13728 15972
rect 13219 15932 13728 15960
rect 13219 15929 13231 15932
rect 13173 15923 13231 15929
rect 13722 15920 13728 15932
rect 13780 15920 13786 15972
rect 14918 15892 14924 15904
rect 11532 15864 14924 15892
rect 10873 15855 10931 15861
rect 14918 15852 14924 15864
rect 14976 15852 14982 15904
rect 1104 15802 15824 15824
rect 1104 15750 5912 15802
rect 5964 15750 5976 15802
rect 6028 15750 6040 15802
rect 6092 15750 6104 15802
rect 6156 15750 10843 15802
rect 10895 15750 10907 15802
rect 10959 15750 10971 15802
rect 11023 15750 11035 15802
rect 11087 15750 15824 15802
rect 1104 15728 15824 15750
rect 2774 15648 2780 15700
rect 2832 15688 2838 15700
rect 3145 15691 3203 15697
rect 2832 15660 2877 15688
rect 2832 15648 2838 15660
rect 3145 15657 3157 15691
rect 3191 15688 3203 15691
rect 5534 15688 5540 15700
rect 3191 15660 5540 15688
rect 3191 15657 3203 15660
rect 3145 15651 3203 15657
rect 5534 15648 5540 15660
rect 5592 15648 5598 15700
rect 5721 15691 5779 15697
rect 5721 15657 5733 15691
rect 5767 15688 5779 15691
rect 5767 15660 7144 15688
rect 5767 15657 5779 15660
rect 5721 15651 5779 15657
rect 934 15580 940 15632
rect 992 15620 998 15632
rect 6822 15620 6828 15632
rect 992 15592 6828 15620
rect 992 15580 998 15592
rect 6822 15580 6828 15592
rect 6880 15580 6886 15632
rect 6917 15623 6975 15629
rect 6917 15589 6929 15623
rect 6963 15620 6975 15623
rect 7006 15620 7012 15632
rect 6963 15592 7012 15620
rect 6963 15589 6975 15592
rect 6917 15583 6975 15589
rect 7006 15580 7012 15592
rect 7064 15580 7070 15632
rect 7116 15620 7144 15660
rect 7190 15648 7196 15700
rect 7248 15688 7254 15700
rect 7745 15691 7803 15697
rect 7745 15688 7757 15691
rect 7248 15660 7757 15688
rect 7248 15648 7254 15660
rect 7745 15657 7757 15660
rect 7791 15657 7803 15691
rect 7745 15651 7803 15657
rect 8113 15691 8171 15697
rect 8113 15657 8125 15691
rect 8159 15688 8171 15691
rect 9677 15691 9735 15697
rect 9677 15688 9689 15691
rect 8159 15660 9689 15688
rect 8159 15657 8171 15660
rect 8113 15651 8171 15657
rect 9677 15657 9689 15660
rect 9723 15657 9735 15691
rect 9677 15651 9735 15657
rect 10318 15648 10324 15700
rect 10376 15688 10382 15700
rect 10873 15691 10931 15697
rect 10873 15688 10885 15691
rect 10376 15660 10885 15688
rect 10376 15648 10382 15660
rect 10873 15657 10885 15660
rect 10919 15657 10931 15691
rect 10873 15651 10931 15657
rect 11333 15691 11391 15697
rect 11333 15657 11345 15691
rect 11379 15688 11391 15691
rect 11882 15688 11888 15700
rect 11379 15660 11888 15688
rect 11379 15657 11391 15660
rect 11333 15651 11391 15657
rect 11882 15648 11888 15660
rect 11940 15648 11946 15700
rect 12437 15691 12495 15697
rect 12437 15688 12449 15691
rect 11992 15660 12449 15688
rect 10778 15620 10784 15632
rect 7116 15592 10784 15620
rect 10778 15580 10784 15592
rect 10836 15580 10842 15632
rect 10962 15580 10968 15632
rect 11020 15620 11026 15632
rect 11992 15620 12020 15660
rect 12437 15657 12449 15660
rect 12483 15657 12495 15691
rect 12437 15651 12495 15657
rect 12802 15648 12808 15700
rect 12860 15688 12866 15700
rect 13449 15691 13507 15697
rect 13449 15688 13461 15691
rect 12860 15660 13461 15688
rect 12860 15648 12866 15660
rect 13449 15657 13461 15660
rect 13495 15657 13507 15691
rect 13449 15651 13507 15657
rect 11020 15592 12020 15620
rect 11020 15580 11026 15592
rect 12066 15580 12072 15632
rect 12124 15620 12130 15632
rect 12710 15620 12716 15632
rect 12124 15592 12716 15620
rect 12124 15580 12130 15592
rect 12710 15580 12716 15592
rect 12768 15580 12774 15632
rect 1857 15555 1915 15561
rect 1857 15521 1869 15555
rect 1903 15552 1915 15555
rect 2314 15552 2320 15564
rect 1903 15524 2320 15552
rect 1903 15521 1915 15524
rect 1857 15515 1915 15521
rect 2314 15512 2320 15524
rect 2372 15512 2378 15564
rect 3237 15555 3295 15561
rect 3237 15521 3249 15555
rect 3283 15552 3295 15555
rect 3418 15552 3424 15564
rect 3283 15524 3424 15552
rect 3283 15521 3295 15524
rect 3237 15515 3295 15521
rect 3418 15512 3424 15524
rect 3476 15512 3482 15564
rect 4525 15555 4583 15561
rect 4525 15521 4537 15555
rect 4571 15552 4583 15555
rect 5442 15552 5448 15564
rect 4571 15524 5448 15552
rect 4571 15521 4583 15524
rect 4525 15515 4583 15521
rect 5442 15512 5448 15524
rect 5500 15512 5506 15564
rect 5813 15555 5871 15561
rect 5813 15521 5825 15555
rect 5859 15552 5871 15555
rect 7650 15552 7656 15564
rect 5859 15524 7656 15552
rect 5859 15521 5871 15524
rect 5813 15515 5871 15521
rect 7650 15512 7656 15524
rect 7708 15512 7714 15564
rect 8754 15512 8760 15564
rect 8812 15552 8818 15564
rect 10045 15555 10103 15561
rect 10045 15552 10057 15555
rect 8812 15524 10057 15552
rect 8812 15512 8818 15524
rect 10045 15521 10057 15524
rect 10091 15521 10103 15555
rect 10045 15515 10103 15521
rect 10137 15555 10195 15561
rect 10137 15521 10149 15555
rect 10183 15552 10195 15555
rect 10502 15552 10508 15564
rect 10183 15524 10508 15552
rect 10183 15521 10195 15524
rect 10137 15515 10195 15521
rect 10502 15512 10508 15524
rect 10560 15512 10566 15564
rect 11241 15555 11299 15561
rect 11241 15521 11253 15555
rect 11287 15521 11299 15555
rect 11241 15515 11299 15521
rect 12360 15524 12756 15552
rect 2133 15487 2191 15493
rect 2133 15453 2145 15487
rect 2179 15453 2191 15487
rect 2133 15447 2191 15453
rect 3329 15487 3387 15493
rect 3329 15453 3341 15487
rect 3375 15453 3387 15487
rect 3329 15447 3387 15453
rect 2148 15348 2176 15447
rect 2774 15376 2780 15428
rect 2832 15416 2838 15428
rect 3344 15416 3372 15447
rect 3786 15444 3792 15496
rect 3844 15484 3850 15496
rect 4062 15484 4068 15496
rect 3844 15456 4068 15484
rect 3844 15444 3850 15456
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 4614 15484 4620 15496
rect 4575 15456 4620 15484
rect 4614 15444 4620 15456
rect 4672 15444 4678 15496
rect 4706 15444 4712 15496
rect 4764 15484 4770 15496
rect 4764 15456 4809 15484
rect 4764 15444 4770 15456
rect 4890 15444 4896 15496
rect 4948 15484 4954 15496
rect 5905 15487 5963 15493
rect 5905 15484 5917 15487
rect 4948 15456 5917 15484
rect 4948 15444 4954 15456
rect 5905 15453 5917 15456
rect 5951 15453 5963 15487
rect 5905 15447 5963 15453
rect 7009 15487 7067 15493
rect 7009 15453 7021 15487
rect 7055 15453 7067 15487
rect 7190 15484 7196 15496
rect 7151 15456 7196 15484
rect 7009 15447 7067 15453
rect 2832 15388 3372 15416
rect 2832 15376 2838 15388
rect 5442 15376 5448 15428
rect 5500 15416 5506 15428
rect 6822 15416 6828 15428
rect 5500 15388 6828 15416
rect 5500 15376 5506 15388
rect 6822 15376 6828 15388
rect 6880 15376 6886 15428
rect 7024 15416 7052 15447
rect 7190 15444 7196 15456
rect 7248 15444 7254 15496
rect 8110 15444 8116 15496
rect 8168 15484 8174 15496
rect 8205 15487 8263 15493
rect 8205 15484 8217 15487
rect 8168 15456 8217 15484
rect 8168 15444 8174 15456
rect 8205 15453 8217 15456
rect 8251 15453 8263 15487
rect 8205 15447 8263 15453
rect 8297 15487 8355 15493
rect 8297 15453 8309 15487
rect 8343 15453 8355 15487
rect 8297 15447 8355 15453
rect 8941 15487 8999 15493
rect 8941 15453 8953 15487
rect 8987 15484 8999 15487
rect 9398 15484 9404 15496
rect 8987 15456 9404 15484
rect 8987 15453 8999 15456
rect 8941 15447 8999 15453
rect 7834 15416 7840 15428
rect 7024 15388 7840 15416
rect 7834 15376 7840 15388
rect 7892 15376 7898 15428
rect 8018 15376 8024 15428
rect 8076 15416 8082 15428
rect 8312 15416 8340 15447
rect 9398 15444 9404 15456
rect 9456 15444 9462 15496
rect 9674 15444 9680 15496
rect 9732 15484 9738 15496
rect 10229 15487 10287 15493
rect 10229 15484 10241 15487
rect 9732 15456 10241 15484
rect 9732 15444 9738 15456
rect 10229 15453 10241 15456
rect 10275 15453 10287 15487
rect 10229 15447 10287 15453
rect 10318 15444 10324 15496
rect 10376 15484 10382 15496
rect 10686 15484 10692 15496
rect 10376 15456 10692 15484
rect 10376 15444 10382 15456
rect 10686 15444 10692 15456
rect 10744 15444 10750 15496
rect 8076 15388 8340 15416
rect 8076 15376 8082 15388
rect 9122 15376 9128 15428
rect 9180 15416 9186 15428
rect 10502 15416 10508 15428
rect 9180 15388 10508 15416
rect 9180 15376 9186 15388
rect 10502 15376 10508 15388
rect 10560 15416 10566 15428
rect 11256 15416 11284 15515
rect 12360 15496 12388 15524
rect 11330 15444 11336 15496
rect 11388 15484 11394 15496
rect 11517 15487 11575 15493
rect 11517 15484 11529 15487
rect 11388 15456 11529 15484
rect 11388 15444 11394 15456
rect 11517 15453 11529 15456
rect 11563 15453 11575 15487
rect 11974 15484 11980 15496
rect 11517 15447 11575 15453
rect 11624 15456 11980 15484
rect 10560 15388 11284 15416
rect 10560 15376 10566 15388
rect 3142 15348 3148 15360
rect 2148 15320 3148 15348
rect 3142 15308 3148 15320
rect 3200 15308 3206 15360
rect 4062 15308 4068 15360
rect 4120 15348 4126 15360
rect 4157 15351 4215 15357
rect 4157 15348 4169 15351
rect 4120 15320 4169 15348
rect 4120 15308 4126 15320
rect 4157 15317 4169 15320
rect 4203 15317 4215 15351
rect 4157 15311 4215 15317
rect 5350 15308 5356 15360
rect 5408 15348 5414 15360
rect 5408 15320 5453 15348
rect 5408 15308 5414 15320
rect 5534 15308 5540 15360
rect 5592 15348 5598 15360
rect 6549 15351 6607 15357
rect 6549 15348 6561 15351
rect 5592 15320 6561 15348
rect 5592 15308 5598 15320
rect 6549 15317 6561 15320
rect 6595 15317 6607 15351
rect 6549 15311 6607 15317
rect 7374 15308 7380 15360
rect 7432 15348 7438 15360
rect 7926 15348 7932 15360
rect 7432 15320 7932 15348
rect 7432 15308 7438 15320
rect 7926 15308 7932 15320
rect 7984 15308 7990 15360
rect 8938 15308 8944 15360
rect 8996 15348 9002 15360
rect 9674 15348 9680 15360
rect 8996 15320 9680 15348
rect 8996 15308 9002 15320
rect 9674 15308 9680 15320
rect 9732 15308 9738 15360
rect 10042 15308 10048 15360
rect 10100 15348 10106 15360
rect 11624 15348 11652 15456
rect 11974 15444 11980 15456
rect 12032 15444 12038 15496
rect 12342 15444 12348 15496
rect 12400 15444 12406 15496
rect 12529 15487 12587 15493
rect 12529 15453 12541 15487
rect 12575 15484 12587 15487
rect 12618 15484 12624 15496
rect 12575 15456 12624 15484
rect 12575 15453 12587 15456
rect 12529 15447 12587 15453
rect 12618 15444 12624 15456
rect 12676 15444 12682 15496
rect 12728 15493 12756 15524
rect 13078 15512 13084 15564
rect 13136 15552 13142 15564
rect 13265 15555 13323 15561
rect 13265 15552 13277 15555
rect 13136 15524 13277 15552
rect 13136 15512 13142 15524
rect 13265 15521 13277 15524
rect 13311 15521 13323 15555
rect 13265 15515 13323 15521
rect 14001 15555 14059 15561
rect 14001 15521 14013 15555
rect 14047 15552 14059 15555
rect 15010 15552 15016 15564
rect 14047 15524 15016 15552
rect 14047 15521 14059 15524
rect 14001 15515 14059 15521
rect 15010 15512 15016 15524
rect 15068 15512 15074 15564
rect 12713 15487 12771 15493
rect 12713 15453 12725 15487
rect 12759 15484 12771 15487
rect 13170 15484 13176 15496
rect 12759 15456 13176 15484
rect 12759 15453 12771 15456
rect 12713 15447 12771 15453
rect 13170 15444 13176 15456
rect 13228 15444 13234 15496
rect 13722 15444 13728 15496
rect 13780 15484 13786 15496
rect 15470 15484 15476 15496
rect 13780 15456 15476 15484
rect 13780 15444 13786 15456
rect 15470 15444 15476 15456
rect 15528 15444 15534 15496
rect 11790 15376 11796 15428
rect 11848 15416 11854 15428
rect 14185 15419 14243 15425
rect 14185 15416 14197 15419
rect 11848 15388 14197 15416
rect 11848 15376 11854 15388
rect 14185 15385 14197 15388
rect 14231 15385 14243 15419
rect 14185 15379 14243 15385
rect 10100 15320 11652 15348
rect 10100 15308 10106 15320
rect 11974 15308 11980 15360
rect 12032 15348 12038 15360
rect 12069 15351 12127 15357
rect 12069 15348 12081 15351
rect 12032 15320 12081 15348
rect 12032 15308 12038 15320
rect 12069 15317 12081 15320
rect 12115 15317 12127 15351
rect 12069 15311 12127 15317
rect 13722 15308 13728 15360
rect 13780 15348 13786 15360
rect 14366 15348 14372 15360
rect 13780 15320 14372 15348
rect 13780 15308 13786 15320
rect 14366 15308 14372 15320
rect 14424 15308 14430 15360
rect 1104 15258 15824 15280
rect 1104 15206 3447 15258
rect 3499 15206 3511 15258
rect 3563 15206 3575 15258
rect 3627 15206 3639 15258
rect 3691 15206 8378 15258
rect 8430 15206 8442 15258
rect 8494 15206 8506 15258
rect 8558 15206 8570 15258
rect 8622 15206 13308 15258
rect 13360 15206 13372 15258
rect 13424 15206 13436 15258
rect 13488 15206 13500 15258
rect 13552 15206 15824 15258
rect 1104 15184 15824 15206
rect 3786 15144 3792 15156
rect 2424 15116 3792 15144
rect 2424 15017 2452 15116
rect 3786 15104 3792 15116
rect 3844 15104 3850 15156
rect 4338 15104 4344 15156
rect 4396 15144 4402 15156
rect 5258 15144 5264 15156
rect 4396 15116 5264 15144
rect 4396 15104 4402 15116
rect 5258 15104 5264 15116
rect 5316 15144 5322 15156
rect 5442 15144 5448 15156
rect 5316 15116 5448 15144
rect 5316 15104 5322 15116
rect 5442 15104 5448 15116
rect 5500 15104 5506 15156
rect 5537 15147 5595 15153
rect 5537 15113 5549 15147
rect 5583 15144 5595 15147
rect 5626 15144 5632 15156
rect 5583 15116 5632 15144
rect 5583 15113 5595 15116
rect 5537 15107 5595 15113
rect 5626 15104 5632 15116
rect 5684 15104 5690 15156
rect 7926 15104 7932 15156
rect 7984 15144 7990 15156
rect 13170 15144 13176 15156
rect 7984 15116 13176 15144
rect 7984 15104 7990 15116
rect 13170 15104 13176 15116
rect 13228 15104 13234 15156
rect 13906 15144 13912 15156
rect 13280 15116 13912 15144
rect 2774 15076 2780 15088
rect 2608 15048 2780 15076
rect 2608 15017 2636 15048
rect 2774 15036 2780 15048
rect 2832 15076 2838 15088
rect 5350 15076 5356 15088
rect 2832 15048 5356 15076
rect 2832 15036 2838 15048
rect 5350 15036 5356 15048
rect 5408 15036 5414 15088
rect 2409 15011 2467 15017
rect 2409 14977 2421 15011
rect 2455 14977 2467 15011
rect 2409 14971 2467 14977
rect 2593 15011 2651 15017
rect 2593 14977 2605 15011
rect 2639 14977 2651 15011
rect 2593 14971 2651 14977
rect 3234 14968 3240 15020
rect 3292 15008 3298 15020
rect 3697 15011 3755 15017
rect 3697 15008 3709 15011
rect 3292 14980 3709 15008
rect 3292 14968 3298 14980
rect 3697 14977 3709 14980
rect 3743 14977 3755 15011
rect 3697 14971 3755 14977
rect 4706 14968 4712 15020
rect 4764 15008 4770 15020
rect 4893 15011 4951 15017
rect 4893 15008 4905 15011
rect 4764 14980 4905 15008
rect 4764 14968 4770 14980
rect 4893 14977 4905 14980
rect 4939 14977 4951 15011
rect 5644 15008 5672 15104
rect 13280 15088 13308 15116
rect 13906 15104 13912 15116
rect 13964 15104 13970 15156
rect 8662 15076 8668 15088
rect 8623 15048 8668 15076
rect 8662 15036 8668 15048
rect 8720 15036 8726 15088
rect 12437 15079 12495 15085
rect 12437 15076 12449 15079
rect 8772 15048 12449 15076
rect 8772 15008 8800 15048
rect 12437 15045 12449 15048
rect 12483 15045 12495 15079
rect 12437 15039 12495 15045
rect 13262 15036 13268 15088
rect 13320 15036 13326 15088
rect 13814 15036 13820 15088
rect 13872 15076 13878 15088
rect 14553 15079 14611 15085
rect 14553 15076 14565 15079
rect 13872 15048 14565 15076
rect 13872 15036 13878 15048
rect 14553 15045 14565 15048
rect 14599 15045 14611 15079
rect 14553 15039 14611 15045
rect 5644 14980 6408 15008
rect 4893 14971 4951 14977
rect 2958 14900 2964 14952
rect 3016 14940 3022 14952
rect 5534 14940 5540 14952
rect 3016 14912 5540 14940
rect 3016 14900 3022 14912
rect 5534 14900 5540 14912
rect 5592 14900 5598 14952
rect 5626 14900 5632 14952
rect 5684 14940 5690 14952
rect 6380 14949 6408 14980
rect 7852 14980 8800 15008
rect 9217 15011 9275 15017
rect 5721 14943 5779 14949
rect 5721 14940 5733 14943
rect 5684 14912 5733 14940
rect 5684 14900 5690 14912
rect 5721 14909 5733 14912
rect 5767 14909 5779 14943
rect 5721 14903 5779 14909
rect 6365 14943 6423 14949
rect 6365 14909 6377 14943
rect 6411 14909 6423 14943
rect 6822 14940 6828 14952
rect 6783 14912 6828 14940
rect 6365 14903 6423 14909
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 7852 14940 7880 14980
rect 9217 14977 9229 15011
rect 9263 14977 9275 15011
rect 9217 14971 9275 14977
rect 6932 14912 7880 14940
rect 2774 14832 2780 14884
rect 2832 14872 2838 14884
rect 3605 14875 3663 14881
rect 3605 14872 3617 14875
rect 2832 14844 3617 14872
rect 2832 14832 2838 14844
rect 3605 14841 3617 14844
rect 3651 14841 3663 14875
rect 4430 14872 4436 14884
rect 3605 14835 3663 14841
rect 3712 14844 4436 14872
rect 1946 14804 1952 14816
rect 1907 14776 1952 14804
rect 1946 14764 1952 14776
rect 2004 14764 2010 14816
rect 2314 14804 2320 14816
rect 2275 14776 2320 14804
rect 2314 14764 2320 14776
rect 2372 14764 2378 14816
rect 3145 14807 3203 14813
rect 3145 14773 3157 14807
rect 3191 14804 3203 14807
rect 3234 14804 3240 14816
rect 3191 14776 3240 14804
rect 3191 14773 3203 14776
rect 3145 14767 3203 14773
rect 3234 14764 3240 14776
rect 3292 14764 3298 14816
rect 3513 14807 3571 14813
rect 3513 14773 3525 14807
rect 3559 14804 3571 14807
rect 3712 14804 3740 14844
rect 4430 14832 4436 14844
rect 4488 14832 4494 14884
rect 4709 14875 4767 14881
rect 4709 14841 4721 14875
rect 4755 14872 4767 14875
rect 5074 14872 5080 14884
rect 4755 14844 5080 14872
rect 4755 14841 4767 14844
rect 4709 14835 4767 14841
rect 5074 14832 5080 14844
rect 5132 14832 5138 14884
rect 5258 14832 5264 14884
rect 5316 14872 5322 14884
rect 6932 14872 6960 14912
rect 8570 14900 8576 14952
rect 8628 14940 8634 14952
rect 9232 14940 9260 14971
rect 9306 14968 9312 15020
rect 9364 15008 9370 15020
rect 9582 15008 9588 15020
rect 9364 14980 9588 15008
rect 9364 14968 9370 14980
rect 9582 14968 9588 14980
rect 9640 15008 9646 15020
rect 11701 15011 11759 15017
rect 11701 15008 11713 15011
rect 9640 14980 11713 15008
rect 9640 14968 9646 14980
rect 11701 14977 11713 14980
rect 11747 15008 11759 15011
rect 12710 15008 12716 15020
rect 11747 14980 12716 15008
rect 11747 14977 11759 14980
rect 11701 14971 11759 14977
rect 12710 14968 12716 14980
rect 12768 14968 12774 15020
rect 12802 14968 12808 15020
rect 12860 15008 12866 15020
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 12860 14980 13001 15008
rect 12860 14968 12866 14980
rect 12989 14977 13001 14980
rect 13035 14977 13047 15011
rect 15378 15008 15384 15020
rect 12989 14971 13047 14977
rect 13096 14980 15384 15008
rect 9490 14940 9496 14952
rect 8628 14912 9496 14940
rect 8628 14900 8634 14912
rect 9490 14900 9496 14912
rect 9548 14900 9554 14952
rect 9766 14900 9772 14952
rect 9824 14940 9830 14952
rect 10045 14943 10103 14949
rect 10045 14940 10057 14943
rect 9824 14912 10057 14940
rect 9824 14900 9830 14912
rect 10045 14909 10057 14912
rect 10091 14940 10103 14943
rect 11790 14940 11796 14952
rect 10091 14912 11796 14940
rect 10091 14909 10103 14912
rect 10045 14903 10103 14909
rect 11790 14900 11796 14912
rect 11848 14900 11854 14952
rect 13096 14940 13124 14980
rect 15378 14968 15384 14980
rect 15436 14968 15442 15020
rect 12636 14912 13124 14940
rect 13633 14943 13691 14949
rect 5316 14844 6960 14872
rect 7092 14875 7150 14881
rect 5316 14832 5322 14844
rect 7092 14841 7104 14875
rect 7138 14872 7150 14875
rect 7190 14872 7196 14884
rect 7138 14844 7196 14872
rect 7138 14841 7150 14844
rect 7092 14835 7150 14841
rect 7190 14832 7196 14844
rect 7248 14832 7254 14884
rect 7558 14832 7564 14884
rect 7616 14872 7622 14884
rect 8588 14872 8616 14900
rect 7616 14844 8616 14872
rect 7616 14832 7622 14844
rect 8662 14832 8668 14884
rect 8720 14872 8726 14884
rect 9125 14875 9183 14881
rect 9125 14872 9137 14875
rect 8720 14844 9137 14872
rect 8720 14832 8726 14844
rect 9125 14841 9137 14844
rect 9171 14872 9183 14875
rect 10870 14872 10876 14884
rect 9171 14844 10876 14872
rect 9171 14841 9183 14844
rect 9125 14835 9183 14841
rect 10870 14832 10876 14844
rect 10928 14832 10934 14884
rect 11517 14875 11575 14881
rect 11517 14841 11529 14875
rect 11563 14872 11575 14875
rect 11974 14872 11980 14884
rect 11563 14844 11980 14872
rect 11563 14841 11575 14844
rect 11517 14835 11575 14841
rect 11974 14832 11980 14844
rect 12032 14872 12038 14884
rect 12250 14872 12256 14884
rect 12032 14844 12256 14872
rect 12032 14832 12038 14844
rect 12250 14832 12256 14844
rect 12308 14832 12314 14884
rect 4338 14804 4344 14816
rect 3559 14776 3740 14804
rect 4299 14776 4344 14804
rect 3559 14773 3571 14776
rect 3513 14767 3571 14773
rect 4338 14764 4344 14776
rect 4396 14764 4402 14816
rect 4801 14807 4859 14813
rect 4801 14773 4813 14807
rect 4847 14804 4859 14807
rect 5810 14804 5816 14816
rect 4847 14776 5816 14804
rect 4847 14773 4859 14776
rect 4801 14767 4859 14773
rect 5810 14764 5816 14776
rect 5868 14764 5874 14816
rect 6181 14807 6239 14813
rect 6181 14773 6193 14807
rect 6227 14804 6239 14807
rect 6270 14804 6276 14816
rect 6227 14776 6276 14804
rect 6227 14773 6239 14776
rect 6181 14767 6239 14773
rect 6270 14764 6276 14776
rect 6328 14764 6334 14816
rect 6362 14764 6368 14816
rect 6420 14804 6426 14816
rect 8205 14807 8263 14813
rect 8205 14804 8217 14807
rect 6420 14776 8217 14804
rect 6420 14764 6426 14776
rect 8205 14773 8217 14776
rect 8251 14773 8263 14807
rect 8205 14767 8263 14773
rect 8938 14764 8944 14816
rect 8996 14804 9002 14816
rect 9033 14807 9091 14813
rect 9033 14804 9045 14807
rect 8996 14776 9045 14804
rect 8996 14764 9002 14776
rect 9033 14773 9045 14776
rect 9079 14773 9091 14807
rect 9033 14767 9091 14773
rect 9861 14807 9919 14813
rect 9861 14773 9873 14807
rect 9907 14804 9919 14807
rect 10318 14804 10324 14816
rect 9907 14776 10324 14804
rect 9907 14773 9919 14776
rect 9861 14767 9919 14773
rect 10318 14764 10324 14776
rect 10376 14764 10382 14816
rect 11057 14807 11115 14813
rect 11057 14773 11069 14807
rect 11103 14804 11115 14807
rect 11146 14804 11152 14816
rect 11103 14776 11152 14804
rect 11103 14773 11115 14776
rect 11057 14767 11115 14773
rect 11146 14764 11152 14776
rect 11204 14764 11210 14816
rect 11425 14807 11483 14813
rect 11425 14773 11437 14807
rect 11471 14804 11483 14807
rect 12158 14804 12164 14816
rect 11471 14776 12164 14804
rect 11471 14773 11483 14776
rect 11425 14767 11483 14773
rect 12158 14764 12164 14776
rect 12216 14804 12222 14816
rect 12636 14804 12664 14912
rect 13633 14909 13645 14943
rect 13679 14940 13691 14943
rect 13998 14940 14004 14952
rect 13679 14912 14004 14940
rect 13679 14909 13691 14912
rect 13633 14903 13691 14909
rect 13998 14900 14004 14912
rect 14056 14900 14062 14952
rect 14366 14940 14372 14952
rect 14327 14912 14372 14940
rect 14366 14900 14372 14912
rect 14424 14900 14430 14952
rect 12897 14875 12955 14881
rect 12897 14841 12909 14875
rect 12943 14872 12955 14875
rect 14826 14872 14832 14884
rect 12943 14844 14832 14872
rect 12943 14841 12955 14844
rect 12897 14835 12955 14841
rect 14826 14832 14832 14844
rect 14884 14872 14890 14884
rect 16390 14872 16396 14884
rect 14884 14844 16396 14872
rect 14884 14832 14890 14844
rect 16390 14832 16396 14844
rect 16448 14832 16454 14884
rect 12802 14804 12808 14816
rect 12216 14776 12664 14804
rect 12763 14776 12808 14804
rect 12216 14764 12222 14776
rect 12802 14764 12808 14776
rect 12860 14764 12866 14816
rect 13814 14804 13820 14816
rect 13775 14776 13820 14804
rect 13814 14764 13820 14776
rect 13872 14764 13878 14816
rect 1104 14714 15824 14736
rect 1104 14662 5912 14714
rect 5964 14662 5976 14714
rect 6028 14662 6040 14714
rect 6092 14662 6104 14714
rect 6156 14662 10843 14714
rect 10895 14662 10907 14714
rect 10959 14662 10971 14714
rect 11023 14662 11035 14714
rect 11087 14662 15824 14714
rect 1104 14640 15824 14662
rect 1578 14600 1584 14612
rect 1539 14572 1584 14600
rect 1578 14560 1584 14572
rect 1636 14560 1642 14612
rect 4157 14603 4215 14609
rect 4157 14569 4169 14603
rect 4203 14600 4215 14603
rect 4798 14600 4804 14612
rect 4203 14572 4804 14600
rect 4203 14569 4215 14572
rect 4157 14563 4215 14569
rect 4798 14560 4804 14572
rect 4856 14560 4862 14612
rect 5718 14600 5724 14612
rect 5092 14572 5724 14600
rect 2041 14535 2099 14541
rect 2041 14501 2053 14535
rect 2087 14532 2099 14535
rect 2682 14532 2688 14544
rect 2087 14504 2688 14532
rect 2087 14501 2099 14504
rect 2041 14495 2099 14501
rect 2682 14492 2688 14504
rect 2740 14492 2746 14544
rect 4430 14492 4436 14544
rect 4488 14532 4494 14544
rect 4525 14535 4583 14541
rect 4525 14532 4537 14535
rect 4488 14504 4537 14532
rect 4488 14492 4494 14504
rect 4525 14501 4537 14504
rect 4571 14501 4583 14535
rect 4525 14495 4583 14501
rect 4614 14492 4620 14544
rect 4672 14532 4678 14544
rect 5092 14532 5120 14572
rect 5718 14560 5724 14572
rect 5776 14560 5782 14612
rect 5810 14560 5816 14612
rect 5868 14600 5874 14612
rect 7926 14600 7932 14612
rect 5868 14572 7932 14600
rect 5868 14560 5874 14572
rect 7926 14560 7932 14572
rect 7984 14560 7990 14612
rect 8110 14560 8116 14612
rect 8168 14600 8174 14612
rect 10873 14603 10931 14609
rect 10873 14600 10885 14603
rect 8168 14572 9628 14600
rect 8168 14560 8174 14572
rect 4672 14504 5120 14532
rect 5629 14535 5687 14541
rect 4672 14492 4678 14504
rect 5629 14501 5641 14535
rect 5675 14532 5687 14535
rect 5902 14532 5908 14544
rect 5675 14504 5908 14532
rect 5675 14501 5687 14504
rect 5629 14495 5687 14501
rect 5902 14492 5908 14504
rect 5960 14492 5966 14544
rect 9306 14532 9312 14544
rect 6656 14504 9312 14532
rect 1949 14467 2007 14473
rect 1949 14433 1961 14467
rect 1995 14464 2007 14467
rect 2958 14464 2964 14476
rect 1995 14436 2964 14464
rect 1995 14433 2007 14436
rect 1949 14427 2007 14433
rect 2958 14424 2964 14436
rect 3016 14424 3022 14476
rect 3145 14467 3203 14473
rect 3145 14433 3157 14467
rect 3191 14464 3203 14467
rect 4246 14464 4252 14476
rect 3191 14436 4252 14464
rect 3191 14433 3203 14436
rect 3145 14427 3203 14433
rect 4246 14424 4252 14436
rect 4304 14424 4310 14476
rect 4632 14464 4660 14492
rect 4632 14436 4752 14464
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14396 2283 14399
rect 2590 14396 2596 14408
rect 2271 14368 2596 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 2590 14356 2596 14368
rect 2648 14356 2654 14408
rect 3050 14356 3056 14408
rect 3108 14396 3114 14408
rect 3237 14399 3295 14405
rect 3237 14396 3249 14399
rect 3108 14368 3249 14396
rect 3108 14356 3114 14368
rect 3237 14365 3249 14368
rect 3283 14365 3295 14399
rect 3237 14359 3295 14365
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14396 3479 14399
rect 4430 14396 4436 14408
rect 3467 14368 4436 14396
rect 3467 14365 3479 14368
rect 3421 14359 3479 14365
rect 4430 14356 4436 14368
rect 4488 14356 4494 14408
rect 4724 14405 4752 14436
rect 5074 14424 5080 14476
rect 5132 14464 5138 14476
rect 5353 14467 5411 14473
rect 5353 14464 5365 14467
rect 5132 14436 5365 14464
rect 5132 14424 5138 14436
rect 5353 14433 5365 14436
rect 5399 14433 5411 14467
rect 5353 14427 5411 14433
rect 5718 14424 5724 14476
rect 5776 14464 5782 14476
rect 6457 14467 6515 14473
rect 6457 14464 6469 14467
rect 5776 14436 6469 14464
rect 5776 14424 5782 14436
rect 6457 14433 6469 14436
rect 6503 14433 6515 14467
rect 6457 14427 6515 14433
rect 4617 14399 4675 14405
rect 4617 14365 4629 14399
rect 4663 14365 4675 14399
rect 4617 14359 4675 14365
rect 4709 14399 4767 14405
rect 4709 14365 4721 14399
rect 4755 14365 4767 14399
rect 6656 14396 6684 14504
rect 9306 14492 9312 14504
rect 9364 14492 9370 14544
rect 9600 14532 9628 14572
rect 9699 14572 10885 14600
rect 9699 14532 9727 14572
rect 10873 14569 10885 14572
rect 10919 14569 10931 14603
rect 10873 14563 10931 14569
rect 11146 14560 11152 14612
rect 11204 14600 11210 14612
rect 12529 14603 12587 14609
rect 12529 14600 12541 14603
rect 11204 14572 12541 14600
rect 11204 14560 11210 14572
rect 12529 14569 12541 14572
rect 12575 14569 12587 14603
rect 12529 14563 12587 14569
rect 13170 14560 13176 14612
rect 13228 14600 13234 14612
rect 14645 14603 14703 14609
rect 14645 14600 14657 14603
rect 13228 14572 14657 14600
rect 13228 14560 13234 14572
rect 14645 14569 14657 14572
rect 14691 14569 14703 14603
rect 14645 14563 14703 14569
rect 9600 14504 9727 14532
rect 9858 14492 9864 14544
rect 9916 14532 9922 14544
rect 10502 14532 10508 14544
rect 9916 14504 10508 14532
rect 9916 14492 9922 14504
rect 10502 14492 10508 14504
rect 10560 14492 10566 14544
rect 11241 14535 11299 14541
rect 11241 14501 11253 14535
rect 11287 14532 11299 14535
rect 13262 14532 13268 14544
rect 11287 14504 13268 14532
rect 11287 14501 11299 14504
rect 11241 14495 11299 14501
rect 7098 14473 7104 14476
rect 7092 14464 7104 14473
rect 7059 14436 7104 14464
rect 7092 14427 7104 14436
rect 7098 14424 7104 14427
rect 7156 14424 7162 14476
rect 7926 14424 7932 14476
rect 7984 14464 7990 14476
rect 9493 14467 9551 14473
rect 7984 14436 9343 14464
rect 7984 14424 7990 14436
rect 6822 14396 6828 14408
rect 4709 14359 4767 14365
rect 5552 14368 6684 14396
rect 6783 14368 6828 14396
rect 4632 14328 4660 14359
rect 5552 14328 5580 14368
rect 6822 14356 6828 14368
rect 6880 14356 6886 14408
rect 8478 14356 8484 14408
rect 8536 14396 8542 14408
rect 8665 14399 8723 14405
rect 8665 14396 8677 14399
rect 8536 14368 8677 14396
rect 8536 14356 8542 14368
rect 8665 14365 8677 14368
rect 8711 14365 8723 14399
rect 8665 14359 8723 14365
rect 4632 14300 5580 14328
rect 5626 14288 5632 14340
rect 5684 14328 5690 14340
rect 6454 14328 6460 14340
rect 5684 14300 6460 14328
rect 5684 14288 5690 14300
rect 6454 14288 6460 14300
rect 6512 14288 6518 14340
rect 8110 14288 8116 14340
rect 8168 14328 8174 14340
rect 9214 14328 9220 14340
rect 8168 14300 9220 14328
rect 8168 14288 8174 14300
rect 9214 14288 9220 14300
rect 9272 14288 9278 14340
rect 9315 14328 9343 14436
rect 9493 14433 9505 14467
rect 9539 14464 9551 14467
rect 9539 14436 9996 14464
rect 9539 14433 9551 14436
rect 9493 14427 9551 14433
rect 9968 14396 9996 14436
rect 10134 14424 10140 14476
rect 10192 14464 10198 14476
rect 10264 14467 10322 14473
rect 10264 14464 10276 14467
rect 10192 14436 10276 14464
rect 10192 14424 10198 14436
rect 10264 14433 10276 14436
rect 10310 14433 10322 14467
rect 10264 14427 10322 14433
rect 10367 14467 10425 14473
rect 10367 14433 10379 14467
rect 10413 14464 10425 14467
rect 10594 14464 10600 14476
rect 10413 14436 10600 14464
rect 10413 14433 10425 14436
rect 10367 14427 10425 14433
rect 10594 14424 10600 14436
rect 10652 14424 10658 14476
rect 11054 14464 11060 14476
rect 10704 14436 11060 14464
rect 10704 14396 10732 14436
rect 11054 14424 11060 14436
rect 11112 14424 11118 14476
rect 11146 14424 11152 14476
rect 11204 14464 11210 14476
rect 11256 14464 11284 14495
rect 13262 14492 13268 14504
rect 13320 14492 13326 14544
rect 13722 14532 13728 14544
rect 13683 14504 13728 14532
rect 13722 14492 13728 14504
rect 13780 14492 13786 14544
rect 11204 14436 11284 14464
rect 11333 14467 11391 14473
rect 11204 14424 11210 14436
rect 11333 14433 11345 14467
rect 11379 14464 11391 14467
rect 12066 14464 12072 14476
rect 11379 14436 12072 14464
rect 11379 14433 11391 14436
rect 11333 14427 11391 14433
rect 12066 14424 12072 14436
rect 12124 14464 12130 14476
rect 12250 14464 12256 14476
rect 12124 14436 12256 14464
rect 12124 14424 12130 14436
rect 12250 14424 12256 14436
rect 12308 14424 12314 14476
rect 12434 14464 12440 14476
rect 12395 14436 12440 14464
rect 12434 14424 12440 14436
rect 12492 14424 12498 14476
rect 13173 14467 13231 14473
rect 13173 14433 13185 14467
rect 13219 14464 13231 14467
rect 13630 14464 13636 14476
rect 13219 14436 13636 14464
rect 13219 14433 13231 14436
rect 13173 14427 13231 14433
rect 13630 14424 13636 14436
rect 13688 14424 13694 14476
rect 14461 14467 14519 14473
rect 14461 14433 14473 14467
rect 14507 14464 14519 14467
rect 15286 14464 15292 14476
rect 14507 14436 15292 14464
rect 14507 14433 14519 14436
rect 14461 14427 14519 14433
rect 15286 14424 15292 14436
rect 15344 14424 15350 14476
rect 11425 14399 11483 14405
rect 11425 14396 11437 14399
rect 9968 14368 10732 14396
rect 10787 14368 11437 14396
rect 9315 14300 9435 14328
rect 2777 14263 2835 14269
rect 2777 14229 2789 14263
rect 2823 14260 2835 14263
rect 5074 14260 5080 14272
rect 2823 14232 5080 14260
rect 2823 14229 2835 14232
rect 2777 14223 2835 14229
rect 5074 14220 5080 14232
rect 5132 14220 5138 14272
rect 5810 14220 5816 14272
rect 5868 14260 5874 14272
rect 6273 14263 6331 14269
rect 6273 14260 6285 14263
rect 5868 14232 6285 14260
rect 5868 14220 5874 14232
rect 6273 14229 6285 14232
rect 6319 14229 6331 14263
rect 6273 14223 6331 14229
rect 7558 14220 7564 14272
rect 7616 14260 7622 14272
rect 8018 14260 8024 14272
rect 7616 14232 8024 14260
rect 7616 14220 7622 14232
rect 8018 14220 8024 14232
rect 8076 14260 8082 14272
rect 8205 14263 8263 14269
rect 8205 14260 8217 14263
rect 8076 14232 8217 14260
rect 8076 14220 8082 14232
rect 8205 14229 8217 14232
rect 8251 14229 8263 14263
rect 8205 14223 8263 14229
rect 9122 14220 9128 14272
rect 9180 14260 9186 14272
rect 9309 14263 9367 14269
rect 9309 14260 9321 14263
rect 9180 14232 9321 14260
rect 9180 14220 9186 14232
rect 9309 14229 9321 14232
rect 9355 14229 9367 14263
rect 9407 14260 9435 14300
rect 9490 14288 9496 14340
rect 9548 14328 9554 14340
rect 10134 14328 10140 14340
rect 9548 14300 10140 14328
rect 9548 14288 9554 14300
rect 10134 14288 10140 14300
rect 10192 14288 10198 14340
rect 10410 14288 10416 14340
rect 10468 14328 10474 14340
rect 10468 14300 10640 14328
rect 10468 14288 10474 14300
rect 10502 14260 10508 14272
rect 9407 14232 10508 14260
rect 9309 14223 9367 14229
rect 10502 14220 10508 14232
rect 10560 14220 10566 14272
rect 10612 14260 10640 14300
rect 10686 14288 10692 14340
rect 10744 14328 10750 14340
rect 10787 14328 10815 14368
rect 11425 14365 11437 14368
rect 11471 14365 11483 14399
rect 11425 14359 11483 14365
rect 12621 14399 12679 14405
rect 12621 14365 12633 14399
rect 12667 14365 12679 14399
rect 12621 14359 12679 14365
rect 12636 14328 12664 14359
rect 12986 14356 12992 14408
rect 13044 14396 13050 14408
rect 13909 14399 13967 14405
rect 13909 14396 13921 14399
rect 13044 14368 13921 14396
rect 13044 14356 13050 14368
rect 13909 14365 13921 14368
rect 13955 14365 13967 14399
rect 13909 14359 13967 14365
rect 10744 14300 10815 14328
rect 10888 14300 12664 14328
rect 10744 14288 10750 14300
rect 10888 14260 10916 14300
rect 10612 14232 10916 14260
rect 10962 14220 10968 14272
rect 11020 14260 11026 14272
rect 12069 14263 12127 14269
rect 12069 14260 12081 14263
rect 11020 14232 12081 14260
rect 11020 14220 11026 14232
rect 12069 14229 12081 14232
rect 12115 14229 12127 14263
rect 12069 14223 12127 14229
rect 13170 14220 13176 14272
rect 13228 14260 13234 14272
rect 13265 14263 13323 14269
rect 13265 14260 13277 14263
rect 13228 14232 13277 14260
rect 13228 14220 13234 14232
rect 13265 14229 13277 14232
rect 13311 14229 13323 14263
rect 13265 14223 13323 14229
rect 1104 14170 15824 14192
rect 1104 14118 3447 14170
rect 3499 14118 3511 14170
rect 3563 14118 3575 14170
rect 3627 14118 3639 14170
rect 3691 14118 8378 14170
rect 8430 14118 8442 14170
rect 8494 14118 8506 14170
rect 8558 14118 8570 14170
rect 8622 14118 13308 14170
rect 13360 14118 13372 14170
rect 13424 14118 13436 14170
rect 13488 14118 13500 14170
rect 13552 14118 15824 14170
rect 1104 14096 15824 14118
rect 2406 14016 2412 14068
rect 2464 14056 2470 14068
rect 3697 14059 3755 14065
rect 3697 14056 3709 14059
rect 2464 14028 3709 14056
rect 2464 14016 2470 14028
rect 3697 14025 3709 14028
rect 3743 14025 3755 14059
rect 3697 14019 3755 14025
rect 4246 14016 4252 14068
rect 4304 14056 4310 14068
rect 7285 14059 7343 14065
rect 4304 14028 7236 14056
rect 4304 14016 4310 14028
rect 2501 13991 2559 13997
rect 2501 13957 2513 13991
rect 2547 13988 2559 13991
rect 4522 13988 4528 14000
rect 2547 13960 4528 13988
rect 2547 13957 2559 13960
rect 2501 13951 2559 13957
rect 4522 13948 4528 13960
rect 4580 13948 4586 14000
rect 7208 13988 7236 14028
rect 7285 14025 7297 14059
rect 7331 14056 7343 14059
rect 8846 14056 8852 14068
rect 7331 14028 8852 14056
rect 7331 14025 7343 14028
rect 7285 14019 7343 14025
rect 8846 14016 8852 14028
rect 8904 14016 8910 14068
rect 9140 14028 10088 14056
rect 9140 13988 9168 14028
rect 7208 13960 9168 13988
rect 10060 13988 10088 14028
rect 10226 14016 10232 14068
rect 10284 14056 10290 14068
rect 11057 14059 11115 14065
rect 11057 14056 11069 14059
rect 10284 14028 11069 14056
rect 10284 14016 10290 14028
rect 11057 14025 11069 14028
rect 11103 14025 11115 14059
rect 12434 14056 12440 14068
rect 12395 14028 12440 14056
rect 11057 14019 11115 14025
rect 12434 14016 12440 14028
rect 12492 14016 12498 14068
rect 10686 13988 10692 14000
rect 10060 13960 10692 13988
rect 10686 13948 10692 13960
rect 10744 13948 10750 14000
rect 10965 13991 11023 13997
rect 10965 13957 10977 13991
rect 11011 13988 11023 13991
rect 12802 13988 12808 14000
rect 11011 13960 12808 13988
rect 11011 13957 11023 13960
rect 10965 13951 11023 13957
rect 12802 13948 12808 13960
rect 12860 13948 12866 14000
rect 13446 13948 13452 14000
rect 13504 13988 13510 14000
rect 15562 13988 15568 14000
rect 13504 13960 15568 13988
rect 13504 13948 13510 13960
rect 15562 13948 15568 13960
rect 15620 13948 15626 14000
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13920 3203 13923
rect 3418 13920 3424 13932
rect 3191 13892 3424 13920
rect 3191 13889 3203 13892
rect 3145 13883 3203 13889
rect 3418 13880 3424 13892
rect 3476 13880 3482 13932
rect 4246 13920 4252 13932
rect 4207 13892 4252 13920
rect 4246 13880 4252 13892
rect 4304 13880 4310 13932
rect 7466 13880 7472 13932
rect 7524 13920 7530 13932
rect 7745 13923 7803 13929
rect 7745 13920 7757 13923
rect 7524 13892 7757 13920
rect 7524 13880 7530 13892
rect 7745 13889 7757 13892
rect 7791 13889 7803 13923
rect 7745 13883 7803 13889
rect 7837 13923 7895 13929
rect 7837 13889 7849 13923
rect 7883 13889 7895 13923
rect 11609 13923 11667 13929
rect 11609 13920 11621 13923
rect 7837 13883 7895 13889
rect 10152 13892 11621 13920
rect 1486 13812 1492 13864
rect 1544 13852 1550 13864
rect 1581 13855 1639 13861
rect 1581 13852 1593 13855
rect 1544 13824 1593 13852
rect 1544 13812 1550 13824
rect 1581 13821 1593 13824
rect 1627 13821 1639 13855
rect 1581 13815 1639 13821
rect 2222 13812 2228 13864
rect 2280 13852 2286 13864
rect 2869 13855 2927 13861
rect 2869 13852 2881 13855
rect 2280 13824 2881 13852
rect 2280 13812 2286 13824
rect 2869 13821 2881 13824
rect 2915 13821 2927 13855
rect 4798 13852 4804 13864
rect 2869 13815 2927 13821
rect 3896 13824 4804 13852
rect 566 13744 572 13796
rect 624 13784 630 13796
rect 1857 13787 1915 13793
rect 1857 13784 1869 13787
rect 624 13756 1869 13784
rect 624 13744 630 13756
rect 1857 13753 1869 13756
rect 1903 13753 1915 13787
rect 1857 13747 1915 13753
rect 3896 13728 3924 13824
rect 4798 13812 4804 13824
rect 4856 13812 4862 13864
rect 4893 13855 4951 13861
rect 4893 13821 4905 13855
rect 4939 13852 4951 13855
rect 4982 13852 4988 13864
rect 4939 13824 4988 13852
rect 4939 13821 4951 13824
rect 4893 13815 4951 13821
rect 4982 13812 4988 13824
rect 5040 13852 5046 13864
rect 6270 13852 6276 13864
rect 5040 13824 6276 13852
rect 5040 13812 5046 13824
rect 6270 13812 6276 13824
rect 6328 13812 6334 13864
rect 7098 13812 7104 13864
rect 7156 13852 7162 13864
rect 7852 13852 7880 13883
rect 10152 13864 10180 13892
rect 11609 13889 11621 13892
rect 11655 13889 11667 13923
rect 11609 13883 11667 13889
rect 12710 13880 12716 13932
rect 12768 13920 12774 13932
rect 13081 13923 13139 13929
rect 13081 13920 13093 13923
rect 12768 13892 13093 13920
rect 12768 13880 12774 13892
rect 13081 13889 13093 13892
rect 13127 13920 13139 13923
rect 13354 13920 13360 13932
rect 13127 13892 13360 13920
rect 13127 13889 13139 13892
rect 13081 13883 13139 13889
rect 13354 13880 13360 13892
rect 13412 13880 13418 13932
rect 13630 13880 13636 13932
rect 13688 13920 13694 13932
rect 13817 13923 13875 13929
rect 13817 13920 13829 13923
rect 13688 13892 13829 13920
rect 13688 13880 13694 13892
rect 13817 13889 13829 13892
rect 13863 13889 13875 13923
rect 14090 13920 14096 13932
rect 14051 13892 14096 13920
rect 13817 13883 13875 13889
rect 14090 13880 14096 13892
rect 14148 13880 14154 13932
rect 9030 13852 9036 13864
rect 7156 13824 7880 13852
rect 7944 13824 9036 13852
rect 7156 13812 7162 13824
rect 4154 13784 4160 13796
rect 4115 13756 4160 13784
rect 4154 13744 4160 13756
rect 4212 13744 4218 13796
rect 4816 13784 4844 13812
rect 5138 13787 5196 13793
rect 5138 13784 5150 13787
rect 4816 13756 5150 13784
rect 5138 13753 5150 13756
rect 5184 13753 5196 13787
rect 5138 13747 5196 13753
rect 6104 13756 6776 13784
rect 2498 13676 2504 13728
rect 2556 13716 2562 13728
rect 2961 13719 3019 13725
rect 2961 13716 2973 13719
rect 2556 13688 2973 13716
rect 2556 13676 2562 13688
rect 2961 13685 2973 13688
rect 3007 13685 3019 13719
rect 2961 13679 3019 13685
rect 3878 13676 3884 13728
rect 3936 13676 3942 13728
rect 4065 13719 4123 13725
rect 4065 13685 4077 13719
rect 4111 13716 4123 13719
rect 6104 13716 6132 13756
rect 6270 13716 6276 13728
rect 4111 13688 6132 13716
rect 6231 13688 6276 13716
rect 4111 13685 4123 13688
rect 4065 13679 4123 13685
rect 6270 13676 6276 13688
rect 6328 13676 6334 13728
rect 6748 13716 6776 13756
rect 6822 13744 6828 13796
rect 6880 13784 6886 13796
rect 7944 13784 7972 13824
rect 9030 13812 9036 13824
rect 9088 13852 9094 13864
rect 9125 13855 9183 13861
rect 9125 13852 9137 13855
rect 9088 13824 9137 13852
rect 9088 13812 9094 13824
rect 9125 13821 9137 13824
rect 9171 13821 9183 13855
rect 10134 13852 10140 13864
rect 9125 13815 9183 13821
rect 9784 13824 10140 13852
rect 6880 13756 7972 13784
rect 8481 13787 8539 13793
rect 6880 13744 6886 13756
rect 8481 13753 8493 13787
rect 8527 13784 8539 13787
rect 8754 13784 8760 13796
rect 8527 13756 8760 13784
rect 8527 13753 8539 13756
rect 8481 13747 8539 13753
rect 8754 13744 8760 13756
rect 8812 13744 8818 13796
rect 8846 13744 8852 13796
rect 8904 13784 8910 13796
rect 9392 13787 9450 13793
rect 8904 13756 9343 13784
rect 8904 13744 8910 13756
rect 7098 13716 7104 13728
rect 6748 13688 7104 13716
rect 7098 13676 7104 13688
rect 7156 13676 7162 13728
rect 7653 13719 7711 13725
rect 7653 13685 7665 13719
rect 7699 13716 7711 13719
rect 7742 13716 7748 13728
rect 7699 13688 7748 13716
rect 7699 13685 7711 13688
rect 7653 13679 7711 13685
rect 7742 13676 7748 13688
rect 7800 13716 7806 13728
rect 7926 13716 7932 13728
rect 7800 13688 7932 13716
rect 7800 13676 7806 13688
rect 7926 13676 7932 13688
rect 7984 13676 7990 13728
rect 9315 13716 9343 13756
rect 9392 13753 9404 13787
rect 9438 13784 9450 13787
rect 9784 13784 9812 13824
rect 10134 13812 10140 13824
rect 10192 13812 10198 13864
rect 10778 13812 10784 13864
rect 10836 13852 10842 13864
rect 10836 13824 13676 13852
rect 10836 13812 10842 13824
rect 9438 13756 9812 13784
rect 9438 13753 9450 13756
rect 9392 13747 9450 13753
rect 10042 13744 10048 13796
rect 10100 13784 10106 13796
rect 10965 13787 11023 13793
rect 10965 13784 10977 13787
rect 10100 13756 10977 13784
rect 10100 13744 10106 13756
rect 10965 13753 10977 13756
rect 11011 13753 11023 13787
rect 10965 13747 11023 13753
rect 11054 13744 11060 13796
rect 11112 13784 11118 13796
rect 12158 13784 12164 13796
rect 11112 13756 12164 13784
rect 11112 13744 11118 13756
rect 12158 13744 12164 13756
rect 12216 13744 12222 13796
rect 12618 13744 12624 13796
rect 12676 13784 12682 13796
rect 13648 13784 13676 13824
rect 13909 13787 13967 13793
rect 13909 13784 13921 13787
rect 12676 13756 13584 13784
rect 13648 13756 13921 13784
rect 12676 13744 12682 13756
rect 9582 13716 9588 13728
rect 9315 13688 9588 13716
rect 9582 13676 9588 13688
rect 9640 13676 9646 13728
rect 9674 13676 9680 13728
rect 9732 13716 9738 13728
rect 10226 13716 10232 13728
rect 9732 13688 10232 13716
rect 9732 13676 9738 13688
rect 10226 13676 10232 13688
rect 10284 13676 10290 13728
rect 10505 13719 10563 13725
rect 10505 13685 10517 13719
rect 10551 13716 10563 13719
rect 10594 13716 10600 13728
rect 10551 13688 10600 13716
rect 10551 13685 10563 13688
rect 10505 13679 10563 13685
rect 10594 13676 10600 13688
rect 10652 13676 10658 13728
rect 11330 13676 11336 13728
rect 11388 13716 11394 13728
rect 11425 13719 11483 13725
rect 11425 13716 11437 13719
rect 11388 13688 11437 13716
rect 11388 13676 11394 13688
rect 11425 13685 11437 13688
rect 11471 13685 11483 13719
rect 11425 13679 11483 13685
rect 11517 13719 11575 13725
rect 11517 13685 11529 13719
rect 11563 13716 11575 13719
rect 11882 13716 11888 13728
rect 11563 13688 11888 13716
rect 11563 13685 11575 13688
rect 11517 13679 11575 13685
rect 11882 13676 11888 13688
rect 11940 13676 11946 13728
rect 12802 13716 12808 13728
rect 12763 13688 12808 13716
rect 12802 13676 12808 13688
rect 12860 13676 12866 13728
rect 12897 13719 12955 13725
rect 12897 13685 12909 13719
rect 12943 13716 12955 13719
rect 13446 13716 13452 13728
rect 12943 13688 13452 13716
rect 12943 13685 12955 13688
rect 12897 13679 12955 13685
rect 13446 13676 13452 13688
rect 13504 13676 13510 13728
rect 13556 13716 13584 13756
rect 13909 13753 13921 13756
rect 13955 13753 13967 13787
rect 13909 13747 13967 13753
rect 13998 13716 14004 13728
rect 13556 13688 14004 13716
rect 13998 13676 14004 13688
rect 14056 13676 14062 13728
rect 1104 13626 15824 13648
rect 1104 13574 5912 13626
rect 5964 13574 5976 13626
rect 6028 13574 6040 13626
rect 6092 13574 6104 13626
rect 6156 13574 10843 13626
rect 10895 13574 10907 13626
rect 10959 13574 10971 13626
rect 11023 13574 11035 13626
rect 11087 13574 15824 13626
rect 1104 13552 15824 13574
rect 2774 13472 2780 13524
rect 2832 13512 2838 13524
rect 6362 13512 6368 13524
rect 2832 13484 2877 13512
rect 3068 13484 6368 13512
rect 2832 13472 2838 13484
rect 2590 13404 2596 13456
rect 2648 13444 2654 13456
rect 3068 13444 3096 13484
rect 6362 13472 6368 13484
rect 6420 13472 6426 13524
rect 7190 13512 7196 13524
rect 7151 13484 7196 13512
rect 7190 13472 7196 13484
rect 7248 13472 7254 13524
rect 7650 13512 7656 13524
rect 7611 13484 7656 13512
rect 7650 13472 7656 13484
rect 7708 13472 7714 13524
rect 8113 13515 8171 13521
rect 8113 13481 8125 13515
rect 8159 13512 8171 13515
rect 8159 13484 10180 13512
rect 8159 13481 8171 13484
rect 8113 13475 8171 13481
rect 2648 13416 3096 13444
rect 3237 13447 3295 13453
rect 2648 13404 2654 13416
rect 3237 13413 3249 13447
rect 3283 13444 3295 13447
rect 3786 13444 3792 13456
rect 3283 13416 3792 13444
rect 3283 13413 3295 13416
rect 3237 13407 3295 13413
rect 3786 13404 3792 13416
rect 3844 13404 3850 13456
rect 6270 13444 6276 13456
rect 3988 13416 6276 13444
rect 1949 13379 2007 13385
rect 1949 13345 1961 13379
rect 1995 13345 2007 13379
rect 1949 13339 2007 13345
rect 1578 13240 1584 13252
rect 1539 13212 1584 13240
rect 1578 13200 1584 13212
rect 1636 13200 1642 13252
rect 1964 13172 1992 13339
rect 2958 13336 2964 13388
rect 3016 13376 3022 13388
rect 3145 13379 3203 13385
rect 3145 13376 3157 13379
rect 3016 13348 3157 13376
rect 3016 13336 3022 13348
rect 3145 13345 3157 13348
rect 3191 13345 3203 13379
rect 3145 13339 3203 13345
rect 2041 13311 2099 13317
rect 2041 13277 2053 13311
rect 2087 13277 2099 13311
rect 2041 13271 2099 13277
rect 2225 13311 2283 13317
rect 2225 13277 2237 13311
rect 2271 13308 2283 13311
rect 3421 13311 3479 13317
rect 2271 13280 3280 13308
rect 2271 13277 2283 13280
rect 2225 13271 2283 13277
rect 2056 13240 2084 13271
rect 2590 13240 2596 13252
rect 2056 13212 2596 13240
rect 2590 13200 2596 13212
rect 2648 13200 2654 13252
rect 3252 13240 3280 13280
rect 3421 13277 3433 13311
rect 3467 13308 3479 13311
rect 3988 13308 4016 13416
rect 6270 13404 6276 13416
rect 6328 13404 6334 13456
rect 7558 13404 7564 13456
rect 7616 13444 7622 13456
rect 8570 13444 8576 13456
rect 7616 13416 8576 13444
rect 7616 13404 7622 13416
rect 8570 13404 8576 13416
rect 8628 13404 8634 13456
rect 9306 13404 9312 13456
rect 9364 13444 9370 13456
rect 10042 13444 10048 13456
rect 9364 13416 10048 13444
rect 9364 13404 9370 13416
rect 10042 13404 10048 13416
rect 10100 13404 10106 13456
rect 10152 13444 10180 13484
rect 10226 13472 10232 13524
rect 10284 13512 10290 13524
rect 12802 13512 12808 13524
rect 10284 13484 12808 13512
rect 10284 13472 10290 13484
rect 12802 13472 12808 13484
rect 12860 13472 12866 13524
rect 12710 13444 12716 13456
rect 10152 13416 10307 13444
rect 4065 13379 4123 13385
rect 4065 13345 4077 13379
rect 4111 13376 4123 13379
rect 5442 13376 5448 13388
rect 4111 13348 5448 13376
rect 4111 13345 4123 13348
rect 4065 13339 4123 13345
rect 5442 13336 5448 13348
rect 5500 13336 5506 13388
rect 6080 13379 6138 13385
rect 6080 13345 6092 13379
rect 6126 13376 6138 13379
rect 6362 13376 6368 13388
rect 6126 13348 6368 13376
rect 6126 13345 6138 13348
rect 6080 13339 6138 13345
rect 6362 13336 6368 13348
rect 6420 13336 6426 13388
rect 6638 13336 6644 13388
rect 6696 13376 6702 13388
rect 7282 13376 7288 13388
rect 6696 13348 7288 13376
rect 6696 13336 6702 13348
rect 7282 13336 7288 13348
rect 7340 13336 7346 13388
rect 8021 13379 8079 13385
rect 8021 13345 8033 13379
rect 8067 13376 8079 13379
rect 8110 13376 8116 13388
rect 8067 13348 8116 13376
rect 8067 13345 8079 13348
rect 8021 13339 8079 13345
rect 8110 13336 8116 13348
rect 8168 13336 8174 13388
rect 8849 13379 8907 13385
rect 8849 13345 8861 13379
rect 8895 13376 8907 13379
rect 9490 13376 9496 13388
rect 8895 13348 9496 13376
rect 8895 13345 8907 13348
rect 8849 13339 8907 13345
rect 9490 13336 9496 13348
rect 9548 13336 9554 13388
rect 9585 13379 9643 13385
rect 9585 13345 9597 13379
rect 9631 13376 9643 13379
rect 9933 13379 9991 13385
rect 9933 13376 9945 13379
rect 9631 13348 9945 13376
rect 9631 13345 9643 13348
rect 9585 13339 9643 13345
rect 9933 13345 9945 13348
rect 9979 13345 9991 13379
rect 10279 13376 10307 13416
rect 10520 13416 12716 13444
rect 10520 13376 10548 13416
rect 12710 13404 12716 13416
rect 12768 13404 12774 13456
rect 13081 13447 13139 13453
rect 13081 13413 13093 13447
rect 13127 13444 13139 13447
rect 13262 13444 13268 13456
rect 13127 13416 13268 13444
rect 13127 13413 13139 13416
rect 13081 13407 13139 13413
rect 13262 13404 13268 13416
rect 13320 13404 13326 13456
rect 13538 13404 13544 13456
rect 13596 13444 13602 13456
rect 13998 13444 14004 13456
rect 13596 13416 14004 13444
rect 13596 13404 13602 13416
rect 13998 13404 14004 13416
rect 14056 13444 14062 13456
rect 14277 13447 14335 13453
rect 14277 13444 14289 13447
rect 14056 13416 14289 13444
rect 14056 13404 14062 13416
rect 14277 13413 14289 13416
rect 14323 13413 14335 13447
rect 14277 13407 14335 13413
rect 10279 13348 10548 13376
rect 9933 13339 9991 13345
rect 10870 13336 10876 13388
rect 10928 13376 10934 13388
rect 11882 13376 11888 13388
rect 10928 13348 11744 13376
rect 11843 13348 11888 13376
rect 10928 13336 10934 13348
rect 4246 13308 4252 13320
rect 3467 13280 4016 13308
rect 4207 13280 4252 13308
rect 3467 13277 3479 13280
rect 3421 13271 3479 13277
rect 4246 13268 4252 13280
rect 4304 13268 4310 13320
rect 5074 13268 5080 13320
rect 5132 13308 5138 13320
rect 5169 13311 5227 13317
rect 5169 13308 5181 13311
rect 5132 13280 5181 13308
rect 5132 13268 5138 13280
rect 5169 13277 5181 13280
rect 5215 13277 5227 13311
rect 5169 13271 5227 13277
rect 5813 13311 5871 13317
rect 5813 13277 5825 13311
rect 5859 13277 5871 13311
rect 5813 13271 5871 13277
rect 4522 13240 4528 13252
rect 3252 13212 4528 13240
rect 4522 13200 4528 13212
rect 4580 13200 4586 13252
rect 4798 13200 4804 13252
rect 4856 13240 4862 13252
rect 4982 13240 4988 13252
rect 4856 13212 4988 13240
rect 4856 13200 4862 13212
rect 4982 13200 4988 13212
rect 5040 13240 5046 13252
rect 5828 13240 5856 13271
rect 7742 13268 7748 13320
rect 7800 13308 7806 13320
rect 8297 13311 8355 13317
rect 8297 13308 8309 13311
rect 7800 13280 8309 13308
rect 7800 13268 7806 13280
rect 8297 13277 8309 13280
rect 8343 13308 8355 13311
rect 8754 13308 8760 13320
rect 8343 13280 8760 13308
rect 8343 13277 8355 13280
rect 8297 13271 8355 13277
rect 8754 13268 8760 13280
rect 8812 13268 8818 13320
rect 9030 13268 9036 13320
rect 9088 13308 9094 13320
rect 9684 13311 9742 13317
rect 9088 13280 9628 13308
rect 9088 13268 9094 13280
rect 8110 13240 8116 13252
rect 5040 13212 5856 13240
rect 6748 13212 8116 13240
rect 5040 13200 5046 13212
rect 2222 13172 2228 13184
rect 1964 13144 2228 13172
rect 2222 13132 2228 13144
rect 2280 13172 2286 13184
rect 6748 13172 6776 13212
rect 8110 13200 8116 13212
rect 8168 13200 8174 13252
rect 8386 13200 8392 13252
rect 8444 13240 8450 13252
rect 9493 13243 9551 13249
rect 9493 13240 9505 13243
rect 8444 13212 9505 13240
rect 8444 13200 8450 13212
rect 9493 13209 9505 13212
rect 9539 13209 9551 13243
rect 9600 13240 9628 13280
rect 9684 13277 9696 13311
rect 9730 13277 9742 13311
rect 9684 13271 9742 13277
rect 9692 13240 9720 13271
rect 11238 13268 11244 13320
rect 11296 13308 11302 13320
rect 11296 13280 11652 13308
rect 11296 13268 11302 13280
rect 9600 13212 9720 13240
rect 9493 13203 9551 13209
rect 10778 13200 10784 13252
rect 10836 13240 10842 13252
rect 11517 13243 11575 13249
rect 11517 13240 11529 13243
rect 10836 13212 11529 13240
rect 10836 13200 10842 13212
rect 11517 13209 11529 13212
rect 11563 13209 11575 13243
rect 11517 13203 11575 13209
rect 2280 13144 6776 13172
rect 2280 13132 2286 13144
rect 7006 13132 7012 13184
rect 7064 13172 7070 13184
rect 7650 13172 7656 13184
rect 7064 13144 7656 13172
rect 7064 13132 7070 13144
rect 7650 13132 7656 13144
rect 7708 13172 7714 13184
rect 10870 13172 10876 13184
rect 7708 13144 10876 13172
rect 7708 13132 7714 13144
rect 10870 13132 10876 13144
rect 10928 13132 10934 13184
rect 11057 13175 11115 13181
rect 11057 13141 11069 13175
rect 11103 13172 11115 13175
rect 11238 13172 11244 13184
rect 11103 13144 11244 13172
rect 11103 13141 11115 13144
rect 11057 13135 11115 13141
rect 11238 13132 11244 13144
rect 11296 13132 11302 13184
rect 11624 13172 11652 13280
rect 11716 13240 11744 13348
rect 11882 13336 11888 13348
rect 11940 13336 11946 13388
rect 12986 13336 12992 13388
rect 13044 13376 13050 13388
rect 13044 13348 13400 13376
rect 13044 13336 13050 13348
rect 11974 13308 11980 13320
rect 11935 13280 11980 13308
rect 11974 13268 11980 13280
rect 12032 13268 12038 13320
rect 12069 13311 12127 13317
rect 12069 13277 12081 13311
rect 12115 13277 12127 13311
rect 12069 13271 12127 13277
rect 12084 13240 12112 13271
rect 12158 13268 12164 13320
rect 12216 13308 12222 13320
rect 13078 13308 13084 13320
rect 12216 13280 13084 13308
rect 12216 13268 12222 13280
rect 13078 13268 13084 13280
rect 13136 13308 13142 13320
rect 13173 13311 13231 13317
rect 13173 13308 13185 13311
rect 13136 13280 13185 13308
rect 13136 13268 13142 13280
rect 13173 13277 13185 13280
rect 13219 13277 13231 13311
rect 13173 13271 13231 13277
rect 13265 13311 13323 13317
rect 13265 13277 13277 13311
rect 13311 13277 13323 13311
rect 13372 13308 13400 13348
rect 13906 13336 13912 13388
rect 13964 13376 13970 13388
rect 14369 13379 14427 13385
rect 14369 13376 14381 13379
rect 13964 13348 14381 13376
rect 13964 13336 13970 13348
rect 14369 13345 14381 13348
rect 14415 13345 14427 13379
rect 14369 13339 14427 13345
rect 14461 13311 14519 13317
rect 14461 13308 14473 13311
rect 13372 13280 14473 13308
rect 13265 13271 13323 13277
rect 14461 13277 14473 13280
rect 14507 13277 14519 13311
rect 14461 13271 14519 13277
rect 11716 13212 12112 13240
rect 12986 13200 12992 13252
rect 13044 13240 13050 13252
rect 13280 13240 13308 13271
rect 13044 13212 13308 13240
rect 13044 13200 13050 13212
rect 12713 13175 12771 13181
rect 12713 13172 12725 13175
rect 11624 13144 12725 13172
rect 12713 13141 12725 13144
rect 12759 13141 12771 13175
rect 12713 13135 12771 13141
rect 13078 13132 13084 13184
rect 13136 13172 13142 13184
rect 13909 13175 13967 13181
rect 13909 13172 13921 13175
rect 13136 13144 13921 13172
rect 13136 13132 13142 13144
rect 13909 13141 13921 13144
rect 13955 13141 13967 13175
rect 13909 13135 13967 13141
rect 1104 13082 15824 13104
rect 1104 13030 3447 13082
rect 3499 13030 3511 13082
rect 3563 13030 3575 13082
rect 3627 13030 3639 13082
rect 3691 13030 8378 13082
rect 8430 13030 8442 13082
rect 8494 13030 8506 13082
rect 8558 13030 8570 13082
rect 8622 13030 13308 13082
rect 13360 13030 13372 13082
rect 13424 13030 13436 13082
rect 13488 13030 13500 13082
rect 13552 13030 15824 13082
rect 1104 13008 15824 13030
rect 1857 12971 1915 12977
rect 1857 12937 1869 12971
rect 1903 12968 1915 12971
rect 3050 12968 3056 12980
rect 1903 12940 3056 12968
rect 1903 12937 1915 12940
rect 1857 12931 1915 12937
rect 3050 12928 3056 12940
rect 3108 12928 3114 12980
rect 4430 12968 4436 12980
rect 4391 12940 4436 12968
rect 4430 12928 4436 12940
rect 4488 12928 4494 12980
rect 4522 12928 4528 12980
rect 4580 12968 4586 12980
rect 6273 12971 6331 12977
rect 6273 12968 6285 12971
rect 4580 12940 6285 12968
rect 4580 12928 4586 12940
rect 6273 12937 6285 12940
rect 6319 12937 6331 12971
rect 6273 12931 6331 12937
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12801 2559 12835
rect 4448 12832 4476 12928
rect 4448 12804 5028 12832
rect 2501 12795 2559 12801
rect 1486 12656 1492 12708
rect 1544 12696 1550 12708
rect 2225 12699 2283 12705
rect 2225 12696 2237 12699
rect 1544 12668 2237 12696
rect 1544 12656 1550 12668
rect 2225 12665 2237 12668
rect 2271 12665 2283 12699
rect 2516 12696 2544 12795
rect 3053 12767 3111 12773
rect 3053 12733 3065 12767
rect 3099 12764 3111 12767
rect 4798 12764 4804 12776
rect 3099 12736 4804 12764
rect 3099 12733 3111 12736
rect 3053 12727 3111 12733
rect 4798 12724 4804 12736
rect 4856 12764 4862 12776
rect 4893 12767 4951 12773
rect 4893 12764 4905 12767
rect 4856 12736 4905 12764
rect 4856 12724 4862 12736
rect 4893 12733 4905 12736
rect 4939 12733 4951 12767
rect 5000 12764 5028 12804
rect 5149 12767 5207 12773
rect 5149 12764 5161 12767
rect 5000 12736 5161 12764
rect 4893 12727 4951 12733
rect 5149 12733 5161 12736
rect 5195 12733 5207 12767
rect 6288 12764 6316 12931
rect 7098 12928 7104 12980
rect 7156 12968 7162 12980
rect 7156 12940 7871 12968
rect 7156 12928 7162 12940
rect 7843 12900 7871 12940
rect 8110 12928 8116 12980
rect 8168 12968 8174 12980
rect 8662 12968 8668 12980
rect 8168 12940 8668 12968
rect 8168 12928 8174 12940
rect 8662 12928 8668 12940
rect 8720 12928 8726 12980
rect 8757 12971 8815 12977
rect 8757 12937 8769 12971
rect 8803 12968 8815 12971
rect 10226 12968 10232 12980
rect 8803 12940 10232 12968
rect 8803 12937 8815 12940
rect 8757 12931 8815 12937
rect 10226 12928 10232 12940
rect 10284 12928 10290 12980
rect 10597 12971 10655 12977
rect 10597 12968 10609 12971
rect 10520 12940 10609 12968
rect 10520 12900 10548 12940
rect 10597 12937 10609 12940
rect 10643 12937 10655 12971
rect 10597 12931 10655 12937
rect 10870 12928 10876 12980
rect 10928 12968 10934 12980
rect 11974 12968 11980 12980
rect 10928 12940 11980 12968
rect 10928 12928 10934 12940
rect 11974 12928 11980 12940
rect 12032 12928 12038 12980
rect 12710 12928 12716 12980
rect 12768 12968 12774 12980
rect 13633 12971 13691 12977
rect 13633 12968 13645 12971
rect 12768 12940 13645 12968
rect 12768 12928 12774 12940
rect 13633 12937 13645 12940
rect 13679 12937 13691 12971
rect 13633 12931 13691 12937
rect 13814 12928 13820 12980
rect 13872 12968 13878 12980
rect 15013 12971 15071 12977
rect 15013 12968 15025 12971
rect 13872 12940 15025 12968
rect 13872 12928 13878 12940
rect 15013 12937 15025 12940
rect 15059 12937 15071 12971
rect 15013 12931 15071 12937
rect 7843 12872 10548 12900
rect 10612 12872 11560 12900
rect 6822 12792 6828 12844
rect 6880 12832 6886 12844
rect 6917 12835 6975 12841
rect 6917 12832 6929 12835
rect 6880 12804 6929 12832
rect 6880 12792 6886 12804
rect 6917 12801 6929 12804
rect 6963 12801 6975 12835
rect 6917 12795 6975 12801
rect 8294 12792 8300 12844
rect 8352 12832 8358 12844
rect 9309 12835 9367 12841
rect 9309 12832 9321 12835
rect 8352 12804 9321 12832
rect 8352 12792 8358 12804
rect 9309 12801 9321 12804
rect 9355 12801 9367 12835
rect 10612 12832 10640 12872
rect 10870 12832 10876 12844
rect 9309 12795 9367 12801
rect 9600 12804 10640 12832
rect 10704 12804 10876 12832
rect 7184 12767 7242 12773
rect 7184 12764 7196 12767
rect 6288 12736 7196 12764
rect 5149 12727 5207 12733
rect 7184 12733 7196 12736
rect 7230 12764 7242 12767
rect 9600 12764 9628 12804
rect 7230 12736 9628 12764
rect 7230 12733 7242 12736
rect 7184 12727 7242 12733
rect 10226 12724 10232 12776
rect 10284 12764 10290 12776
rect 10704 12764 10732 12804
rect 10870 12792 10876 12804
rect 10928 12792 10934 12844
rect 11241 12835 11299 12841
rect 11241 12801 11253 12835
rect 11287 12832 11299 12835
rect 11422 12832 11428 12844
rect 11287 12804 11428 12832
rect 11287 12801 11299 12804
rect 11241 12795 11299 12801
rect 11422 12792 11428 12804
rect 11480 12792 11486 12844
rect 11532 12832 11560 12872
rect 11790 12860 11796 12912
rect 11848 12900 11854 12912
rect 11848 12872 11893 12900
rect 11848 12860 11854 12872
rect 13262 12860 13268 12912
rect 13320 12900 13326 12912
rect 14734 12900 14740 12912
rect 13320 12872 14740 12900
rect 13320 12860 13326 12872
rect 14734 12860 14740 12872
rect 14792 12860 14798 12912
rect 12986 12832 12992 12844
rect 11532 12804 12992 12832
rect 12986 12792 12992 12804
rect 13044 12792 13050 12844
rect 13630 12792 13636 12844
rect 13688 12832 13694 12844
rect 14185 12835 14243 12841
rect 14185 12832 14197 12835
rect 13688 12804 14197 12832
rect 13688 12792 13694 12804
rect 14185 12801 14197 12804
rect 14231 12801 14243 12835
rect 14185 12795 14243 12801
rect 10284 12736 10732 12764
rect 10284 12724 10290 12736
rect 10778 12724 10784 12776
rect 10836 12764 10842 12776
rect 11057 12767 11115 12773
rect 11057 12764 11069 12767
rect 10836 12736 11069 12764
rect 10836 12724 10842 12736
rect 11057 12733 11069 12736
rect 11103 12733 11115 12767
rect 11057 12727 11115 12733
rect 11790 12724 11796 12776
rect 11848 12764 11854 12776
rect 11977 12767 12035 12773
rect 11977 12764 11989 12767
rect 11848 12736 11989 12764
rect 11848 12724 11854 12736
rect 11977 12733 11989 12736
rect 12023 12733 12035 12767
rect 14829 12767 14887 12773
rect 14829 12764 14841 12767
rect 11977 12727 12035 12733
rect 12268 12736 14841 12764
rect 3320 12699 3378 12705
rect 3320 12696 3332 12699
rect 2516 12668 3332 12696
rect 2225 12659 2283 12665
rect 3320 12665 3332 12668
rect 3366 12696 3378 12699
rect 7006 12696 7012 12708
rect 3366 12668 7012 12696
rect 3366 12665 3378 12668
rect 3320 12659 3378 12665
rect 7006 12656 7012 12668
rect 7064 12656 7070 12708
rect 8754 12696 8760 12708
rect 7107 12668 8760 12696
rect 2317 12631 2375 12637
rect 2317 12597 2329 12631
rect 2363 12628 2375 12631
rect 4338 12628 4344 12640
rect 2363 12600 4344 12628
rect 2363 12597 2375 12600
rect 2317 12591 2375 12597
rect 4338 12588 4344 12600
rect 4396 12588 4402 12640
rect 5626 12588 5632 12640
rect 5684 12628 5690 12640
rect 7107 12628 7135 12668
rect 8754 12656 8760 12668
rect 8812 12656 8818 12708
rect 9214 12696 9220 12708
rect 9175 12668 9220 12696
rect 9214 12656 9220 12668
rect 9272 12656 9278 12708
rect 10410 12696 10416 12708
rect 9876 12668 10416 12696
rect 5684 12600 7135 12628
rect 5684 12588 5690 12600
rect 7374 12588 7380 12640
rect 7432 12628 7438 12640
rect 8297 12631 8355 12637
rect 8297 12628 8309 12631
rect 7432 12600 8309 12628
rect 7432 12588 7438 12600
rect 8297 12597 8309 12600
rect 8343 12628 8355 12631
rect 8846 12628 8852 12640
rect 8343 12600 8852 12628
rect 8343 12597 8355 12600
rect 8297 12591 8355 12597
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 9125 12631 9183 12637
rect 9125 12597 9137 12631
rect 9171 12628 9183 12631
rect 9876 12628 9904 12668
rect 10410 12656 10416 12668
rect 10468 12656 10474 12708
rect 10594 12656 10600 12708
rect 10652 12696 10658 12708
rect 10652 12668 11100 12696
rect 10652 12656 10658 12668
rect 9171 12600 9904 12628
rect 9953 12631 10011 12637
rect 9171 12597 9183 12600
rect 9125 12591 9183 12597
rect 9953 12597 9965 12631
rect 9999 12628 10011 12631
rect 10134 12628 10140 12640
rect 9999 12600 10140 12628
rect 9999 12597 10011 12600
rect 9953 12591 10011 12597
rect 10134 12588 10140 12600
rect 10192 12588 10198 12640
rect 10226 12588 10232 12640
rect 10284 12628 10290 12640
rect 10965 12631 11023 12637
rect 10965 12628 10977 12631
rect 10284 12600 10977 12628
rect 10284 12588 10290 12600
rect 10965 12597 10977 12600
rect 11011 12597 11023 12631
rect 11072 12628 11100 12668
rect 11606 12656 11612 12708
rect 11664 12696 11670 12708
rect 12158 12696 12164 12708
rect 11664 12668 12164 12696
rect 11664 12656 11670 12668
rect 12158 12656 12164 12668
rect 12216 12656 12222 12708
rect 12268 12628 12296 12736
rect 14829 12733 14841 12736
rect 14875 12733 14887 12767
rect 14829 12727 14887 12733
rect 14093 12699 14151 12705
rect 14093 12696 14105 12699
rect 12452 12668 14105 12696
rect 12452 12637 12480 12668
rect 14093 12665 14105 12668
rect 14139 12665 14151 12699
rect 14093 12659 14151 12665
rect 11072 12600 12296 12628
rect 12437 12631 12495 12637
rect 10965 12591 11023 12597
rect 12437 12597 12449 12631
rect 12483 12597 12495 12631
rect 12437 12591 12495 12597
rect 12710 12588 12716 12640
rect 12768 12628 12774 12640
rect 12805 12631 12863 12637
rect 12805 12628 12817 12631
rect 12768 12600 12817 12628
rect 12768 12588 12774 12600
rect 12805 12597 12817 12600
rect 12851 12597 12863 12631
rect 12805 12591 12863 12597
rect 12897 12631 12955 12637
rect 12897 12597 12909 12631
rect 12943 12628 12955 12631
rect 13078 12628 13084 12640
rect 12943 12600 13084 12628
rect 12943 12597 12955 12600
rect 12897 12591 12955 12597
rect 13078 12588 13084 12600
rect 13136 12588 13142 12640
rect 13998 12628 14004 12640
rect 13959 12600 14004 12628
rect 13998 12588 14004 12600
rect 14056 12588 14062 12640
rect 1104 12538 15824 12560
rect 1104 12486 5912 12538
rect 5964 12486 5976 12538
rect 6028 12486 6040 12538
rect 6092 12486 6104 12538
rect 6156 12486 10843 12538
rect 10895 12486 10907 12538
rect 10959 12486 10971 12538
rect 11023 12486 11035 12538
rect 11087 12486 15824 12538
rect 1104 12464 15824 12486
rect 1578 12384 1584 12436
rect 1636 12424 1642 12436
rect 1673 12427 1731 12433
rect 1673 12424 1685 12427
rect 1636 12396 1685 12424
rect 1636 12384 1642 12396
rect 1673 12393 1685 12396
rect 1719 12393 1731 12427
rect 1673 12387 1731 12393
rect 4890 12384 4896 12436
rect 4948 12424 4954 12436
rect 5169 12427 5227 12433
rect 5169 12424 5181 12427
rect 4948 12396 5181 12424
rect 4948 12384 4954 12396
rect 5169 12393 5181 12396
rect 5215 12393 5227 12427
rect 5169 12387 5227 12393
rect 5626 12384 5632 12436
rect 5684 12424 5690 12436
rect 5905 12427 5963 12433
rect 5905 12424 5917 12427
rect 5684 12396 5917 12424
rect 5684 12384 5690 12396
rect 5905 12393 5917 12396
rect 5951 12393 5963 12427
rect 5905 12387 5963 12393
rect 6273 12427 6331 12433
rect 6273 12393 6285 12427
rect 6319 12424 6331 12427
rect 6454 12424 6460 12436
rect 6319 12396 6460 12424
rect 6319 12393 6331 12396
rect 6273 12387 6331 12393
rect 6454 12384 6460 12396
rect 6512 12384 6518 12436
rect 6638 12384 6644 12436
rect 6696 12424 6702 12436
rect 7098 12424 7104 12436
rect 6696 12396 7104 12424
rect 6696 12384 6702 12396
rect 7098 12384 7104 12396
rect 7156 12424 7162 12436
rect 7156 12396 8064 12424
rect 7156 12384 7162 12396
rect 2041 12359 2099 12365
rect 2041 12325 2053 12359
rect 2087 12356 2099 12359
rect 2682 12356 2688 12368
rect 2087 12328 2688 12356
rect 2087 12325 2099 12328
rect 2041 12319 2099 12325
rect 2682 12316 2688 12328
rect 2740 12316 2746 12368
rect 4154 12316 4160 12368
rect 4212 12356 4218 12368
rect 5077 12359 5135 12365
rect 5077 12356 5089 12359
rect 4212 12328 5089 12356
rect 4212 12316 4218 12328
rect 5077 12325 5089 12328
rect 5123 12325 5135 12359
rect 5077 12319 5135 12325
rect 5350 12316 5356 12368
rect 5408 12356 5414 12368
rect 6365 12359 6423 12365
rect 6365 12356 6377 12359
rect 5408 12328 6377 12356
rect 5408 12316 5414 12328
rect 6365 12325 6377 12328
rect 6411 12356 6423 12359
rect 6546 12356 6552 12368
rect 6411 12328 6552 12356
rect 6411 12325 6423 12328
rect 6365 12319 6423 12325
rect 6546 12316 6552 12328
rect 6604 12316 6610 12368
rect 7466 12356 7472 12368
rect 7427 12328 7472 12356
rect 7466 12316 7472 12328
rect 7524 12316 7530 12368
rect 8036 12356 8064 12396
rect 8754 12384 8760 12436
rect 8812 12424 8818 12436
rect 9306 12424 9312 12436
rect 8812 12396 9312 12424
rect 8812 12384 8818 12396
rect 9306 12384 9312 12396
rect 9364 12384 9370 12436
rect 9582 12384 9588 12436
rect 9640 12424 9646 12436
rect 9677 12427 9735 12433
rect 9677 12424 9689 12427
rect 9640 12396 9689 12424
rect 9640 12384 9646 12396
rect 9677 12393 9689 12396
rect 9723 12393 9735 12427
rect 9677 12387 9735 12393
rect 10045 12427 10103 12433
rect 10045 12393 10057 12427
rect 10091 12424 10103 12427
rect 10091 12396 10640 12424
rect 10091 12393 10103 12396
rect 10045 12387 10103 12393
rect 8036 12328 8156 12356
rect 2593 12291 2651 12297
rect 2593 12257 2605 12291
rect 2639 12288 2651 12291
rect 2774 12288 2780 12300
rect 2639 12260 2780 12288
rect 2639 12257 2651 12260
rect 2593 12251 2651 12257
rect 2774 12248 2780 12260
rect 2832 12248 2838 12300
rect 3329 12291 3387 12297
rect 3329 12257 3341 12291
rect 3375 12288 3387 12291
rect 7190 12288 7196 12300
rect 3375 12260 7196 12288
rect 3375 12257 3387 12260
rect 3329 12251 3387 12257
rect 7190 12248 7196 12260
rect 7248 12248 7254 12300
rect 7561 12291 7619 12297
rect 7561 12257 7573 12291
rect 7607 12288 7619 12291
rect 8018 12288 8024 12300
rect 7607 12260 8024 12288
rect 7607 12257 7619 12260
rect 7561 12251 7619 12257
rect 8018 12248 8024 12260
rect 8076 12248 8082 12300
rect 8128 12288 8156 12328
rect 8662 12316 8668 12368
rect 8720 12356 8726 12368
rect 9858 12356 9864 12368
rect 8720 12328 9864 12356
rect 8720 12316 8726 12328
rect 9858 12316 9864 12328
rect 9916 12356 9922 12368
rect 10137 12359 10195 12365
rect 10137 12356 10149 12359
rect 9916 12328 10149 12356
rect 9916 12316 9922 12328
rect 10137 12325 10149 12328
rect 10183 12325 10195 12359
rect 10612 12356 10640 12396
rect 10686 12384 10692 12436
rect 10744 12424 10750 12436
rect 10873 12427 10931 12433
rect 10873 12424 10885 12427
rect 10744 12396 10885 12424
rect 10744 12384 10750 12396
rect 10873 12393 10885 12396
rect 10919 12393 10931 12427
rect 10873 12387 10931 12393
rect 11241 12427 11299 12433
rect 11241 12393 11253 12427
rect 11287 12424 11299 12427
rect 11287 12396 12296 12424
rect 11287 12393 11299 12396
rect 11241 12387 11299 12393
rect 11606 12356 11612 12368
rect 10612 12328 11612 12356
rect 10137 12319 10195 12325
rect 11606 12316 11612 12328
rect 11664 12316 11670 12368
rect 12268 12356 12296 12396
rect 12342 12384 12348 12436
rect 12400 12424 12406 12436
rect 12529 12427 12587 12433
rect 12529 12424 12541 12427
rect 12400 12396 12541 12424
rect 12400 12384 12406 12396
rect 12529 12393 12541 12396
rect 12575 12393 12587 12427
rect 12529 12387 12587 12393
rect 13170 12384 13176 12436
rect 13228 12424 13234 12436
rect 13633 12427 13691 12433
rect 13633 12424 13645 12427
rect 13228 12396 13645 12424
rect 13228 12384 13234 12396
rect 13633 12393 13645 12396
rect 13679 12393 13691 12427
rect 13633 12387 13691 12393
rect 14458 12384 14464 12436
rect 14516 12424 14522 12436
rect 14645 12427 14703 12433
rect 14645 12424 14657 12427
rect 14516 12396 14657 12424
rect 14516 12384 14522 12396
rect 14645 12393 14657 12396
rect 14691 12393 14703 12427
rect 14645 12387 14703 12393
rect 14734 12384 14740 12436
rect 14792 12424 14798 12436
rect 15102 12424 15108 12436
rect 14792 12396 15108 12424
rect 14792 12384 14798 12396
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 15286 12356 15292 12368
rect 12268 12328 15292 12356
rect 15286 12316 15292 12328
rect 15344 12316 15350 12368
rect 10410 12288 10416 12300
rect 8128 12260 10416 12288
rect 10410 12248 10416 12260
rect 10468 12248 10474 12300
rect 11146 12248 11152 12300
rect 11204 12288 11210 12300
rect 11333 12291 11391 12297
rect 11333 12288 11345 12291
rect 11204 12260 11345 12288
rect 11204 12248 11210 12260
rect 11333 12257 11345 12260
rect 11379 12257 11391 12291
rect 11333 12251 11391 12257
rect 12158 12248 12164 12300
rect 12216 12288 12222 12300
rect 12434 12288 12440 12300
rect 12216 12260 12440 12288
rect 12216 12248 12222 12260
rect 12434 12248 12440 12260
rect 12492 12248 12498 12300
rect 13262 12288 13268 12300
rect 12544 12260 13268 12288
rect 2130 12220 2136 12232
rect 2091 12192 2136 12220
rect 2130 12180 2136 12192
rect 2188 12180 2194 12232
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12220 2375 12223
rect 4065 12223 4123 12229
rect 2363 12192 3004 12220
rect 2363 12189 2375 12192
rect 2317 12183 2375 12189
rect 2976 12084 3004 12192
rect 4065 12189 4077 12223
rect 4111 12220 4123 12223
rect 4433 12223 4491 12229
rect 4433 12220 4445 12223
rect 4111 12192 4445 12220
rect 4111 12189 4123 12192
rect 4065 12183 4123 12189
rect 4433 12189 4445 12192
rect 4479 12220 4491 12223
rect 4890 12220 4896 12232
rect 4479 12192 4896 12220
rect 4479 12189 4491 12192
rect 4433 12183 4491 12189
rect 4890 12180 4896 12192
rect 4948 12180 4954 12232
rect 5350 12220 5356 12232
rect 5311 12192 5356 12220
rect 5350 12180 5356 12192
rect 5408 12180 5414 12232
rect 5718 12180 5724 12232
rect 5776 12220 5782 12232
rect 6454 12220 6460 12232
rect 5776 12192 6460 12220
rect 5776 12180 5782 12192
rect 6454 12180 6460 12192
rect 6512 12180 6518 12232
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12220 6607 12223
rect 6638 12220 6644 12232
rect 6595 12192 6644 12220
rect 6595 12189 6607 12192
rect 6549 12183 6607 12189
rect 6638 12180 6644 12192
rect 6696 12180 6702 12232
rect 6914 12180 6920 12232
rect 6972 12220 6978 12232
rect 7653 12223 7711 12229
rect 7653 12220 7665 12223
rect 6972 12192 7665 12220
rect 6972 12180 6978 12192
rect 7653 12189 7665 12192
rect 7699 12189 7711 12223
rect 7653 12183 7711 12189
rect 8297 12223 8355 12229
rect 8297 12189 8309 12223
rect 8343 12220 8355 12223
rect 8846 12220 8852 12232
rect 8343 12192 8852 12220
rect 8343 12189 8355 12192
rect 8297 12183 8355 12189
rect 8846 12180 8852 12192
rect 8904 12180 8910 12232
rect 8941 12223 8999 12229
rect 8941 12189 8953 12223
rect 8987 12220 8999 12223
rect 9490 12220 9496 12232
rect 8987 12192 9496 12220
rect 8987 12189 8999 12192
rect 8941 12183 8999 12189
rect 9490 12180 9496 12192
rect 9548 12180 9554 12232
rect 9674 12180 9680 12232
rect 9732 12220 9738 12232
rect 10134 12220 10140 12232
rect 9732 12192 10140 12220
rect 9732 12180 9738 12192
rect 10134 12180 10140 12192
rect 10192 12180 10198 12232
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12189 10287 12223
rect 11425 12223 11483 12229
rect 11425 12220 11437 12223
rect 10229 12183 10287 12189
rect 10382 12192 11437 12220
rect 4338 12112 4344 12164
rect 4396 12152 4402 12164
rect 6730 12152 6736 12164
rect 4396 12124 6736 12152
rect 4396 12112 4402 12124
rect 6730 12112 6736 12124
rect 6788 12112 6794 12164
rect 7101 12155 7159 12161
rect 7101 12121 7113 12155
rect 7147 12152 7159 12155
rect 7834 12152 7840 12164
rect 7147 12124 7840 12152
rect 7147 12121 7159 12124
rect 7101 12115 7159 12121
rect 7834 12112 7840 12124
rect 7892 12112 7898 12164
rect 9030 12152 9036 12164
rect 7944 12124 9036 12152
rect 3786 12084 3792 12096
rect 2976 12056 3792 12084
rect 3786 12044 3792 12056
rect 3844 12044 3850 12096
rect 4709 12087 4767 12093
rect 4709 12053 4721 12087
rect 4755 12084 4767 12087
rect 7944 12084 7972 12124
rect 9030 12112 9036 12124
rect 9088 12112 9094 12164
rect 9306 12112 9312 12164
rect 9364 12152 9370 12164
rect 10244 12152 10272 12183
rect 10382 12152 10410 12192
rect 11425 12189 11437 12192
rect 11471 12189 11483 12223
rect 12544 12220 12572 12260
rect 13262 12248 13268 12260
rect 13320 12248 13326 12300
rect 13722 12288 13728 12300
rect 13683 12260 13728 12288
rect 13722 12248 13728 12260
rect 13780 12248 13786 12300
rect 14461 12291 14519 12297
rect 14461 12257 14473 12291
rect 14507 12288 14519 12291
rect 14734 12288 14740 12300
rect 14507 12260 14740 12288
rect 14507 12257 14519 12260
rect 14461 12251 14519 12257
rect 14734 12248 14740 12260
rect 14792 12288 14798 12300
rect 14918 12288 14924 12300
rect 14792 12260 14924 12288
rect 14792 12248 14798 12260
rect 14918 12248 14924 12260
rect 14976 12248 14982 12300
rect 11425 12183 11483 12189
rect 12176 12192 12572 12220
rect 12621 12223 12679 12229
rect 9364 12124 10410 12152
rect 9364 12112 9370 12124
rect 10502 12112 10508 12164
rect 10560 12152 10566 12164
rect 12069 12155 12127 12161
rect 12069 12152 12081 12155
rect 10560 12124 12081 12152
rect 10560 12112 10566 12124
rect 12069 12121 12081 12124
rect 12115 12121 12127 12155
rect 12069 12115 12127 12121
rect 4755 12056 7972 12084
rect 4755 12053 4767 12056
rect 4709 12047 4767 12053
rect 8018 12044 8024 12096
rect 8076 12084 8082 12096
rect 12176 12084 12204 12192
rect 12621 12189 12633 12223
rect 12667 12189 12679 12223
rect 13814 12220 13820 12232
rect 13775 12192 13820 12220
rect 12621 12183 12679 12189
rect 12434 12112 12440 12164
rect 12492 12152 12498 12164
rect 12636 12152 12664 12183
rect 13814 12180 13820 12192
rect 13872 12180 13878 12232
rect 12492 12124 12664 12152
rect 12492 12112 12498 12124
rect 13722 12112 13728 12164
rect 13780 12152 13786 12164
rect 13906 12152 13912 12164
rect 13780 12124 13912 12152
rect 13780 12112 13786 12124
rect 13906 12112 13912 12124
rect 13964 12112 13970 12164
rect 8076 12056 12204 12084
rect 8076 12044 8082 12056
rect 12342 12044 12348 12096
rect 12400 12084 12406 12096
rect 12526 12084 12532 12096
rect 12400 12056 12532 12084
rect 12400 12044 12406 12056
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 13265 12087 13323 12093
rect 13265 12053 13277 12087
rect 13311 12084 13323 12087
rect 13998 12084 14004 12096
rect 13311 12056 14004 12084
rect 13311 12053 13323 12056
rect 13265 12047 13323 12053
rect 13998 12044 14004 12056
rect 14056 12044 14062 12096
rect 1104 11994 15824 12016
rect 1104 11942 3447 11994
rect 3499 11942 3511 11994
rect 3563 11942 3575 11994
rect 3627 11942 3639 11994
rect 3691 11942 8378 11994
rect 8430 11942 8442 11994
rect 8494 11942 8506 11994
rect 8558 11942 8570 11994
rect 8622 11942 13308 11994
rect 13360 11942 13372 11994
rect 13424 11942 13436 11994
rect 13488 11942 13500 11994
rect 13552 11942 15824 11994
rect 1104 11920 15824 11942
rect 3326 11880 3332 11892
rect 3068 11852 3332 11880
rect 2774 11772 2780 11824
rect 2832 11812 2838 11824
rect 3068 11812 3096 11852
rect 3326 11840 3332 11852
rect 3384 11840 3390 11892
rect 6273 11883 6331 11889
rect 6273 11849 6285 11883
rect 6319 11880 6331 11883
rect 7558 11880 7564 11892
rect 6319 11852 7564 11880
rect 6319 11849 6331 11852
rect 6273 11843 6331 11849
rect 7558 11840 7564 11852
rect 7616 11840 7622 11892
rect 7834 11840 7840 11892
rect 7892 11880 7898 11892
rect 8205 11883 8263 11889
rect 8205 11880 8217 11883
rect 7892 11852 8217 11880
rect 7892 11840 7898 11852
rect 8205 11849 8217 11852
rect 8251 11880 8263 11883
rect 10042 11880 10048 11892
rect 8251 11852 8432 11880
rect 8251 11849 8263 11852
rect 8205 11843 8263 11849
rect 2832 11784 3096 11812
rect 2832 11772 2838 11784
rect 2501 11747 2559 11753
rect 2501 11713 2513 11747
rect 2547 11744 2559 11747
rect 2958 11744 2964 11756
rect 2547 11716 2964 11744
rect 2547 11713 2559 11716
rect 2501 11707 2559 11713
rect 2958 11704 2964 11716
rect 3016 11704 3022 11756
rect 3068 11753 3096 11784
rect 6362 11772 6368 11824
rect 6420 11812 6426 11824
rect 6420 11784 6868 11812
rect 6420 11772 6426 11784
rect 6840 11756 6868 11784
rect 3053 11747 3111 11753
rect 3053 11713 3065 11747
rect 3099 11713 3111 11747
rect 4522 11744 4528 11756
rect 3053 11707 3111 11713
rect 4264 11716 4528 11744
rect 2314 11676 2320 11688
rect 2275 11648 2320 11676
rect 2314 11636 2320 11648
rect 2372 11636 2378 11688
rect 3320 11679 3378 11685
rect 3320 11645 3332 11679
rect 3366 11676 3378 11679
rect 4062 11676 4068 11688
rect 3366 11648 4068 11676
rect 3366 11645 3378 11648
rect 3320 11639 3378 11645
rect 4062 11636 4068 11648
rect 4120 11636 4126 11688
rect 2406 11568 2412 11620
rect 2464 11608 2470 11620
rect 4264 11608 4292 11716
rect 4522 11704 4528 11716
rect 4580 11704 4586 11756
rect 4798 11704 4804 11756
rect 4856 11744 4862 11756
rect 4893 11747 4951 11753
rect 4893 11744 4905 11747
rect 4856 11716 4905 11744
rect 4856 11704 4862 11716
rect 4893 11713 4905 11716
rect 4939 11713 4951 11747
rect 6638 11744 6644 11756
rect 4893 11707 4951 11713
rect 5920 11716 6644 11744
rect 5920 11676 5948 11716
rect 6638 11704 6644 11716
rect 6696 11704 6702 11756
rect 6822 11744 6828 11756
rect 6783 11716 6828 11744
rect 6822 11704 6828 11716
rect 6880 11704 6886 11756
rect 8404 11744 8432 11852
rect 8496 11852 9628 11880
rect 10003 11852 10048 11880
rect 8496 11824 8524 11852
rect 8478 11772 8484 11824
rect 8536 11772 8542 11824
rect 9600 11812 9628 11852
rect 10042 11840 10048 11852
rect 10100 11840 10106 11892
rect 11146 11880 11152 11892
rect 10152 11852 11152 11880
rect 10152 11812 10180 11852
rect 11146 11840 11152 11852
rect 11204 11840 11210 11892
rect 11238 11840 11244 11892
rect 11296 11880 11302 11892
rect 11974 11880 11980 11892
rect 11296 11852 11980 11880
rect 11296 11840 11302 11852
rect 11974 11840 11980 11852
rect 12032 11880 12038 11892
rect 13078 11880 13084 11892
rect 12032 11852 13084 11880
rect 12032 11840 12038 11852
rect 13078 11840 13084 11852
rect 13136 11840 13142 11892
rect 10502 11812 10508 11824
rect 9600 11784 10180 11812
rect 10463 11784 10508 11812
rect 10502 11772 10508 11784
rect 10560 11772 10566 11824
rect 10962 11772 10968 11824
rect 11020 11812 11026 11824
rect 12437 11815 12495 11821
rect 12437 11812 12449 11815
rect 11020 11784 12449 11812
rect 11020 11772 11026 11784
rect 12437 11781 12449 11784
rect 12483 11781 12495 11815
rect 12437 11775 12495 11781
rect 12544 11784 13124 11812
rect 8404 11716 8800 11744
rect 2464 11580 4292 11608
rect 4356 11648 5948 11676
rect 2464 11568 2470 11580
rect 1578 11500 1584 11552
rect 1636 11540 1642 11552
rect 1857 11543 1915 11549
rect 1857 11540 1869 11543
rect 1636 11512 1869 11540
rect 1636 11500 1642 11512
rect 1857 11509 1869 11512
rect 1903 11509 1915 11543
rect 1857 11503 1915 11509
rect 2225 11543 2283 11549
rect 2225 11509 2237 11543
rect 2271 11540 2283 11543
rect 4356 11540 4384 11648
rect 6270 11636 6276 11688
rect 6328 11676 6334 11688
rect 7081 11679 7139 11685
rect 7081 11676 7093 11679
rect 6328 11648 7093 11676
rect 6328 11636 6334 11648
rect 7081 11645 7093 11648
rect 7127 11645 7139 11679
rect 7081 11639 7139 11645
rect 8110 11636 8116 11688
rect 8168 11676 8174 11688
rect 8478 11676 8484 11688
rect 8168 11648 8484 11676
rect 8168 11636 8174 11648
rect 8478 11636 8484 11648
rect 8536 11636 8542 11688
rect 8665 11679 8723 11685
rect 8665 11645 8677 11679
rect 8711 11645 8723 11679
rect 8772 11676 8800 11716
rect 9674 11704 9680 11756
rect 9732 11744 9738 11756
rect 11057 11747 11115 11753
rect 11057 11744 11069 11747
rect 9732 11716 11069 11744
rect 9732 11704 9738 11716
rect 11057 11713 11069 11716
rect 11103 11713 11115 11747
rect 11057 11707 11115 11713
rect 11146 11704 11152 11756
rect 11204 11744 11210 11756
rect 12544 11744 12572 11784
rect 12986 11744 12992 11756
rect 11204 11716 12572 11744
rect 12947 11716 12992 11744
rect 11204 11704 11210 11716
rect 12986 11704 12992 11716
rect 13044 11704 13050 11756
rect 13096 11744 13124 11784
rect 14185 11747 14243 11753
rect 14185 11744 14197 11747
rect 13096 11716 14197 11744
rect 14185 11713 14197 11716
rect 14231 11713 14243 11747
rect 14185 11707 14243 11713
rect 8938 11685 8944 11688
rect 8921 11679 8944 11685
rect 8921 11676 8933 11679
rect 8772 11648 8933 11676
rect 8665 11639 8723 11645
rect 8921 11645 8933 11648
rect 8996 11676 9002 11688
rect 8996 11648 9069 11676
rect 8921 11639 8944 11645
rect 4798 11568 4804 11620
rect 4856 11608 4862 11620
rect 5166 11617 5172 11620
rect 5138 11611 5172 11617
rect 5138 11608 5150 11611
rect 4856 11580 5150 11608
rect 4856 11568 4862 11580
rect 5138 11577 5150 11580
rect 5224 11608 5230 11620
rect 5224 11580 5286 11608
rect 5138 11571 5172 11577
rect 5166 11568 5172 11571
rect 5224 11568 5230 11580
rect 7926 11568 7932 11620
rect 7984 11608 7990 11620
rect 8680 11608 8708 11639
rect 8938 11636 8944 11639
rect 8996 11636 9002 11648
rect 10226 11636 10232 11688
rect 10284 11676 10290 11688
rect 10284 11648 11008 11676
rect 10284 11636 10290 11648
rect 9582 11608 9588 11620
rect 7984 11580 9588 11608
rect 7984 11568 7990 11580
rect 9582 11568 9588 11580
rect 9640 11608 9646 11620
rect 10318 11608 10324 11620
rect 9640 11580 10324 11608
rect 9640 11568 9646 11580
rect 10318 11568 10324 11580
rect 10376 11568 10382 11620
rect 10870 11608 10876 11620
rect 10831 11580 10876 11608
rect 10870 11568 10876 11580
rect 10928 11568 10934 11620
rect 10980 11608 11008 11648
rect 11422 11636 11428 11688
rect 11480 11676 11486 11688
rect 12897 11679 12955 11685
rect 12897 11676 12909 11679
rect 11480 11648 12909 11676
rect 11480 11636 11486 11648
rect 12897 11645 12909 11648
rect 12943 11645 12955 11679
rect 13998 11676 14004 11688
rect 13959 11648 14004 11676
rect 12897 11639 12955 11645
rect 13998 11636 14004 11648
rect 14056 11636 14062 11688
rect 14826 11676 14832 11688
rect 14787 11648 14832 11676
rect 14826 11636 14832 11648
rect 14884 11636 14890 11688
rect 14366 11608 14372 11620
rect 10980 11580 14372 11608
rect 14366 11568 14372 11580
rect 14424 11568 14430 11620
rect 2271 11512 4384 11540
rect 4433 11543 4491 11549
rect 2271 11509 2283 11512
rect 2225 11503 2283 11509
rect 4433 11509 4445 11543
rect 4479 11540 4491 11543
rect 8110 11540 8116 11552
rect 4479 11512 8116 11540
rect 4479 11509 4491 11512
rect 4433 11503 4491 11509
rect 8110 11500 8116 11512
rect 8168 11540 8174 11552
rect 9674 11540 9680 11552
rect 8168 11512 9680 11540
rect 8168 11500 8174 11512
rect 9674 11500 9680 11512
rect 9732 11500 9738 11552
rect 10965 11543 11023 11549
rect 10965 11509 10977 11543
rect 11011 11540 11023 11543
rect 11238 11540 11244 11552
rect 11011 11512 11244 11540
rect 11011 11509 11023 11512
rect 10965 11503 11023 11509
rect 11238 11500 11244 11512
rect 11296 11500 11302 11552
rect 11701 11543 11759 11549
rect 11701 11509 11713 11543
rect 11747 11540 11759 11543
rect 12618 11540 12624 11552
rect 11747 11512 12624 11540
rect 11747 11509 11759 11512
rect 11701 11503 11759 11509
rect 12618 11500 12624 11512
rect 12676 11500 12682 11552
rect 12805 11543 12863 11549
rect 12805 11509 12817 11543
rect 12851 11540 12863 11543
rect 13170 11540 13176 11552
rect 12851 11512 13176 11540
rect 12851 11509 12863 11512
rect 12805 11503 12863 11509
rect 13170 11500 13176 11512
rect 13228 11500 13234 11552
rect 13630 11540 13636 11552
rect 13591 11512 13636 11540
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 14090 11500 14096 11552
rect 14148 11540 14154 11552
rect 14148 11512 14193 11540
rect 14148 11500 14154 11512
rect 14458 11500 14464 11552
rect 14516 11540 14522 11552
rect 15013 11543 15071 11549
rect 15013 11540 15025 11543
rect 14516 11512 15025 11540
rect 14516 11500 14522 11512
rect 15013 11509 15025 11512
rect 15059 11509 15071 11543
rect 15013 11503 15071 11509
rect 1104 11450 15824 11472
rect 1104 11398 5912 11450
rect 5964 11398 5976 11450
rect 6028 11398 6040 11450
rect 6092 11398 6104 11450
rect 6156 11398 10843 11450
rect 10895 11398 10907 11450
rect 10959 11398 10971 11450
rect 11023 11398 11035 11450
rect 11087 11398 15824 11450
rect 1104 11376 15824 11398
rect 1596 11308 5203 11336
rect 1596 11209 1624 11308
rect 1854 11268 1860 11280
rect 1815 11240 1860 11268
rect 1854 11228 1860 11240
rect 1912 11228 1918 11280
rect 2774 11268 2780 11280
rect 2148 11240 2780 11268
rect 2148 11209 2176 11240
rect 2774 11228 2780 11240
rect 2832 11268 2838 11280
rect 2832 11240 3280 11268
rect 2832 11228 2838 11240
rect 2406 11209 2412 11212
rect 1581 11203 1639 11209
rect 1581 11169 1593 11203
rect 1627 11169 1639 11203
rect 1581 11163 1639 11169
rect 2133 11203 2191 11209
rect 2133 11169 2145 11203
rect 2179 11169 2191 11203
rect 2133 11163 2191 11169
rect 2400 11163 2412 11209
rect 2464 11200 2470 11212
rect 2464 11172 2500 11200
rect 2406 11160 2412 11163
rect 2464 11160 2470 11172
rect 2958 11160 2964 11212
rect 3016 11200 3022 11212
rect 3016 11172 3188 11200
rect 3016 11160 3022 11172
rect 3160 11064 3188 11172
rect 3252 11132 3280 11240
rect 4430 11228 4436 11280
rect 4488 11228 4494 11280
rect 5175 11268 5203 11308
rect 5258 11296 5264 11348
rect 5316 11336 5322 11348
rect 5442 11336 5448 11348
rect 5316 11308 5448 11336
rect 5316 11296 5322 11308
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 5810 11296 5816 11348
rect 5868 11336 5874 11348
rect 6089 11339 6147 11345
rect 6089 11336 6101 11339
rect 5868 11308 6101 11336
rect 5868 11296 5874 11308
rect 6089 11305 6101 11308
rect 6135 11305 6147 11339
rect 6089 11299 6147 11305
rect 7650 11296 7656 11348
rect 7708 11336 7714 11348
rect 7745 11339 7803 11345
rect 7745 11336 7757 11339
rect 7708 11308 7757 11336
rect 7708 11296 7714 11308
rect 7745 11305 7757 11308
rect 7791 11305 7803 11339
rect 7745 11299 7803 11305
rect 8018 11296 8024 11348
rect 8076 11336 8082 11348
rect 8205 11339 8263 11345
rect 8205 11336 8217 11339
rect 8076 11308 8217 11336
rect 8076 11296 8082 11308
rect 8205 11305 8217 11308
rect 8251 11305 8263 11339
rect 8205 11299 8263 11305
rect 8754 11296 8760 11348
rect 8812 11336 8818 11348
rect 8849 11339 8907 11345
rect 8849 11336 8861 11339
rect 8812 11308 8861 11336
rect 8812 11296 8818 11308
rect 8849 11305 8861 11308
rect 8895 11305 8907 11339
rect 11517 11339 11575 11345
rect 8849 11299 8907 11305
rect 9140 11308 11008 11336
rect 5994 11268 6000 11280
rect 5175 11240 6000 11268
rect 5994 11228 6000 11240
rect 6052 11228 6058 11280
rect 6610 11271 6668 11277
rect 6610 11268 6622 11271
rect 6095 11240 6622 11268
rect 3694 11160 3700 11212
rect 3752 11200 3758 11212
rect 4321 11203 4379 11209
rect 4321 11200 4333 11203
rect 3752 11172 4333 11200
rect 3752 11160 3758 11172
rect 4321 11169 4333 11172
rect 4367 11169 4379 11203
rect 4448 11200 4476 11228
rect 4614 11200 4620 11212
rect 4448 11172 4620 11200
rect 4321 11163 4379 11169
rect 4614 11160 4620 11172
rect 4672 11200 4678 11212
rect 6095 11200 6123 11240
rect 6610 11237 6622 11240
rect 6656 11268 6668 11271
rect 6730 11268 6736 11280
rect 6656 11240 6736 11268
rect 6656 11237 6668 11240
rect 6610 11231 6668 11237
rect 6730 11228 6736 11240
rect 6788 11228 6794 11280
rect 8294 11228 8300 11280
rect 8352 11268 8358 11280
rect 9140 11268 9168 11308
rect 10980 11280 11008 11308
rect 11517 11305 11529 11339
rect 11563 11336 11575 11339
rect 11790 11336 11796 11348
rect 11563 11308 11796 11336
rect 11563 11305 11575 11308
rect 11517 11299 11575 11305
rect 11790 11296 11796 11308
rect 11848 11296 11854 11348
rect 12342 11296 12348 11348
rect 12400 11336 12406 11348
rect 12713 11339 12771 11345
rect 12713 11336 12725 11339
rect 12400 11308 12725 11336
rect 12400 11296 12406 11308
rect 12713 11305 12725 11308
rect 12759 11305 12771 11339
rect 12713 11299 12771 11305
rect 12894 11296 12900 11348
rect 12952 11336 12958 11348
rect 13081 11339 13139 11345
rect 13081 11336 13093 11339
rect 12952 11308 13093 11336
rect 12952 11296 12958 11308
rect 13081 11305 13093 11308
rect 13127 11305 13139 11339
rect 13081 11299 13139 11305
rect 13909 11339 13967 11345
rect 13909 11305 13921 11339
rect 13955 11336 13967 11339
rect 14090 11336 14096 11348
rect 13955 11308 14096 11336
rect 13955 11305 13967 11308
rect 13909 11299 13967 11305
rect 14090 11296 14096 11308
rect 14148 11296 14154 11348
rect 14366 11336 14372 11348
rect 14327 11308 14372 11336
rect 14366 11296 14372 11308
rect 14424 11296 14430 11348
rect 8352 11240 9168 11268
rect 8352 11228 8358 11240
rect 9214 11228 9220 11280
rect 9272 11268 9278 11280
rect 9674 11268 9680 11280
rect 9272 11240 9680 11268
rect 9272 11228 9278 11240
rect 9674 11228 9680 11240
rect 9732 11228 9738 11280
rect 10042 11268 10048 11280
rect 9784 11240 10048 11268
rect 4672 11172 6123 11200
rect 6273 11203 6331 11209
rect 4672 11160 4678 11172
rect 6273 11169 6285 11203
rect 6319 11200 6331 11203
rect 8662 11200 8668 11212
rect 6319 11172 8668 11200
rect 6319 11169 6331 11172
rect 6273 11163 6331 11169
rect 8662 11160 8668 11172
rect 8720 11160 8726 11212
rect 9784 11200 9812 11240
rect 10042 11228 10048 11240
rect 10100 11228 10106 11280
rect 10962 11228 10968 11280
rect 11020 11228 11026 11280
rect 11054 11228 11060 11280
rect 11112 11268 11118 11280
rect 11885 11271 11943 11277
rect 11885 11268 11897 11271
rect 11112 11240 11897 11268
rect 11112 11228 11118 11240
rect 11885 11237 11897 11240
rect 11931 11237 11943 11271
rect 11885 11231 11943 11237
rect 11977 11271 12035 11277
rect 11977 11237 11989 11271
rect 12023 11268 12035 11271
rect 15194 11268 15200 11280
rect 12023 11240 15200 11268
rect 12023 11237 12035 11240
rect 11977 11231 12035 11237
rect 14384 11212 14412 11240
rect 15194 11228 15200 11240
rect 15252 11228 15258 11280
rect 8864 11172 9812 11200
rect 9944 11203 10002 11209
rect 4062 11132 4068 11144
rect 3252 11104 4068 11132
rect 4062 11092 4068 11104
rect 4120 11092 4126 11144
rect 6362 11132 6368 11144
rect 6323 11104 6368 11132
rect 6362 11092 6368 11104
rect 6420 11092 6426 11144
rect 7466 11092 7472 11144
rect 7524 11132 7530 11144
rect 8864 11132 8892 11172
rect 9944 11169 9956 11203
rect 9990 11200 10002 11203
rect 10410 11200 10416 11212
rect 9990 11172 10416 11200
rect 9990 11169 10002 11172
rect 9944 11163 10002 11169
rect 10410 11160 10416 11172
rect 10468 11200 10474 11212
rect 12434 11200 12440 11212
rect 10468 11172 12440 11200
rect 10468 11160 10474 11172
rect 12434 11160 12440 11172
rect 12492 11160 12498 11212
rect 13078 11160 13084 11212
rect 13136 11200 13142 11212
rect 13173 11203 13231 11209
rect 13173 11200 13185 11203
rect 13136 11172 13185 11200
rect 13136 11160 13142 11172
rect 13173 11169 13185 11172
rect 13219 11169 13231 11203
rect 14274 11200 14280 11212
rect 14235 11172 14280 11200
rect 13173 11163 13231 11169
rect 14274 11160 14280 11172
rect 14332 11160 14338 11212
rect 14366 11160 14372 11212
rect 14424 11160 14430 11212
rect 7524 11104 8892 11132
rect 7524 11092 7530 11104
rect 9582 11092 9588 11144
rect 9640 11132 9646 11144
rect 9677 11135 9735 11141
rect 9677 11132 9689 11135
rect 9640 11104 9689 11132
rect 9640 11092 9646 11104
rect 9677 11101 9689 11104
rect 9723 11101 9735 11135
rect 9677 11095 9735 11101
rect 10962 11092 10968 11144
rect 11020 11132 11026 11144
rect 12069 11135 12127 11141
rect 12069 11132 12081 11135
rect 11020 11104 12081 11132
rect 11020 11092 11026 11104
rect 12069 11101 12081 11104
rect 12115 11101 12127 11135
rect 12069 11095 12127 11101
rect 12342 11092 12348 11144
rect 12400 11132 12406 11144
rect 13265 11135 13323 11141
rect 13265 11132 13277 11135
rect 12400 11104 13277 11132
rect 12400 11092 12406 11104
rect 13265 11101 13277 11104
rect 13311 11101 13323 11135
rect 13265 11095 13323 11101
rect 14461 11135 14519 11141
rect 14461 11101 14473 11135
rect 14507 11101 14519 11135
rect 14461 11095 14519 11101
rect 3326 11064 3332 11076
rect 3160 11036 3332 11064
rect 3326 11024 3332 11036
rect 3384 11064 3390 11076
rect 3513 11067 3571 11073
rect 3513 11064 3525 11067
rect 3384 11036 3525 11064
rect 3384 11024 3390 11036
rect 3513 11033 3525 11036
rect 3559 11033 3571 11067
rect 3513 11027 3571 11033
rect 5074 11024 5080 11076
rect 5132 11064 5138 11076
rect 5350 11064 5356 11076
rect 5132 11036 5356 11064
rect 5132 11024 5138 11036
rect 5350 11024 5356 11036
rect 5408 11024 5414 11076
rect 13814 11064 13820 11076
rect 7484 11036 9720 11064
rect 3970 10956 3976 11008
rect 4028 10996 4034 11008
rect 5166 10996 5172 11008
rect 4028 10968 5172 10996
rect 4028 10956 4034 10968
rect 5166 10956 5172 10968
rect 5224 10956 5230 11008
rect 5442 10956 5448 11008
rect 5500 10996 5506 11008
rect 7484 10996 7512 11036
rect 5500 10968 7512 10996
rect 5500 10956 5506 10968
rect 8018 10956 8024 11008
rect 8076 10996 8082 11008
rect 9214 10996 9220 11008
rect 8076 10968 9220 10996
rect 8076 10956 8082 10968
rect 9214 10956 9220 10968
rect 9272 10956 9278 11008
rect 9692 10996 9720 11036
rect 10888 11036 13820 11064
rect 10888 10996 10916 11036
rect 13814 11024 13820 11036
rect 13872 11064 13878 11076
rect 14476 11064 14504 11095
rect 13872 11036 14504 11064
rect 13872 11024 13878 11036
rect 9692 10968 10916 10996
rect 10962 10956 10968 11008
rect 11020 10996 11026 11008
rect 11057 10999 11115 11005
rect 11057 10996 11069 10999
rect 11020 10968 11069 10996
rect 11020 10956 11026 10968
rect 11057 10965 11069 10968
rect 11103 10965 11115 10999
rect 11057 10959 11115 10965
rect 11146 10956 11152 11008
rect 11204 10996 11210 11008
rect 11790 10996 11796 11008
rect 11204 10968 11796 10996
rect 11204 10956 11210 10968
rect 11790 10956 11796 10968
rect 11848 10956 11854 11008
rect 13722 10956 13728 11008
rect 13780 10996 13786 11008
rect 14550 10996 14556 11008
rect 13780 10968 14556 10996
rect 13780 10956 13786 10968
rect 14550 10956 14556 10968
rect 14608 10956 14614 11008
rect 1104 10906 15824 10928
rect 1104 10854 3447 10906
rect 3499 10854 3511 10906
rect 3563 10854 3575 10906
rect 3627 10854 3639 10906
rect 3691 10854 8378 10906
rect 8430 10854 8442 10906
rect 8494 10854 8506 10906
rect 8558 10854 8570 10906
rect 8622 10854 13308 10906
rect 13360 10854 13372 10906
rect 13424 10854 13436 10906
rect 13488 10854 13500 10906
rect 13552 10854 15824 10906
rect 1104 10832 15824 10854
rect 1581 10795 1639 10801
rect 1581 10761 1593 10795
rect 1627 10792 1639 10795
rect 1670 10792 1676 10804
rect 1627 10764 1676 10792
rect 1627 10761 1639 10764
rect 1581 10755 1639 10761
rect 1670 10752 1676 10764
rect 1728 10752 1734 10804
rect 1857 10795 1915 10801
rect 1857 10761 1869 10795
rect 1903 10792 1915 10795
rect 2130 10792 2136 10804
rect 1903 10764 2136 10792
rect 1903 10761 1915 10764
rect 1857 10755 1915 10761
rect 2130 10752 2136 10764
rect 2188 10752 2194 10804
rect 2958 10752 2964 10804
rect 3016 10792 3022 10804
rect 4433 10795 4491 10801
rect 3016 10764 4384 10792
rect 3016 10752 3022 10764
rect 4356 10724 4384 10764
rect 4433 10761 4445 10795
rect 4479 10792 4491 10795
rect 5166 10792 5172 10804
rect 4479 10764 5172 10792
rect 4479 10761 4491 10764
rect 4433 10755 4491 10761
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 6270 10792 6276 10804
rect 5592 10764 6276 10792
rect 5592 10752 5598 10764
rect 6270 10752 6276 10764
rect 6328 10752 6334 10804
rect 6362 10752 6368 10804
rect 6420 10792 6426 10804
rect 12986 10792 12992 10804
rect 6420 10764 12992 10792
rect 6420 10752 6426 10764
rect 12986 10752 12992 10764
rect 13044 10752 13050 10804
rect 4522 10724 4528 10736
rect 4356 10696 4528 10724
rect 4522 10684 4528 10696
rect 4580 10684 4586 10736
rect 7834 10684 7840 10736
rect 7892 10724 7898 10736
rect 8205 10727 8263 10733
rect 8205 10724 8217 10727
rect 7892 10696 8217 10724
rect 7892 10684 7898 10696
rect 8205 10693 8217 10696
rect 8251 10693 8263 10727
rect 8205 10687 8263 10693
rect 9674 10684 9680 10736
rect 9732 10724 9738 10736
rect 10045 10727 10103 10733
rect 10045 10724 10057 10727
rect 9732 10696 10057 10724
rect 9732 10684 9738 10696
rect 10045 10693 10057 10696
rect 10091 10724 10103 10727
rect 10502 10724 10508 10736
rect 10091 10696 10508 10724
rect 10091 10693 10103 10696
rect 10045 10687 10103 10693
rect 10502 10684 10508 10696
rect 10560 10684 10566 10736
rect 11885 10727 11943 10733
rect 11885 10693 11897 10727
rect 11931 10724 11943 10727
rect 12066 10724 12072 10736
rect 11931 10696 12072 10724
rect 11931 10693 11943 10696
rect 11885 10687 11943 10693
rect 12066 10684 12072 10696
rect 12124 10684 12130 10736
rect 15013 10727 15071 10733
rect 15013 10724 15025 10727
rect 12176 10696 15025 10724
rect 2498 10656 2504 10668
rect 2459 10628 2504 10656
rect 2498 10616 2504 10628
rect 2556 10616 2562 10668
rect 2774 10616 2780 10668
rect 2832 10656 2838 10668
rect 3053 10659 3111 10665
rect 3053 10656 3065 10659
rect 2832 10628 3065 10656
rect 2832 10616 2838 10628
rect 3053 10625 3065 10628
rect 3099 10625 3111 10659
rect 3053 10619 3111 10625
rect 4062 10616 4068 10668
rect 4120 10656 4126 10668
rect 4893 10659 4951 10665
rect 4893 10656 4905 10659
rect 4120 10628 4905 10656
rect 4120 10616 4126 10628
rect 4893 10625 4905 10628
rect 4939 10625 4951 10659
rect 6822 10656 6828 10668
rect 6783 10628 6828 10656
rect 4893 10619 4951 10625
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 7926 10616 7932 10668
rect 7984 10656 7990 10668
rect 8665 10659 8723 10665
rect 8665 10656 8677 10659
rect 7984 10628 8677 10656
rect 7984 10616 7990 10628
rect 8665 10625 8677 10628
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 11606 10616 11612 10668
rect 11664 10656 11670 10668
rect 11974 10656 11980 10668
rect 11664 10628 11980 10656
rect 11664 10616 11670 10628
rect 11974 10616 11980 10628
rect 12032 10616 12038 10668
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 1670 10588 1676 10600
rect 1443 10560 1676 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 1670 10548 1676 10560
rect 1728 10548 1734 10600
rect 2225 10591 2283 10597
rect 2225 10557 2237 10591
rect 2271 10588 2283 10591
rect 8202 10588 8208 10600
rect 2271 10560 8208 10588
rect 2271 10557 2283 10560
rect 2225 10551 2283 10557
rect 8202 10548 8208 10560
rect 8260 10548 8266 10600
rect 10318 10548 10324 10600
rect 10376 10588 10382 10600
rect 10505 10591 10563 10597
rect 10505 10588 10517 10591
rect 10376 10560 10517 10588
rect 10376 10548 10382 10560
rect 10505 10557 10517 10560
rect 10551 10557 10563 10591
rect 12176 10588 12204 10696
rect 15013 10693 15025 10696
rect 15059 10693 15071 10727
rect 15013 10687 15071 10693
rect 12986 10656 12992 10668
rect 12947 10628 12992 10656
rect 12986 10616 12992 10628
rect 13044 10616 13050 10668
rect 13078 10616 13084 10668
rect 13136 10656 13142 10668
rect 13354 10656 13360 10668
rect 13136 10628 13360 10656
rect 13136 10616 13142 10628
rect 13354 10616 13360 10628
rect 13412 10616 13418 10668
rect 13814 10616 13820 10668
rect 13872 10656 13878 10668
rect 14185 10659 14243 10665
rect 14185 10656 14197 10659
rect 13872 10628 14197 10656
rect 13872 10616 13878 10628
rect 14185 10625 14197 10628
rect 14231 10625 14243 10659
rect 14185 10619 14243 10625
rect 10505 10551 10563 10557
rect 10704 10560 12204 10588
rect 3320 10523 3378 10529
rect 3320 10489 3332 10523
rect 3366 10520 3378 10523
rect 5160 10523 5218 10529
rect 3366 10492 4476 10520
rect 3366 10489 3378 10492
rect 3320 10483 3378 10489
rect 4448 10464 4476 10492
rect 5160 10489 5172 10523
rect 5206 10520 5218 10523
rect 5258 10520 5264 10532
rect 5206 10492 5264 10520
rect 5206 10489 5218 10492
rect 5160 10483 5218 10489
rect 5258 10480 5264 10492
rect 5316 10480 5322 10532
rect 5350 10480 5356 10532
rect 5408 10520 5414 10532
rect 7092 10523 7150 10529
rect 5408 10492 6500 10520
rect 5408 10480 5414 10492
rect 2314 10412 2320 10464
rect 2372 10452 2378 10464
rect 2372 10424 2417 10452
rect 2372 10412 2378 10424
rect 4430 10412 4436 10464
rect 4488 10452 4494 10464
rect 6362 10452 6368 10464
rect 4488 10424 6368 10452
rect 4488 10412 4494 10424
rect 6362 10412 6368 10424
rect 6420 10412 6426 10464
rect 6472 10452 6500 10492
rect 7092 10489 7104 10523
rect 7138 10520 7150 10523
rect 7374 10520 7380 10532
rect 7138 10492 7380 10520
rect 7138 10489 7150 10492
rect 7092 10483 7150 10489
rect 7374 10480 7380 10492
rect 7432 10480 7438 10532
rect 8910 10523 8968 10529
rect 8910 10489 8922 10523
rect 8956 10489 8968 10523
rect 8910 10483 8968 10489
rect 8925 10452 8953 10483
rect 9766 10480 9772 10532
rect 9824 10520 9830 10532
rect 10594 10520 10600 10532
rect 9824 10492 10600 10520
rect 9824 10480 9830 10492
rect 10594 10480 10600 10492
rect 10652 10480 10658 10532
rect 6472 10424 8953 10452
rect 9214 10412 9220 10464
rect 9272 10452 9278 10464
rect 10704 10452 10732 10560
rect 12894 10548 12900 10600
rect 12952 10588 12958 10600
rect 14001 10591 14059 10597
rect 14001 10588 14013 10591
rect 12952 10560 14013 10588
rect 12952 10548 12958 10560
rect 14001 10557 14013 10560
rect 14047 10557 14059 10591
rect 14001 10551 14059 10557
rect 14274 10548 14280 10600
rect 14332 10588 14338 10600
rect 14829 10591 14887 10597
rect 14829 10588 14841 10591
rect 14332 10560 14841 10588
rect 14332 10548 14338 10560
rect 14829 10557 14841 10560
rect 14875 10588 14887 10591
rect 15930 10588 15936 10600
rect 14875 10560 15936 10588
rect 14875 10557 14887 10560
rect 14829 10551 14887 10557
rect 15930 10548 15936 10560
rect 15988 10548 15994 10600
rect 10778 10529 10784 10532
rect 10772 10483 10784 10529
rect 10836 10520 10842 10532
rect 12342 10520 12348 10532
rect 10836 10492 12348 10520
rect 10778 10480 10784 10483
rect 10836 10480 10842 10492
rect 12342 10480 12348 10492
rect 12400 10480 12406 10532
rect 12805 10523 12863 10529
rect 12805 10489 12817 10523
rect 12851 10520 12863 10523
rect 13262 10520 13268 10532
rect 12851 10492 13268 10520
rect 12851 10489 12863 10492
rect 12805 10483 12863 10489
rect 13262 10480 13268 10492
rect 13320 10480 13326 10532
rect 13354 10480 13360 10532
rect 13412 10520 13418 10532
rect 14093 10523 14151 10529
rect 14093 10520 14105 10523
rect 13412 10492 14105 10520
rect 13412 10480 13418 10492
rect 14093 10489 14105 10492
rect 14139 10489 14151 10523
rect 14093 10483 14151 10489
rect 9272 10424 10732 10452
rect 9272 10412 9278 10424
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12894 10452 12900 10464
rect 12492 10424 12537 10452
rect 12855 10424 12900 10452
rect 12492 10412 12498 10424
rect 12894 10412 12900 10424
rect 12952 10412 12958 10464
rect 13633 10455 13691 10461
rect 13633 10421 13645 10455
rect 13679 10452 13691 10455
rect 13906 10452 13912 10464
rect 13679 10424 13912 10452
rect 13679 10421 13691 10424
rect 13633 10415 13691 10421
rect 13906 10412 13912 10424
rect 13964 10412 13970 10464
rect 1104 10362 15824 10384
rect 1104 10310 5912 10362
rect 5964 10310 5976 10362
rect 6028 10310 6040 10362
rect 6092 10310 6104 10362
rect 6156 10310 10843 10362
rect 10895 10310 10907 10362
rect 10959 10310 10971 10362
rect 11023 10310 11035 10362
rect 11087 10310 15824 10362
rect 1104 10288 15824 10310
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10248 1639 10251
rect 4522 10248 4528 10260
rect 1627 10220 4528 10248
rect 1627 10217 1639 10220
rect 1581 10211 1639 10217
rect 4522 10208 4528 10220
rect 4580 10208 4586 10260
rect 5442 10248 5448 10260
rect 5403 10220 5448 10248
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 10502 10248 10508 10260
rect 6104 10220 10508 10248
rect 2400 10183 2458 10189
rect 2400 10149 2412 10183
rect 2446 10180 2458 10183
rect 2498 10180 2504 10192
rect 2446 10152 2504 10180
rect 2446 10149 2458 10152
rect 2400 10143 2458 10149
rect 2498 10140 2504 10152
rect 2556 10140 2562 10192
rect 2682 10140 2688 10192
rect 2740 10180 2746 10192
rect 6104 10180 6132 10220
rect 10502 10208 10508 10220
rect 10560 10208 10566 10260
rect 10686 10208 10692 10260
rect 10744 10248 10750 10260
rect 11057 10251 11115 10257
rect 11057 10248 11069 10251
rect 10744 10220 11069 10248
rect 10744 10208 10750 10220
rect 11057 10217 11069 10220
rect 11103 10217 11115 10251
rect 11057 10211 11115 10217
rect 11517 10251 11575 10257
rect 11517 10217 11529 10251
rect 11563 10217 11575 10251
rect 11517 10211 11575 10217
rect 11885 10251 11943 10257
rect 11885 10217 11897 10251
rect 11931 10248 11943 10251
rect 12158 10248 12164 10260
rect 11931 10220 12164 10248
rect 11931 10217 11943 10220
rect 11885 10211 11943 10217
rect 2740 10152 6132 10180
rect 6172 10183 6230 10189
rect 2740 10140 2746 10152
rect 6172 10149 6184 10183
rect 6218 10180 6230 10183
rect 6270 10180 6276 10192
rect 6218 10152 6276 10180
rect 6218 10149 6230 10152
rect 6172 10143 6230 10149
rect 6270 10140 6276 10152
rect 6328 10140 6334 10192
rect 8012 10183 8070 10189
rect 8012 10149 8024 10183
rect 8058 10180 8070 10183
rect 8110 10180 8116 10192
rect 8058 10152 8116 10180
rect 8058 10149 8070 10152
rect 8012 10143 8070 10149
rect 8110 10140 8116 10152
rect 8168 10140 8174 10192
rect 8662 10140 8668 10192
rect 8720 10180 8726 10192
rect 11532 10180 11560 10211
rect 12158 10208 12164 10220
rect 12216 10248 12222 10260
rect 12342 10248 12348 10260
rect 12216 10220 12348 10248
rect 12216 10208 12222 10220
rect 12342 10208 12348 10220
rect 12400 10208 12406 10260
rect 12434 10208 12440 10260
rect 12492 10248 12498 10260
rect 13173 10251 13231 10257
rect 13173 10248 13185 10251
rect 12492 10220 13185 10248
rect 12492 10208 12498 10220
rect 13173 10217 13185 10220
rect 13219 10217 13231 10251
rect 13173 10211 13231 10217
rect 13909 10251 13967 10257
rect 13909 10217 13921 10251
rect 13955 10248 13967 10251
rect 13998 10248 14004 10260
rect 13955 10220 14004 10248
rect 13955 10217 13967 10220
rect 13909 10211 13967 10217
rect 13998 10208 14004 10220
rect 14056 10208 14062 10260
rect 14277 10183 14335 10189
rect 14277 10180 14289 10183
rect 8720 10152 11560 10180
rect 11624 10152 14289 10180
rect 8720 10140 8726 10152
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10072 1458 10124
rect 2133 10115 2191 10121
rect 2133 10081 2145 10115
rect 2179 10112 2191 10115
rect 2774 10112 2780 10124
rect 2179 10084 2780 10112
rect 2179 10081 2191 10084
rect 2133 10075 2191 10081
rect 2774 10072 2780 10084
rect 2832 10072 2838 10124
rect 4332 10115 4390 10121
rect 4332 10081 4344 10115
rect 4378 10112 4390 10115
rect 5074 10112 5080 10124
rect 4378 10084 5080 10112
rect 4378 10081 4390 10084
rect 4332 10075 4390 10081
rect 5074 10072 5080 10084
rect 5132 10072 5138 10124
rect 9933 10115 9991 10121
rect 9933 10112 9945 10115
rect 5368 10084 9945 10112
rect 4062 10044 4068 10056
rect 4023 10016 4068 10044
rect 4062 10004 4068 10016
rect 4120 10004 4126 10056
rect 3513 9911 3571 9917
rect 3513 9877 3525 9911
rect 3559 9908 3571 9911
rect 3786 9908 3792 9920
rect 3559 9880 3792 9908
rect 3559 9877 3571 9880
rect 3513 9871 3571 9877
rect 3786 9868 3792 9880
rect 3844 9908 3850 9920
rect 5368 9908 5396 10084
rect 9933 10081 9945 10084
rect 9979 10081 9991 10115
rect 9933 10075 9991 10081
rect 10502 10072 10508 10124
rect 10560 10112 10566 10124
rect 10560 10084 10732 10112
rect 10560 10072 10566 10084
rect 5902 10044 5908 10056
rect 5863 10016 5908 10044
rect 5902 10004 5908 10016
rect 5960 10004 5966 10056
rect 7742 10044 7748 10056
rect 7703 10016 7748 10044
rect 7742 10004 7748 10016
rect 7800 10004 7806 10056
rect 9582 10004 9588 10056
rect 9640 10044 9646 10056
rect 9677 10047 9735 10053
rect 9677 10044 9689 10047
rect 9640 10016 9689 10044
rect 9640 10004 9646 10016
rect 9677 10013 9689 10016
rect 9723 10013 9735 10047
rect 9677 10007 9735 10013
rect 7098 9936 7104 9988
rect 7156 9976 7162 9988
rect 7285 9979 7343 9985
rect 7285 9976 7297 9979
rect 7156 9948 7297 9976
rect 7156 9936 7162 9948
rect 7285 9945 7297 9948
rect 7331 9945 7343 9979
rect 7285 9939 7343 9945
rect 3844 9880 5396 9908
rect 3844 9868 3850 9880
rect 5902 9868 5908 9920
rect 5960 9908 5966 9920
rect 7760 9908 7788 10004
rect 9125 9979 9183 9985
rect 9125 9945 9137 9979
rect 9171 9976 9183 9979
rect 9306 9976 9312 9988
rect 9171 9948 9312 9976
rect 9171 9945 9183 9948
rect 9125 9939 9183 9945
rect 9306 9936 9312 9948
rect 9364 9936 9370 9988
rect 10704 9976 10732 10084
rect 10778 10072 10784 10124
rect 10836 10112 10842 10124
rect 11624 10112 11652 10152
rect 14277 10149 14289 10152
rect 14323 10149 14335 10183
rect 14277 10143 14335 10149
rect 14366 10140 14372 10192
rect 14424 10140 14430 10192
rect 10836 10084 11652 10112
rect 11977 10115 12035 10121
rect 10836 10072 10842 10084
rect 11977 10081 11989 10115
rect 12023 10112 12035 10115
rect 12250 10112 12256 10124
rect 12023 10084 12256 10112
rect 12023 10081 12035 10084
rect 11977 10075 12035 10081
rect 12250 10072 12256 10084
rect 12308 10112 12314 10124
rect 12434 10112 12440 10124
rect 12308 10084 12440 10112
rect 12308 10072 12314 10084
rect 12434 10072 12440 10084
rect 12492 10072 12498 10124
rect 13078 10112 13084 10124
rect 13039 10084 13084 10112
rect 13078 10072 13084 10084
rect 13136 10072 13142 10124
rect 13998 10072 14004 10124
rect 14056 10112 14062 10124
rect 14384 10112 14412 10140
rect 14056 10084 14412 10112
rect 14056 10072 14062 10084
rect 12158 10044 12164 10056
rect 12119 10016 12164 10044
rect 12158 10004 12164 10016
rect 12216 10004 12222 10056
rect 13265 10047 13323 10053
rect 13265 10013 13277 10047
rect 13311 10013 13323 10047
rect 14366 10044 14372 10056
rect 14327 10016 14372 10044
rect 13265 10007 13323 10013
rect 12713 9979 12771 9985
rect 12713 9976 12725 9979
rect 10704 9948 12725 9976
rect 12713 9945 12725 9948
rect 12759 9945 12771 9979
rect 12713 9939 12771 9945
rect 5960 9880 7788 9908
rect 5960 9868 5966 9880
rect 10594 9868 10600 9920
rect 10652 9908 10658 9920
rect 10778 9908 10784 9920
rect 10652 9880 10784 9908
rect 10652 9868 10658 9880
rect 10778 9868 10784 9880
rect 10836 9868 10842 9920
rect 11238 9868 11244 9920
rect 11296 9908 11302 9920
rect 13280 9908 13308 10007
rect 14366 10004 14372 10016
rect 14424 10004 14430 10056
rect 14461 10047 14519 10053
rect 14461 10013 14473 10047
rect 14507 10013 14519 10047
rect 14461 10007 14519 10013
rect 14182 9936 14188 9988
rect 14240 9976 14246 9988
rect 14476 9976 14504 10007
rect 14240 9948 14504 9976
rect 14240 9936 14246 9948
rect 11296 9880 13308 9908
rect 11296 9868 11302 9880
rect 1104 9818 15824 9840
rect 1104 9766 3447 9818
rect 3499 9766 3511 9818
rect 3563 9766 3575 9818
rect 3627 9766 3639 9818
rect 3691 9766 8378 9818
rect 8430 9766 8442 9818
rect 8494 9766 8506 9818
rect 8558 9766 8570 9818
rect 8622 9766 13308 9818
rect 13360 9766 13372 9818
rect 13424 9766 13436 9818
rect 13488 9766 13500 9818
rect 13552 9766 15824 9818
rect 1104 9744 15824 9766
rect 1857 9707 1915 9713
rect 1857 9673 1869 9707
rect 1903 9704 1915 9707
rect 2314 9704 2320 9716
rect 1903 9676 2320 9704
rect 1903 9673 1915 9676
rect 1857 9667 1915 9673
rect 2314 9664 2320 9676
rect 2372 9664 2378 9716
rect 2590 9664 2596 9716
rect 2648 9704 2654 9716
rect 2958 9704 2964 9716
rect 2648 9676 2964 9704
rect 2648 9664 2654 9676
rect 2958 9664 2964 9676
rect 3016 9664 3022 9716
rect 4062 9704 4068 9716
rect 3068 9676 4068 9704
rect 2498 9568 2504 9580
rect 2459 9540 2504 9568
rect 2498 9528 2504 9540
rect 2556 9528 2562 9580
rect 3068 9577 3096 9676
rect 4062 9664 4068 9676
rect 4120 9664 4126 9716
rect 5902 9704 5908 9716
rect 5276 9676 5908 9704
rect 4430 9636 4436 9648
rect 4391 9608 4436 9636
rect 4430 9596 4436 9608
rect 4488 9596 4494 9648
rect 5276 9577 5304 9676
rect 5902 9664 5908 9676
rect 5960 9664 5966 9716
rect 5994 9664 6000 9716
rect 6052 9704 6058 9716
rect 8110 9704 8116 9716
rect 6052 9676 8116 9704
rect 6052 9664 6058 9676
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 12437 9707 12495 9713
rect 9048 9676 11468 9704
rect 6270 9596 6276 9648
rect 6328 9636 6334 9648
rect 8662 9636 8668 9648
rect 6328 9608 8668 9636
rect 6328 9596 6334 9608
rect 8662 9596 8668 9608
rect 8720 9596 8726 9648
rect 3053 9571 3111 9577
rect 3053 9537 3065 9571
rect 3099 9537 3111 9571
rect 3053 9531 3111 9537
rect 5261 9571 5319 9577
rect 5261 9537 5273 9571
rect 5307 9537 5319 9571
rect 5261 9531 5319 9537
rect 8202 9528 8208 9580
rect 8260 9568 8266 9580
rect 9048 9568 9076 9676
rect 10226 9596 10232 9648
rect 10284 9636 10290 9648
rect 10413 9639 10471 9645
rect 10413 9636 10425 9639
rect 10284 9608 10425 9636
rect 10284 9596 10290 9608
rect 10413 9605 10425 9608
rect 10459 9605 10471 9639
rect 11440 9636 11468 9676
rect 12437 9673 12449 9707
rect 12483 9704 12495 9707
rect 13078 9704 13084 9716
rect 12483 9676 13084 9704
rect 12483 9673 12495 9676
rect 12437 9667 12495 9673
rect 13078 9664 13084 9676
rect 13136 9664 13142 9716
rect 13633 9639 13691 9645
rect 13633 9636 13645 9639
rect 11440 9608 13645 9636
rect 10413 9599 10471 9605
rect 13633 9605 13645 9608
rect 13679 9605 13691 9639
rect 13633 9599 13691 9605
rect 13998 9596 14004 9648
rect 14056 9636 14062 9648
rect 14056 9608 14872 9636
rect 14056 9596 14062 9608
rect 12986 9568 12992 9580
rect 8260 9540 9076 9568
rect 12360 9540 12992 9568
rect 8260 9528 8266 9540
rect 2317 9503 2375 9509
rect 2317 9469 2329 9503
rect 2363 9500 2375 9503
rect 3602 9500 3608 9512
rect 2363 9472 3608 9500
rect 2363 9469 2375 9472
rect 2317 9463 2375 9469
rect 3602 9460 3608 9472
rect 3660 9460 3666 9512
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9500 5135 9503
rect 5169 9503 5227 9509
rect 5169 9500 5181 9503
rect 5123 9472 5181 9500
rect 5123 9469 5135 9472
rect 5077 9463 5135 9469
rect 5169 9469 5181 9472
rect 5215 9469 5227 9503
rect 8570 9500 8576 9512
rect 5169 9463 5227 9469
rect 5460 9472 8576 9500
rect 2225 9435 2283 9441
rect 2225 9401 2237 9435
rect 2271 9432 2283 9435
rect 2958 9432 2964 9444
rect 2271 9404 2964 9432
rect 2271 9401 2283 9404
rect 2225 9395 2283 9401
rect 2958 9392 2964 9404
rect 3016 9392 3022 9444
rect 3320 9435 3378 9441
rect 3320 9401 3332 9435
rect 3366 9432 3378 9435
rect 5460 9432 5488 9472
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 9033 9503 9091 9509
rect 9033 9469 9045 9503
rect 9079 9500 9091 9503
rect 9122 9500 9128 9512
rect 9079 9472 9128 9500
rect 9079 9469 9091 9472
rect 9033 9463 9091 9469
rect 9122 9460 9128 9472
rect 9180 9460 9186 9512
rect 9582 9460 9588 9512
rect 9640 9500 9646 9512
rect 10505 9503 10563 9509
rect 10505 9500 10517 9503
rect 9640 9472 10517 9500
rect 9640 9460 9646 9472
rect 10505 9469 10517 9472
rect 10551 9469 10563 9503
rect 12066 9500 12072 9512
rect 10505 9463 10563 9469
rect 10704 9472 12072 9500
rect 5534 9441 5540 9444
rect 3366 9404 5488 9432
rect 3366 9401 3378 9404
rect 3320 9395 3378 9401
rect 5528 9395 5540 9441
rect 5592 9432 5598 9444
rect 5592 9404 5628 9432
rect 5534 9392 5540 9395
rect 5592 9392 5598 9404
rect 5810 9392 5816 9444
rect 5868 9432 5874 9444
rect 6270 9432 6276 9444
rect 5868 9404 6276 9432
rect 5868 9392 5874 9404
rect 6270 9392 6276 9404
rect 6328 9392 6334 9444
rect 7190 9432 7196 9444
rect 6564 9404 7113 9432
rect 7151 9404 7196 9432
rect 4890 9364 4896 9376
rect 4851 9336 4896 9364
rect 4890 9324 4896 9336
rect 4948 9324 4954 9376
rect 5169 9367 5227 9373
rect 5169 9333 5181 9367
rect 5215 9364 5227 9367
rect 6564 9364 6592 9404
rect 5215 9336 6592 9364
rect 6641 9367 6699 9373
rect 5215 9333 5227 9336
rect 5169 9327 5227 9333
rect 6641 9333 6653 9367
rect 6687 9364 6699 9367
rect 6914 9364 6920 9376
rect 6687 9336 6920 9364
rect 6687 9333 6699 9336
rect 6641 9327 6699 9333
rect 6914 9324 6920 9336
rect 6972 9324 6978 9376
rect 7085 9364 7113 9404
rect 7190 9392 7196 9404
rect 7248 9392 7254 9444
rect 8754 9432 8760 9444
rect 8715 9404 8760 9432
rect 8754 9392 8760 9404
rect 8812 9392 8818 9444
rect 9300 9435 9358 9441
rect 9300 9401 9312 9435
rect 9346 9432 9358 9435
rect 10704 9432 10732 9472
rect 12066 9460 12072 9472
rect 12124 9460 12130 9512
rect 12360 9500 12388 9540
rect 12986 9528 12992 9540
rect 13044 9568 13050 9580
rect 14185 9571 14243 9577
rect 14185 9568 14197 9571
rect 13044 9540 14197 9568
rect 13044 9528 13050 9540
rect 14185 9537 14197 9540
rect 14231 9537 14243 9571
rect 14185 9531 14243 9537
rect 12268 9472 12388 9500
rect 9346 9404 10732 9432
rect 10772 9435 10830 9441
rect 9346 9401 9358 9404
rect 9300 9395 9358 9401
rect 10772 9401 10784 9435
rect 10818 9432 10830 9435
rect 11146 9432 11152 9444
rect 10818 9404 11152 9432
rect 10818 9401 10830 9404
rect 10772 9395 10830 9401
rect 11146 9392 11152 9404
rect 11204 9432 11210 9444
rect 12158 9432 12164 9444
rect 11204 9404 12164 9432
rect 11204 9392 11210 9404
rect 12158 9392 12164 9404
rect 12216 9392 12222 9444
rect 9122 9364 9128 9376
rect 7085 9336 9128 9364
rect 9122 9324 9128 9336
rect 9180 9324 9186 9376
rect 9582 9324 9588 9376
rect 9640 9364 9646 9376
rect 11606 9364 11612 9376
rect 9640 9336 11612 9364
rect 9640 9324 9646 9336
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 11882 9364 11888 9376
rect 11843 9336 11888 9364
rect 11882 9324 11888 9336
rect 11940 9364 11946 9376
rect 12268 9364 12296 9472
rect 12618 9460 12624 9512
rect 12676 9500 12682 9512
rect 12805 9503 12863 9509
rect 12805 9500 12817 9503
rect 12676 9472 12817 9500
rect 12676 9460 12682 9472
rect 12805 9469 12817 9472
rect 12851 9469 12863 9503
rect 12805 9463 12863 9469
rect 13446 9460 13452 9512
rect 13504 9500 13510 9512
rect 14844 9509 14872 9608
rect 14001 9503 14059 9509
rect 14001 9500 14013 9503
rect 13504 9472 14013 9500
rect 13504 9460 13510 9472
rect 14001 9469 14013 9472
rect 14047 9469 14059 9503
rect 14001 9463 14059 9469
rect 14829 9503 14887 9509
rect 14829 9469 14841 9503
rect 14875 9469 14887 9503
rect 14829 9463 14887 9469
rect 12897 9435 12955 9441
rect 12897 9401 12909 9435
rect 12943 9432 12955 9435
rect 14274 9432 14280 9444
rect 12943 9404 14280 9432
rect 12943 9401 12955 9404
rect 12897 9395 12955 9401
rect 14274 9392 14280 9404
rect 14332 9392 14338 9444
rect 14090 9364 14096 9376
rect 11940 9336 12296 9364
rect 14051 9336 14096 9364
rect 11940 9324 11946 9336
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 15010 9364 15016 9376
rect 14971 9336 15016 9364
rect 15010 9324 15016 9336
rect 15068 9324 15074 9376
rect 1104 9274 15824 9296
rect 1104 9222 5912 9274
rect 5964 9222 5976 9274
rect 6028 9222 6040 9274
rect 6092 9222 6104 9274
rect 6156 9222 10843 9274
rect 10895 9222 10907 9274
rect 10959 9222 10971 9274
rect 11023 9222 11035 9274
rect 11087 9222 15824 9274
rect 1104 9200 15824 9222
rect 2958 9120 2964 9172
rect 3016 9160 3022 9172
rect 13357 9163 13415 9169
rect 13357 9160 13369 9163
rect 3016 9132 13369 9160
rect 3016 9120 3022 9132
rect 13357 9129 13369 9132
rect 13403 9129 13415 9163
rect 13357 9123 13415 9129
rect 2498 9052 2504 9104
rect 2556 9092 2562 9104
rect 5810 9092 5816 9104
rect 2556 9064 5816 9092
rect 2556 9052 2562 9064
rect 5810 9052 5816 9064
rect 5868 9052 5874 9104
rect 5994 9101 6000 9104
rect 5988 9055 6000 9101
rect 6052 9092 6058 9104
rect 6052 9064 6088 9092
rect 5994 9052 6000 9055
rect 6052 9052 6058 9064
rect 6270 9052 6276 9104
rect 6328 9092 6334 9104
rect 9922 9095 9980 9101
rect 9922 9092 9934 9095
rect 6328 9064 9934 9092
rect 6328 9052 6334 9064
rect 9922 9061 9934 9064
rect 9968 9092 9980 9095
rect 11882 9092 11888 9104
rect 9968 9064 11888 9092
rect 9968 9061 9980 9064
rect 9922 9055 9980 9061
rect 11882 9052 11888 9064
rect 11940 9052 11946 9104
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 2038 9024 2044 9036
rect 1443 8996 2044 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2038 8984 2044 8996
rect 2096 8984 2102 9036
rect 2400 9027 2458 9033
rect 2400 8993 2412 9027
rect 2446 9024 2458 9027
rect 4154 9024 4160 9036
rect 2446 8996 4160 9024
rect 2446 8993 2458 8996
rect 2400 8987 2458 8993
rect 4154 8984 4160 8996
rect 4212 8984 4218 9036
rect 4516 9027 4574 9033
rect 4516 8993 4528 9027
rect 4562 9024 4574 9027
rect 5442 9024 5448 9036
rect 4562 8996 5448 9024
rect 4562 8993 4574 8996
rect 4516 8987 4574 8993
rect 5442 8984 5448 8996
rect 5500 8984 5506 9036
rect 5721 9027 5779 9033
rect 5721 8993 5733 9027
rect 5767 9024 5779 9027
rect 5767 8996 7236 9024
rect 5767 8993 5779 8996
rect 5721 8987 5779 8993
rect 2130 8956 2136 8968
rect 2091 8928 2136 8956
rect 2130 8916 2136 8928
rect 2188 8916 2194 8968
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 4249 8959 4307 8965
rect 4249 8956 4261 8959
rect 4120 8928 4261 8956
rect 4120 8916 4126 8928
rect 4249 8925 4261 8928
rect 4295 8925 4307 8959
rect 7208 8956 7236 8996
rect 7282 8984 7288 9036
rect 7340 9024 7346 9036
rect 7817 9027 7875 9033
rect 7817 9024 7829 9027
rect 7340 8996 7829 9024
rect 7340 8984 7346 8996
rect 7817 8993 7829 8996
rect 7863 8993 7875 9027
rect 7817 8987 7875 8993
rect 8846 8984 8852 9036
rect 8904 9024 8910 9036
rect 9030 9024 9036 9036
rect 8904 8996 9036 9024
rect 8904 8984 8910 8996
rect 9030 8984 9036 8996
rect 9088 8984 9094 9036
rect 9214 8984 9220 9036
rect 9272 9024 9278 9036
rect 9677 9027 9735 9033
rect 9677 9024 9689 9027
rect 9272 8996 9689 9024
rect 9272 8984 9278 8996
rect 9677 8993 9689 8996
rect 9723 8993 9735 9027
rect 10226 9024 10232 9036
rect 9677 8987 9735 8993
rect 9784 8996 10232 9024
rect 7561 8959 7619 8965
rect 7561 8956 7573 8959
rect 7208 8928 7573 8956
rect 4249 8919 4307 8925
rect 7561 8925 7573 8928
rect 7607 8925 7619 8959
rect 7561 8919 7619 8925
rect 5629 8891 5687 8897
rect 5629 8857 5641 8891
rect 5675 8888 5687 8891
rect 5718 8888 5724 8900
rect 5675 8860 5724 8888
rect 5675 8857 5687 8860
rect 5629 8851 5687 8857
rect 5718 8848 5724 8860
rect 5776 8848 5782 8900
rect 937 8823 995 8829
rect 937 8789 949 8823
rect 983 8820 995 8823
rect 1581 8823 1639 8829
rect 1581 8820 1593 8823
rect 983 8792 1593 8820
rect 983 8789 995 8792
rect 937 8783 995 8789
rect 1581 8789 1593 8792
rect 1627 8789 1639 8823
rect 1581 8783 1639 8789
rect 3513 8823 3571 8829
rect 3513 8789 3525 8823
rect 3559 8820 3571 8823
rect 3786 8820 3792 8832
rect 3559 8792 3792 8820
rect 3559 8789 3571 8792
rect 3513 8783 3571 8789
rect 3786 8780 3792 8792
rect 3844 8780 3850 8832
rect 4890 8780 4896 8832
rect 4948 8820 4954 8832
rect 6454 8820 6460 8832
rect 4948 8792 6460 8820
rect 4948 8780 4954 8792
rect 6454 8780 6460 8792
rect 6512 8780 6518 8832
rect 7101 8823 7159 8829
rect 7101 8789 7113 8823
rect 7147 8820 7159 8823
rect 7282 8820 7288 8832
rect 7147 8792 7288 8820
rect 7147 8789 7159 8792
rect 7101 8783 7159 8789
rect 7282 8780 7288 8792
rect 7340 8780 7346 8832
rect 7576 8820 7604 8919
rect 8570 8916 8576 8968
rect 8628 8956 8634 8968
rect 9582 8956 9588 8968
rect 8628 8928 9588 8956
rect 8628 8916 8634 8928
rect 9582 8916 9588 8928
rect 9640 8956 9646 8968
rect 9784 8956 9812 8996
rect 10226 8984 10232 8996
rect 10284 8984 10290 9036
rect 10502 8984 10508 9036
rect 10560 9024 10566 9036
rect 11784 9027 11842 9033
rect 10560 8996 10732 9024
rect 10560 8984 10566 8996
rect 9640 8928 9812 8956
rect 9640 8916 9646 8928
rect 10704 8888 10732 8996
rect 11784 8993 11796 9027
rect 11830 9024 11842 9027
rect 12250 9024 12256 9036
rect 11830 8996 12256 9024
rect 11830 8993 11842 8996
rect 11784 8987 11842 8993
rect 12250 8984 12256 8996
rect 12308 9024 12314 9036
rect 13538 9024 13544 9036
rect 12308 8996 13544 9024
rect 12308 8984 12314 8996
rect 13538 8984 13544 8996
rect 13596 8984 13602 9036
rect 13630 8984 13636 9036
rect 13688 9024 13694 9036
rect 13725 9027 13783 9033
rect 13725 9024 13737 9027
rect 13688 8996 13737 9024
rect 13688 8984 13694 8996
rect 13725 8993 13737 8996
rect 13771 8993 13783 9027
rect 13725 8987 13783 8993
rect 10962 8916 10968 8968
rect 11020 8956 11026 8968
rect 11517 8959 11575 8965
rect 11517 8956 11529 8959
rect 11020 8928 11529 8956
rect 11020 8916 11026 8928
rect 11517 8925 11529 8928
rect 11563 8925 11575 8959
rect 11517 8919 11575 8925
rect 12526 8916 12532 8968
rect 12584 8956 12590 8968
rect 13817 8959 13875 8965
rect 13817 8956 13829 8959
rect 12584 8928 13829 8956
rect 12584 8916 12590 8928
rect 13817 8925 13829 8928
rect 13863 8925 13875 8959
rect 13817 8919 13875 8925
rect 14001 8959 14059 8965
rect 14001 8925 14013 8959
rect 14047 8956 14059 8959
rect 14458 8956 14464 8968
rect 14047 8928 14464 8956
rect 14047 8925 14059 8928
rect 14001 8919 14059 8925
rect 14458 8916 14464 8928
rect 14516 8916 14522 8968
rect 14553 8959 14611 8965
rect 14553 8925 14565 8959
rect 14599 8956 14611 8959
rect 15562 8956 15568 8968
rect 14599 8928 15568 8956
rect 14599 8925 14611 8928
rect 14553 8919 14611 8925
rect 15562 8916 15568 8928
rect 15620 8916 15626 8968
rect 11057 8891 11115 8897
rect 11057 8888 11069 8891
rect 10704 8860 11069 8888
rect 11057 8857 11069 8860
rect 11103 8888 11115 8891
rect 11238 8888 11244 8900
rect 11103 8860 11244 8888
rect 11103 8857 11115 8860
rect 11057 8851 11115 8857
rect 11238 8848 11244 8860
rect 11296 8848 11302 8900
rect 12710 8848 12716 8900
rect 12768 8888 12774 8900
rect 12768 8860 14044 8888
rect 12768 8848 12774 8860
rect 14016 8832 14044 8860
rect 7834 8820 7840 8832
rect 7576 8792 7840 8820
rect 7834 8780 7840 8792
rect 7892 8780 7898 8832
rect 8202 8780 8208 8832
rect 8260 8820 8266 8832
rect 8941 8823 8999 8829
rect 8941 8820 8953 8823
rect 8260 8792 8953 8820
rect 8260 8780 8266 8792
rect 8941 8789 8953 8792
rect 8987 8820 8999 8823
rect 10318 8820 10324 8832
rect 8987 8792 10324 8820
rect 8987 8789 8999 8792
rect 8941 8783 8999 8789
rect 10318 8780 10324 8792
rect 10376 8780 10382 8832
rect 10594 8780 10600 8832
rect 10652 8820 10658 8832
rect 12434 8820 12440 8832
rect 10652 8792 12440 8820
rect 10652 8780 10658 8792
rect 12434 8780 12440 8792
rect 12492 8780 12498 8832
rect 12897 8823 12955 8829
rect 12897 8789 12909 8823
rect 12943 8820 12955 8823
rect 13078 8820 13084 8832
rect 12943 8792 13084 8820
rect 12943 8789 12955 8792
rect 12897 8783 12955 8789
rect 13078 8780 13084 8792
rect 13136 8780 13142 8832
rect 13998 8780 14004 8832
rect 14056 8780 14062 8832
rect 1104 8730 15824 8752
rect 1104 8678 3447 8730
rect 3499 8678 3511 8730
rect 3563 8678 3575 8730
rect 3627 8678 3639 8730
rect 3691 8678 8378 8730
rect 8430 8678 8442 8730
rect 8494 8678 8506 8730
rect 8558 8678 8570 8730
rect 8622 8678 13308 8730
rect 13360 8678 13372 8730
rect 13424 8678 13436 8730
rect 13488 8678 13500 8730
rect 13552 8678 15824 8730
rect 1104 8656 15824 8678
rect 2225 8619 2283 8625
rect 2225 8585 2237 8619
rect 2271 8616 2283 8619
rect 2958 8616 2964 8628
rect 2271 8588 2964 8616
rect 2271 8585 2283 8588
rect 2225 8579 2283 8585
rect 2958 8576 2964 8588
rect 3016 8576 3022 8628
rect 4062 8616 4068 8628
rect 3068 8588 4068 8616
rect 2130 8508 2136 8560
rect 2188 8548 2194 8560
rect 3068 8548 3096 8588
rect 4062 8576 4068 8588
rect 4120 8576 4126 8628
rect 4433 8619 4491 8625
rect 4433 8585 4445 8619
rect 4479 8616 4491 8619
rect 11146 8616 11152 8628
rect 4479 8588 11152 8616
rect 4479 8585 4491 8588
rect 4433 8579 4491 8585
rect 11146 8576 11152 8588
rect 11204 8616 11210 8628
rect 11204 8588 11836 8616
rect 11204 8576 11210 8588
rect 2188 8520 3096 8548
rect 2188 8508 2194 8520
rect 3068 8489 3096 8520
rect 5994 8508 6000 8560
rect 6052 8548 6058 8560
rect 6270 8548 6276 8560
rect 6052 8520 6276 8548
rect 6052 8508 6058 8520
rect 6270 8508 6276 8520
rect 6328 8508 6334 8560
rect 9674 8508 9680 8560
rect 9732 8548 9738 8560
rect 9858 8548 9864 8560
rect 9732 8520 9864 8548
rect 9732 8508 9738 8520
rect 9858 8508 9864 8520
rect 9916 8508 9922 8560
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8480 2099 8483
rect 2869 8483 2927 8489
rect 2087 8452 2820 8480
rect 2087 8449 2099 8452
rect 2041 8443 2099 8449
rect 2682 8412 2688 8424
rect 2643 8384 2688 8412
rect 2682 8372 2688 8384
rect 2740 8372 2746 8424
rect 1762 8344 1768 8356
rect 1723 8316 1768 8344
rect 1762 8304 1768 8316
rect 1820 8304 1826 8356
rect 1857 8347 1915 8353
rect 1857 8313 1869 8347
rect 1903 8344 1915 8347
rect 2314 8344 2320 8356
rect 1903 8316 2320 8344
rect 1903 8313 1915 8316
rect 1857 8307 1915 8313
rect 2314 8304 2320 8316
rect 2372 8304 2378 8356
rect 1026 8236 1032 8288
rect 1084 8276 1090 8288
rect 1397 8279 1455 8285
rect 1397 8276 1409 8279
rect 1084 8248 1409 8276
rect 1084 8236 1090 8248
rect 1397 8245 1409 8248
rect 1443 8245 1455 8279
rect 1397 8239 1455 8245
rect 2222 8236 2228 8288
rect 2280 8276 2286 8288
rect 2593 8279 2651 8285
rect 2593 8276 2605 8279
rect 2280 8248 2605 8276
rect 2280 8236 2286 8248
rect 2593 8245 2605 8248
rect 2639 8245 2651 8279
rect 2792 8276 2820 8452
rect 2869 8449 2881 8483
rect 2915 8449 2927 8483
rect 2869 8443 2927 8449
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8449 3111 8483
rect 3053 8443 3111 8449
rect 2884 8412 2912 8443
rect 4062 8440 4068 8492
rect 4120 8480 4126 8492
rect 4890 8480 4896 8492
rect 4120 8452 4896 8480
rect 4120 8440 4126 8452
rect 4890 8440 4896 8452
rect 4948 8440 4954 8492
rect 7834 8440 7840 8492
rect 7892 8480 7898 8492
rect 7892 8452 8708 8480
rect 7892 8440 7898 8452
rect 8680 8424 8708 8452
rect 10042 8440 10048 8492
rect 10100 8480 10106 8492
rect 11808 8480 11836 8588
rect 11882 8576 11888 8628
rect 11940 8616 11946 8628
rect 12437 8619 12495 8625
rect 11940 8588 11985 8616
rect 11940 8576 11946 8588
rect 12437 8585 12449 8619
rect 12483 8616 12495 8619
rect 14090 8616 14096 8628
rect 12483 8588 14096 8616
rect 12483 8585 12495 8588
rect 12437 8579 12495 8585
rect 14090 8576 14096 8588
rect 14148 8576 14154 8628
rect 12342 8508 12348 8560
rect 12400 8548 12406 8560
rect 12618 8548 12624 8560
rect 12400 8520 12624 8548
rect 12400 8508 12406 8520
rect 12618 8508 12624 8520
rect 12676 8508 12682 8560
rect 13633 8551 13691 8557
rect 13633 8517 13645 8551
rect 13679 8548 13691 8551
rect 13814 8548 13820 8560
rect 13679 8520 13820 8548
rect 13679 8517 13691 8520
rect 13633 8511 13691 8517
rect 13814 8508 13820 8520
rect 13872 8508 13878 8560
rect 14458 8548 14464 8560
rect 14016 8520 14464 8548
rect 12989 8483 13047 8489
rect 12989 8480 13001 8483
rect 10100 8452 10640 8480
rect 11808 8452 13001 8480
rect 10100 8440 10106 8452
rect 3326 8421 3332 8424
rect 2884 8384 3280 8412
rect 3252 8344 3280 8384
rect 3320 8375 3332 8421
rect 3384 8412 3390 8424
rect 5534 8412 5540 8424
rect 3384 8384 3420 8412
rect 5000 8384 5540 8412
rect 3326 8372 3332 8375
rect 3384 8372 3390 8384
rect 5000 8344 5028 8384
rect 5534 8372 5540 8384
rect 5592 8372 5598 8424
rect 6730 8372 6736 8424
rect 6788 8412 6794 8424
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 6788 8384 6837 8412
rect 6788 8372 6794 8384
rect 6825 8381 6837 8384
rect 6871 8381 6883 8415
rect 6825 8375 6883 8381
rect 6914 8372 6920 8424
rect 6972 8412 6978 8424
rect 7926 8412 7932 8424
rect 6972 8384 7932 8412
rect 6972 8372 6978 8384
rect 7926 8372 7932 8384
rect 7984 8412 7990 8424
rect 8662 8412 8668 8424
rect 7984 8384 8432 8412
rect 8575 8384 8668 8412
rect 7984 8372 7990 8384
rect 5166 8353 5172 8356
rect 5160 8344 5172 8353
rect 3252 8316 5028 8344
rect 5127 8316 5172 8344
rect 5160 8307 5172 8316
rect 5166 8304 5172 8307
rect 5224 8304 5230 8356
rect 5810 8304 5816 8356
rect 5868 8344 5874 8356
rect 7070 8347 7128 8353
rect 7070 8344 7082 8347
rect 5868 8316 7082 8344
rect 5868 8304 5874 8316
rect 7070 8313 7082 8316
rect 7116 8344 7128 8347
rect 7282 8344 7288 8356
rect 7116 8316 7288 8344
rect 7116 8313 7128 8316
rect 7070 8307 7128 8313
rect 7282 8304 7288 8316
rect 7340 8304 7346 8356
rect 8404 8344 8432 8384
rect 8662 8372 8668 8384
rect 8720 8412 8726 8424
rect 9214 8412 9220 8424
rect 8720 8384 9220 8412
rect 8720 8372 8726 8384
rect 9214 8372 9220 8384
rect 9272 8412 9278 8424
rect 10505 8415 10563 8421
rect 10505 8412 10517 8415
rect 9272 8384 10517 8412
rect 9272 8372 9278 8384
rect 10505 8381 10517 8384
rect 10551 8381 10563 8415
rect 10612 8412 10640 8452
rect 12989 8449 13001 8452
rect 13035 8480 13047 8483
rect 14016 8480 14044 8520
rect 14458 8508 14464 8520
rect 14516 8508 14522 8560
rect 14182 8480 14188 8492
rect 13035 8452 14044 8480
rect 14143 8452 14188 8480
rect 13035 8449 13047 8452
rect 12989 8443 13047 8449
rect 14182 8440 14188 8452
rect 14240 8440 14246 8492
rect 14093 8415 14151 8421
rect 14093 8412 14105 8415
rect 10612 8384 14105 8412
rect 10505 8375 10563 8381
rect 14093 8381 14105 8384
rect 14139 8381 14151 8415
rect 14093 8375 14151 8381
rect 14829 8415 14887 8421
rect 14829 8381 14841 8415
rect 14875 8412 14887 8415
rect 15102 8412 15108 8424
rect 14875 8384 15108 8412
rect 14875 8381 14887 8384
rect 14829 8375 14887 8381
rect 8910 8347 8968 8353
rect 8910 8344 8922 8347
rect 8036 8316 8340 8344
rect 8404 8316 8922 8344
rect 3326 8276 3332 8288
rect 2792 8248 3332 8276
rect 2593 8239 2651 8245
rect 3326 8236 3332 8248
rect 3384 8276 3390 8288
rect 3786 8276 3792 8288
rect 3384 8248 3792 8276
rect 3384 8236 3390 8248
rect 3786 8236 3792 8248
rect 3844 8236 3850 8288
rect 4154 8236 4160 8288
rect 4212 8276 4218 8288
rect 8036 8276 8064 8316
rect 8202 8276 8208 8288
rect 4212 8248 8064 8276
rect 8163 8248 8208 8276
rect 4212 8236 4218 8248
rect 8202 8236 8208 8248
rect 8260 8236 8266 8288
rect 8312 8276 8340 8316
rect 8910 8313 8922 8316
rect 8956 8313 8968 8347
rect 8910 8307 8968 8313
rect 8386 8276 8392 8288
rect 8312 8248 8392 8276
rect 8386 8236 8392 8248
rect 8444 8236 8450 8288
rect 9858 8236 9864 8288
rect 9916 8276 9922 8288
rect 10045 8279 10103 8285
rect 10045 8276 10057 8279
rect 9916 8248 10057 8276
rect 9916 8236 9922 8248
rect 10045 8245 10057 8248
rect 10091 8245 10103 8279
rect 10520 8276 10548 8375
rect 15102 8372 15108 8384
rect 15160 8372 15166 8424
rect 10686 8304 10692 8356
rect 10744 8353 10750 8356
rect 10744 8347 10808 8353
rect 10744 8313 10762 8347
rect 10796 8313 10808 8347
rect 10744 8307 10808 8313
rect 10744 8304 10750 8307
rect 10962 8304 10968 8356
rect 11020 8304 11026 8356
rect 11330 8304 11336 8356
rect 11388 8344 11394 8356
rect 11388 8316 11744 8344
rect 11388 8304 11394 8316
rect 10980 8276 11008 8304
rect 10520 8248 11008 8276
rect 10045 8239 10103 8245
rect 11146 8236 11152 8288
rect 11204 8276 11210 8288
rect 11606 8276 11612 8288
rect 11204 8248 11612 8276
rect 11204 8236 11210 8248
rect 11606 8236 11612 8248
rect 11664 8236 11670 8288
rect 11716 8276 11744 8316
rect 12066 8304 12072 8356
rect 12124 8344 12130 8356
rect 12710 8344 12716 8356
rect 12124 8316 12716 8344
rect 12124 8304 12130 8316
rect 12710 8304 12716 8316
rect 12768 8344 12774 8356
rect 12897 8347 12955 8353
rect 12897 8344 12909 8347
rect 12768 8316 12909 8344
rect 12768 8304 12774 8316
rect 12897 8313 12909 8316
rect 12943 8313 12955 8347
rect 14458 8344 14464 8356
rect 12897 8307 12955 8313
rect 13004 8316 14464 8344
rect 12805 8279 12863 8285
rect 12805 8276 12817 8279
rect 11716 8248 12817 8276
rect 12805 8245 12817 8248
rect 12851 8276 12863 8279
rect 13004 8276 13032 8316
rect 14458 8304 14464 8316
rect 14516 8304 14522 8356
rect 13998 8276 14004 8288
rect 12851 8248 13032 8276
rect 13959 8248 14004 8276
rect 12851 8245 12863 8248
rect 12805 8239 12863 8245
rect 13998 8236 14004 8248
rect 14056 8236 14062 8288
rect 15010 8276 15016 8288
rect 14971 8248 15016 8276
rect 15010 8236 15016 8248
rect 15068 8236 15074 8288
rect 1104 8186 15824 8208
rect 1104 8134 5912 8186
rect 5964 8134 5976 8186
rect 6028 8134 6040 8186
rect 6092 8134 6104 8186
rect 6156 8134 10843 8186
rect 10895 8134 10907 8186
rect 10959 8134 10971 8186
rect 11023 8134 11035 8186
rect 11087 8134 15824 8186
rect 1104 8112 15824 8134
rect 3513 8075 3571 8081
rect 3513 8041 3525 8075
rect 3559 8072 3571 8075
rect 4154 8072 4160 8084
rect 3559 8044 4160 8072
rect 3559 8041 3571 8044
rect 3513 8035 3571 8041
rect 4154 8032 4160 8044
rect 4212 8032 4218 8084
rect 4893 8075 4951 8081
rect 4893 8041 4905 8075
rect 4939 8072 4951 8075
rect 11517 8075 11575 8081
rect 11517 8072 11529 8075
rect 4939 8044 11529 8072
rect 4939 8041 4951 8044
rect 4893 8035 4951 8041
rect 11517 8041 11529 8044
rect 11563 8041 11575 8075
rect 11517 8035 11575 8041
rect 11606 8032 11612 8084
rect 11664 8072 11670 8084
rect 11977 8075 12035 8081
rect 11977 8072 11989 8075
rect 11664 8044 11989 8072
rect 11664 8032 11670 8044
rect 11977 8041 11989 8044
rect 12023 8072 12035 8075
rect 12526 8072 12532 8084
rect 12023 8044 12532 8072
rect 12023 8041 12035 8044
rect 11977 8035 12035 8041
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 12710 8072 12716 8084
rect 12671 8044 12716 8072
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 13909 8075 13967 8081
rect 13909 8041 13921 8075
rect 13955 8072 13967 8075
rect 13998 8072 14004 8084
rect 13955 8044 14004 8072
rect 13955 8041 13967 8044
rect 13909 8035 13967 8041
rect 13998 8032 14004 8044
rect 14056 8032 14062 8084
rect 2682 7964 2688 8016
rect 2740 8004 2746 8016
rect 3050 8004 3056 8016
rect 2740 7976 3056 8004
rect 2740 7964 2746 7976
rect 3050 7964 3056 7976
rect 3108 7964 3114 8016
rect 4062 7964 4068 8016
rect 4120 8004 4126 8016
rect 5166 8004 5172 8016
rect 4120 7976 5172 8004
rect 4120 7964 4126 7976
rect 5166 7964 5172 7976
rect 5224 8004 5230 8016
rect 5224 7976 8340 8004
rect 5224 7964 5230 7976
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 1946 7936 1952 7948
rect 1443 7908 1952 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 1946 7896 1952 7908
rect 2004 7896 2010 7948
rect 2130 7936 2136 7948
rect 2091 7908 2136 7936
rect 2130 7896 2136 7908
rect 2188 7896 2194 7948
rect 2400 7939 2458 7945
rect 2400 7905 2412 7939
rect 2446 7936 2458 7939
rect 2446 7908 3924 7936
rect 2446 7905 2458 7908
rect 2400 7899 2458 7905
rect 3896 7868 3924 7908
rect 5534 7896 5540 7948
rect 5592 7936 5598 7948
rect 5701 7939 5759 7945
rect 5701 7936 5713 7939
rect 5592 7908 5713 7936
rect 5592 7896 5598 7908
rect 5701 7905 5713 7908
rect 5747 7905 5759 7939
rect 5701 7899 5759 7905
rect 6822 7896 6828 7948
rect 6880 7936 6886 7948
rect 7374 7936 7380 7948
rect 6880 7908 7380 7936
rect 6880 7896 6886 7908
rect 7374 7896 7380 7908
rect 7432 7936 7438 7948
rect 7541 7939 7599 7945
rect 7541 7936 7553 7939
rect 7432 7908 7553 7936
rect 7432 7896 7438 7908
rect 7541 7905 7553 7908
rect 7587 7905 7599 7939
rect 7541 7899 7599 7905
rect 4246 7868 4252 7880
rect 3896 7840 4252 7868
rect 4246 7828 4252 7840
rect 4304 7828 4310 7880
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7837 5043 7871
rect 4985 7831 5043 7837
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7868 5227 7871
rect 5215 7840 5396 7868
rect 5215 7837 5227 7840
rect 5169 7831 5227 7837
rect 5000 7800 5028 7831
rect 5258 7800 5264 7812
rect 5000 7772 5264 7800
rect 5258 7760 5264 7772
rect 5316 7760 5322 7812
rect 1486 7692 1492 7744
rect 1544 7732 1550 7744
rect 1581 7735 1639 7741
rect 1581 7732 1593 7735
rect 1544 7704 1593 7732
rect 1544 7692 1550 7704
rect 1581 7701 1593 7704
rect 1627 7701 1639 7735
rect 4522 7732 4528 7744
rect 4483 7704 4528 7732
rect 1581 7695 1639 7701
rect 4522 7692 4528 7704
rect 4580 7692 4586 7744
rect 4614 7692 4620 7744
rect 4672 7732 4678 7744
rect 5368 7732 5396 7840
rect 5442 7828 5448 7880
rect 5500 7868 5506 7880
rect 5500 7840 5545 7868
rect 5500 7828 5506 7840
rect 6730 7828 6736 7880
rect 6788 7868 6794 7880
rect 7285 7871 7343 7877
rect 7285 7868 7297 7871
rect 6788 7840 7297 7868
rect 6788 7828 6794 7840
rect 7285 7837 7297 7840
rect 7331 7837 7343 7871
rect 8312 7868 8340 7976
rect 8386 7964 8392 8016
rect 8444 8004 8450 8016
rect 9922 8007 9980 8013
rect 9922 8004 9934 8007
rect 8444 7976 9934 8004
rect 8444 7964 8450 7976
rect 9922 7973 9934 7976
rect 9968 7973 9980 8007
rect 9922 7967 9980 7973
rect 10410 7964 10416 8016
rect 10468 8004 10474 8016
rect 11885 8007 11943 8013
rect 11885 8004 11897 8007
rect 10468 7976 11897 8004
rect 10468 7964 10474 7976
rect 11885 7973 11897 7976
rect 11931 7973 11943 8007
rect 11885 7967 11943 7973
rect 12342 7964 12348 8016
rect 12400 8004 12406 8016
rect 13081 8007 13139 8013
rect 13081 8004 13093 8007
rect 12400 7976 13093 8004
rect 12400 7964 12406 7976
rect 13081 7973 13093 7976
rect 13127 7973 13139 8007
rect 13081 7967 13139 7973
rect 8754 7896 8760 7948
rect 8812 7936 8818 7948
rect 9309 7939 9367 7945
rect 9309 7936 9321 7939
rect 8812 7908 9321 7936
rect 8812 7896 8818 7908
rect 9309 7905 9321 7908
rect 9355 7905 9367 7939
rect 9309 7899 9367 7905
rect 10318 7896 10324 7948
rect 10376 7936 10382 7948
rect 10376 7908 13308 7936
rect 10376 7896 10382 7908
rect 8312 7840 8892 7868
rect 7285 7831 7343 7837
rect 6086 7732 6092 7744
rect 4672 7704 6092 7732
rect 4672 7692 4678 7704
rect 6086 7692 6092 7704
rect 6144 7692 6150 7744
rect 6178 7692 6184 7744
rect 6236 7732 6242 7744
rect 6825 7735 6883 7741
rect 6825 7732 6837 7735
rect 6236 7704 6837 7732
rect 6236 7692 6242 7704
rect 6825 7701 6837 7704
rect 6871 7732 6883 7735
rect 7558 7732 7564 7744
rect 6871 7704 7564 7732
rect 6871 7701 6883 7704
rect 6825 7695 6883 7701
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 8665 7735 8723 7741
rect 8665 7701 8677 7735
rect 8711 7732 8723 7735
rect 8864 7732 8892 7840
rect 9214 7828 9220 7880
rect 9272 7868 9278 7880
rect 9677 7871 9735 7877
rect 9677 7868 9689 7871
rect 9272 7840 9689 7868
rect 9272 7828 9278 7840
rect 9677 7837 9689 7840
rect 9723 7837 9735 7871
rect 9677 7831 9735 7837
rect 11054 7828 11060 7880
rect 11112 7868 11118 7880
rect 12069 7871 12127 7877
rect 12069 7868 12081 7871
rect 11112 7840 12081 7868
rect 11112 7828 11118 7840
rect 12069 7837 12081 7840
rect 12115 7837 12127 7871
rect 12069 7831 12127 7837
rect 12526 7828 12532 7880
rect 12584 7868 12590 7880
rect 13280 7877 13308 7908
rect 13722 7896 13728 7948
rect 13780 7936 13786 7948
rect 14277 7939 14335 7945
rect 14277 7936 14289 7939
rect 13780 7908 14289 7936
rect 13780 7896 13786 7908
rect 14277 7905 14289 7908
rect 14323 7905 14335 7939
rect 14826 7936 14832 7948
rect 14277 7899 14335 7905
rect 14384 7908 14832 7936
rect 13173 7871 13231 7877
rect 13173 7868 13185 7871
rect 12584 7840 13185 7868
rect 12584 7828 12590 7840
rect 13173 7837 13185 7840
rect 13219 7837 13231 7871
rect 13173 7831 13231 7837
rect 13265 7871 13323 7877
rect 13265 7837 13277 7871
rect 13311 7837 13323 7871
rect 13265 7831 13323 7837
rect 13814 7828 13820 7880
rect 13872 7868 13878 7880
rect 14384 7877 14412 7908
rect 14826 7896 14832 7908
rect 14884 7896 14890 7948
rect 14369 7871 14427 7877
rect 14369 7868 14381 7871
rect 13872 7840 14381 7868
rect 13872 7828 13878 7840
rect 14369 7837 14381 7840
rect 14415 7837 14427 7871
rect 14369 7831 14427 7837
rect 14461 7871 14519 7877
rect 14461 7837 14473 7871
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 10778 7760 10784 7812
rect 10836 7800 10842 7812
rect 12342 7800 12348 7812
rect 10836 7772 12348 7800
rect 10836 7760 10842 7772
rect 12342 7760 12348 7772
rect 12400 7760 12406 7812
rect 13078 7760 13084 7812
rect 13136 7800 13142 7812
rect 14182 7800 14188 7812
rect 13136 7772 14188 7800
rect 13136 7760 13142 7772
rect 14182 7760 14188 7772
rect 14240 7800 14246 7812
rect 14476 7800 14504 7831
rect 14240 7772 14504 7800
rect 14240 7760 14246 7772
rect 9122 7732 9128 7744
rect 8711 7704 8892 7732
rect 9083 7704 9128 7732
rect 8711 7701 8723 7704
rect 8665 7695 8723 7701
rect 9122 7692 9128 7704
rect 9180 7692 9186 7744
rect 9214 7692 9220 7744
rect 9272 7732 9278 7744
rect 9490 7732 9496 7744
rect 9272 7704 9496 7732
rect 9272 7692 9278 7704
rect 9490 7692 9496 7704
rect 9548 7692 9554 7744
rect 9858 7692 9864 7744
rect 9916 7732 9922 7744
rect 10686 7732 10692 7744
rect 9916 7704 10692 7732
rect 9916 7692 9922 7704
rect 10686 7692 10692 7704
rect 10744 7732 10750 7744
rect 11057 7735 11115 7741
rect 11057 7732 11069 7735
rect 10744 7704 11069 7732
rect 10744 7692 10750 7704
rect 11057 7701 11069 7704
rect 11103 7701 11115 7735
rect 11057 7695 11115 7701
rect 11606 7692 11612 7744
rect 11664 7732 11670 7744
rect 13998 7732 14004 7744
rect 11664 7704 14004 7732
rect 11664 7692 11670 7704
rect 13998 7692 14004 7704
rect 14056 7692 14062 7744
rect 1104 7642 15824 7664
rect 1104 7590 3447 7642
rect 3499 7590 3511 7642
rect 3563 7590 3575 7642
rect 3627 7590 3639 7642
rect 3691 7590 8378 7642
rect 8430 7590 8442 7642
rect 8494 7590 8506 7642
rect 8558 7590 8570 7642
rect 8622 7590 13308 7642
rect 13360 7590 13372 7642
rect 13424 7590 13436 7642
rect 13488 7590 13500 7642
rect 13552 7590 15824 7642
rect 1104 7568 15824 7590
rect 4433 7531 4491 7537
rect 4433 7528 4445 7531
rect 3068 7500 4445 7528
rect 1857 7463 1915 7469
rect 1857 7429 1869 7463
rect 1903 7460 1915 7463
rect 2958 7460 2964 7472
rect 1903 7432 2964 7460
rect 1903 7429 1915 7432
rect 1857 7423 1915 7429
rect 2958 7420 2964 7432
rect 3016 7420 3022 7472
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 3068 7392 3096 7500
rect 4433 7497 4445 7500
rect 4479 7528 4491 7531
rect 4614 7528 4620 7540
rect 4479 7500 4620 7528
rect 4479 7497 4491 7500
rect 4433 7491 4491 7497
rect 4614 7488 4620 7500
rect 4672 7488 4678 7540
rect 5166 7528 5172 7540
rect 4908 7500 5172 7528
rect 4908 7460 4936 7500
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 5258 7488 5264 7540
rect 5316 7528 5322 7540
rect 10505 7531 10563 7537
rect 10505 7528 10517 7531
rect 5316 7500 10517 7528
rect 5316 7488 5322 7500
rect 10505 7497 10517 7500
rect 10551 7497 10563 7531
rect 11606 7528 11612 7540
rect 10505 7491 10563 7497
rect 10888 7500 11612 7528
rect 10888 7472 10916 7500
rect 11606 7488 11612 7500
rect 11664 7488 11670 7540
rect 11790 7488 11796 7540
rect 11848 7528 11854 7540
rect 12250 7528 12256 7540
rect 11848 7500 12256 7528
rect 11848 7488 11854 7500
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 12437 7531 12495 7537
rect 12437 7528 12449 7531
rect 12360 7500 12449 7528
rect 2547 7364 3096 7392
rect 4172 7432 4936 7460
rect 6273 7463 6331 7469
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 2130 7284 2136 7336
rect 2188 7324 2194 7336
rect 3053 7327 3111 7333
rect 3053 7324 3065 7327
rect 2188 7296 3065 7324
rect 2188 7284 2194 7296
rect 3053 7293 3065 7296
rect 3099 7293 3111 7327
rect 3053 7287 3111 7293
rect 2225 7259 2283 7265
rect 2225 7225 2237 7259
rect 2271 7256 2283 7259
rect 2498 7256 2504 7268
rect 2271 7228 2504 7256
rect 2271 7225 2283 7228
rect 2225 7219 2283 7225
rect 2498 7216 2504 7228
rect 2556 7216 2562 7268
rect 3320 7259 3378 7265
rect 3320 7225 3332 7259
rect 3366 7256 3378 7259
rect 4172 7256 4200 7432
rect 6273 7429 6285 7463
rect 6319 7460 6331 7463
rect 6822 7460 6828 7472
rect 6319 7432 6828 7460
rect 6319 7429 6331 7432
rect 6273 7423 6331 7429
rect 6822 7420 6828 7432
rect 6880 7420 6886 7472
rect 8205 7463 8263 7469
rect 8205 7429 8217 7463
rect 8251 7429 8263 7463
rect 8205 7423 8263 7429
rect 4246 7352 4252 7404
rect 4304 7392 4310 7404
rect 4614 7392 4620 7404
rect 4304 7364 4620 7392
rect 4304 7352 4310 7364
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 6086 7352 6092 7404
rect 6144 7392 6150 7404
rect 6144 7364 6960 7392
rect 6144 7352 6150 7364
rect 4893 7327 4951 7333
rect 4893 7293 4905 7327
rect 4939 7324 4951 7327
rect 4982 7324 4988 7336
rect 4939 7296 4988 7324
rect 4939 7293 4951 7296
rect 4893 7287 4951 7293
rect 4982 7284 4988 7296
rect 5040 7284 5046 7336
rect 5994 7324 6000 7336
rect 5092 7296 6000 7324
rect 5092 7256 5120 7296
rect 5994 7284 6000 7296
rect 6052 7284 6058 7336
rect 6730 7284 6736 7336
rect 6788 7324 6794 7336
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 6788 7296 6837 7324
rect 6788 7284 6794 7296
rect 6825 7293 6837 7296
rect 6871 7293 6883 7327
rect 6932 7324 6960 7364
rect 6932 7296 7227 7324
rect 6825 7287 6883 7293
rect 3366 7228 4200 7256
rect 4356 7228 5120 7256
rect 5160 7259 5218 7265
rect 3366 7225 3378 7228
rect 3320 7219 3378 7225
rect 2317 7191 2375 7197
rect 2317 7157 2329 7191
rect 2363 7188 2375 7191
rect 4356 7188 4384 7228
rect 5160 7225 5172 7259
rect 5206 7256 5218 7259
rect 6178 7256 6184 7268
rect 5206 7228 6184 7256
rect 5206 7225 5218 7228
rect 5160 7219 5218 7225
rect 6178 7216 6184 7228
rect 6236 7216 6242 7268
rect 7006 7216 7012 7268
rect 7064 7265 7070 7268
rect 7064 7259 7128 7265
rect 7064 7225 7082 7259
rect 7116 7225 7128 7259
rect 7199 7256 7227 7296
rect 7650 7284 7656 7336
rect 7708 7324 7714 7336
rect 8220 7324 8248 7423
rect 9766 7420 9772 7472
rect 9824 7460 9830 7472
rect 10226 7460 10232 7472
rect 9824 7432 10232 7460
rect 9824 7420 9830 7432
rect 10226 7420 10232 7432
rect 10284 7460 10290 7472
rect 10870 7460 10876 7472
rect 10284 7432 10876 7460
rect 10284 7420 10290 7432
rect 10870 7420 10876 7432
rect 10928 7420 10934 7472
rect 10962 7420 10968 7472
rect 11020 7460 11026 7472
rect 12360 7460 12388 7500
rect 12437 7497 12449 7500
rect 12483 7497 12495 7531
rect 12437 7491 12495 7497
rect 13633 7531 13691 7537
rect 13633 7497 13645 7531
rect 13679 7528 13691 7531
rect 14366 7528 14372 7540
rect 13679 7500 14372 7528
rect 13679 7497 13691 7500
rect 13633 7491 13691 7497
rect 14366 7488 14372 7500
rect 14424 7488 14430 7540
rect 11020 7432 12388 7460
rect 11020 7420 11026 7432
rect 8294 7352 8300 7404
rect 8352 7392 8358 7404
rect 10778 7392 10784 7404
rect 8352 7364 8800 7392
rect 8352 7352 8358 7364
rect 8662 7324 8668 7336
rect 7708 7296 8248 7324
rect 8623 7296 8668 7324
rect 7708 7284 7714 7296
rect 8662 7284 8668 7296
rect 8720 7284 8726 7336
rect 8772 7324 8800 7364
rect 10060 7364 10784 7392
rect 10060 7324 10088 7364
rect 10778 7352 10784 7364
rect 10836 7352 10842 7404
rect 11054 7392 11060 7404
rect 11015 7364 11060 7392
rect 11054 7352 11060 7364
rect 11112 7392 11118 7404
rect 11701 7395 11759 7401
rect 11112 7364 11652 7392
rect 11112 7352 11118 7364
rect 11624 7336 11652 7364
rect 11701 7361 11713 7395
rect 11747 7392 11759 7395
rect 12250 7392 12256 7404
rect 11747 7364 12256 7392
rect 11747 7361 11759 7364
rect 11701 7355 11759 7361
rect 12250 7352 12256 7364
rect 12308 7352 12314 7404
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 12360 7364 13001 7392
rect 8772 7296 10088 7324
rect 10134 7284 10140 7336
rect 10192 7324 10198 7336
rect 10870 7324 10876 7336
rect 10192 7296 10793 7324
rect 10831 7296 10876 7324
rect 10192 7284 10198 7296
rect 8910 7259 8968 7265
rect 8910 7256 8922 7259
rect 7199 7228 8922 7256
rect 7064 7219 7128 7225
rect 8910 7225 8922 7228
rect 8956 7225 8968 7259
rect 8910 7219 8968 7225
rect 7064 7216 7070 7219
rect 9306 7216 9312 7268
rect 9364 7256 9370 7268
rect 10765 7256 10793 7296
rect 10870 7284 10876 7296
rect 10928 7284 10934 7336
rect 10965 7327 11023 7333
rect 10965 7293 10977 7327
rect 11011 7324 11023 7327
rect 11330 7324 11336 7336
rect 11011 7296 11336 7324
rect 11011 7293 11023 7296
rect 10965 7287 11023 7293
rect 11330 7284 11336 7296
rect 11388 7284 11394 7336
rect 11606 7324 11612 7336
rect 11519 7296 11612 7324
rect 11606 7284 11612 7296
rect 11664 7324 11670 7336
rect 12360 7324 12388 7364
rect 12989 7361 13001 7364
rect 13035 7361 13047 7395
rect 12989 7355 13047 7361
rect 13906 7352 13912 7404
rect 13964 7392 13970 7404
rect 14093 7395 14151 7401
rect 14093 7392 14105 7395
rect 13964 7364 14105 7392
rect 13964 7352 13970 7364
rect 14093 7361 14105 7364
rect 14139 7361 14151 7395
rect 14093 7355 14151 7361
rect 14182 7352 14188 7404
rect 14240 7392 14246 7404
rect 14277 7395 14335 7401
rect 14277 7392 14289 7395
rect 14240 7364 14289 7392
rect 14240 7352 14246 7364
rect 14277 7361 14289 7364
rect 14323 7361 14335 7395
rect 14277 7355 14335 7361
rect 12805 7327 12863 7333
rect 12805 7324 12817 7327
rect 11664 7296 12388 7324
rect 12636 7296 12817 7324
rect 11664 7284 11670 7296
rect 11698 7256 11704 7268
rect 9364 7228 10180 7256
rect 10765 7228 11704 7256
rect 9364 7216 9370 7228
rect 2363 7160 4384 7188
rect 2363 7157 2375 7160
rect 2317 7151 2375 7157
rect 5258 7148 5264 7200
rect 5316 7188 5322 7200
rect 5810 7188 5816 7200
rect 5316 7160 5816 7188
rect 5316 7148 5322 7160
rect 5810 7148 5816 7160
rect 5868 7148 5874 7200
rect 7190 7148 7196 7200
rect 7248 7188 7254 7200
rect 10045 7191 10103 7197
rect 10045 7188 10057 7191
rect 7248 7160 10057 7188
rect 7248 7148 7254 7160
rect 10045 7157 10057 7160
rect 10091 7157 10103 7191
rect 10152 7188 10180 7228
rect 11698 7216 11704 7228
rect 11756 7216 11762 7268
rect 12636 7200 12664 7296
rect 12805 7293 12817 7296
rect 12851 7293 12863 7327
rect 12805 7287 12863 7293
rect 12894 7284 12900 7336
rect 12952 7324 12958 7336
rect 14001 7327 14059 7333
rect 14001 7324 14013 7327
rect 12952 7296 14013 7324
rect 12952 7284 12958 7296
rect 14001 7293 14013 7296
rect 14047 7293 14059 7327
rect 14001 7287 14059 7293
rect 14642 7284 14648 7336
rect 14700 7324 14706 7336
rect 14829 7327 14887 7333
rect 14829 7324 14841 7327
rect 14700 7296 14841 7324
rect 14700 7284 14706 7296
rect 14829 7293 14841 7296
rect 14875 7293 14887 7327
rect 14829 7287 14887 7293
rect 12250 7188 12256 7200
rect 10152 7160 12256 7188
rect 10045 7151 10103 7157
rect 12250 7148 12256 7160
rect 12308 7148 12314 7200
rect 12618 7148 12624 7200
rect 12676 7148 12682 7200
rect 12894 7188 12900 7200
rect 12855 7160 12900 7188
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 13998 7148 14004 7200
rect 14056 7188 14062 7200
rect 14366 7188 14372 7200
rect 14056 7160 14372 7188
rect 14056 7148 14062 7160
rect 14366 7148 14372 7160
rect 14424 7148 14430 7200
rect 15010 7188 15016 7200
rect 14971 7160 15016 7188
rect 15010 7148 15016 7160
rect 15068 7148 15074 7200
rect 1104 7098 15824 7120
rect 1104 7046 5912 7098
rect 5964 7046 5976 7098
rect 6028 7046 6040 7098
rect 6092 7046 6104 7098
rect 6156 7046 10843 7098
rect 10895 7046 10907 7098
rect 10959 7046 10971 7098
rect 11023 7046 11035 7098
rect 11087 7046 15824 7098
rect 1104 7024 15824 7046
rect 4982 6944 4988 6996
rect 5040 6984 5046 6996
rect 5442 6984 5448 6996
rect 5040 6956 5448 6984
rect 5040 6944 5046 6956
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 7006 6944 7012 6996
rect 7064 6984 7070 6996
rect 8941 6987 8999 6993
rect 8941 6984 8953 6987
rect 7064 6956 8953 6984
rect 7064 6944 7070 6956
rect 8941 6953 8953 6956
rect 8987 6984 8999 6987
rect 9490 6984 9496 6996
rect 8987 6956 9496 6984
rect 8987 6953 8999 6956
rect 8941 6947 8999 6953
rect 9490 6944 9496 6956
rect 9548 6944 9554 6996
rect 10045 6987 10103 6993
rect 10045 6953 10057 6987
rect 10091 6984 10103 6987
rect 11514 6984 11520 6996
rect 10091 6956 11520 6984
rect 10091 6953 10103 6956
rect 10045 6947 10103 6953
rect 11514 6944 11520 6956
rect 11572 6944 11578 6996
rect 11698 6944 11704 6996
rect 11756 6984 11762 6996
rect 12437 6987 12495 6993
rect 12437 6984 12449 6987
rect 11756 6956 12449 6984
rect 11756 6944 11762 6956
rect 12437 6953 12449 6956
rect 12483 6953 12495 6987
rect 12437 6947 12495 6953
rect 1857 6919 1915 6925
rect 1857 6885 1869 6919
rect 1903 6916 1915 6919
rect 2774 6916 2780 6928
rect 1903 6888 2780 6916
rect 1903 6885 1915 6888
rect 1857 6879 1915 6885
rect 2774 6876 2780 6888
rect 2832 6876 2838 6928
rect 4893 6919 4951 6925
rect 4893 6885 4905 6919
rect 4939 6916 4951 6919
rect 10502 6916 10508 6928
rect 4939 6888 10508 6916
rect 4939 6885 4951 6888
rect 4893 6879 4951 6885
rect 10502 6876 10508 6888
rect 10560 6876 10566 6928
rect 10686 6876 10692 6928
rect 10744 6916 10750 6928
rect 11241 6919 11299 6925
rect 11241 6916 11253 6919
rect 10744 6888 11253 6916
rect 10744 6876 10750 6888
rect 11241 6885 11253 6888
rect 11287 6885 11299 6919
rect 12452 6916 12480 6947
rect 13170 6944 13176 6996
rect 13228 6984 13234 6996
rect 13265 6987 13323 6993
rect 13265 6984 13277 6987
rect 13228 6956 13277 6984
rect 13228 6944 13234 6956
rect 13265 6953 13277 6956
rect 13311 6953 13323 6987
rect 13265 6947 13323 6953
rect 13630 6944 13636 6996
rect 13688 6984 13694 6996
rect 14826 6984 14832 6996
rect 13688 6956 14832 6984
rect 13688 6944 13694 6956
rect 14826 6944 14832 6956
rect 14884 6944 14890 6996
rect 14090 6916 14096 6928
rect 12452 6888 14096 6916
rect 11241 6879 11299 6885
rect 14090 6876 14096 6888
rect 14148 6876 14154 6928
rect 1578 6848 1584 6860
rect 1539 6820 1584 6848
rect 1578 6808 1584 6820
rect 1636 6808 1642 6860
rect 2400 6851 2458 6857
rect 2400 6817 2412 6851
rect 2446 6848 2458 6851
rect 4430 6848 4436 6860
rect 2446 6820 4436 6848
rect 2446 6817 2458 6820
rect 2400 6811 2458 6817
rect 4430 6808 4436 6820
rect 4488 6808 4494 6860
rect 5442 6808 5448 6860
rect 5500 6848 5506 6860
rect 5721 6851 5779 6857
rect 5721 6848 5733 6851
rect 5500 6820 5733 6848
rect 5500 6808 5506 6820
rect 5721 6817 5733 6820
rect 5767 6817 5779 6851
rect 5721 6811 5779 6817
rect 5988 6851 6046 6857
rect 5988 6817 6000 6851
rect 6034 6848 6046 6851
rect 6546 6848 6552 6860
rect 6034 6820 6552 6848
rect 6034 6817 6046 6820
rect 5988 6811 6046 6817
rect 6546 6808 6552 6820
rect 6604 6808 6610 6860
rect 6730 6808 6736 6860
rect 6788 6848 6794 6860
rect 7558 6848 7564 6860
rect 6788 6820 7564 6848
rect 6788 6808 6794 6820
rect 7558 6808 7564 6820
rect 7616 6808 7622 6860
rect 7834 6857 7840 6860
rect 7828 6848 7840 6857
rect 7795 6820 7840 6848
rect 7828 6811 7840 6820
rect 7834 6808 7840 6811
rect 7892 6808 7898 6860
rect 8110 6808 8116 6860
rect 8168 6848 8174 6860
rect 8168 6820 10548 6848
rect 8168 6808 8174 6820
rect 2130 6780 2136 6792
rect 2091 6752 2136 6780
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 4985 6783 5043 6789
rect 4985 6749 4997 6783
rect 5031 6749 5043 6783
rect 4985 6743 5043 6749
rect 5169 6783 5227 6789
rect 5169 6749 5181 6783
rect 5215 6780 5227 6783
rect 5626 6780 5632 6792
rect 5215 6752 5632 6780
rect 5215 6749 5227 6752
rect 5169 6743 5227 6749
rect 3513 6715 3571 6721
rect 3513 6681 3525 6715
rect 3559 6712 3571 6715
rect 3786 6712 3792 6724
rect 3559 6684 3792 6712
rect 3559 6681 3571 6684
rect 3513 6675 3571 6681
rect 3786 6672 3792 6684
rect 3844 6672 3850 6724
rect 4525 6647 4583 6653
rect 4525 6613 4537 6647
rect 4571 6644 4583 6647
rect 4890 6644 4896 6656
rect 4571 6616 4896 6644
rect 4571 6613 4583 6616
rect 4525 6607 4583 6613
rect 4890 6604 4896 6616
rect 4948 6604 4954 6656
rect 5000 6644 5028 6743
rect 5626 6740 5632 6752
rect 5684 6740 5690 6792
rect 10134 6780 10140 6792
rect 10095 6752 10140 6780
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 10318 6740 10324 6792
rect 10376 6780 10382 6792
rect 10520 6780 10548 6820
rect 11146 6808 11152 6860
rect 11204 6848 11210 6860
rect 11330 6848 11336 6860
rect 11204 6820 11336 6848
rect 11204 6808 11210 6820
rect 11330 6808 11336 6820
rect 11388 6808 11394 6860
rect 11698 6808 11704 6860
rect 11756 6848 11762 6860
rect 11882 6848 11888 6860
rect 11756 6820 11888 6848
rect 11756 6808 11762 6820
rect 11882 6808 11888 6820
rect 11940 6848 11946 6860
rect 13630 6848 13636 6860
rect 11940 6820 12756 6848
rect 13591 6820 13636 6848
rect 11940 6808 11946 6820
rect 11425 6783 11483 6789
rect 11425 6780 11437 6783
rect 10376 6752 10421 6780
rect 10520 6752 11437 6780
rect 10376 6740 10382 6752
rect 11425 6749 11437 6752
rect 11471 6749 11483 6783
rect 12526 6780 12532 6792
rect 12487 6752 12532 6780
rect 11425 6743 11483 6749
rect 12526 6740 12532 6752
rect 12584 6740 12590 6792
rect 12621 6783 12679 6789
rect 12621 6749 12633 6783
rect 12667 6749 12679 6783
rect 12728 6780 12756 6820
rect 13630 6808 13636 6820
rect 13688 6808 13694 6860
rect 13722 6808 13728 6860
rect 13780 6848 13786 6860
rect 13780 6820 13825 6848
rect 13780 6808 13786 6820
rect 14182 6808 14188 6860
rect 14240 6848 14246 6860
rect 14461 6851 14519 6857
rect 14461 6848 14473 6851
rect 14240 6820 14473 6848
rect 14240 6808 14246 6820
rect 14461 6817 14473 6820
rect 14507 6817 14519 6851
rect 14461 6811 14519 6817
rect 13817 6783 13875 6789
rect 13817 6780 13829 6783
rect 12728 6752 13829 6780
rect 12621 6743 12679 6749
rect 13817 6749 13829 6752
rect 13863 6749 13875 6783
rect 13817 6743 13875 6749
rect 6840 6684 7604 6712
rect 6840 6644 6868 6684
rect 5000 6616 6868 6644
rect 6914 6604 6920 6656
rect 6972 6644 6978 6656
rect 7101 6647 7159 6653
rect 7101 6644 7113 6647
rect 6972 6616 7113 6644
rect 6972 6604 6978 6616
rect 7101 6613 7113 6616
rect 7147 6613 7159 6647
rect 7576 6644 7604 6684
rect 8662 6672 8668 6724
rect 8720 6712 8726 6724
rect 12636 6712 12664 6743
rect 14734 6712 14740 6724
rect 8720 6684 12664 6712
rect 12728 6684 14740 6712
rect 8720 6672 8726 6684
rect 8846 6644 8852 6656
rect 7576 6616 8852 6644
rect 7101 6607 7159 6613
rect 8846 6604 8852 6616
rect 8904 6604 8910 6656
rect 9674 6644 9680 6656
rect 9635 6616 9680 6644
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 10318 6604 10324 6656
rect 10376 6644 10382 6656
rect 10594 6644 10600 6656
rect 10376 6616 10600 6644
rect 10376 6604 10382 6616
rect 10594 6604 10600 6616
rect 10652 6604 10658 6656
rect 10686 6604 10692 6656
rect 10744 6644 10750 6656
rect 10873 6647 10931 6653
rect 10873 6644 10885 6647
rect 10744 6616 10885 6644
rect 10744 6604 10750 6616
rect 10873 6613 10885 6616
rect 10919 6613 10931 6647
rect 10873 6607 10931 6613
rect 11330 6604 11336 6656
rect 11388 6644 11394 6656
rect 12069 6647 12127 6653
rect 12069 6644 12081 6647
rect 11388 6616 12081 6644
rect 11388 6604 11394 6616
rect 12069 6613 12081 6616
rect 12115 6613 12127 6647
rect 12069 6607 12127 6613
rect 12526 6604 12532 6656
rect 12584 6644 12590 6656
rect 12728 6644 12756 6684
rect 14734 6672 14740 6684
rect 14792 6672 14798 6724
rect 12584 6616 12756 6644
rect 12584 6604 12590 6616
rect 13170 6604 13176 6656
rect 13228 6644 13234 6656
rect 14645 6647 14703 6653
rect 14645 6644 14657 6647
rect 13228 6616 14657 6644
rect 13228 6604 13234 6616
rect 14645 6613 14657 6616
rect 14691 6613 14703 6647
rect 14645 6607 14703 6613
rect 1104 6554 15824 6576
rect 1104 6502 3447 6554
rect 3499 6502 3511 6554
rect 3563 6502 3575 6554
rect 3627 6502 3639 6554
rect 3691 6502 8378 6554
rect 8430 6502 8442 6554
rect 8494 6502 8506 6554
rect 8558 6502 8570 6554
rect 8622 6502 13308 6554
rect 13360 6502 13372 6554
rect 13424 6502 13436 6554
rect 13488 6502 13500 6554
rect 13552 6502 15824 6554
rect 1104 6480 15824 6502
rect 5258 6440 5264 6452
rect 2516 6412 5264 6440
rect 1946 6332 1952 6384
rect 2004 6372 2010 6384
rect 2314 6372 2320 6384
rect 2004 6344 2320 6372
rect 2004 6332 2010 6344
rect 2314 6332 2320 6344
rect 2372 6332 2378 6384
rect 1302 6264 1308 6316
rect 1360 6304 1366 6316
rect 2130 6304 2136 6316
rect 1360 6276 2136 6304
rect 1360 6264 1366 6276
rect 2130 6264 2136 6276
rect 2188 6264 2194 6316
rect 2516 6313 2544 6412
rect 5258 6400 5264 6412
rect 5316 6400 5322 6452
rect 5626 6400 5632 6452
rect 5684 6440 5690 6452
rect 6273 6443 6331 6449
rect 6273 6440 6285 6443
rect 5684 6412 6285 6440
rect 5684 6400 5690 6412
rect 6273 6409 6285 6412
rect 6319 6409 6331 6443
rect 6273 6403 6331 6409
rect 6454 6400 6460 6452
rect 6512 6440 6518 6452
rect 10502 6440 10508 6452
rect 6512 6412 9720 6440
rect 10463 6412 10508 6440
rect 6512 6400 6518 6412
rect 2501 6307 2559 6313
rect 2501 6273 2513 6307
rect 2547 6273 2559 6307
rect 9692 6304 9720 6412
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 10594 6400 10600 6452
rect 10652 6440 10658 6452
rect 10778 6440 10784 6452
rect 10652 6412 10784 6440
rect 10652 6400 10658 6412
rect 10778 6400 10784 6412
rect 10836 6400 10842 6452
rect 12437 6443 12495 6449
rect 12437 6409 12449 6443
rect 12483 6440 12495 6443
rect 13630 6440 13636 6452
rect 12483 6412 13636 6440
rect 12483 6409 12495 6412
rect 12437 6403 12495 6409
rect 13630 6400 13636 6412
rect 13688 6400 13694 6452
rect 9766 6332 9772 6384
rect 9824 6372 9830 6384
rect 10045 6375 10103 6381
rect 10045 6372 10057 6375
rect 9824 6344 10057 6372
rect 9824 6332 9830 6344
rect 10045 6341 10057 6344
rect 10091 6372 10103 6375
rect 12710 6372 12716 6384
rect 10091 6344 12716 6372
rect 10091 6341 10103 6344
rect 10045 6335 10103 6341
rect 12710 6332 12716 6344
rect 12768 6332 12774 6384
rect 13078 6332 13084 6384
rect 13136 6372 13142 6384
rect 13136 6344 14872 6372
rect 13136 6332 13142 6344
rect 2501 6267 2559 6273
rect 5920 6276 6960 6304
rect 9692 6276 10272 6304
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6205 1455 6239
rect 2148 6236 2176 6264
rect 3053 6239 3111 6245
rect 3053 6236 3065 6239
rect 2148 6208 3065 6236
rect 1397 6199 1455 6205
rect 3053 6205 3065 6208
rect 3099 6236 3111 6239
rect 4893 6239 4951 6245
rect 4893 6236 4905 6239
rect 3099 6208 4905 6236
rect 3099 6205 3111 6208
rect 3053 6199 3111 6205
rect 4893 6205 4905 6208
rect 4939 6236 4951 6239
rect 5442 6236 5448 6248
rect 4939 6208 5448 6236
rect 4939 6205 4951 6208
rect 4893 6199 4951 6205
rect 1412 6168 1440 6199
rect 5442 6196 5448 6208
rect 5500 6196 5506 6248
rect 5718 6196 5724 6248
rect 5776 6236 5782 6248
rect 5920 6236 5948 6276
rect 6822 6236 6828 6248
rect 5776 6208 5948 6236
rect 6783 6208 6828 6236
rect 5776 6196 5782 6208
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 6932 6236 6960 6276
rect 8110 6236 8116 6248
rect 6932 6208 8116 6236
rect 8110 6196 8116 6208
rect 8168 6196 8174 6248
rect 8665 6239 8723 6245
rect 8665 6205 8677 6239
rect 8711 6236 8723 6239
rect 9214 6236 9220 6248
rect 8711 6208 9220 6236
rect 8711 6205 8723 6208
rect 8665 6199 8723 6205
rect 2498 6168 2504 6180
rect 1412 6140 2504 6168
rect 2498 6128 2504 6140
rect 2556 6128 2562 6180
rect 3326 6177 3332 6180
rect 3320 6168 3332 6177
rect 3287 6140 3332 6168
rect 3320 6131 3332 6140
rect 3326 6128 3332 6131
rect 3384 6128 3390 6180
rect 5160 6171 5218 6177
rect 5160 6137 5172 6171
rect 5206 6168 5218 6171
rect 5206 6140 6875 6168
rect 5206 6137 5218 6140
rect 5160 6131 5218 6137
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 1854 6100 1860 6112
rect 1815 6072 1860 6100
rect 1854 6060 1860 6072
rect 1912 6060 1918 6112
rect 2222 6100 2228 6112
rect 2183 6072 2228 6100
rect 2222 6060 2228 6072
rect 2280 6060 2286 6112
rect 2314 6060 2320 6112
rect 2372 6100 2378 6112
rect 4430 6100 4436 6112
rect 2372 6072 2417 6100
rect 4343 6072 4436 6100
rect 2372 6060 2378 6072
rect 4430 6060 4436 6072
rect 4488 6100 4494 6112
rect 5718 6100 5724 6112
rect 4488 6072 5724 6100
rect 4488 6060 4494 6072
rect 5718 6060 5724 6072
rect 5776 6060 5782 6112
rect 6847 6100 6875 6140
rect 6914 6128 6920 6180
rect 6972 6168 6978 6180
rect 7070 6171 7128 6177
rect 7070 6168 7082 6171
rect 6972 6140 7082 6168
rect 6972 6128 6978 6140
rect 7070 6137 7082 6140
rect 7116 6137 7128 6171
rect 7070 6131 7128 6137
rect 7558 6128 7564 6180
rect 7616 6168 7622 6180
rect 8680 6168 8708 6199
rect 9214 6196 9220 6208
rect 9272 6196 9278 6248
rect 9490 6196 9496 6248
rect 9548 6236 9554 6248
rect 10134 6236 10140 6248
rect 9548 6208 10140 6236
rect 9548 6196 9554 6208
rect 10134 6196 10140 6208
rect 10192 6196 10198 6248
rect 10244 6236 10272 6276
rect 10502 6264 10508 6316
rect 10560 6304 10566 6316
rect 11057 6307 11115 6313
rect 11057 6304 11069 6307
rect 10560 6276 11069 6304
rect 10560 6264 10566 6276
rect 11057 6273 11069 6276
rect 11103 6273 11115 6307
rect 11057 6267 11115 6273
rect 12158 6264 12164 6316
rect 12216 6304 12222 6316
rect 12989 6307 13047 6313
rect 12989 6304 13001 6307
rect 12216 6276 13001 6304
rect 12216 6264 12222 6276
rect 12989 6273 13001 6276
rect 13035 6273 13047 6307
rect 12989 6267 13047 6273
rect 13262 6264 13268 6316
rect 13320 6304 13326 6316
rect 14185 6307 14243 6313
rect 14185 6304 14197 6307
rect 13320 6276 14197 6304
rect 13320 6264 13326 6276
rect 14185 6273 14197 6276
rect 14231 6273 14243 6307
rect 14185 6267 14243 6273
rect 10686 6236 10692 6248
rect 10244 6208 10692 6236
rect 10686 6196 10692 6208
rect 10744 6196 10750 6248
rect 10962 6236 10968 6248
rect 10923 6208 10968 6236
rect 10962 6196 10968 6208
rect 11020 6196 11026 6248
rect 14844 6245 14872 6344
rect 14093 6239 14151 6245
rect 14093 6236 14105 6239
rect 11072 6208 14105 6236
rect 7616 6140 8708 6168
rect 8932 6171 8990 6177
rect 7616 6128 7622 6140
rect 8932 6137 8944 6171
rect 8978 6137 8990 6171
rect 8932 6131 8990 6137
rect 7374 6100 7380 6112
rect 6847 6072 7380 6100
rect 7374 6060 7380 6072
rect 7432 6100 7438 6112
rect 8202 6100 8208 6112
rect 7432 6072 8208 6100
rect 7432 6060 7438 6072
rect 8202 6060 8208 6072
rect 8260 6060 8266 6112
rect 8754 6060 8760 6112
rect 8812 6100 8818 6112
rect 8947 6100 8975 6131
rect 9398 6128 9404 6180
rect 9456 6168 9462 6180
rect 10873 6171 10931 6177
rect 10873 6168 10885 6171
rect 9456 6140 10885 6168
rect 9456 6128 9462 6140
rect 10873 6137 10885 6140
rect 10919 6137 10931 6171
rect 10873 6131 10931 6137
rect 9950 6100 9956 6112
rect 8812 6072 9956 6100
rect 8812 6060 8818 6072
rect 9950 6060 9956 6072
rect 10008 6060 10014 6112
rect 10686 6060 10692 6112
rect 10744 6100 10750 6112
rect 11072 6100 11100 6208
rect 14093 6205 14105 6208
rect 14139 6205 14151 6239
rect 14093 6199 14151 6205
rect 14829 6239 14887 6245
rect 14829 6205 14841 6239
rect 14875 6205 14887 6239
rect 14829 6199 14887 6205
rect 11974 6128 11980 6180
rect 12032 6168 12038 6180
rect 12805 6171 12863 6177
rect 12805 6168 12817 6171
rect 12032 6140 12817 6168
rect 12032 6128 12038 6140
rect 12805 6137 12817 6140
rect 12851 6168 12863 6171
rect 13265 6171 13323 6177
rect 13265 6168 13277 6171
rect 12851 6140 13277 6168
rect 12851 6137 12863 6140
rect 12805 6131 12863 6137
rect 13265 6137 13277 6140
rect 13311 6137 13323 6171
rect 13722 6168 13728 6180
rect 13265 6131 13323 6137
rect 13464 6140 13728 6168
rect 10744 6072 11100 6100
rect 11701 6103 11759 6109
rect 10744 6060 10750 6072
rect 11701 6069 11713 6103
rect 11747 6100 11759 6103
rect 12342 6100 12348 6112
rect 11747 6072 12348 6100
rect 11747 6069 11759 6072
rect 11701 6063 11759 6069
rect 12342 6060 12348 6072
rect 12400 6060 12406 6112
rect 12897 6103 12955 6109
rect 12897 6069 12909 6103
rect 12943 6100 12955 6103
rect 13464 6100 13492 6140
rect 13722 6128 13728 6140
rect 13780 6128 13786 6180
rect 14001 6171 14059 6177
rect 14001 6137 14013 6171
rect 14047 6168 14059 6171
rect 14182 6168 14188 6180
rect 14047 6140 14188 6168
rect 14047 6137 14059 6140
rect 14001 6131 14059 6137
rect 14182 6128 14188 6140
rect 14240 6128 14246 6180
rect 13630 6100 13636 6112
rect 12943 6072 13492 6100
rect 13591 6072 13636 6100
rect 12943 6069 12955 6072
rect 12897 6063 12955 6069
rect 13630 6060 13636 6072
rect 13688 6060 13694 6112
rect 13814 6060 13820 6112
rect 13872 6100 13878 6112
rect 15013 6103 15071 6109
rect 15013 6100 15025 6103
rect 13872 6072 15025 6100
rect 13872 6060 13878 6072
rect 15013 6069 15025 6072
rect 15059 6069 15071 6103
rect 15013 6063 15071 6069
rect 1104 6010 15824 6032
rect 1104 5958 5912 6010
rect 5964 5958 5976 6010
rect 6028 5958 6040 6010
rect 6092 5958 6104 6010
rect 6156 5958 10843 6010
rect 10895 5958 10907 6010
rect 10959 5958 10971 6010
rect 11023 5958 11035 6010
rect 11087 5958 15824 6010
rect 1104 5936 15824 5958
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 1854 5896 1860 5908
rect 1627 5868 1860 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 1854 5856 1860 5868
rect 1912 5856 1918 5908
rect 2041 5899 2099 5905
rect 2041 5865 2053 5899
rect 2087 5896 2099 5899
rect 4890 5896 4896 5908
rect 2087 5868 4752 5896
rect 4851 5868 4896 5896
rect 2087 5865 2099 5868
rect 2041 5859 2099 5865
rect 1949 5831 2007 5837
rect 1949 5797 1961 5831
rect 1995 5828 2007 5831
rect 4430 5828 4436 5840
rect 1995 5800 4436 5828
rect 1995 5797 2007 5800
rect 1949 5791 2007 5797
rect 4430 5788 4436 5800
rect 4488 5788 4494 5840
rect 4724 5828 4752 5868
rect 4890 5856 4896 5868
rect 4948 5856 4954 5908
rect 5442 5856 5448 5908
rect 5500 5896 5506 5908
rect 5718 5896 5724 5908
rect 5500 5868 5724 5896
rect 5500 5856 5506 5868
rect 5718 5856 5724 5868
rect 5776 5856 5782 5908
rect 5920 5868 6224 5896
rect 5920 5828 5948 5868
rect 4724 5800 5948 5828
rect 5988 5831 6046 5837
rect 5988 5797 6000 5831
rect 6034 5828 6046 5831
rect 6086 5828 6092 5840
rect 6034 5800 6092 5828
rect 6034 5797 6046 5800
rect 5988 5791 6046 5797
rect 6086 5788 6092 5800
rect 6144 5788 6150 5840
rect 6196 5828 6224 5868
rect 6546 5856 6552 5908
rect 6604 5896 6610 5908
rect 7101 5899 7159 5905
rect 7101 5896 7113 5899
rect 6604 5868 7113 5896
rect 6604 5856 6610 5868
rect 7101 5865 7113 5868
rect 7147 5865 7159 5899
rect 10226 5896 10232 5908
rect 7101 5859 7159 5865
rect 10152 5868 10232 5896
rect 9674 5828 9680 5840
rect 6196 5800 9680 5828
rect 9674 5788 9680 5800
rect 9732 5788 9738 5840
rect 10045 5831 10103 5837
rect 10045 5797 10057 5831
rect 10091 5828 10103 5831
rect 10152 5828 10180 5868
rect 10226 5856 10232 5868
rect 10284 5856 10290 5908
rect 11241 5899 11299 5905
rect 11241 5865 11253 5899
rect 11287 5896 11299 5899
rect 11974 5896 11980 5908
rect 11287 5868 11980 5896
rect 11287 5865 11299 5868
rect 11241 5859 11299 5865
rect 11974 5856 11980 5868
rect 12032 5856 12038 5908
rect 12069 5899 12127 5905
rect 12069 5865 12081 5899
rect 12115 5896 12127 5899
rect 12342 5896 12348 5908
rect 12115 5868 12348 5896
rect 12115 5865 12127 5868
rect 12069 5859 12127 5865
rect 12342 5856 12348 5868
rect 12400 5856 12406 5908
rect 13446 5856 13452 5908
rect 13504 5896 13510 5908
rect 13633 5899 13691 5905
rect 13633 5896 13645 5899
rect 13504 5868 13645 5896
rect 13504 5856 13510 5868
rect 13633 5865 13645 5868
rect 13679 5865 13691 5899
rect 13633 5859 13691 5865
rect 11330 5828 11336 5840
rect 10091 5800 10180 5828
rect 11291 5800 11336 5828
rect 10091 5797 10103 5800
rect 10045 5791 10103 5797
rect 11330 5788 11336 5800
rect 11388 5788 11394 5840
rect 12437 5831 12495 5837
rect 12437 5797 12449 5831
rect 12483 5828 12495 5831
rect 12526 5828 12532 5840
rect 12483 5800 12532 5828
rect 12483 5797 12495 5800
rect 12437 5791 12495 5797
rect 12526 5788 12532 5800
rect 12584 5788 12590 5840
rect 12710 5788 12716 5840
rect 12768 5828 12774 5840
rect 12986 5828 12992 5840
rect 12768 5800 12992 5828
rect 12768 5788 12774 5800
rect 12986 5788 12992 5800
rect 13044 5788 13050 5840
rect 13538 5788 13544 5840
rect 13596 5828 13602 5840
rect 13725 5831 13783 5837
rect 13725 5828 13737 5831
rect 13596 5800 13737 5828
rect 13596 5788 13602 5800
rect 13725 5797 13737 5800
rect 13771 5797 13783 5831
rect 13725 5791 13783 5797
rect 3145 5763 3203 5769
rect 3145 5729 3157 5763
rect 3191 5729 3203 5763
rect 3145 5723 3203 5729
rect 3237 5763 3295 5769
rect 3237 5729 3249 5763
rect 3283 5760 3295 5763
rect 6822 5760 6828 5772
rect 3283 5732 6828 5760
rect 3283 5729 3295 5732
rect 3237 5723 3295 5729
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5692 2283 5695
rect 2774 5692 2780 5704
rect 2271 5664 2780 5692
rect 2271 5661 2283 5664
rect 2225 5655 2283 5661
rect 2774 5652 2780 5664
rect 2832 5652 2838 5704
rect 3160 5624 3188 5723
rect 6822 5720 6828 5732
rect 6880 5720 6886 5772
rect 7558 5720 7564 5772
rect 7616 5760 7622 5772
rect 7653 5763 7711 5769
rect 7653 5760 7665 5763
rect 7616 5732 7665 5760
rect 7616 5720 7622 5732
rect 7653 5729 7665 5732
rect 7699 5729 7711 5763
rect 7653 5723 7711 5729
rect 7920 5763 7978 5769
rect 7920 5729 7932 5763
rect 7966 5760 7978 5763
rect 9766 5760 9772 5772
rect 7966 5732 9772 5760
rect 7966 5729 7978 5732
rect 7920 5723 7978 5729
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 9950 5720 9956 5772
rect 10008 5760 10014 5772
rect 13262 5760 13268 5772
rect 10008 5732 13268 5760
rect 10008 5720 10014 5732
rect 13262 5720 13268 5732
rect 13320 5720 13326 5772
rect 14461 5763 14519 5769
rect 14461 5729 14473 5763
rect 14507 5760 14519 5763
rect 14550 5760 14556 5772
rect 14507 5732 14556 5760
rect 14507 5729 14519 5732
rect 14461 5723 14519 5729
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5692 3479 5695
rect 4062 5692 4068 5704
rect 3467 5664 4068 5692
rect 3467 5661 3479 5664
rect 3421 5655 3479 5661
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 4982 5692 4988 5704
rect 4943 5664 4988 5692
rect 4982 5652 4988 5664
rect 5040 5652 5046 5704
rect 5169 5695 5227 5701
rect 5169 5661 5181 5695
rect 5215 5692 5227 5695
rect 5534 5692 5540 5704
rect 5215 5664 5540 5692
rect 5215 5661 5227 5664
rect 5169 5655 5227 5661
rect 5534 5652 5540 5664
rect 5592 5652 5598 5704
rect 5718 5692 5724 5704
rect 5679 5664 5724 5692
rect 5718 5652 5724 5664
rect 5776 5652 5782 5704
rect 10137 5695 10195 5701
rect 8680 5664 9812 5692
rect 3160 5596 5580 5624
rect 2777 5559 2835 5565
rect 2777 5525 2789 5559
rect 2823 5556 2835 5559
rect 4430 5556 4436 5568
rect 2823 5528 4436 5556
rect 2823 5525 2835 5528
rect 2777 5519 2835 5525
rect 4430 5516 4436 5528
rect 4488 5516 4494 5568
rect 4525 5559 4583 5565
rect 4525 5525 4537 5559
rect 4571 5556 4583 5559
rect 4890 5556 4896 5568
rect 4571 5528 4896 5556
rect 4571 5525 4583 5528
rect 4525 5519 4583 5525
rect 4890 5516 4896 5528
rect 4948 5516 4954 5568
rect 5552 5556 5580 5596
rect 6730 5584 6736 5636
rect 6788 5624 6794 5636
rect 6788 5596 7696 5624
rect 6788 5584 6794 5596
rect 7006 5556 7012 5568
rect 5552 5528 7012 5556
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 7668 5556 7696 5596
rect 8680 5556 8708 5664
rect 8846 5584 8852 5636
rect 8904 5624 8910 5636
rect 9677 5627 9735 5633
rect 9677 5624 9689 5627
rect 8904 5596 9689 5624
rect 8904 5584 8910 5596
rect 9677 5593 9689 5596
rect 9723 5593 9735 5627
rect 9784 5624 9812 5664
rect 10137 5661 10149 5695
rect 10183 5692 10195 5695
rect 10226 5692 10232 5704
rect 10183 5664 10232 5692
rect 10183 5661 10195 5664
rect 10137 5655 10195 5661
rect 10226 5652 10232 5664
rect 10284 5652 10290 5704
rect 10321 5695 10379 5701
rect 10321 5661 10333 5695
rect 10367 5692 10379 5695
rect 10502 5692 10508 5704
rect 10367 5664 10508 5692
rect 10367 5661 10379 5664
rect 10321 5655 10379 5661
rect 10502 5652 10508 5664
rect 10560 5652 10566 5704
rect 11517 5695 11575 5701
rect 11517 5661 11529 5695
rect 11563 5692 11575 5695
rect 11606 5692 11612 5704
rect 11563 5664 11612 5692
rect 11563 5661 11575 5664
rect 11517 5655 11575 5661
rect 11606 5652 11612 5664
rect 11664 5652 11670 5704
rect 12526 5692 12532 5704
rect 12487 5664 12532 5692
rect 12526 5652 12532 5664
rect 12584 5652 12590 5704
rect 12621 5695 12679 5701
rect 12621 5661 12633 5695
rect 12667 5661 12679 5695
rect 12621 5655 12679 5661
rect 10873 5627 10931 5633
rect 10873 5624 10885 5627
rect 9784 5596 10885 5624
rect 9677 5587 9735 5593
rect 10873 5593 10885 5596
rect 10919 5593 10931 5627
rect 10873 5587 10931 5593
rect 11330 5584 11336 5636
rect 11388 5624 11394 5636
rect 11882 5624 11888 5636
rect 11388 5596 11888 5624
rect 11388 5584 11394 5596
rect 11882 5584 11888 5596
rect 11940 5584 11946 5636
rect 12158 5584 12164 5636
rect 12216 5624 12222 5636
rect 12636 5624 12664 5655
rect 12802 5652 12808 5704
rect 12860 5692 12866 5704
rect 13817 5695 13875 5701
rect 13817 5692 13829 5695
rect 12860 5664 13829 5692
rect 12860 5652 12866 5664
rect 13817 5661 13829 5664
rect 13863 5661 13875 5695
rect 13817 5655 13875 5661
rect 12216 5596 12664 5624
rect 12216 5584 12222 5596
rect 13170 5584 13176 5636
rect 13228 5624 13234 5636
rect 14476 5624 14504 5723
rect 14550 5720 14556 5732
rect 14608 5720 14614 5772
rect 13228 5596 14504 5624
rect 13228 5584 13234 5596
rect 7668 5528 8708 5556
rect 9033 5559 9091 5565
rect 9033 5525 9045 5559
rect 9079 5556 9091 5559
rect 9122 5556 9128 5568
rect 9079 5528 9128 5556
rect 9079 5525 9091 5528
rect 9033 5519 9091 5525
rect 9122 5516 9128 5528
rect 9180 5516 9186 5568
rect 9398 5516 9404 5568
rect 9456 5556 9462 5568
rect 13265 5559 13323 5565
rect 13265 5556 13277 5559
rect 9456 5528 13277 5556
rect 9456 5516 9462 5528
rect 13265 5525 13277 5528
rect 13311 5525 13323 5559
rect 13265 5519 13323 5525
rect 13722 5516 13728 5568
rect 13780 5556 13786 5568
rect 14645 5559 14703 5565
rect 14645 5556 14657 5559
rect 13780 5528 14657 5556
rect 13780 5516 13786 5528
rect 14645 5525 14657 5528
rect 14691 5525 14703 5559
rect 14645 5519 14703 5525
rect 1104 5466 15824 5488
rect 1104 5414 3447 5466
rect 3499 5414 3511 5466
rect 3563 5414 3575 5466
rect 3627 5414 3639 5466
rect 3691 5414 8378 5466
rect 8430 5414 8442 5466
rect 8494 5414 8506 5466
rect 8558 5414 8570 5466
rect 8622 5414 13308 5466
rect 13360 5414 13372 5466
rect 13424 5414 13436 5466
rect 13488 5414 13500 5466
rect 13552 5414 15824 5466
rect 1104 5392 15824 5414
rect 1394 5352 1400 5364
rect 1355 5324 1400 5352
rect 1394 5312 1400 5324
rect 1452 5312 1458 5364
rect 5258 5352 5264 5364
rect 3160 5324 5264 5352
rect 2590 5284 2596 5296
rect 1872 5256 2596 5284
rect 1872 5225 1900 5256
rect 2590 5244 2596 5256
rect 2648 5244 2654 5296
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5185 1915 5219
rect 1857 5179 1915 5185
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5216 2099 5219
rect 2682 5216 2688 5228
rect 2087 5188 2688 5216
rect 2087 5185 2099 5188
rect 2041 5179 2099 5185
rect 2682 5176 2688 5188
rect 2740 5176 2746 5228
rect 2958 5216 2964 5228
rect 2919 5188 2964 5216
rect 2958 5176 2964 5188
rect 3016 5176 3022 5228
rect 3160 5225 3188 5324
rect 5258 5312 5264 5324
rect 5316 5312 5322 5364
rect 5534 5312 5540 5364
rect 5592 5352 5598 5364
rect 6273 5355 6331 5361
rect 6273 5352 6285 5355
rect 5592 5324 6285 5352
rect 5592 5312 5598 5324
rect 6273 5321 6285 5324
rect 6319 5321 6331 5355
rect 6273 5315 6331 5321
rect 7006 5312 7012 5364
rect 7064 5352 7070 5364
rect 9217 5355 9275 5361
rect 9217 5352 9229 5355
rect 7064 5324 8800 5352
rect 7064 5312 7070 5324
rect 3418 5244 3424 5296
rect 3476 5284 3482 5296
rect 4798 5284 4804 5296
rect 3476 5256 4804 5284
rect 3476 5244 3482 5256
rect 4798 5244 4804 5256
rect 4856 5244 4862 5296
rect 8772 5284 8800 5324
rect 8956 5324 9229 5352
rect 8956 5284 8984 5324
rect 9217 5321 9229 5324
rect 9263 5321 9275 5355
rect 9217 5315 9275 5321
rect 9674 5312 9680 5364
rect 9732 5352 9738 5364
rect 12250 5352 12256 5364
rect 9732 5324 12256 5352
rect 9732 5312 9738 5324
rect 12250 5312 12256 5324
rect 12308 5312 12314 5364
rect 12342 5312 12348 5364
rect 12400 5352 12406 5364
rect 12400 5324 14872 5352
rect 12400 5312 12406 5324
rect 8772 5256 8984 5284
rect 9122 5244 9128 5296
rect 9180 5284 9186 5296
rect 9582 5284 9588 5296
rect 9180 5256 9588 5284
rect 9180 5244 9186 5256
rect 9582 5244 9588 5256
rect 9640 5244 9646 5296
rect 9766 5244 9772 5296
rect 9824 5284 9830 5296
rect 10226 5284 10232 5296
rect 9824 5256 10232 5284
rect 9824 5244 9830 5256
rect 10226 5244 10232 5256
rect 10284 5244 10290 5296
rect 10318 5244 10324 5296
rect 10376 5284 10382 5296
rect 10413 5287 10471 5293
rect 10413 5284 10425 5287
rect 10376 5256 10425 5284
rect 10376 5244 10382 5256
rect 10413 5253 10425 5256
rect 10459 5253 10471 5287
rect 13633 5287 13691 5293
rect 13633 5284 13645 5287
rect 10413 5247 10471 5253
rect 10612 5256 13645 5284
rect 3145 5219 3203 5225
rect 3145 5185 3157 5219
rect 3191 5185 3203 5219
rect 3145 5179 3203 5185
rect 4062 5176 4068 5228
rect 4120 5216 4126 5228
rect 4249 5219 4307 5225
rect 4249 5216 4261 5219
rect 4120 5188 4261 5216
rect 4120 5176 4126 5188
rect 4249 5185 4261 5188
rect 4295 5185 4307 5219
rect 4249 5179 4307 5185
rect 6638 5176 6644 5228
rect 6696 5216 6702 5228
rect 6696 5188 7512 5216
rect 6696 5176 6702 5188
rect 1670 5108 1676 5160
rect 1728 5148 1734 5160
rect 1765 5151 1823 5157
rect 1765 5148 1777 5151
rect 1728 5120 1777 5148
rect 1728 5108 1734 5120
rect 1765 5117 1777 5120
rect 1811 5117 1823 5151
rect 1765 5111 1823 5117
rect 2869 5151 2927 5157
rect 2869 5117 2881 5151
rect 2915 5148 2927 5151
rect 4522 5148 4528 5160
rect 2915 5120 4528 5148
rect 2915 5117 2927 5120
rect 2869 5111 2927 5117
rect 4522 5108 4528 5120
rect 4580 5108 4586 5160
rect 4798 5108 4804 5160
rect 4856 5148 4862 5160
rect 4893 5151 4951 5157
rect 4893 5148 4905 5151
rect 4856 5120 4905 5148
rect 4856 5108 4862 5120
rect 4893 5117 4905 5120
rect 4939 5117 4951 5151
rect 4893 5111 4951 5117
rect 5160 5151 5218 5157
rect 5160 5117 5172 5151
rect 5206 5148 5218 5151
rect 5626 5148 5632 5160
rect 5206 5120 5632 5148
rect 5206 5117 5218 5120
rect 5160 5111 5218 5117
rect 5626 5108 5632 5120
rect 5684 5108 5690 5160
rect 6086 5108 6092 5160
rect 6144 5148 6150 5160
rect 6362 5148 6368 5160
rect 6144 5120 6368 5148
rect 6144 5108 6150 5120
rect 6362 5108 6368 5120
rect 6420 5108 6426 5160
rect 7006 5108 7012 5160
rect 7064 5148 7070 5160
rect 7377 5151 7435 5157
rect 7377 5148 7389 5151
rect 7064 5120 7389 5148
rect 7064 5108 7070 5120
rect 7377 5117 7389 5120
rect 7423 5117 7435 5151
rect 7484 5148 7512 5188
rect 8570 5176 8576 5228
rect 8628 5216 8634 5228
rect 9861 5219 9919 5225
rect 9861 5216 9873 5219
rect 8628 5188 9873 5216
rect 8628 5176 8634 5188
rect 9861 5185 9873 5188
rect 9907 5185 9919 5219
rect 9861 5179 9919 5185
rect 9950 5176 9956 5228
rect 10008 5216 10014 5228
rect 10612 5216 10640 5256
rect 13633 5253 13645 5256
rect 13679 5253 13691 5287
rect 13633 5247 13691 5253
rect 10008 5188 10640 5216
rect 10008 5176 10014 5188
rect 10870 5176 10876 5228
rect 10928 5216 10934 5228
rect 10965 5219 11023 5225
rect 10965 5216 10977 5219
rect 10928 5188 10977 5216
rect 10928 5176 10934 5188
rect 10965 5185 10977 5188
rect 11011 5185 11023 5219
rect 10965 5179 11023 5185
rect 11164 5188 11744 5216
rect 8386 5148 8392 5160
rect 7484 5120 8392 5148
rect 7377 5111 7435 5117
rect 8386 5108 8392 5120
rect 8444 5148 8450 5160
rect 10778 5148 10784 5160
rect 8444 5120 10180 5148
rect 10739 5120 10784 5148
rect 8444 5108 8450 5120
rect 4065 5083 4123 5089
rect 4065 5049 4077 5083
rect 4111 5080 4123 5083
rect 7466 5080 7472 5092
rect 4111 5052 7472 5080
rect 4111 5049 4123 5052
rect 4065 5043 4123 5049
rect 7466 5040 7472 5052
rect 7524 5040 7530 5092
rect 7644 5083 7702 5089
rect 7644 5049 7656 5083
rect 7690 5080 7702 5083
rect 7834 5080 7840 5092
rect 7690 5052 7840 5080
rect 7690 5049 7702 5052
rect 7644 5043 7702 5049
rect 7834 5040 7840 5052
rect 7892 5040 7898 5092
rect 9122 5080 9128 5092
rect 8588 5052 9128 5080
rect 2501 5015 2559 5021
rect 2501 4981 2513 5015
rect 2547 5012 2559 5015
rect 3510 5012 3516 5024
rect 2547 4984 3516 5012
rect 2547 4981 2559 4984
rect 2501 4975 2559 4981
rect 3510 4972 3516 4984
rect 3568 4972 3574 5024
rect 3694 5012 3700 5024
rect 3655 4984 3700 5012
rect 3694 4972 3700 4984
rect 3752 4972 3758 5024
rect 4157 5015 4215 5021
rect 4157 4981 4169 5015
rect 4203 5012 4215 5015
rect 5534 5012 5540 5024
rect 4203 4984 5540 5012
rect 4203 4981 4215 4984
rect 4157 4975 4215 4981
rect 5534 4972 5540 4984
rect 5592 4972 5598 5024
rect 5718 4972 5724 5024
rect 5776 5012 5782 5024
rect 7926 5012 7932 5024
rect 5776 4984 7932 5012
rect 5776 4972 5782 4984
rect 7926 4972 7932 4984
rect 7984 5012 7990 5024
rect 8588 5012 8616 5052
rect 9122 5040 9128 5052
rect 9180 5040 9186 5092
rect 9214 5040 9220 5092
rect 9272 5080 9278 5092
rect 10152 5080 10180 5120
rect 10778 5108 10784 5120
rect 10836 5108 10842 5160
rect 10873 5083 10931 5089
rect 10873 5080 10885 5083
rect 9272 5052 10088 5080
rect 10152 5052 10885 5080
rect 9272 5040 9278 5052
rect 8754 5012 8760 5024
rect 7984 4984 8616 5012
rect 8715 4984 8760 5012
rect 7984 4972 7990 4984
rect 8754 4972 8760 4984
rect 8812 4972 8818 5024
rect 9490 4972 9496 5024
rect 9548 5012 9554 5024
rect 9585 5015 9643 5021
rect 9585 5012 9597 5015
rect 9548 4984 9597 5012
rect 9548 4972 9554 4984
rect 9585 4981 9597 4984
rect 9631 4981 9643 5015
rect 9585 4975 9643 4981
rect 9677 5015 9735 5021
rect 9677 4981 9689 5015
rect 9723 5012 9735 5015
rect 9766 5012 9772 5024
rect 9723 4984 9772 5012
rect 9723 4981 9735 4984
rect 9677 4975 9735 4981
rect 9766 4972 9772 4984
rect 9824 4972 9830 5024
rect 10060 5012 10088 5052
rect 10873 5049 10885 5052
rect 10919 5080 10931 5083
rect 11164 5080 11192 5188
rect 11514 5108 11520 5160
rect 11572 5148 11578 5160
rect 11609 5151 11667 5157
rect 11609 5148 11621 5151
rect 11572 5120 11621 5148
rect 11572 5108 11578 5120
rect 11609 5117 11621 5120
rect 11655 5117 11667 5151
rect 11716 5148 11744 5188
rect 11790 5176 11796 5228
rect 11848 5216 11854 5228
rect 12342 5216 12348 5228
rect 11848 5188 12348 5216
rect 11848 5176 11854 5188
rect 12342 5176 12348 5188
rect 12400 5176 12406 5228
rect 12434 5176 12440 5228
rect 12492 5216 12498 5228
rect 12618 5216 12624 5228
rect 12492 5188 12624 5216
rect 12492 5176 12498 5188
rect 12618 5176 12624 5188
rect 12676 5176 12682 5228
rect 12710 5176 12716 5228
rect 12768 5216 12774 5228
rect 12897 5219 12955 5225
rect 12897 5216 12909 5219
rect 12768 5188 12909 5216
rect 12768 5176 12774 5188
rect 12897 5185 12909 5188
rect 12943 5185 12955 5219
rect 12897 5179 12955 5185
rect 12986 5176 12992 5228
rect 13044 5216 13050 5228
rect 13044 5188 13089 5216
rect 13044 5176 13050 5188
rect 13354 5176 13360 5228
rect 13412 5216 13418 5228
rect 14185 5219 14243 5225
rect 14185 5216 14197 5219
rect 13412 5188 14197 5216
rect 13412 5176 13418 5188
rect 14185 5185 14197 5188
rect 14231 5185 14243 5219
rect 14185 5179 14243 5185
rect 11882 5148 11888 5160
rect 11716 5120 11888 5148
rect 11609 5111 11667 5117
rect 11882 5108 11888 5120
rect 11940 5108 11946 5160
rect 12250 5108 12256 5160
rect 12308 5148 12314 5160
rect 12308 5120 13032 5148
rect 12308 5108 12314 5120
rect 12805 5083 12863 5089
rect 12805 5080 12817 5083
rect 10919 5052 11192 5080
rect 11256 5052 12817 5080
rect 10919 5049 10931 5052
rect 10873 5043 10931 5049
rect 11256 5012 11284 5052
rect 12805 5049 12817 5052
rect 12851 5049 12863 5083
rect 13004 5080 13032 5120
rect 13078 5108 13084 5160
rect 13136 5148 13142 5160
rect 13630 5148 13636 5160
rect 13136 5120 13636 5148
rect 13136 5108 13142 5120
rect 13630 5108 13636 5120
rect 13688 5148 13694 5160
rect 14844 5157 14872 5324
rect 14001 5151 14059 5157
rect 14001 5148 14013 5151
rect 13688 5120 14013 5148
rect 13688 5108 13694 5120
rect 14001 5117 14013 5120
rect 14047 5117 14059 5151
rect 14001 5111 14059 5117
rect 14829 5151 14887 5157
rect 14829 5117 14841 5151
rect 14875 5117 14887 5151
rect 14829 5111 14887 5117
rect 13538 5080 13544 5092
rect 13004 5052 13544 5080
rect 12805 5043 12863 5049
rect 13538 5040 13544 5052
rect 13596 5080 13602 5092
rect 13596 5052 14872 5080
rect 13596 5040 13602 5052
rect 14844 5024 14872 5052
rect 11790 5012 11796 5024
rect 10060 4984 11284 5012
rect 11751 4984 11796 5012
rect 11790 4972 11796 4984
rect 11848 4972 11854 5024
rect 12437 5015 12495 5021
rect 12437 4981 12449 5015
rect 12483 5012 12495 5015
rect 12986 5012 12992 5024
rect 12483 4984 12992 5012
rect 12483 4981 12495 4984
rect 12437 4975 12495 4981
rect 12986 4972 12992 4984
rect 13044 4972 13050 5024
rect 13722 4972 13728 5024
rect 13780 5012 13786 5024
rect 14093 5015 14151 5021
rect 14093 5012 14105 5015
rect 13780 4984 14105 5012
rect 13780 4972 13786 4984
rect 14093 4981 14105 4984
rect 14139 4981 14151 5015
rect 14093 4975 14151 4981
rect 14826 4972 14832 5024
rect 14884 4972 14890 5024
rect 15010 5012 15016 5024
rect 14971 4984 15016 5012
rect 15010 4972 15016 4984
rect 15068 4972 15074 5024
rect 1104 4922 15824 4944
rect 1104 4870 5912 4922
rect 5964 4870 5976 4922
rect 6028 4870 6040 4922
rect 6092 4870 6104 4922
rect 6156 4870 10843 4922
rect 10895 4870 10907 4922
rect 10959 4870 10971 4922
rect 11023 4870 11035 4922
rect 11087 4870 15824 4922
rect 1104 4848 15824 4870
rect 2777 4811 2835 4817
rect 2777 4777 2789 4811
rect 2823 4808 2835 4811
rect 3418 4808 3424 4820
rect 2823 4780 3424 4808
rect 2823 4777 2835 4780
rect 2777 4771 2835 4777
rect 3418 4768 3424 4780
rect 3476 4768 3482 4820
rect 3694 4768 3700 4820
rect 3752 4808 3758 4820
rect 4525 4811 4583 4817
rect 4525 4808 4537 4811
rect 3752 4780 4537 4808
rect 3752 4768 3758 4780
rect 4525 4777 4537 4780
rect 4571 4777 4583 4811
rect 4525 4771 4583 4777
rect 4982 4768 4988 4820
rect 5040 4808 5046 4820
rect 5261 4811 5319 4817
rect 5261 4808 5273 4811
rect 5040 4780 5273 4808
rect 5040 4768 5046 4780
rect 5261 4777 5273 4780
rect 5307 4777 5319 4811
rect 5261 4771 5319 4777
rect 5350 4768 5356 4820
rect 5408 4808 5414 4820
rect 7190 4808 7196 4820
rect 5408 4780 7196 4808
rect 5408 4768 5414 4780
rect 7190 4768 7196 4780
rect 7248 4768 7254 4820
rect 7466 4768 7472 4820
rect 7524 4808 7530 4820
rect 8297 4811 8355 4817
rect 8297 4808 8309 4811
rect 7524 4780 8309 4808
rect 7524 4768 7530 4780
rect 8297 4777 8309 4780
rect 8343 4777 8355 4811
rect 8297 4771 8355 4777
rect 8386 4768 8392 4820
rect 8444 4808 8450 4820
rect 8757 4811 8815 4817
rect 8757 4808 8769 4811
rect 8444 4780 8769 4808
rect 8444 4768 8450 4780
rect 8757 4777 8769 4780
rect 8803 4808 8815 4811
rect 9122 4808 9128 4820
rect 8803 4780 9128 4808
rect 8803 4777 8815 4780
rect 8757 4771 8815 4777
rect 9122 4768 9128 4780
rect 9180 4768 9186 4820
rect 9306 4768 9312 4820
rect 9364 4808 9370 4820
rect 9490 4808 9496 4820
rect 9364 4780 9496 4808
rect 9364 4768 9370 4780
rect 9490 4768 9496 4780
rect 9548 4768 9554 4820
rect 9677 4811 9735 4817
rect 9677 4777 9689 4811
rect 9723 4808 9735 4811
rect 9950 4808 9956 4820
rect 9723 4780 9956 4808
rect 9723 4777 9735 4780
rect 9677 4771 9735 4777
rect 9950 4768 9956 4780
rect 10008 4768 10014 4820
rect 10045 4811 10103 4817
rect 10045 4777 10057 4811
rect 10091 4808 10103 4811
rect 10410 4808 10416 4820
rect 10091 4780 10416 4808
rect 10091 4777 10103 4780
rect 10045 4771 10103 4777
rect 10410 4768 10416 4780
rect 10468 4768 10474 4820
rect 11330 4808 11336 4820
rect 10704 4780 11336 4808
rect 1664 4743 1722 4749
rect 1664 4709 1676 4743
rect 1710 4740 1722 4743
rect 3970 4740 3976 4752
rect 1710 4712 3976 4740
rect 1710 4709 1722 4712
rect 1664 4703 1722 4709
rect 3970 4700 3976 4712
rect 4028 4700 4034 4752
rect 4430 4740 4436 4752
rect 4391 4712 4436 4740
rect 4430 4700 4436 4712
rect 4488 4700 4494 4752
rect 6270 4740 6276 4752
rect 4724 4712 6276 4740
rect 2130 4632 2136 4684
rect 2188 4672 2194 4684
rect 3237 4675 3295 4681
rect 3237 4672 3249 4675
rect 2188 4644 3249 4672
rect 2188 4632 2194 4644
rect 3237 4641 3249 4644
rect 3283 4672 3295 4675
rect 4062 4672 4068 4684
rect 3283 4644 4068 4672
rect 3283 4641 3295 4644
rect 3237 4635 3295 4641
rect 4062 4632 4068 4644
rect 4120 4632 4126 4684
rect 3050 4564 3056 4616
rect 3108 4604 3114 4616
rect 3326 4604 3332 4616
rect 3108 4576 3332 4604
rect 3108 4564 3114 4576
rect 3326 4564 3332 4576
rect 3384 4564 3390 4616
rect 3510 4604 3516 4616
rect 3471 4576 3516 4604
rect 3510 4564 3516 4576
rect 3568 4564 3574 4616
rect 4724 4613 4752 4712
rect 6270 4700 6276 4712
rect 6328 4700 6334 4752
rect 6702 4743 6760 4749
rect 6702 4740 6714 4743
rect 6380 4712 6714 4740
rect 4798 4632 4804 4684
rect 4856 4672 4862 4684
rect 5258 4672 5264 4684
rect 4856 4644 5264 4672
rect 4856 4632 4862 4644
rect 5258 4632 5264 4644
rect 5316 4632 5322 4684
rect 5626 4672 5632 4684
rect 5587 4644 5632 4672
rect 5626 4632 5632 4644
rect 5684 4632 5690 4684
rect 6178 4632 6184 4684
rect 6236 4672 6242 4684
rect 6380 4672 6408 4712
rect 6702 4709 6714 4712
rect 6748 4709 6760 4743
rect 6702 4703 6760 4709
rect 7558 4700 7564 4752
rect 7616 4740 7622 4752
rect 7926 4740 7932 4752
rect 7616 4712 7932 4740
rect 7616 4700 7622 4712
rect 7926 4700 7932 4712
rect 7984 4740 7990 4752
rect 8570 4740 8576 4752
rect 7984 4712 8576 4740
rect 7984 4700 7990 4712
rect 8570 4700 8576 4712
rect 8628 4700 8634 4752
rect 10704 4740 10732 4780
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 13078 4808 13084 4820
rect 11808 4780 13084 4808
rect 11808 4740 11836 4780
rect 13078 4768 13084 4780
rect 13136 4768 13142 4820
rect 13262 4808 13268 4820
rect 13223 4780 13268 4808
rect 13262 4768 13268 4780
rect 13320 4768 13326 4820
rect 13538 4768 13544 4820
rect 13596 4808 13602 4820
rect 13725 4811 13783 4817
rect 13725 4808 13737 4811
rect 13596 4780 13737 4808
rect 13596 4768 13602 4780
rect 13725 4777 13737 4780
rect 13771 4777 13783 4811
rect 14642 4808 14648 4820
rect 14603 4780 14648 4808
rect 13725 4771 13783 4777
rect 14642 4768 14648 4780
rect 14700 4768 14706 4820
rect 12802 4740 12808 4752
rect 9968 4712 10732 4740
rect 11348 4712 11836 4740
rect 11900 4712 12808 4740
rect 6236 4644 6408 4672
rect 6457 4675 6515 4681
rect 6236 4632 6242 4644
rect 6457 4641 6469 4675
rect 6503 4672 6515 4675
rect 7006 4672 7012 4684
rect 6503 4644 7012 4672
rect 6503 4641 6515 4644
rect 6457 4635 6515 4641
rect 7006 4632 7012 4644
rect 7064 4632 7070 4684
rect 8665 4675 8723 4681
rect 8665 4641 8677 4675
rect 8711 4672 8723 4675
rect 9968 4672 9996 4712
rect 10134 4672 10140 4684
rect 8711 4644 9996 4672
rect 10095 4644 10140 4672
rect 8711 4641 8723 4644
rect 8665 4635 8723 4641
rect 10134 4632 10140 4644
rect 10192 4632 10198 4684
rect 10686 4672 10692 4684
rect 10244 4644 10692 4672
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4573 4767 4607
rect 5718 4604 5724 4616
rect 5679 4576 5724 4604
rect 4709 4567 4767 4573
rect 5718 4564 5724 4576
rect 5776 4564 5782 4616
rect 5810 4564 5816 4616
rect 5868 4604 5874 4616
rect 5868 4576 5913 4604
rect 5868 4564 5874 4576
rect 7466 4564 7472 4616
rect 7524 4604 7530 4616
rect 8110 4604 8116 4616
rect 7524 4576 8116 4604
rect 7524 4564 7530 4576
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 8570 4564 8576 4616
rect 8628 4604 8634 4616
rect 8849 4607 8907 4613
rect 8849 4604 8861 4607
rect 8628 4576 8861 4604
rect 8628 4564 8634 4576
rect 8849 4573 8861 4576
rect 8895 4573 8907 4607
rect 8849 4567 8907 4573
rect 10042 4564 10048 4616
rect 10100 4604 10106 4616
rect 10244 4613 10272 4644
rect 10686 4632 10692 4644
rect 10744 4632 10750 4684
rect 10778 4632 10784 4684
rect 10836 4672 10842 4684
rect 11348 4681 11376 4712
rect 11241 4675 11299 4681
rect 11241 4672 11253 4675
rect 10836 4644 11253 4672
rect 10836 4632 10842 4644
rect 11241 4641 11253 4644
rect 11287 4641 11299 4675
rect 11241 4635 11299 4641
rect 11333 4675 11391 4681
rect 11333 4641 11345 4675
rect 11379 4641 11391 4675
rect 11333 4635 11391 4641
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 10100 4576 10241 4604
rect 10100 4564 10106 4576
rect 10229 4573 10241 4576
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 10318 4564 10324 4616
rect 10376 4604 10382 4616
rect 10962 4604 10968 4616
rect 10376 4576 10968 4604
rect 10376 4564 10382 4576
rect 10962 4564 10968 4576
rect 11020 4604 11026 4616
rect 11517 4607 11575 4613
rect 11517 4604 11529 4607
rect 11020 4576 11529 4604
rect 11020 4564 11026 4576
rect 11517 4573 11529 4576
rect 11563 4604 11575 4607
rect 11900 4604 11928 4712
rect 12802 4700 12808 4712
rect 12860 4700 12866 4752
rect 13446 4700 13452 4752
rect 13504 4740 13510 4752
rect 13633 4743 13691 4749
rect 13633 4740 13645 4743
rect 13504 4712 13645 4740
rect 13504 4700 13510 4712
rect 13633 4709 13645 4712
rect 13679 4709 13691 4743
rect 13633 4703 13691 4709
rect 12437 4675 12495 4681
rect 12437 4672 12449 4675
rect 11563 4576 11928 4604
rect 11992 4644 12449 4672
rect 11563 4573 11575 4576
rect 11517 4567 11575 4573
rect 2869 4539 2927 4545
rect 2869 4505 2881 4539
rect 2915 4536 2927 4539
rect 2958 4536 2964 4548
rect 2915 4508 2964 4536
rect 2915 4505 2927 4508
rect 2869 4499 2927 4505
rect 2958 4496 2964 4508
rect 3016 4496 3022 4548
rect 3602 4496 3608 4548
rect 3660 4536 3666 4548
rect 5350 4536 5356 4548
rect 3660 4508 5356 4536
rect 3660 4496 3666 4508
rect 5350 4496 5356 4508
rect 5408 4496 5414 4548
rect 5442 4496 5448 4548
rect 5500 4536 5506 4548
rect 6270 4536 6276 4548
rect 5500 4508 6276 4536
rect 5500 4496 5506 4508
rect 6270 4496 6276 4508
rect 6328 4496 6334 4548
rect 8478 4496 8484 4548
rect 8536 4536 8542 4548
rect 11146 4536 11152 4548
rect 8536 4508 11152 4536
rect 8536 4496 8542 4508
rect 11146 4496 11152 4508
rect 11204 4496 11210 4548
rect 11992 4536 12020 4644
rect 12437 4641 12449 4644
rect 12483 4641 12495 4675
rect 14458 4672 14464 4684
rect 14419 4644 14464 4672
rect 12437 4635 12495 4641
rect 14458 4632 14464 4644
rect 14516 4632 14522 4684
rect 12250 4564 12256 4616
rect 12308 4604 12314 4616
rect 12529 4607 12587 4613
rect 12529 4604 12541 4607
rect 12308 4576 12541 4604
rect 12308 4564 12314 4576
rect 12529 4573 12541 4576
rect 12575 4573 12587 4607
rect 12710 4604 12716 4616
rect 12671 4576 12716 4604
rect 12529 4567 12587 4573
rect 12710 4564 12716 4576
rect 12768 4604 12774 4616
rect 13354 4604 13360 4616
rect 12768 4576 13360 4604
rect 12768 4564 12774 4576
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 13817 4607 13875 4613
rect 13817 4604 13829 4607
rect 13648 4576 13829 4604
rect 11256 4508 12020 4536
rect 4062 4468 4068 4480
rect 4023 4440 4068 4468
rect 4062 4428 4068 4440
rect 4120 4428 4126 4480
rect 4798 4428 4804 4480
rect 4856 4468 4862 4480
rect 6362 4468 6368 4480
rect 4856 4440 6368 4468
rect 4856 4428 4862 4440
rect 6362 4428 6368 4440
rect 6420 4428 6426 4480
rect 6822 4428 6828 4480
rect 6880 4468 6886 4480
rect 7466 4468 7472 4480
rect 6880 4440 7472 4468
rect 6880 4428 6886 4440
rect 7466 4428 7472 4440
rect 7524 4428 7530 4480
rect 7834 4468 7840 4480
rect 7747 4440 7840 4468
rect 7834 4428 7840 4440
rect 7892 4468 7898 4480
rect 8754 4468 8760 4480
rect 7892 4440 8760 4468
rect 7892 4428 7898 4440
rect 8754 4428 8760 4440
rect 8812 4468 8818 4480
rect 9306 4468 9312 4480
rect 8812 4440 9312 4468
rect 8812 4428 8818 4440
rect 9306 4428 9312 4440
rect 9364 4428 9370 4480
rect 9582 4428 9588 4480
rect 9640 4468 9646 4480
rect 10134 4468 10140 4480
rect 9640 4440 10140 4468
rect 9640 4428 9646 4440
rect 10134 4428 10140 4440
rect 10192 4428 10198 4480
rect 10594 4428 10600 4480
rect 10652 4468 10658 4480
rect 10873 4471 10931 4477
rect 10873 4468 10885 4471
rect 10652 4440 10885 4468
rect 10652 4428 10658 4440
rect 10873 4437 10885 4440
rect 10919 4437 10931 4471
rect 10873 4431 10931 4437
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 11256 4468 11284 4508
rect 11112 4440 11284 4468
rect 11112 4428 11118 4440
rect 11514 4428 11520 4480
rect 11572 4468 11578 4480
rect 12069 4471 12127 4477
rect 12069 4468 12081 4471
rect 11572 4440 12081 4468
rect 11572 4428 11578 4440
rect 12069 4437 12081 4440
rect 12115 4437 12127 4471
rect 12069 4431 12127 4437
rect 12710 4428 12716 4480
rect 12768 4468 12774 4480
rect 13648 4468 13676 4576
rect 13817 4573 13829 4576
rect 13863 4573 13875 4607
rect 13817 4567 13875 4573
rect 12768 4440 13676 4468
rect 12768 4428 12774 4440
rect 1104 4378 15824 4400
rect 1104 4326 3447 4378
rect 3499 4326 3511 4378
rect 3563 4326 3575 4378
rect 3627 4326 3639 4378
rect 3691 4326 8378 4378
rect 8430 4326 8442 4378
rect 8494 4326 8506 4378
rect 8558 4326 8570 4378
rect 8622 4326 13308 4378
rect 13360 4326 13372 4378
rect 13424 4326 13436 4378
rect 13488 4326 13500 4378
rect 13552 4326 15824 4378
rect 1104 4304 15824 4326
rect 5350 4264 5356 4276
rect 2608 4236 5356 4264
rect 2225 4131 2283 4137
rect 2225 4097 2237 4131
rect 2271 4128 2283 4131
rect 2608 4128 2636 4236
rect 5350 4224 5356 4236
rect 5408 4224 5414 4276
rect 5534 4264 5540 4276
rect 5495 4236 5540 4264
rect 5534 4224 5540 4236
rect 5592 4224 5598 4276
rect 5626 4224 5632 4276
rect 5684 4264 5690 4276
rect 6825 4267 6883 4273
rect 6825 4264 6837 4267
rect 5684 4236 6837 4264
rect 5684 4224 5690 4236
rect 6825 4233 6837 4236
rect 6871 4233 6883 4267
rect 6825 4227 6883 4233
rect 7466 4224 7472 4276
rect 7524 4264 7530 4276
rect 8021 4267 8079 4273
rect 8021 4264 8033 4267
rect 7524 4236 8033 4264
rect 7524 4224 7530 4236
rect 8021 4233 8033 4236
rect 8067 4233 8079 4267
rect 8021 4227 8079 4233
rect 8849 4267 8907 4273
rect 8849 4233 8861 4267
rect 8895 4264 8907 4267
rect 9030 4264 9036 4276
rect 8895 4236 9036 4264
rect 8895 4233 8907 4236
rect 8849 4227 8907 4233
rect 9030 4224 9036 4236
rect 9088 4224 9094 4276
rect 9306 4224 9312 4276
rect 9364 4264 9370 4276
rect 10318 4264 10324 4276
rect 9364 4236 10324 4264
rect 9364 4224 9370 4236
rect 10318 4224 10324 4236
rect 10376 4224 10382 4276
rect 10962 4224 10968 4276
rect 11020 4224 11026 4276
rect 11241 4267 11299 4273
rect 11241 4233 11253 4267
rect 11287 4264 11299 4267
rect 11422 4264 11428 4276
rect 11287 4236 11428 4264
rect 11287 4233 11299 4236
rect 11241 4227 11299 4233
rect 11422 4224 11428 4236
rect 11480 4224 11486 4276
rect 11514 4224 11520 4276
rect 11572 4264 11578 4276
rect 11882 4264 11888 4276
rect 11572 4236 11888 4264
rect 11572 4224 11578 4236
rect 11882 4224 11888 4236
rect 11940 4224 11946 4276
rect 12710 4224 12716 4276
rect 12768 4264 12774 4276
rect 12768 4236 13032 4264
rect 12768 4224 12774 4236
rect 3973 4199 4031 4205
rect 3973 4165 3985 4199
rect 4019 4165 4031 4199
rect 3973 4159 4031 4165
rect 2271 4100 2636 4128
rect 3988 4128 4016 4159
rect 4246 4156 4252 4208
rect 4304 4196 4310 4208
rect 6454 4196 6460 4208
rect 4304 4168 4660 4196
rect 4304 4156 4310 4168
rect 4522 4128 4528 4140
rect 3988 4100 4528 4128
rect 2271 4097 2283 4100
rect 2225 4091 2283 4097
rect 4522 4088 4528 4100
rect 4580 4088 4586 4140
rect 4632 4137 4660 4168
rect 6012 4168 6460 4196
rect 6012 4137 6040 4168
rect 6454 4156 6460 4168
rect 6512 4156 6518 4208
rect 6840 4168 8708 4196
rect 6840 4140 6868 4168
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4097 4675 4131
rect 4617 4091 4675 4097
rect 5997 4131 6055 4137
rect 5997 4097 6009 4131
rect 6043 4097 6055 4131
rect 5997 4091 6055 4097
rect 6089 4131 6147 4137
rect 6089 4097 6101 4131
rect 6135 4097 6147 4131
rect 6089 4091 6147 4097
rect 1302 4020 1308 4072
rect 1360 4060 1366 4072
rect 2593 4063 2651 4069
rect 2593 4060 2605 4063
rect 1360 4032 2605 4060
rect 1360 4020 1366 4032
rect 2593 4029 2605 4032
rect 2639 4029 2651 4063
rect 2593 4023 2651 4029
rect 3326 4020 3332 4072
rect 3384 4060 3390 4072
rect 4798 4060 4804 4072
rect 3384 4032 4804 4060
rect 3384 4020 3390 4032
rect 4798 4020 4804 4032
rect 4856 4020 4862 4072
rect 4893 4063 4951 4069
rect 4893 4029 4905 4063
rect 4939 4060 4951 4063
rect 5534 4060 5540 4072
rect 4939 4032 5540 4060
rect 4939 4029 4951 4032
rect 4893 4023 4951 4029
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 5902 4020 5908 4072
rect 5960 4060 5966 4072
rect 6104 4060 6132 4091
rect 6822 4088 6828 4140
rect 6880 4088 6886 4140
rect 7374 4128 7380 4140
rect 7335 4100 7380 4128
rect 7374 4088 7380 4100
rect 7432 4088 7438 4140
rect 7926 4088 7932 4140
rect 7984 4128 7990 4140
rect 8573 4131 8631 4137
rect 8573 4128 8585 4131
rect 7984 4100 8585 4128
rect 7984 4088 7990 4100
rect 8573 4097 8585 4100
rect 8619 4097 8631 4131
rect 8680 4128 8708 4168
rect 9674 4156 9680 4208
rect 9732 4196 9738 4208
rect 9858 4196 9864 4208
rect 9732 4168 9864 4196
rect 9732 4156 9738 4168
rect 9858 4156 9864 4168
rect 9916 4156 9922 4208
rect 10870 4196 10876 4208
rect 10704 4168 10876 4196
rect 9401 4131 9459 4137
rect 8680 4100 9352 4128
rect 8573 4091 8631 4097
rect 9324 4072 9352 4100
rect 9401 4097 9413 4131
rect 9447 4128 9459 4131
rect 10704 4128 10732 4168
rect 10870 4156 10876 4168
rect 10928 4156 10934 4208
rect 10980 4137 11008 4224
rect 12250 4196 12256 4208
rect 11532 4168 12256 4196
rect 9447 4100 10732 4128
rect 10965 4131 11023 4137
rect 9447 4097 9459 4100
rect 9401 4091 9459 4097
rect 10965 4097 10977 4131
rect 11011 4097 11023 4131
rect 11330 4128 11336 4140
rect 10965 4091 11023 4097
rect 11072 4100 11336 4128
rect 5960 4032 6132 4060
rect 5960 4020 5966 4032
rect 6362 4020 6368 4072
rect 6420 4060 6426 4072
rect 7190 4060 7196 4072
rect 6420 4032 7196 4060
rect 6420 4020 6426 4032
rect 7190 4020 7196 4032
rect 7248 4060 7254 4072
rect 7285 4063 7343 4069
rect 7285 4060 7297 4063
rect 7248 4032 7297 4060
rect 7248 4020 7254 4032
rect 7285 4029 7297 4032
rect 7331 4029 7343 4063
rect 7285 4023 7343 4029
rect 7834 4020 7840 4072
rect 7892 4060 7898 4072
rect 9030 4060 9036 4072
rect 7892 4032 9036 4060
rect 7892 4020 7898 4032
rect 9030 4020 9036 4032
rect 9088 4020 9094 4072
rect 9122 4020 9128 4072
rect 9180 4060 9186 4072
rect 9217 4063 9275 4069
rect 9217 4060 9229 4063
rect 9180 4032 9229 4060
rect 9180 4020 9186 4032
rect 9217 4029 9229 4032
rect 9263 4029 9275 4063
rect 9217 4023 9275 4029
rect 9306 4020 9312 4072
rect 9364 4060 9370 4072
rect 9364 4032 9409 4060
rect 9364 4020 9370 4032
rect 9490 4020 9496 4072
rect 9548 4060 9554 4072
rect 10229 4063 10287 4069
rect 10229 4060 10241 4063
rect 9548 4032 10241 4060
rect 9548 4020 9554 4032
rect 10229 4029 10241 4032
rect 10275 4029 10287 4063
rect 10229 4023 10287 4029
rect 10873 4063 10931 4069
rect 10873 4029 10885 4063
rect 10919 4060 10931 4063
rect 11072 4060 11100 4100
rect 11330 4088 11336 4100
rect 11388 4088 11394 4140
rect 11422 4060 11428 4072
rect 10919 4032 11100 4060
rect 11164 4032 11428 4060
rect 10919 4029 10931 4032
rect 10873 4023 10931 4029
rect 1949 3995 2007 4001
rect 1949 3961 1961 3995
rect 1995 3992 2007 3995
rect 2130 3992 2136 4004
rect 1995 3964 2136 3992
rect 1995 3961 2007 3964
rect 1949 3955 2007 3961
rect 2130 3952 2136 3964
rect 2188 3952 2194 4004
rect 2774 3952 2780 4004
rect 2832 4001 2838 4004
rect 2832 3995 2896 4001
rect 2832 3961 2850 3995
rect 2884 3961 2896 3995
rect 2832 3955 2896 3961
rect 2832 3952 2838 3955
rect 3050 3952 3056 4004
rect 3108 3992 3114 4004
rect 5169 3995 5227 4001
rect 5169 3992 5181 3995
rect 3108 3964 5181 3992
rect 3108 3952 3114 3964
rect 5169 3961 5181 3964
rect 5215 3961 5227 3995
rect 5169 3955 5227 3961
rect 5626 3952 5632 4004
rect 5684 3992 5690 4004
rect 6178 3992 6184 4004
rect 5684 3964 6184 3992
rect 5684 3952 5690 3964
rect 6178 3952 6184 3964
rect 6236 3952 6242 4004
rect 6270 3952 6276 4004
rect 6328 3992 6334 4004
rect 6454 3992 6460 4004
rect 6328 3964 6460 3992
rect 6328 3952 6334 3964
rect 6454 3952 6460 3964
rect 6512 3952 6518 4004
rect 6822 3992 6828 4004
rect 6748 3964 6828 3992
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 1670 3924 1676 3936
rect 1627 3896 1676 3924
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 1670 3884 1676 3896
rect 1728 3884 1734 3936
rect 2041 3927 2099 3933
rect 2041 3893 2053 3927
rect 2087 3924 2099 3927
rect 2958 3924 2964 3936
rect 2087 3896 2964 3924
rect 2087 3893 2099 3896
rect 2041 3887 2099 3893
rect 2958 3884 2964 3896
rect 3016 3884 3022 3936
rect 4065 3927 4123 3933
rect 4065 3893 4077 3927
rect 4111 3924 4123 3927
rect 4246 3924 4252 3936
rect 4111 3896 4252 3924
rect 4111 3893 4123 3896
rect 4065 3887 4123 3893
rect 4246 3884 4252 3896
rect 4304 3884 4310 3936
rect 4430 3924 4436 3936
rect 4391 3896 4436 3924
rect 4430 3884 4436 3896
rect 4488 3884 4494 3936
rect 4522 3884 4528 3936
rect 4580 3924 4586 3936
rect 4580 3896 4625 3924
rect 4580 3884 4586 3896
rect 4798 3884 4804 3936
rect 4856 3924 4862 3936
rect 5905 3927 5963 3933
rect 5905 3924 5917 3927
rect 4856 3896 5917 3924
rect 4856 3884 4862 3896
rect 5905 3893 5917 3896
rect 5951 3924 5963 3927
rect 6748 3924 6776 3964
rect 6822 3952 6828 3964
rect 6880 3952 6886 4004
rect 7006 3952 7012 4004
rect 7064 3992 7070 4004
rect 8110 3992 8116 4004
rect 7064 3964 8116 3992
rect 7064 3952 7070 3964
rect 8110 3952 8116 3964
rect 8168 3952 8174 4004
rect 8389 3995 8447 4001
rect 8389 3961 8401 3995
rect 8435 3992 8447 3995
rect 9858 3992 9864 4004
rect 8435 3964 9864 3992
rect 8435 3961 8447 3964
rect 8389 3955 8447 3961
rect 9858 3952 9864 3964
rect 9916 3952 9922 4004
rect 10781 3995 10839 4001
rect 10781 3961 10793 3995
rect 10827 3992 10839 3995
rect 11164 3992 11192 4032
rect 11422 4020 11428 4032
rect 11480 4020 11486 4072
rect 11532 3992 11560 4168
rect 12250 4156 12256 4168
rect 12308 4156 12314 4208
rect 11698 4088 11704 4140
rect 11756 4128 11762 4140
rect 13004 4137 13032 4236
rect 13078 4224 13084 4276
rect 13136 4224 13142 4276
rect 13096 4196 13124 4224
rect 13262 4196 13268 4208
rect 13096 4168 13268 4196
rect 13262 4156 13268 4168
rect 13320 4156 13326 4208
rect 11793 4131 11851 4137
rect 11793 4128 11805 4131
rect 11756 4100 11805 4128
rect 11756 4088 11762 4100
rect 11793 4097 11805 4100
rect 11839 4097 11851 4131
rect 11793 4091 11851 4097
rect 12989 4131 13047 4137
rect 12989 4097 13001 4131
rect 13035 4097 13047 4131
rect 12989 4091 13047 4097
rect 13078 4088 13084 4140
rect 13136 4128 13142 4140
rect 14185 4131 14243 4137
rect 14185 4128 14197 4131
rect 13136 4100 14197 4128
rect 13136 4088 13142 4100
rect 14185 4097 14197 4100
rect 14231 4097 14243 4131
rect 14185 4091 14243 4097
rect 11609 4063 11667 4069
rect 11609 4029 11621 4063
rect 11655 4060 11667 4063
rect 12066 4060 12072 4072
rect 11655 4032 12072 4060
rect 11655 4029 11667 4032
rect 11609 4023 11667 4029
rect 12066 4020 12072 4032
rect 12124 4020 12130 4072
rect 12526 4020 12532 4072
rect 12584 4060 12590 4072
rect 13354 4060 13360 4072
rect 12584 4032 13360 4060
rect 12584 4020 12590 4032
rect 13354 4020 13360 4032
rect 13412 4060 13418 4072
rect 14829 4063 14887 4069
rect 14829 4060 14841 4063
rect 13412 4032 14841 4060
rect 13412 4020 13418 4032
rect 14829 4029 14841 4032
rect 14875 4029 14887 4063
rect 14829 4023 14887 4029
rect 10827 3964 11192 3992
rect 11256 3964 11560 3992
rect 11701 3995 11759 4001
rect 10827 3961 10839 3964
rect 10781 3955 10839 3961
rect 5951 3896 6776 3924
rect 7193 3927 7251 3933
rect 5951 3893 5963 3896
rect 5905 3887 5963 3893
rect 7193 3893 7205 3927
rect 7239 3924 7251 3927
rect 7282 3924 7288 3936
rect 7239 3896 7288 3924
rect 7239 3893 7251 3896
rect 7193 3887 7251 3893
rect 7282 3884 7288 3896
rect 7340 3884 7346 3936
rect 8481 3927 8539 3933
rect 8481 3893 8493 3927
rect 8527 3924 8539 3927
rect 9030 3924 9036 3936
rect 8527 3896 9036 3924
rect 8527 3893 8539 3896
rect 8481 3887 8539 3893
rect 9030 3884 9036 3896
rect 9088 3884 9094 3936
rect 10045 3927 10103 3933
rect 10045 3893 10057 3927
rect 10091 3924 10103 3927
rect 10226 3924 10232 3936
rect 10091 3896 10232 3924
rect 10091 3893 10103 3896
rect 10045 3887 10103 3893
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 10410 3924 10416 3936
rect 10371 3896 10416 3924
rect 10410 3884 10416 3896
rect 10468 3884 10474 3936
rect 10686 3884 10692 3936
rect 10744 3924 10750 3936
rect 11256 3924 11284 3964
rect 11701 3961 11713 3995
rect 11747 3992 11759 3995
rect 11882 3992 11888 4004
rect 11747 3964 11888 3992
rect 11747 3961 11759 3964
rect 11701 3955 11759 3961
rect 11882 3952 11888 3964
rect 11940 3952 11946 4004
rect 12802 3992 12808 4004
rect 12763 3964 12808 3992
rect 12802 3952 12808 3964
rect 12860 3952 12866 4004
rect 13998 3992 14004 4004
rect 13464 3964 13768 3992
rect 13959 3964 14004 3992
rect 10744 3896 11284 3924
rect 10744 3884 10750 3896
rect 11330 3884 11336 3936
rect 11388 3924 11394 3936
rect 11790 3924 11796 3936
rect 11388 3896 11796 3924
rect 11388 3884 11394 3896
rect 11790 3884 11796 3896
rect 11848 3884 11854 3936
rect 12250 3884 12256 3936
rect 12308 3924 12314 3936
rect 12437 3927 12495 3933
rect 12437 3924 12449 3927
rect 12308 3896 12449 3924
rect 12308 3884 12314 3896
rect 12437 3893 12449 3896
rect 12483 3893 12495 3927
rect 12437 3887 12495 3893
rect 12897 3927 12955 3933
rect 12897 3893 12909 3927
rect 12943 3924 12955 3927
rect 13464 3924 13492 3964
rect 13630 3924 13636 3936
rect 12943 3896 13492 3924
rect 13591 3896 13636 3924
rect 12943 3893 12955 3896
rect 12897 3887 12955 3893
rect 13630 3884 13636 3896
rect 13688 3884 13694 3936
rect 13740 3924 13768 3964
rect 13998 3952 14004 3964
rect 14056 3952 14062 4004
rect 14093 3995 14151 4001
rect 14093 3961 14105 3995
rect 14139 3992 14151 3995
rect 15102 3992 15108 4004
rect 14139 3964 15108 3992
rect 14139 3961 14151 3964
rect 14093 3955 14151 3961
rect 15102 3952 15108 3964
rect 15160 3952 15166 4004
rect 14274 3924 14280 3936
rect 13740 3896 14280 3924
rect 14274 3884 14280 3896
rect 14332 3884 14338 3936
rect 15010 3884 15016 3936
rect 15068 3924 15074 3936
rect 15068 3896 15113 3924
rect 15068 3884 15074 3896
rect 1104 3834 15824 3856
rect 1104 3782 5912 3834
rect 5964 3782 5976 3834
rect 6028 3782 6040 3834
rect 6092 3782 6104 3834
rect 6156 3782 10843 3834
rect 10895 3782 10907 3834
rect 10959 3782 10971 3834
rect 11023 3782 11035 3834
rect 11087 3782 15824 3834
rect 1104 3760 15824 3782
rect 2777 3723 2835 3729
rect 2777 3689 2789 3723
rect 2823 3689 2835 3723
rect 2777 3683 2835 3689
rect 1664 3655 1722 3661
rect 1664 3621 1676 3655
rect 1710 3652 1722 3655
rect 2406 3652 2412 3664
rect 1710 3624 2412 3652
rect 1710 3621 1722 3624
rect 1664 3615 1722 3621
rect 2406 3612 2412 3624
rect 2464 3612 2470 3664
rect 2792 3652 2820 3683
rect 2866 3680 2872 3732
rect 2924 3720 2930 3732
rect 2924 3692 2969 3720
rect 2924 3680 2930 3692
rect 3234 3680 3240 3732
rect 3292 3720 3298 3732
rect 3329 3723 3387 3729
rect 3329 3720 3341 3723
rect 3292 3692 3341 3720
rect 3292 3680 3298 3692
rect 3329 3689 3341 3692
rect 3375 3689 3387 3723
rect 3329 3683 3387 3689
rect 4065 3723 4123 3729
rect 4065 3689 4077 3723
rect 4111 3720 4123 3723
rect 4522 3720 4528 3732
rect 4111 3692 4528 3720
rect 4111 3689 4123 3692
rect 4065 3683 4123 3689
rect 4522 3680 4528 3692
rect 4580 3680 4586 3732
rect 4893 3723 4951 3729
rect 4893 3689 4905 3723
rect 4939 3720 4951 3723
rect 5813 3723 5871 3729
rect 4939 3692 5771 3720
rect 4939 3689 4951 3692
rect 4893 3683 4951 3689
rect 3970 3652 3976 3664
rect 2792 3624 3976 3652
rect 3970 3612 3976 3624
rect 4028 3612 4034 3664
rect 4154 3612 4160 3664
rect 4212 3652 4218 3664
rect 4433 3655 4491 3661
rect 4433 3652 4445 3655
rect 4212 3624 4445 3652
rect 4212 3612 4218 3624
rect 4433 3621 4445 3624
rect 4479 3621 4491 3655
rect 4433 3615 4491 3621
rect 566 3544 572 3596
rect 624 3584 630 3596
rect 1486 3584 1492 3596
rect 624 3556 1492 3584
rect 624 3544 630 3556
rect 1486 3544 1492 3556
rect 1544 3544 1550 3596
rect 2130 3544 2136 3596
rect 2188 3584 2194 3596
rect 3234 3584 3240 3596
rect 2188 3556 2636 3584
rect 3195 3556 3240 3584
rect 2188 3544 2194 3556
rect 1302 3476 1308 3528
rect 1360 3516 1366 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 1360 3488 1409 3516
rect 1360 3476 1366 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 2608 3516 2636 3556
rect 3234 3544 3240 3556
rect 3292 3544 3298 3596
rect 3602 3584 3608 3596
rect 3528 3556 3608 3584
rect 3528 3525 3556 3556
rect 3602 3544 3608 3556
rect 3660 3544 3666 3596
rect 5350 3584 5356 3596
rect 5311 3556 5356 3584
rect 5350 3544 5356 3556
rect 5408 3544 5414 3596
rect 5743 3584 5771 3692
rect 5813 3689 5825 3723
rect 5859 3720 5871 3723
rect 7101 3723 7159 3729
rect 7101 3720 7113 3723
rect 5859 3692 7113 3720
rect 5859 3689 5871 3692
rect 5813 3683 5871 3689
rect 7101 3689 7113 3692
rect 7147 3689 7159 3723
rect 7101 3683 7159 3689
rect 7469 3723 7527 3729
rect 7469 3689 7481 3723
rect 7515 3720 7527 3723
rect 7742 3720 7748 3732
rect 7515 3692 7748 3720
rect 7515 3689 7527 3692
rect 7469 3683 7527 3689
rect 7742 3680 7748 3692
rect 7800 3680 7806 3732
rect 8294 3720 8300 3732
rect 8255 3692 8300 3720
rect 8294 3680 8300 3692
rect 8352 3680 8358 3732
rect 8478 3680 8484 3732
rect 8536 3720 8542 3732
rect 8757 3723 8815 3729
rect 8757 3720 8769 3723
rect 8536 3692 8769 3720
rect 8536 3680 8542 3692
rect 8757 3689 8769 3692
rect 8803 3689 8815 3723
rect 8757 3683 8815 3689
rect 9677 3723 9735 3729
rect 9677 3689 9689 3723
rect 9723 3720 9735 3723
rect 10686 3720 10692 3732
rect 9723 3692 10692 3720
rect 9723 3689 9735 3692
rect 9677 3683 9735 3689
rect 10686 3680 10692 3692
rect 10744 3680 10750 3732
rect 11790 3680 11796 3732
rect 11848 3680 11854 3732
rect 12066 3680 12072 3732
rect 12124 3720 12130 3732
rect 12618 3720 12624 3732
rect 12124 3692 12624 3720
rect 12124 3680 12130 3692
rect 12618 3680 12624 3692
rect 12676 3680 12682 3732
rect 13262 3720 13268 3732
rect 13223 3692 13268 3720
rect 13262 3680 13268 3692
rect 13320 3680 13326 3732
rect 13633 3723 13691 3729
rect 13633 3689 13645 3723
rect 13679 3720 13691 3723
rect 13906 3720 13912 3732
rect 13679 3692 13912 3720
rect 13679 3689 13691 3692
rect 13633 3683 13691 3689
rect 13906 3680 13912 3692
rect 13964 3680 13970 3732
rect 14642 3720 14648 3732
rect 14603 3692 14648 3720
rect 14642 3680 14648 3692
rect 14700 3680 14706 3732
rect 6178 3612 6184 3664
rect 6236 3652 6242 3664
rect 7009 3655 7067 3661
rect 6236 3624 6281 3652
rect 6236 3612 6242 3624
rect 7009 3621 7021 3655
rect 7055 3652 7067 3655
rect 7929 3655 7987 3661
rect 7929 3652 7941 3655
rect 7055 3624 7941 3652
rect 7055 3621 7067 3624
rect 7009 3615 7067 3621
rect 7929 3621 7941 3624
rect 7975 3652 7987 3655
rect 8386 3652 8392 3664
rect 7975 3624 8392 3652
rect 7975 3621 7987 3624
rect 7929 3615 7987 3621
rect 8386 3612 8392 3624
rect 8444 3652 8450 3664
rect 8444 3624 9076 3652
rect 8444 3612 8450 3624
rect 6270 3584 6276 3596
rect 5743 3556 6276 3584
rect 6270 3544 6276 3556
rect 6328 3544 6334 3596
rect 7190 3544 7196 3596
rect 7248 3584 7254 3596
rect 7834 3584 7840 3596
rect 7248 3556 7840 3584
rect 7248 3544 7254 3556
rect 7834 3544 7840 3556
rect 7892 3544 7898 3596
rect 8570 3584 8576 3596
rect 8128 3556 8576 3584
rect 3513 3519 3571 3525
rect 2608 3488 3464 3516
rect 1397 3479 1455 3485
rect 3436 3448 3464 3488
rect 3513 3485 3525 3519
rect 3559 3485 3571 3519
rect 4522 3516 4528 3528
rect 4483 3488 4528 3516
rect 3513 3479 3571 3485
rect 4522 3476 4528 3488
rect 4580 3476 4586 3528
rect 4709 3519 4767 3525
rect 4709 3485 4721 3519
rect 4755 3516 4767 3519
rect 4982 3516 4988 3528
rect 4755 3488 4988 3516
rect 4755 3485 4767 3488
rect 4709 3479 4767 3485
rect 4982 3476 4988 3488
rect 5040 3476 5046 3528
rect 5442 3516 5448 3528
rect 5403 3488 5448 3516
rect 5442 3476 5448 3488
rect 5500 3476 5506 3528
rect 5629 3519 5687 3525
rect 5629 3485 5641 3519
rect 5675 3485 5687 3519
rect 5629 3479 5687 3485
rect 4798 3448 4804 3460
rect 3436 3420 4804 3448
rect 4798 3408 4804 3420
rect 4856 3408 4862 3460
rect 5644 3392 5672 3479
rect 5810 3476 5816 3528
rect 5868 3516 5874 3528
rect 6178 3516 6184 3528
rect 5868 3488 6184 3516
rect 5868 3476 5874 3488
rect 6178 3476 6184 3488
rect 6236 3476 6242 3528
rect 6457 3519 6515 3525
rect 6457 3485 6469 3519
rect 6503 3516 6515 3519
rect 6914 3516 6920 3528
rect 6503 3488 6920 3516
rect 6503 3485 6515 3488
rect 6457 3479 6515 3485
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 7285 3519 7343 3525
rect 7285 3485 7297 3519
rect 7331 3516 7343 3519
rect 7374 3516 7380 3528
rect 7331 3488 7380 3516
rect 7331 3485 7343 3488
rect 7285 3479 7343 3485
rect 7374 3476 7380 3488
rect 7432 3476 7438 3528
rect 8128 3525 8156 3556
rect 8570 3544 8576 3556
rect 8628 3544 8634 3596
rect 8665 3587 8723 3593
rect 8665 3553 8677 3587
rect 8711 3584 8723 3587
rect 8711 3556 8975 3584
rect 8711 3553 8723 3556
rect 8665 3547 8723 3553
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3485 8171 3519
rect 8113 3479 8171 3485
rect 8202 3476 8208 3528
rect 8260 3516 8266 3528
rect 8849 3519 8907 3525
rect 8849 3516 8861 3519
rect 8260 3488 8861 3516
rect 8260 3476 8266 3488
rect 8849 3485 8861 3488
rect 8895 3485 8907 3519
rect 8849 3479 8907 3485
rect 5718 3408 5724 3460
rect 5776 3448 5782 3460
rect 6641 3451 6699 3457
rect 6641 3448 6653 3451
rect 5776 3420 6653 3448
rect 5776 3408 5782 3420
rect 6641 3417 6653 3420
rect 6687 3417 6699 3451
rect 6641 3411 6699 3417
rect 8662 3408 8668 3460
rect 8720 3448 8726 3460
rect 8947 3448 8975 3556
rect 9048 3516 9076 3624
rect 9306 3612 9312 3664
rect 9364 3652 9370 3664
rect 10137 3655 10195 3661
rect 10137 3652 10149 3655
rect 9364 3624 9720 3652
rect 9364 3612 9370 3624
rect 9692 3596 9720 3624
rect 9876 3624 10149 3652
rect 9674 3544 9680 3596
rect 9732 3544 9738 3596
rect 9876 3528 9904 3624
rect 10137 3621 10149 3624
rect 10183 3621 10195 3655
rect 10137 3615 10195 3621
rect 11514 3612 11520 3664
rect 11572 3652 11578 3664
rect 11808 3652 11836 3680
rect 12437 3655 12495 3661
rect 11572 3624 11744 3652
rect 11808 3624 12204 3652
rect 11572 3612 11578 3624
rect 10045 3587 10103 3593
rect 10045 3553 10057 3587
rect 10091 3584 10103 3587
rect 10226 3584 10232 3596
rect 10091 3556 10232 3584
rect 10091 3553 10103 3556
rect 10045 3547 10103 3553
rect 10226 3544 10232 3556
rect 10284 3544 10290 3596
rect 10502 3544 10508 3596
rect 10560 3584 10566 3596
rect 10962 3584 10968 3596
rect 10560 3556 10968 3584
rect 10560 3544 10566 3556
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 11238 3584 11244 3596
rect 11199 3556 11244 3584
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 11716 3593 11744 3624
rect 11333 3587 11391 3593
rect 11333 3553 11345 3587
rect 11379 3584 11391 3587
rect 11701 3587 11759 3593
rect 11379 3556 11560 3584
rect 11379 3553 11391 3556
rect 11333 3547 11391 3553
rect 9122 3516 9128 3528
rect 9048 3488 9128 3516
rect 9122 3476 9128 3488
rect 9180 3476 9186 3528
rect 9582 3476 9588 3528
rect 9640 3516 9646 3528
rect 9858 3516 9864 3528
rect 9640 3488 9864 3516
rect 9640 3476 9646 3488
rect 9858 3476 9864 3488
rect 9916 3476 9922 3528
rect 10134 3476 10140 3528
rect 10192 3516 10198 3528
rect 10321 3519 10379 3525
rect 10321 3516 10333 3519
rect 10192 3488 10333 3516
rect 10192 3476 10198 3488
rect 10321 3485 10333 3488
rect 10367 3516 10379 3519
rect 11425 3519 11483 3525
rect 11425 3516 11437 3519
rect 10367 3488 11437 3516
rect 10367 3485 10379 3488
rect 10321 3479 10379 3485
rect 11425 3485 11437 3488
rect 11471 3485 11483 3519
rect 11532 3516 11560 3556
rect 11701 3553 11713 3587
rect 11747 3553 11759 3587
rect 12176 3584 12204 3624
rect 12437 3621 12449 3655
rect 12483 3652 12495 3655
rect 15194 3652 15200 3664
rect 12483 3624 15200 3652
rect 12483 3621 12495 3624
rect 12437 3615 12495 3621
rect 15194 3612 15200 3624
rect 15252 3652 15258 3664
rect 15930 3652 15936 3664
rect 15252 3624 15936 3652
rect 15252 3612 15258 3624
rect 15930 3612 15936 3624
rect 15988 3612 15994 3664
rect 12529 3587 12587 3593
rect 12529 3584 12541 3587
rect 12176 3556 12541 3584
rect 11701 3547 11759 3553
rect 12529 3553 12541 3556
rect 12575 3584 12587 3587
rect 13170 3584 13176 3596
rect 12575 3556 13176 3584
rect 12575 3553 12587 3556
rect 12529 3547 12587 3553
rect 13170 3544 13176 3556
rect 13228 3544 13234 3596
rect 13262 3544 13268 3596
rect 13320 3584 13326 3596
rect 13725 3587 13783 3593
rect 13725 3584 13737 3587
rect 13320 3556 13737 3584
rect 13320 3544 13326 3556
rect 13725 3553 13737 3556
rect 13771 3553 13783 3587
rect 14458 3584 14464 3596
rect 14419 3556 14464 3584
rect 13725 3547 13783 3553
rect 14458 3544 14464 3556
rect 14516 3544 14522 3596
rect 11606 3516 11612 3528
rect 11519 3488 11612 3516
rect 11425 3479 11483 3485
rect 11606 3476 11612 3488
rect 11664 3516 11670 3528
rect 12066 3516 12072 3528
rect 11664 3488 12072 3516
rect 11664 3476 11670 3488
rect 12066 3476 12072 3488
rect 12124 3476 12130 3528
rect 12618 3516 12624 3528
rect 12579 3488 12624 3516
rect 12618 3476 12624 3488
rect 12676 3476 12682 3528
rect 13817 3519 13875 3525
rect 13817 3485 13829 3519
rect 13863 3485 13875 3519
rect 13817 3479 13875 3485
rect 8720 3420 8975 3448
rect 8720 3408 8726 3420
rect 9030 3408 9036 3460
rect 9088 3448 9094 3460
rect 10686 3448 10692 3460
rect 9088 3420 10692 3448
rect 9088 3408 9094 3420
rect 10686 3408 10692 3420
rect 10744 3408 10750 3460
rect 10870 3448 10876 3460
rect 10831 3420 10876 3448
rect 10870 3408 10876 3420
rect 10928 3408 10934 3460
rect 13832 3448 13860 3479
rect 11072 3420 12572 3448
rect 2314 3340 2320 3392
rect 2372 3380 2378 3392
rect 4893 3383 4951 3389
rect 4893 3380 4905 3383
rect 2372 3352 4905 3380
rect 2372 3340 2378 3352
rect 4893 3349 4905 3352
rect 4939 3349 4951 3383
rect 4893 3343 4951 3349
rect 4982 3340 4988 3392
rect 5040 3380 5046 3392
rect 5626 3380 5632 3392
rect 5040 3352 5085 3380
rect 5539 3352 5632 3380
rect 5040 3340 5046 3352
rect 5626 3340 5632 3352
rect 5684 3380 5690 3392
rect 11072 3380 11100 3420
rect 5684 3352 11100 3380
rect 5684 3340 5690 3352
rect 11238 3340 11244 3392
rect 11296 3380 11302 3392
rect 11698 3380 11704 3392
rect 11296 3352 11704 3380
rect 11296 3340 11302 3352
rect 11698 3340 11704 3352
rect 11756 3340 11762 3392
rect 11882 3380 11888 3392
rect 11843 3352 11888 3380
rect 11882 3340 11888 3352
rect 11940 3340 11946 3392
rect 11974 3340 11980 3392
rect 12032 3380 12038 3392
rect 12069 3383 12127 3389
rect 12069 3380 12081 3383
rect 12032 3352 12081 3380
rect 12032 3340 12038 3352
rect 12069 3349 12081 3352
rect 12115 3349 12127 3383
rect 12544 3380 12572 3420
rect 12728 3420 13860 3448
rect 12728 3380 12756 3420
rect 12544 3352 12756 3380
rect 12069 3343 12127 3349
rect 13814 3340 13820 3392
rect 13872 3380 13878 3392
rect 14550 3380 14556 3392
rect 13872 3352 14556 3380
rect 13872 3340 13878 3352
rect 14550 3340 14556 3352
rect 14608 3340 14614 3392
rect 1104 3290 15824 3312
rect 1104 3238 3447 3290
rect 3499 3238 3511 3290
rect 3563 3238 3575 3290
rect 3627 3238 3639 3290
rect 3691 3238 8378 3290
rect 8430 3238 8442 3290
rect 8494 3238 8506 3290
rect 8558 3238 8570 3290
rect 8622 3238 13308 3290
rect 13360 3238 13372 3290
rect 13424 3238 13436 3290
rect 13488 3238 13500 3290
rect 13552 3238 15824 3290
rect 1104 3216 15824 3238
rect 1026 3136 1032 3188
rect 1084 3176 1090 3188
rect 1578 3176 1584 3188
rect 1084 3148 1584 3176
rect 1084 3136 1090 3148
rect 1578 3136 1584 3148
rect 1636 3136 1642 3188
rect 4249 3179 4307 3185
rect 4249 3145 4261 3179
rect 4295 3176 4307 3179
rect 4338 3176 4344 3188
rect 4295 3148 4344 3176
rect 4295 3145 4307 3148
rect 4249 3139 4307 3145
rect 4338 3136 4344 3148
rect 4396 3136 4402 3188
rect 4522 3136 4528 3188
rect 4580 3176 4586 3188
rect 6825 3179 6883 3185
rect 6825 3176 6837 3179
rect 4580 3148 6837 3176
rect 4580 3136 4586 3148
rect 6825 3145 6837 3148
rect 6871 3145 6883 3179
rect 7374 3176 7380 3188
rect 6825 3139 6883 3145
rect 7024 3148 7380 3176
rect 2777 3111 2835 3117
rect 2777 3077 2789 3111
rect 2823 3108 2835 3111
rect 2866 3108 2872 3120
rect 2823 3080 2872 3108
rect 2823 3077 2835 3080
rect 2777 3071 2835 3077
rect 2866 3068 2872 3080
rect 2924 3068 2930 3120
rect 5442 3068 5448 3120
rect 5500 3108 5506 3120
rect 6362 3108 6368 3120
rect 5500 3080 6368 3108
rect 5500 3068 5506 3080
rect 6362 3068 6368 3080
rect 6420 3068 6426 3120
rect 1302 3000 1308 3052
rect 1360 3040 1366 3052
rect 1397 3043 1455 3049
rect 1397 3040 1409 3043
rect 1360 3012 1409 3040
rect 1360 3000 1366 3012
rect 1397 3009 1409 3012
rect 1443 3009 1455 3043
rect 1397 3003 1455 3009
rect 4246 3000 4252 3052
rect 4304 3000 4310 3052
rect 4614 3000 4620 3052
rect 4672 3040 4678 3052
rect 4985 3043 5043 3049
rect 4985 3040 4997 3043
rect 4672 3012 4997 3040
rect 4672 3000 4678 3012
rect 4985 3009 4997 3012
rect 5031 3040 5043 3043
rect 5626 3040 5632 3052
rect 5031 3012 5632 3040
rect 5031 3009 5043 3012
rect 4985 3003 5043 3009
rect 5626 3000 5632 3012
rect 5684 3000 5690 3052
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 5859 3012 6132 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 3136 2975 3194 2981
rect 3136 2941 3148 2975
rect 3182 2972 3194 2975
rect 3694 2972 3700 2984
rect 3182 2944 3700 2972
rect 3182 2941 3194 2944
rect 3136 2935 3194 2941
rect 3694 2932 3700 2944
rect 3752 2932 3758 2984
rect 4264 2972 4292 3000
rect 5986 2975 6044 2981
rect 5986 2972 5998 2975
rect 4264 2944 5998 2972
rect 5986 2941 5998 2944
rect 6032 2941 6044 2975
rect 6104 2972 6132 3012
rect 6178 3000 6184 3052
rect 6236 3040 6242 3052
rect 6236 3012 6281 3040
rect 6236 3000 6242 3012
rect 6454 2972 6460 2984
rect 6104 2944 6460 2972
rect 5986 2935 6044 2941
rect 6454 2932 6460 2944
rect 6512 2932 6518 2984
rect 1664 2907 1722 2913
rect 1664 2873 1676 2907
rect 1710 2904 1722 2907
rect 1762 2904 1768 2916
rect 1710 2876 1768 2904
rect 1710 2873 1722 2876
rect 1664 2867 1722 2873
rect 1762 2864 1768 2876
rect 1820 2864 1826 2916
rect 2498 2864 2504 2916
rect 2556 2904 2562 2916
rect 4706 2904 4712 2916
rect 2556 2876 4712 2904
rect 2556 2864 2562 2876
rect 4706 2864 4712 2876
rect 4764 2864 4770 2916
rect 6086 2864 6092 2916
rect 6144 2904 6150 2916
rect 7024 2904 7052 3148
rect 7374 3136 7380 3148
rect 7432 3136 7438 3188
rect 7653 3179 7711 3185
rect 7653 3145 7665 3179
rect 7699 3176 7711 3179
rect 8662 3176 8668 3188
rect 7699 3148 8668 3176
rect 7699 3145 7711 3148
rect 7653 3139 7711 3145
rect 8662 3136 8668 3148
rect 8720 3136 8726 3188
rect 9214 3176 9220 3188
rect 9175 3148 9220 3176
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 11241 3179 11299 3185
rect 11241 3145 11253 3179
rect 11287 3176 11299 3179
rect 12434 3176 12440 3188
rect 11287 3148 12440 3176
rect 11287 3145 11299 3148
rect 11241 3139 11299 3145
rect 12434 3136 12440 3148
rect 12492 3136 12498 3188
rect 12526 3136 12532 3188
rect 12584 3176 12590 3188
rect 15289 3179 15347 3185
rect 15289 3176 15301 3179
rect 12584 3148 15301 3176
rect 12584 3136 12590 3148
rect 15289 3145 15301 3148
rect 15335 3145 15347 3179
rect 15289 3139 15347 3145
rect 10502 3068 10508 3120
rect 10560 3108 10566 3120
rect 11606 3108 11612 3120
rect 10560 3080 11612 3108
rect 10560 3068 10566 3080
rect 11606 3068 11612 3080
rect 11664 3068 11670 3120
rect 13262 3068 13268 3120
rect 13320 3108 13326 3120
rect 13906 3108 13912 3120
rect 13320 3080 13912 3108
rect 13320 3068 13326 3080
rect 13906 3068 13912 3080
rect 13964 3068 13970 3120
rect 13998 3068 14004 3120
rect 14056 3108 14062 3120
rect 14918 3108 14924 3120
rect 14056 3080 14924 3108
rect 14056 3068 14062 3080
rect 14918 3068 14924 3080
rect 14976 3068 14982 3120
rect 7190 3000 7196 3052
rect 7248 3000 7254 3052
rect 7374 3040 7380 3052
rect 7335 3012 7380 3040
rect 7374 3000 7380 3012
rect 7432 3000 7438 3052
rect 7466 3000 7472 3052
rect 7524 3040 7530 3052
rect 8205 3043 8263 3049
rect 8205 3040 8217 3043
rect 7524 3012 8217 3040
rect 7524 3000 7530 3012
rect 8205 3009 8217 3012
rect 8251 3009 8263 3043
rect 8205 3003 8263 3009
rect 8846 3000 8852 3052
rect 8904 3040 8910 3052
rect 9769 3043 9827 3049
rect 9769 3040 9781 3043
rect 8904 3012 9781 3040
rect 8904 3000 8910 3012
rect 9769 3009 9781 3012
rect 9815 3009 9827 3043
rect 9769 3003 9827 3009
rect 10318 3000 10324 3052
rect 10376 3040 10382 3052
rect 10965 3043 11023 3049
rect 10965 3040 10977 3043
rect 10376 3012 10977 3040
rect 10376 3000 10382 3012
rect 10965 3009 10977 3012
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 11146 3000 11152 3052
rect 11204 3040 11210 3052
rect 11793 3043 11851 3049
rect 11793 3040 11805 3043
rect 11204 3012 11805 3040
rect 11204 3000 11210 3012
rect 11793 3009 11805 3012
rect 11839 3009 11851 3043
rect 12897 3043 12955 3049
rect 12897 3040 12909 3043
rect 11793 3003 11851 3009
rect 12360 3012 12909 3040
rect 7208 2972 7236 3000
rect 12360 2984 12388 3012
rect 12897 3009 12909 3012
rect 12943 3009 12955 3043
rect 13078 3040 13084 3052
rect 13039 3012 13084 3040
rect 12897 3003 12955 3009
rect 13078 3000 13084 3012
rect 13136 3000 13142 3052
rect 13817 3043 13875 3049
rect 13817 3009 13829 3043
rect 13863 3040 13875 3043
rect 14734 3040 14740 3052
rect 13863 3012 14740 3040
rect 13863 3009 13875 3012
rect 13817 3003 13875 3009
rect 14734 3000 14740 3012
rect 14792 3000 14798 3052
rect 8478 2972 8484 2984
rect 7208 2944 8484 2972
rect 8478 2932 8484 2944
rect 8536 2932 8542 2984
rect 8570 2932 8576 2984
rect 8628 2972 8634 2984
rect 9214 2972 9220 2984
rect 8628 2944 8673 2972
rect 8772 2944 9220 2972
rect 8628 2932 8634 2944
rect 6144 2876 7052 2904
rect 6144 2864 6150 2876
rect 7098 2864 7104 2916
rect 7156 2904 7162 2916
rect 7193 2907 7251 2913
rect 7193 2904 7205 2907
rect 7156 2876 7205 2904
rect 7156 2864 7162 2876
rect 7193 2873 7205 2876
rect 7239 2873 7251 2907
rect 7193 2867 7251 2873
rect 7285 2907 7343 2913
rect 7285 2873 7297 2907
rect 7331 2904 7343 2907
rect 7650 2904 7656 2916
rect 7331 2876 7656 2904
rect 7331 2873 7343 2876
rect 7285 2867 7343 2873
rect 7650 2864 7656 2876
rect 7708 2864 7714 2916
rect 8113 2907 8171 2913
rect 8113 2873 8125 2907
rect 8159 2904 8171 2907
rect 8772 2904 8800 2944
rect 9214 2932 9220 2944
rect 9272 2932 9278 2984
rect 9677 2975 9735 2981
rect 9677 2941 9689 2975
rect 9723 2972 9735 2975
rect 10410 2972 10416 2984
rect 9723 2944 10416 2972
rect 9723 2941 9735 2944
rect 9677 2935 9735 2941
rect 10410 2932 10416 2944
rect 10468 2932 10474 2984
rect 10594 2932 10600 2984
rect 10652 2972 10658 2984
rect 10873 2975 10931 2981
rect 10873 2972 10885 2975
rect 10652 2944 10885 2972
rect 10652 2932 10658 2944
rect 10873 2941 10885 2944
rect 10919 2941 10931 2975
rect 10873 2935 10931 2941
rect 11609 2975 11667 2981
rect 11609 2941 11621 2975
rect 11655 2972 11667 2975
rect 12342 2972 12348 2984
rect 11655 2944 12348 2972
rect 11655 2941 11667 2944
rect 11609 2935 11667 2941
rect 12342 2932 12348 2944
rect 12400 2932 12406 2984
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 12492 2944 12848 2972
rect 12492 2932 12498 2944
rect 8159 2876 8800 2904
rect 8849 2907 8907 2913
rect 8159 2873 8171 2876
rect 8113 2867 8171 2873
rect 8849 2873 8861 2907
rect 8895 2904 8907 2907
rect 9122 2904 9128 2916
rect 8895 2876 9128 2904
rect 8895 2873 8907 2876
rect 8849 2867 8907 2873
rect 9122 2864 9128 2876
rect 9180 2864 9186 2916
rect 10781 2907 10839 2913
rect 9416 2876 10548 2904
rect 2866 2796 2872 2848
rect 2924 2836 2930 2848
rect 3878 2836 3884 2848
rect 2924 2808 3884 2836
rect 2924 2796 2930 2808
rect 3878 2796 3884 2808
rect 3936 2796 3942 2848
rect 4338 2836 4344 2848
rect 4299 2808 4344 2836
rect 4338 2796 4344 2808
rect 4396 2796 4402 2848
rect 4798 2836 4804 2848
rect 4759 2808 4804 2836
rect 4798 2796 4804 2808
rect 4856 2796 4862 2848
rect 5169 2839 5227 2845
rect 5169 2805 5181 2839
rect 5215 2836 5227 2839
rect 5350 2836 5356 2848
rect 5215 2808 5356 2836
rect 5215 2805 5227 2808
rect 5169 2799 5227 2805
rect 5350 2796 5356 2808
rect 5408 2796 5414 2848
rect 5442 2796 5448 2848
rect 5500 2836 5506 2848
rect 5537 2839 5595 2845
rect 5537 2836 5549 2839
rect 5500 2808 5549 2836
rect 5500 2796 5506 2808
rect 5537 2805 5549 2808
rect 5583 2805 5595 2839
rect 5537 2799 5595 2805
rect 5629 2839 5687 2845
rect 5629 2805 5641 2839
rect 5675 2836 5687 2839
rect 7834 2836 7840 2848
rect 5675 2808 7840 2836
rect 5675 2805 5687 2808
rect 5629 2799 5687 2805
rect 7834 2796 7840 2808
rect 7892 2796 7898 2848
rect 8021 2839 8079 2845
rect 8021 2805 8033 2839
rect 8067 2836 8079 2839
rect 9416 2836 9444 2876
rect 8067 2808 9444 2836
rect 8067 2805 8079 2808
rect 8021 2799 8079 2805
rect 9490 2796 9496 2848
rect 9548 2836 9554 2848
rect 9585 2839 9643 2845
rect 9585 2836 9597 2839
rect 9548 2808 9597 2836
rect 9548 2796 9554 2808
rect 9585 2805 9597 2808
rect 9631 2805 9643 2839
rect 9585 2799 9643 2805
rect 9766 2796 9772 2848
rect 9824 2836 9830 2848
rect 10413 2839 10471 2845
rect 10413 2836 10425 2839
rect 9824 2808 10425 2836
rect 9824 2796 9830 2808
rect 10413 2805 10425 2808
rect 10459 2805 10471 2839
rect 10520 2836 10548 2876
rect 10781 2873 10793 2907
rect 10827 2904 10839 2907
rect 11238 2904 11244 2916
rect 10827 2876 11244 2904
rect 10827 2873 10839 2876
rect 10781 2867 10839 2873
rect 11238 2864 11244 2876
rect 11296 2864 11302 2916
rect 11701 2907 11759 2913
rect 11701 2873 11713 2907
rect 11747 2904 11759 2907
rect 11882 2904 11888 2916
rect 11747 2876 11888 2904
rect 11747 2873 11759 2876
rect 11701 2867 11759 2873
rect 11882 2864 11888 2876
rect 11940 2904 11946 2916
rect 12820 2913 12848 2944
rect 12986 2932 12992 2984
rect 13044 2972 13050 2984
rect 13633 2975 13691 2981
rect 13633 2972 13645 2975
rect 13044 2944 13645 2972
rect 13044 2932 13050 2944
rect 13633 2941 13645 2944
rect 13679 2941 13691 2975
rect 13633 2935 13691 2941
rect 14090 2932 14096 2984
rect 14148 2972 14154 2984
rect 14550 2972 14556 2984
rect 14148 2944 14556 2972
rect 14148 2932 14154 2944
rect 14550 2932 14556 2944
rect 14608 2932 14614 2984
rect 14826 2932 14832 2984
rect 14884 2972 14890 2984
rect 15473 2975 15531 2981
rect 15473 2972 15485 2975
rect 14884 2944 15485 2972
rect 14884 2932 14890 2944
rect 15473 2941 15485 2944
rect 15519 2941 15531 2975
rect 15473 2935 15531 2941
rect 12805 2907 12863 2913
rect 11940 2876 12572 2904
rect 11940 2864 11946 2876
rect 12158 2836 12164 2848
rect 10520 2808 12164 2836
rect 10413 2799 10471 2805
rect 12158 2796 12164 2808
rect 12216 2796 12222 2848
rect 12342 2796 12348 2848
rect 12400 2836 12406 2848
rect 12437 2839 12495 2845
rect 12437 2836 12449 2839
rect 12400 2808 12449 2836
rect 12400 2796 12406 2808
rect 12437 2805 12449 2808
rect 12483 2805 12495 2839
rect 12544 2836 12572 2876
rect 12805 2873 12817 2907
rect 12851 2904 12863 2907
rect 14642 2904 14648 2916
rect 12851 2876 14648 2904
rect 12851 2873 12863 2876
rect 12805 2867 12863 2873
rect 14642 2864 14648 2876
rect 14700 2904 14706 2916
rect 14700 2876 14872 2904
rect 14700 2864 14706 2876
rect 13998 2836 14004 2848
rect 12544 2808 14004 2836
rect 12437 2799 12495 2805
rect 13998 2796 14004 2808
rect 14056 2796 14062 2848
rect 14734 2836 14740 2848
rect 14695 2808 14740 2836
rect 14734 2796 14740 2808
rect 14792 2796 14798 2848
rect 14844 2836 14872 2876
rect 15102 2864 15108 2916
rect 15160 2904 15166 2916
rect 16758 2904 16764 2916
rect 15160 2876 16764 2904
rect 15160 2864 15166 2876
rect 16758 2864 16764 2876
rect 16816 2864 16822 2916
rect 15286 2836 15292 2848
rect 14844 2808 15292 2836
rect 15286 2796 15292 2808
rect 15344 2796 15350 2848
rect 1104 2746 15824 2768
rect 1104 2694 5912 2746
rect 5964 2694 5976 2746
rect 6028 2694 6040 2746
rect 6092 2694 6104 2746
rect 6156 2694 10843 2746
rect 10895 2694 10907 2746
rect 10959 2694 10971 2746
rect 11023 2694 11035 2746
rect 11087 2694 15824 2746
rect 1104 2672 15824 2694
rect 2041 2635 2099 2641
rect 2041 2601 2053 2635
rect 2087 2632 2099 2635
rect 2314 2632 2320 2644
rect 2087 2604 2320 2632
rect 2087 2601 2099 2604
rect 2041 2595 2099 2601
rect 2314 2592 2320 2604
rect 2372 2592 2378 2644
rect 2866 2632 2872 2644
rect 2827 2604 2872 2632
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 3237 2635 3295 2641
rect 3237 2601 3249 2635
rect 3283 2632 3295 2635
rect 3326 2632 3332 2644
rect 3283 2604 3332 2632
rect 3283 2601 3295 2604
rect 3237 2595 3295 2601
rect 3326 2592 3332 2604
rect 3384 2592 3390 2644
rect 3970 2632 3976 2644
rect 3712 2604 3976 2632
rect 2222 2524 2228 2576
rect 2280 2524 2286 2576
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2496 2007 2499
rect 2240 2496 2268 2524
rect 3712 2496 3740 2604
rect 3970 2592 3976 2604
rect 4028 2592 4034 2644
rect 5534 2632 5540 2644
rect 5495 2604 5540 2632
rect 5534 2592 5540 2604
rect 5592 2592 5598 2644
rect 5810 2592 5816 2644
rect 5868 2632 5874 2644
rect 5997 2635 6055 2641
rect 5997 2632 6009 2635
rect 5868 2604 6009 2632
rect 5868 2592 5874 2604
rect 5997 2601 6009 2604
rect 6043 2601 6055 2635
rect 5997 2595 6055 2601
rect 6730 2592 6736 2644
rect 6788 2632 6794 2644
rect 6788 2604 7512 2632
rect 6788 2592 6794 2604
rect 7377 2567 7435 2573
rect 7377 2564 7389 2567
rect 1995 2468 3740 2496
rect 3804 2536 7389 2564
rect 1995 2465 2007 2468
rect 1949 2459 2007 2465
rect 2222 2428 2228 2440
rect 2183 2400 2228 2428
rect 2222 2388 2228 2400
rect 2280 2388 2286 2440
rect 2777 2431 2835 2437
rect 2777 2397 2789 2431
rect 2823 2428 2835 2431
rect 3234 2428 3240 2440
rect 2823 2400 3240 2428
rect 2823 2397 2835 2400
rect 2777 2391 2835 2397
rect 3234 2388 3240 2400
rect 3292 2428 3298 2440
rect 3329 2431 3387 2437
rect 3329 2428 3341 2431
rect 3292 2400 3341 2428
rect 3292 2388 3298 2400
rect 3329 2397 3341 2400
rect 3375 2397 3387 2431
rect 3329 2391 3387 2397
rect 3418 2388 3424 2440
rect 3476 2428 3482 2440
rect 3694 2428 3700 2440
rect 3476 2400 3521 2428
rect 3655 2400 3700 2428
rect 3476 2388 3482 2400
rect 3694 2388 3700 2400
rect 3752 2388 3758 2440
rect 1581 2363 1639 2369
rect 1581 2329 1593 2363
rect 1627 2360 1639 2363
rect 3804 2360 3832 2536
rect 7377 2533 7389 2536
rect 7423 2533 7435 2567
rect 7484 2564 7512 2604
rect 7834 2592 7840 2644
rect 7892 2632 7898 2644
rect 8665 2635 8723 2641
rect 8665 2632 8677 2635
rect 7892 2604 8677 2632
rect 7892 2592 7898 2604
rect 8665 2601 8677 2604
rect 8711 2601 8723 2635
rect 8665 2595 8723 2601
rect 9582 2592 9588 2644
rect 9640 2632 9646 2644
rect 10965 2635 11023 2641
rect 10965 2632 10977 2635
rect 9640 2604 10977 2632
rect 9640 2592 9646 2604
rect 10965 2601 10977 2604
rect 11011 2601 11023 2635
rect 10965 2595 11023 2601
rect 11425 2635 11483 2641
rect 11425 2601 11437 2635
rect 11471 2632 11483 2635
rect 12250 2632 12256 2644
rect 11471 2604 12256 2632
rect 11471 2601 11483 2604
rect 11425 2595 11483 2601
rect 12250 2592 12256 2604
rect 12308 2592 12314 2644
rect 12342 2592 12348 2644
rect 12400 2632 12406 2644
rect 13262 2632 13268 2644
rect 12400 2604 13268 2632
rect 12400 2592 12406 2604
rect 13262 2592 13268 2604
rect 13320 2592 13326 2644
rect 7484 2536 9628 2564
rect 7377 2527 7435 2533
rect 4332 2499 4390 2505
rect 4332 2465 4344 2499
rect 4378 2496 4390 2499
rect 4378 2468 5488 2496
rect 4378 2465 4390 2468
rect 4332 2459 4390 2465
rect 5460 2428 5488 2468
rect 5534 2456 5540 2508
rect 5592 2496 5598 2508
rect 5905 2499 5963 2505
rect 5905 2496 5917 2499
rect 5592 2468 5917 2496
rect 5592 2456 5598 2468
rect 5905 2465 5917 2468
rect 5951 2465 5963 2499
rect 7006 2496 7012 2508
rect 5905 2459 5963 2465
rect 5992 2468 7012 2496
rect 5992 2428 6020 2468
rect 7006 2456 7012 2468
rect 7064 2456 7070 2508
rect 7098 2456 7104 2508
rect 7156 2496 7162 2508
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 7156 2468 7297 2496
rect 7156 2456 7162 2468
rect 7285 2465 7297 2468
rect 7331 2496 7343 2499
rect 8202 2496 8208 2508
rect 7331 2468 8208 2496
rect 7331 2465 7343 2468
rect 7285 2459 7343 2465
rect 8202 2456 8208 2468
rect 8260 2456 8266 2508
rect 8573 2499 8631 2505
rect 8573 2465 8585 2499
rect 8619 2496 8631 2499
rect 8938 2496 8944 2508
rect 8619 2468 8944 2496
rect 8619 2465 8631 2468
rect 8573 2459 8631 2465
rect 8938 2456 8944 2468
rect 8996 2456 9002 2508
rect 9600 2505 9628 2536
rect 10042 2524 10048 2576
rect 10100 2564 10106 2576
rect 11333 2567 11391 2573
rect 10100 2536 10732 2564
rect 10100 2524 10106 2536
rect 9585 2499 9643 2505
rect 9585 2465 9597 2499
rect 9631 2465 9643 2499
rect 9585 2459 9643 2465
rect 10137 2499 10195 2505
rect 10137 2465 10149 2499
rect 10183 2496 10195 2499
rect 10594 2496 10600 2508
rect 10183 2468 10600 2496
rect 10183 2465 10195 2468
rect 10137 2459 10195 2465
rect 10594 2456 10600 2468
rect 10652 2456 10658 2508
rect 5460 2400 6020 2428
rect 6181 2431 6239 2437
rect 6181 2397 6193 2431
rect 6227 2428 6239 2431
rect 6546 2428 6552 2440
rect 6227 2400 6552 2428
rect 6227 2397 6239 2400
rect 6181 2391 6239 2397
rect 6546 2388 6552 2400
rect 6604 2388 6610 2440
rect 7466 2428 7472 2440
rect 7427 2400 7472 2428
rect 7466 2388 7472 2400
rect 7524 2388 7530 2440
rect 8754 2428 8760 2440
rect 8715 2400 8760 2428
rect 8754 2388 8760 2400
rect 8812 2388 8818 2440
rect 9214 2388 9220 2440
rect 9272 2428 9278 2440
rect 10042 2428 10048 2440
rect 9272 2400 10048 2428
rect 9272 2388 9278 2400
rect 10042 2388 10048 2400
rect 10100 2388 10106 2440
rect 10229 2431 10287 2437
rect 10229 2397 10241 2431
rect 10275 2428 10287 2431
rect 10318 2428 10324 2440
rect 10275 2400 10324 2428
rect 10275 2397 10287 2400
rect 10229 2391 10287 2397
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 10410 2388 10416 2440
rect 10468 2428 10474 2440
rect 10704 2428 10732 2536
rect 11333 2533 11345 2567
rect 11379 2564 11391 2567
rect 13630 2564 13636 2576
rect 11379 2536 13636 2564
rect 11379 2533 11391 2536
rect 11333 2527 11391 2533
rect 13630 2524 13636 2536
rect 13688 2524 13694 2576
rect 14737 2567 14795 2573
rect 14737 2533 14749 2567
rect 14783 2564 14795 2567
rect 15102 2564 15108 2576
rect 14783 2536 15108 2564
rect 14783 2533 14795 2536
rect 14737 2527 14795 2533
rect 15102 2524 15108 2536
rect 15160 2524 15166 2576
rect 11606 2456 11612 2508
rect 11664 2496 11670 2508
rect 11793 2499 11851 2505
rect 11793 2496 11805 2499
rect 11664 2468 11805 2496
rect 11664 2456 11670 2468
rect 11793 2465 11805 2468
rect 11839 2496 11851 2499
rect 12342 2496 12348 2508
rect 11839 2468 12348 2496
rect 11839 2465 11851 2468
rect 11793 2459 11851 2465
rect 12342 2456 12348 2468
rect 12400 2456 12406 2508
rect 12618 2496 12624 2508
rect 12579 2468 12624 2496
rect 12618 2456 12624 2468
rect 12676 2456 12682 2508
rect 12710 2456 12716 2508
rect 12768 2496 12774 2508
rect 13541 2499 13599 2505
rect 13541 2496 13553 2499
rect 12768 2468 13553 2496
rect 12768 2456 12774 2468
rect 13541 2465 13553 2468
rect 13587 2465 13599 2499
rect 14458 2496 14464 2508
rect 14419 2468 14464 2496
rect 13541 2459 13599 2465
rect 14458 2456 14464 2468
rect 14516 2456 14522 2508
rect 11517 2431 11575 2437
rect 11517 2428 11529 2431
rect 10468 2400 10513 2428
rect 10704 2400 11529 2428
rect 10468 2388 10474 2400
rect 11517 2397 11529 2400
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 11698 2388 11704 2440
rect 11756 2428 11762 2440
rect 11974 2428 11980 2440
rect 11756 2400 11980 2428
rect 11756 2388 11762 2400
rect 11974 2388 11980 2400
rect 12032 2388 12038 2440
rect 12802 2428 12808 2440
rect 12763 2400 12808 2428
rect 12802 2388 12808 2400
rect 12860 2388 12866 2440
rect 13722 2428 13728 2440
rect 13683 2400 13728 2428
rect 13722 2388 13728 2400
rect 13780 2388 13786 2440
rect 1627 2332 3832 2360
rect 1627 2329 1639 2332
rect 1581 2323 1639 2329
rect 5350 2320 5356 2372
rect 5408 2360 5414 2372
rect 5810 2360 5816 2372
rect 5408 2332 5816 2360
rect 5408 2320 5414 2332
rect 5810 2320 5816 2332
rect 5868 2320 5874 2372
rect 8205 2363 8263 2369
rect 8205 2329 8217 2363
rect 8251 2360 8263 2363
rect 14182 2360 14188 2372
rect 8251 2332 14188 2360
rect 8251 2329 8263 2332
rect 8205 2323 8263 2329
rect 14182 2320 14188 2332
rect 14240 2320 14246 2372
rect 3605 2295 3663 2301
rect 3605 2261 3617 2295
rect 3651 2292 3663 2295
rect 3786 2292 3792 2304
rect 3651 2264 3792 2292
rect 3651 2261 3663 2264
rect 3605 2255 3663 2261
rect 3786 2252 3792 2264
rect 3844 2292 3850 2304
rect 4062 2292 4068 2304
rect 3844 2264 4068 2292
rect 3844 2252 3850 2264
rect 4062 2252 4068 2264
rect 4120 2252 4126 2304
rect 4246 2252 4252 2304
rect 4304 2292 4310 2304
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 4304 2264 5457 2292
rect 4304 2252 4310 2264
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 6914 2292 6920 2304
rect 6875 2264 6920 2292
rect 5445 2255 5503 2261
rect 6914 2252 6920 2264
rect 6972 2252 6978 2304
rect 7926 2252 7932 2304
rect 7984 2292 7990 2304
rect 9122 2292 9128 2304
rect 7984 2264 9128 2292
rect 7984 2252 7990 2264
rect 9122 2252 9128 2264
rect 9180 2252 9186 2304
rect 9398 2292 9404 2304
rect 9359 2264 9404 2292
rect 9398 2252 9404 2264
rect 9456 2252 9462 2304
rect 9766 2292 9772 2304
rect 9727 2264 9772 2292
rect 9766 2252 9772 2264
rect 9824 2252 9830 2304
rect 10042 2252 10048 2304
rect 10100 2292 10106 2304
rect 11698 2292 11704 2304
rect 10100 2264 11704 2292
rect 10100 2252 10106 2264
rect 11698 2252 11704 2264
rect 11756 2252 11762 2304
rect 11974 2292 11980 2304
rect 11935 2264 11980 2292
rect 11974 2252 11980 2264
rect 12032 2252 12038 2304
rect 1104 2202 15824 2224
rect 1104 2150 3447 2202
rect 3499 2150 3511 2202
rect 3563 2150 3575 2202
rect 3627 2150 3639 2202
rect 3691 2150 8378 2202
rect 8430 2150 8442 2202
rect 8494 2150 8506 2202
rect 8558 2150 8570 2202
rect 8622 2150 13308 2202
rect 13360 2150 13372 2202
rect 13424 2150 13436 2202
rect 13488 2150 13500 2202
rect 13552 2150 15824 2202
rect 1104 2128 15824 2150
rect 5258 2048 5264 2100
rect 5316 2088 5322 2100
rect 9398 2088 9404 2100
rect 5316 2060 9404 2088
rect 5316 2048 5322 2060
rect 9398 2048 9404 2060
rect 9456 2048 9462 2100
rect 10686 2048 10692 2100
rect 10744 2088 10750 2100
rect 13170 2088 13176 2100
rect 10744 2060 13176 2088
rect 10744 2048 10750 2060
rect 13170 2048 13176 2060
rect 13228 2048 13234 2100
rect 14458 2088 14464 2100
rect 14419 2060 14464 2088
rect 14458 2048 14464 2060
rect 14516 2048 14522 2100
rect 2038 1980 2044 2032
rect 2096 2020 2102 2032
rect 12802 2020 12808 2032
rect 2096 1992 12808 2020
rect 2096 1980 2102 1992
rect 12802 1980 12808 1992
rect 12860 1980 12866 2032
rect 198 1912 204 1964
rect 256 1952 262 1964
rect 11974 1952 11980 1964
rect 256 1924 11980 1952
rect 256 1912 262 1924
rect 11974 1912 11980 1924
rect 12032 1912 12038 1964
rect 4154 1844 4160 1896
rect 4212 1884 4218 1896
rect 6733 1887 6791 1893
rect 6733 1884 6745 1887
rect 4212 1856 6745 1884
rect 4212 1844 4218 1856
rect 6733 1853 6745 1856
rect 6779 1853 6791 1887
rect 6733 1847 6791 1853
rect 7006 1844 7012 1896
rect 7064 1884 7070 1896
rect 11606 1884 11612 1896
rect 7064 1856 11612 1884
rect 7064 1844 7070 1856
rect 11606 1844 11612 1856
rect 11664 1844 11670 1896
rect 11701 1887 11759 1893
rect 11701 1853 11713 1887
rect 11747 1884 11759 1887
rect 13722 1884 13728 1896
rect 11747 1856 13728 1884
rect 11747 1853 11759 1856
rect 11701 1847 11759 1853
rect 13722 1844 13728 1856
rect 13780 1844 13786 1896
rect 4890 1776 4896 1828
rect 4948 1816 4954 1828
rect 7101 1819 7159 1825
rect 7101 1816 7113 1819
rect 4948 1788 7113 1816
rect 4948 1776 4954 1788
rect 7101 1785 7113 1788
rect 7147 1785 7159 1819
rect 7101 1779 7159 1785
rect 7282 1776 7288 1828
rect 7340 1816 7346 1828
rect 10962 1816 10968 1828
rect 7340 1788 10968 1816
rect 7340 1776 7346 1788
rect 10962 1776 10968 1788
rect 11020 1776 11026 1828
rect 11057 1819 11115 1825
rect 11057 1785 11069 1819
rect 11103 1816 11115 1819
rect 12618 1816 12624 1828
rect 11103 1788 12624 1816
rect 11103 1785 11115 1788
rect 11057 1779 11115 1785
rect 12618 1776 12624 1788
rect 12676 1776 12682 1828
rect 2958 1708 2964 1760
rect 3016 1748 3022 1760
rect 9766 1748 9772 1760
rect 3016 1720 9772 1748
rect 3016 1708 3022 1720
rect 9766 1708 9772 1720
rect 9824 1708 9830 1760
rect 10594 1708 10600 1760
rect 10652 1748 10658 1760
rect 15470 1748 15476 1760
rect 10652 1720 15476 1748
rect 10652 1708 10658 1720
rect 15470 1708 15476 1720
rect 15528 1708 15534 1760
rect 1946 1640 1952 1692
rect 2004 1680 2010 1692
rect 6914 1680 6920 1692
rect 2004 1652 6920 1680
rect 2004 1640 2010 1652
rect 6914 1640 6920 1652
rect 6972 1640 6978 1692
rect 7101 1683 7159 1689
rect 7101 1649 7113 1683
rect 7147 1680 7159 1683
rect 12710 1680 12716 1692
rect 7147 1652 12716 1680
rect 7147 1649 7159 1652
rect 7101 1643 7159 1649
rect 12710 1640 12716 1652
rect 12768 1640 12774 1692
rect 2222 1572 2228 1624
rect 2280 1612 2286 1624
rect 10226 1612 10232 1624
rect 2280 1584 10232 1612
rect 2280 1572 2286 1584
rect 10226 1572 10232 1584
rect 10284 1572 10290 1624
rect 11146 1572 11152 1624
rect 11204 1612 11210 1624
rect 16298 1612 16304 1624
rect 11204 1584 16304 1612
rect 11204 1572 11210 1584
rect 16298 1572 16304 1584
rect 16356 1572 16362 1624
rect 6270 1504 6276 1556
rect 6328 1544 6334 1556
rect 8478 1544 8484 1556
rect 6328 1516 8484 1544
rect 6328 1504 6334 1516
rect 8478 1504 8484 1516
rect 8536 1504 8542 1556
rect 8846 1504 8852 1556
rect 8904 1544 8910 1556
rect 9858 1544 9864 1556
rect 8904 1516 9864 1544
rect 8904 1504 8910 1516
rect 9858 1504 9864 1516
rect 9916 1504 9922 1556
rect 11422 1504 11428 1556
rect 11480 1544 11486 1556
rect 15102 1544 15108 1556
rect 11480 1516 15108 1544
rect 11480 1504 11486 1516
rect 15102 1504 15108 1516
rect 15160 1504 15166 1556
rect 1394 1436 1400 1488
rect 1452 1476 1458 1488
rect 6638 1476 6644 1488
rect 1452 1448 6644 1476
rect 1452 1436 1458 1448
rect 6638 1436 6644 1448
rect 6696 1436 6702 1488
rect 6733 1479 6791 1485
rect 6733 1445 6745 1479
rect 6779 1476 6791 1479
rect 11057 1479 11115 1485
rect 11057 1476 11069 1479
rect 6779 1448 11069 1476
rect 6779 1445 6791 1448
rect 6733 1439 6791 1445
rect 11057 1445 11069 1448
rect 11103 1445 11115 1479
rect 11057 1439 11115 1445
rect 1118 1368 1124 1420
rect 1176 1408 1182 1420
rect 11701 1411 11759 1417
rect 11701 1408 11713 1411
rect 1176 1380 11713 1408
rect 1176 1368 1182 1380
rect 11701 1377 11713 1380
rect 11747 1377 11759 1411
rect 14461 1411 14519 1417
rect 14461 1408 14473 1411
rect 11701 1371 11759 1377
rect 11808 1380 14473 1408
rect 2222 1300 2228 1352
rect 2280 1340 2286 1352
rect 9490 1340 9496 1352
rect 2280 1312 9496 1340
rect 2280 1300 2286 1312
rect 9490 1300 9496 1312
rect 9548 1300 9554 1352
rect 937 1275 995 1281
rect 937 1241 949 1275
rect 983 1272 995 1275
rect 5994 1272 6000 1284
rect 983 1244 6000 1272
rect 983 1241 995 1244
rect 937 1235 995 1241
rect 5994 1232 6000 1244
rect 6052 1232 6058 1284
rect 6730 1232 6736 1284
rect 6788 1272 6794 1284
rect 11808 1272 11836 1380
rect 14461 1377 14473 1380
rect 14507 1377 14519 1411
rect 14461 1371 14519 1377
rect 6788 1244 11836 1272
rect 6788 1232 6794 1244
rect 1854 1164 1860 1216
rect 1912 1204 1918 1216
rect 7558 1204 7564 1216
rect 1912 1176 7564 1204
rect 1912 1164 1918 1176
rect 7558 1164 7564 1176
rect 7616 1164 7622 1216
rect 4706 1096 4712 1148
rect 4764 1136 4770 1148
rect 9306 1136 9312 1148
rect 4764 1108 9312 1136
rect 4764 1096 4770 1108
rect 9306 1096 9312 1108
rect 9364 1096 9370 1148
rect 7374 1028 7380 1080
rect 7432 1068 7438 1080
rect 13078 1068 13084 1080
rect 7432 1040 13084 1068
rect 7432 1028 7438 1040
rect 13078 1028 13084 1040
rect 13136 1028 13142 1080
rect 8202 960 8208 1012
rect 8260 1000 8266 1012
rect 9306 1000 9312 1012
rect 8260 972 9312 1000
rect 8260 960 8266 972
rect 9306 960 9312 972
rect 9364 960 9370 1012
rect 4430 892 4436 944
rect 4488 932 4494 944
rect 9582 932 9588 944
rect 4488 904 9588 932
rect 4488 892 4494 904
rect 9582 892 9588 904
rect 9640 892 9646 944
rect 8938 620 8944 672
rect 8996 660 9002 672
rect 12618 660 12624 672
rect 8996 632 12624 660
rect 8996 620 9002 632
rect 12618 620 12624 632
rect 12676 620 12682 672
<< via1 >>
rect 12256 18776 12308 18828
rect 13912 18776 13964 18828
rect 10600 18232 10652 18284
rect 11060 18232 11112 18284
rect 8300 18164 8352 18216
rect 9588 18164 9640 18216
rect 10508 18164 10560 18216
rect 15108 18164 15160 18216
rect 3424 18096 3476 18148
rect 8852 18096 8904 18148
rect 10692 18096 10744 18148
rect 11428 18096 11480 18148
rect 7472 18028 7524 18080
rect 11152 18028 11204 18080
rect 3516 17960 3568 18012
rect 12808 17960 12860 18012
rect 6092 17892 6144 17944
rect 8944 17892 8996 17944
rect 7104 17824 7156 17876
rect 9680 17824 9732 17876
rect 7932 17756 7984 17808
rect 10232 17756 10284 17808
rect 11704 17756 11756 17808
rect 12348 17756 12400 17808
rect 1768 17688 1820 17740
rect 12532 17688 12584 17740
rect 7012 17620 7064 17672
rect 14004 17620 14056 17672
rect 572 17552 624 17604
rect 11980 17552 12032 17604
rect 13544 17552 13596 17604
rect 14188 17552 14240 17604
rect 4988 17484 5040 17536
rect 6276 17484 6328 17536
rect 6368 17484 6420 17536
rect 10140 17484 10192 17536
rect 3447 17382 3499 17434
rect 3511 17382 3563 17434
rect 3575 17382 3627 17434
rect 3639 17382 3691 17434
rect 8378 17382 8430 17434
rect 8442 17382 8494 17434
rect 8506 17382 8558 17434
rect 8570 17382 8622 17434
rect 13308 17382 13360 17434
rect 13372 17382 13424 17434
rect 13436 17382 13488 17434
rect 13500 17382 13552 17434
rect 4252 17280 4304 17332
rect 7840 17212 7892 17264
rect 5172 17144 5224 17196
rect 5264 17144 5316 17196
rect 6092 17187 6144 17196
rect 6092 17153 6101 17187
rect 6101 17153 6135 17187
rect 6135 17153 6144 17187
rect 6092 17144 6144 17153
rect 5356 17076 5408 17128
rect 6644 17144 6696 17196
rect 7380 17144 7432 17196
rect 7656 17144 7708 17196
rect 8024 17144 8076 17196
rect 10416 17187 10468 17196
rect 10416 17153 10425 17187
rect 10425 17153 10459 17187
rect 10459 17153 10468 17187
rect 10416 17144 10468 17153
rect 7196 17076 7248 17128
rect 10324 17076 10376 17128
rect 12164 17144 12216 17196
rect 11796 17076 11848 17128
rect 13636 17144 13688 17196
rect 14556 17187 14608 17196
rect 14556 17153 14565 17187
rect 14565 17153 14599 17187
rect 14599 17153 14608 17187
rect 14556 17144 14608 17153
rect 2136 17051 2188 17060
rect 2136 17017 2145 17051
rect 2145 17017 2179 17051
rect 2179 17017 2188 17051
rect 2136 17008 2188 17017
rect 3056 17051 3108 17060
rect 3056 17017 3065 17051
rect 3065 17017 3099 17051
rect 3099 17017 3108 17051
rect 3056 17008 3108 17017
rect 4528 17008 4580 17060
rect 4988 17008 5040 17060
rect 4804 16983 4856 16992
rect 4804 16949 4813 16983
rect 4813 16949 4847 16983
rect 4847 16949 4856 16983
rect 4804 16940 4856 16949
rect 5080 16940 5132 16992
rect 8484 17008 8536 17060
rect 8668 17008 8720 17060
rect 12256 17008 12308 17060
rect 12808 17008 12860 17060
rect 13728 17008 13780 17060
rect 6736 16940 6788 16992
rect 7472 16940 7524 16992
rect 7748 16940 7800 16992
rect 8944 16940 8996 16992
rect 9772 16983 9824 16992
rect 9772 16949 9781 16983
rect 9781 16949 9815 16983
rect 9815 16949 9824 16983
rect 9772 16940 9824 16949
rect 10692 16940 10744 16992
rect 11152 16983 11204 16992
rect 11152 16949 11161 16983
rect 11161 16949 11195 16983
rect 11195 16949 11204 16983
rect 11152 16940 11204 16949
rect 5912 16838 5964 16890
rect 5976 16838 6028 16890
rect 6040 16838 6092 16890
rect 6104 16838 6156 16890
rect 10843 16838 10895 16890
rect 10907 16838 10959 16890
rect 10971 16838 11023 16890
rect 11035 16838 11087 16890
rect 3332 16736 3384 16788
rect 1584 16643 1636 16652
rect 1584 16609 1593 16643
rect 1593 16609 1627 16643
rect 1627 16609 1636 16643
rect 1584 16600 1636 16609
rect 1860 16643 1912 16652
rect 1860 16609 1869 16643
rect 1869 16609 1903 16643
rect 1903 16609 1912 16643
rect 1860 16600 1912 16609
rect 2412 16600 2464 16652
rect 2964 16600 3016 16652
rect 5632 16736 5684 16788
rect 6276 16736 6328 16788
rect 6736 16736 6788 16788
rect 7104 16736 7156 16788
rect 9680 16779 9732 16788
rect 9680 16745 9689 16779
rect 9689 16745 9723 16779
rect 9723 16745 9732 16779
rect 9680 16736 9732 16745
rect 10140 16736 10192 16788
rect 10232 16736 10284 16788
rect 14004 16779 14056 16788
rect 14004 16745 14013 16779
rect 14013 16745 14047 16779
rect 14047 16745 14056 16779
rect 14004 16736 14056 16745
rect 2228 16532 2280 16584
rect 7932 16668 7984 16720
rect 8300 16668 8352 16720
rect 11060 16668 11112 16720
rect 12900 16668 12952 16720
rect 4896 16600 4948 16652
rect 4344 16575 4396 16584
rect 4344 16541 4353 16575
rect 4353 16541 4387 16575
rect 4387 16541 4396 16575
rect 4344 16532 4396 16541
rect 1400 16464 1452 16516
rect 4252 16464 4304 16516
rect 5724 16507 5776 16516
rect 5724 16473 5733 16507
rect 5733 16473 5767 16507
rect 5767 16473 5776 16507
rect 5724 16464 5776 16473
rect 6368 16600 6420 16652
rect 7288 16643 7340 16652
rect 7288 16609 7297 16643
rect 7297 16609 7331 16643
rect 7331 16609 7340 16643
rect 7288 16600 7340 16609
rect 8116 16600 8168 16652
rect 8208 16600 8260 16652
rect 9864 16600 9916 16652
rect 10784 16600 10836 16652
rect 11152 16600 11204 16652
rect 12348 16643 12400 16652
rect 12348 16609 12357 16643
rect 12357 16609 12391 16643
rect 12391 16609 12400 16643
rect 12348 16600 12400 16609
rect 13084 16643 13136 16652
rect 13084 16609 13093 16643
rect 13093 16609 13127 16643
rect 13127 16609 13136 16643
rect 13084 16600 13136 16609
rect 13912 16600 13964 16652
rect 14280 16600 14332 16652
rect 7932 16532 7984 16584
rect 9312 16532 9364 16584
rect 10232 16532 10284 16584
rect 10416 16532 10468 16584
rect 2228 16396 2280 16448
rect 6736 16396 6788 16448
rect 6920 16439 6972 16448
rect 6920 16405 6929 16439
rect 6929 16405 6963 16439
rect 6963 16405 6972 16439
rect 6920 16396 6972 16405
rect 7012 16396 7064 16448
rect 8852 16464 8904 16516
rect 12808 16532 12860 16584
rect 11980 16464 12032 16516
rect 12532 16507 12584 16516
rect 12532 16473 12541 16507
rect 12541 16473 12575 16507
rect 12575 16473 12584 16507
rect 12532 16464 12584 16473
rect 10416 16396 10468 16448
rect 10876 16396 10928 16448
rect 3447 16294 3499 16346
rect 3511 16294 3563 16346
rect 3575 16294 3627 16346
rect 3639 16294 3691 16346
rect 8378 16294 8430 16346
rect 8442 16294 8494 16346
rect 8506 16294 8558 16346
rect 8570 16294 8622 16346
rect 13308 16294 13360 16346
rect 13372 16294 13424 16346
rect 13436 16294 13488 16346
rect 13500 16294 13552 16346
rect 2872 16192 2924 16244
rect 204 16124 256 16176
rect 4068 16124 4120 16176
rect 4620 16192 4672 16244
rect 4712 16124 4764 16176
rect 2780 16056 2832 16108
rect 3976 16056 4028 16108
rect 4160 16056 4212 16108
rect 4988 16124 5040 16176
rect 4896 16099 4948 16108
rect 4896 16065 4905 16099
rect 4905 16065 4939 16099
rect 4939 16065 4948 16099
rect 4896 16056 4948 16065
rect 1676 15988 1728 16040
rect 6736 16056 6788 16108
rect 7104 16056 7156 16108
rect 9588 16192 9640 16244
rect 11244 16192 11296 16244
rect 11336 16192 11388 16244
rect 9680 16124 9732 16176
rect 7748 15988 7800 16040
rect 7840 15988 7892 16040
rect 8852 16056 8904 16108
rect 9312 16056 9364 16108
rect 9956 16056 10008 16108
rect 10324 16056 10376 16108
rect 10416 16056 10468 16108
rect 8944 15988 8996 16040
rect 9496 15988 9548 16040
rect 5448 15920 5500 15972
rect 7196 15920 7248 15972
rect 8668 15920 8720 15972
rect 3148 15852 3200 15904
rect 3516 15895 3568 15904
rect 3516 15861 3525 15895
rect 3525 15861 3559 15895
rect 3559 15861 3568 15895
rect 3516 15852 3568 15861
rect 3884 15852 3936 15904
rect 4344 15895 4396 15904
rect 4344 15861 4353 15895
rect 4353 15861 4387 15895
rect 4387 15861 4396 15895
rect 4344 15852 4396 15861
rect 6276 15852 6328 15904
rect 9036 15852 9088 15904
rect 9220 15895 9272 15904
rect 9220 15861 9229 15895
rect 9229 15861 9263 15895
rect 9263 15861 9272 15895
rect 9220 15852 9272 15861
rect 9588 15852 9640 15904
rect 10048 15920 10100 15972
rect 10784 15963 10836 15972
rect 10784 15929 10793 15963
rect 10793 15929 10827 15963
rect 10827 15929 10836 15963
rect 10784 15920 10836 15929
rect 10232 15852 10284 15904
rect 10416 15895 10468 15904
rect 10416 15861 10425 15895
rect 10425 15861 10459 15895
rect 10459 15861 10468 15895
rect 10416 15852 10468 15861
rect 10692 15852 10744 15904
rect 11060 15920 11112 15972
rect 11888 15988 11940 16040
rect 12072 16056 12124 16108
rect 16764 16056 16816 16108
rect 12532 15988 12584 16040
rect 12900 15988 12952 16040
rect 12992 15988 13044 16040
rect 14556 15988 14608 16040
rect 11980 15920 12032 15972
rect 13728 15920 13780 15972
rect 14924 15852 14976 15904
rect 5912 15750 5964 15802
rect 5976 15750 6028 15802
rect 6040 15750 6092 15802
rect 6104 15750 6156 15802
rect 10843 15750 10895 15802
rect 10907 15750 10959 15802
rect 10971 15750 11023 15802
rect 11035 15750 11087 15802
rect 2780 15691 2832 15700
rect 2780 15657 2789 15691
rect 2789 15657 2823 15691
rect 2823 15657 2832 15691
rect 2780 15648 2832 15657
rect 5540 15648 5592 15700
rect 940 15580 992 15632
rect 6828 15580 6880 15632
rect 7012 15580 7064 15632
rect 7196 15648 7248 15700
rect 10324 15648 10376 15700
rect 11888 15648 11940 15700
rect 10784 15580 10836 15632
rect 10968 15580 11020 15632
rect 12808 15648 12860 15700
rect 12072 15580 12124 15632
rect 12716 15580 12768 15632
rect 2320 15512 2372 15564
rect 3424 15512 3476 15564
rect 5448 15512 5500 15564
rect 7656 15512 7708 15564
rect 8760 15512 8812 15564
rect 10508 15512 10560 15564
rect 2780 15376 2832 15428
rect 3792 15444 3844 15496
rect 4068 15444 4120 15496
rect 4620 15487 4672 15496
rect 4620 15453 4629 15487
rect 4629 15453 4663 15487
rect 4663 15453 4672 15487
rect 4620 15444 4672 15453
rect 4712 15487 4764 15496
rect 4712 15453 4721 15487
rect 4721 15453 4755 15487
rect 4755 15453 4764 15487
rect 4712 15444 4764 15453
rect 4896 15444 4948 15496
rect 7196 15487 7248 15496
rect 5448 15376 5500 15428
rect 6828 15376 6880 15428
rect 7196 15453 7205 15487
rect 7205 15453 7239 15487
rect 7239 15453 7248 15487
rect 7196 15444 7248 15453
rect 8116 15444 8168 15496
rect 7840 15376 7892 15428
rect 8024 15376 8076 15428
rect 9404 15444 9456 15496
rect 9680 15444 9732 15496
rect 10324 15444 10376 15496
rect 10692 15444 10744 15496
rect 9128 15376 9180 15428
rect 10508 15376 10560 15428
rect 11336 15444 11388 15496
rect 3148 15308 3200 15360
rect 4068 15308 4120 15360
rect 5356 15351 5408 15360
rect 5356 15317 5365 15351
rect 5365 15317 5399 15351
rect 5399 15317 5408 15351
rect 5356 15308 5408 15317
rect 5540 15308 5592 15360
rect 7380 15308 7432 15360
rect 7932 15308 7984 15360
rect 8944 15308 8996 15360
rect 9680 15308 9732 15360
rect 10048 15308 10100 15360
rect 11980 15444 12032 15496
rect 12348 15444 12400 15496
rect 12624 15444 12676 15496
rect 13084 15512 13136 15564
rect 15016 15512 15068 15564
rect 13176 15444 13228 15496
rect 13728 15444 13780 15496
rect 15476 15444 15528 15496
rect 11796 15376 11848 15428
rect 11980 15308 12032 15360
rect 13728 15308 13780 15360
rect 14372 15308 14424 15360
rect 3447 15206 3499 15258
rect 3511 15206 3563 15258
rect 3575 15206 3627 15258
rect 3639 15206 3691 15258
rect 8378 15206 8430 15258
rect 8442 15206 8494 15258
rect 8506 15206 8558 15258
rect 8570 15206 8622 15258
rect 13308 15206 13360 15258
rect 13372 15206 13424 15258
rect 13436 15206 13488 15258
rect 13500 15206 13552 15258
rect 3792 15104 3844 15156
rect 4344 15104 4396 15156
rect 5264 15104 5316 15156
rect 5448 15104 5500 15156
rect 5632 15104 5684 15156
rect 7932 15104 7984 15156
rect 13176 15104 13228 15156
rect 2780 15036 2832 15088
rect 5356 15036 5408 15088
rect 3240 14968 3292 15020
rect 4712 14968 4764 15020
rect 13912 15104 13964 15156
rect 8668 15079 8720 15088
rect 8668 15045 8677 15079
rect 8677 15045 8711 15079
rect 8711 15045 8720 15079
rect 8668 15036 8720 15045
rect 13268 15036 13320 15088
rect 13820 15036 13872 15088
rect 2964 14900 3016 14952
rect 5540 14900 5592 14952
rect 5632 14900 5684 14952
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 2780 14832 2832 14884
rect 1952 14807 2004 14816
rect 1952 14773 1961 14807
rect 1961 14773 1995 14807
rect 1995 14773 2004 14807
rect 1952 14764 2004 14773
rect 2320 14807 2372 14816
rect 2320 14773 2329 14807
rect 2329 14773 2363 14807
rect 2363 14773 2372 14807
rect 2320 14764 2372 14773
rect 3240 14764 3292 14816
rect 4436 14832 4488 14884
rect 5080 14832 5132 14884
rect 5264 14832 5316 14884
rect 8576 14900 8628 14952
rect 9312 14968 9364 15020
rect 9588 14968 9640 15020
rect 12716 14968 12768 15020
rect 12808 14968 12860 15020
rect 9496 14900 9548 14952
rect 9772 14900 9824 14952
rect 11796 14900 11848 14952
rect 15384 14968 15436 15020
rect 7196 14832 7248 14884
rect 7564 14832 7616 14884
rect 8668 14832 8720 14884
rect 10876 14832 10928 14884
rect 11980 14832 12032 14884
rect 12256 14832 12308 14884
rect 4344 14807 4396 14816
rect 4344 14773 4353 14807
rect 4353 14773 4387 14807
rect 4387 14773 4396 14807
rect 4344 14764 4396 14773
rect 5816 14764 5868 14816
rect 6276 14764 6328 14816
rect 6368 14764 6420 14816
rect 8944 14764 8996 14816
rect 10324 14764 10376 14816
rect 11152 14764 11204 14816
rect 12164 14764 12216 14816
rect 14004 14900 14056 14952
rect 14372 14943 14424 14952
rect 14372 14909 14381 14943
rect 14381 14909 14415 14943
rect 14415 14909 14424 14943
rect 14372 14900 14424 14909
rect 14832 14832 14884 14884
rect 16396 14832 16448 14884
rect 12808 14807 12860 14816
rect 12808 14773 12817 14807
rect 12817 14773 12851 14807
rect 12851 14773 12860 14807
rect 12808 14764 12860 14773
rect 13820 14807 13872 14816
rect 13820 14773 13829 14807
rect 13829 14773 13863 14807
rect 13863 14773 13872 14807
rect 13820 14764 13872 14773
rect 5912 14662 5964 14714
rect 5976 14662 6028 14714
rect 6040 14662 6092 14714
rect 6104 14662 6156 14714
rect 10843 14662 10895 14714
rect 10907 14662 10959 14714
rect 10971 14662 11023 14714
rect 11035 14662 11087 14714
rect 1584 14603 1636 14612
rect 1584 14569 1593 14603
rect 1593 14569 1627 14603
rect 1627 14569 1636 14603
rect 1584 14560 1636 14569
rect 4804 14560 4856 14612
rect 2688 14492 2740 14544
rect 4436 14492 4488 14544
rect 4620 14492 4672 14544
rect 5724 14560 5776 14612
rect 5816 14560 5868 14612
rect 7932 14560 7984 14612
rect 8116 14560 8168 14612
rect 5908 14492 5960 14544
rect 2964 14424 3016 14476
rect 4252 14424 4304 14476
rect 2596 14356 2648 14408
rect 3056 14356 3108 14408
rect 4436 14356 4488 14408
rect 5080 14424 5132 14476
rect 5724 14424 5776 14476
rect 9312 14492 9364 14544
rect 11152 14560 11204 14612
rect 13176 14560 13228 14612
rect 9864 14492 9916 14544
rect 10508 14492 10560 14544
rect 7104 14467 7156 14476
rect 7104 14433 7138 14467
rect 7138 14433 7156 14467
rect 7104 14424 7156 14433
rect 7932 14424 7984 14476
rect 6828 14399 6880 14408
rect 6828 14365 6837 14399
rect 6837 14365 6871 14399
rect 6871 14365 6880 14399
rect 6828 14356 6880 14365
rect 8484 14356 8536 14408
rect 5632 14288 5684 14340
rect 6460 14288 6512 14340
rect 8116 14288 8168 14340
rect 9220 14288 9272 14340
rect 10140 14424 10192 14476
rect 10600 14424 10652 14476
rect 11060 14424 11112 14476
rect 11152 14424 11204 14476
rect 13268 14492 13320 14544
rect 13728 14535 13780 14544
rect 13728 14501 13737 14535
rect 13737 14501 13771 14535
rect 13771 14501 13780 14535
rect 13728 14492 13780 14501
rect 12072 14424 12124 14476
rect 12256 14424 12308 14476
rect 12440 14467 12492 14476
rect 12440 14433 12449 14467
rect 12449 14433 12483 14467
rect 12483 14433 12492 14467
rect 12440 14424 12492 14433
rect 13636 14467 13688 14476
rect 13636 14433 13645 14467
rect 13645 14433 13679 14467
rect 13679 14433 13688 14467
rect 13636 14424 13688 14433
rect 15292 14424 15344 14476
rect 5080 14220 5132 14272
rect 5816 14220 5868 14272
rect 7564 14220 7616 14272
rect 8024 14220 8076 14272
rect 9128 14220 9180 14272
rect 9496 14288 9548 14340
rect 10140 14288 10192 14340
rect 10416 14288 10468 14340
rect 10508 14220 10560 14272
rect 10692 14288 10744 14340
rect 12992 14356 13044 14408
rect 10968 14220 11020 14272
rect 13176 14220 13228 14272
rect 3447 14118 3499 14170
rect 3511 14118 3563 14170
rect 3575 14118 3627 14170
rect 3639 14118 3691 14170
rect 8378 14118 8430 14170
rect 8442 14118 8494 14170
rect 8506 14118 8558 14170
rect 8570 14118 8622 14170
rect 13308 14118 13360 14170
rect 13372 14118 13424 14170
rect 13436 14118 13488 14170
rect 13500 14118 13552 14170
rect 2412 14016 2464 14068
rect 4252 14016 4304 14068
rect 4528 13948 4580 14000
rect 8852 14016 8904 14068
rect 10232 14016 10284 14068
rect 12440 14059 12492 14068
rect 12440 14025 12449 14059
rect 12449 14025 12483 14059
rect 12483 14025 12492 14059
rect 12440 14016 12492 14025
rect 10692 13948 10744 14000
rect 12808 13948 12860 14000
rect 13452 13948 13504 14000
rect 15568 13948 15620 14000
rect 3424 13880 3476 13932
rect 4252 13923 4304 13932
rect 4252 13889 4261 13923
rect 4261 13889 4295 13923
rect 4295 13889 4304 13923
rect 4252 13880 4304 13889
rect 7472 13880 7524 13932
rect 1492 13812 1544 13864
rect 2228 13812 2280 13864
rect 572 13744 624 13796
rect 4804 13812 4856 13864
rect 4988 13812 5040 13864
rect 6276 13812 6328 13864
rect 7104 13812 7156 13864
rect 12716 13880 12768 13932
rect 13360 13880 13412 13932
rect 13636 13880 13688 13932
rect 14096 13923 14148 13932
rect 14096 13889 14105 13923
rect 14105 13889 14139 13923
rect 14139 13889 14148 13923
rect 14096 13880 14148 13889
rect 4160 13787 4212 13796
rect 4160 13753 4169 13787
rect 4169 13753 4203 13787
rect 4203 13753 4212 13787
rect 4160 13744 4212 13753
rect 2504 13676 2556 13728
rect 3884 13676 3936 13728
rect 6276 13719 6328 13728
rect 6276 13685 6285 13719
rect 6285 13685 6319 13719
rect 6319 13685 6328 13719
rect 6276 13676 6328 13685
rect 6828 13744 6880 13796
rect 9036 13812 9088 13864
rect 8760 13744 8812 13796
rect 8852 13744 8904 13796
rect 7104 13676 7156 13728
rect 7748 13676 7800 13728
rect 7932 13676 7984 13728
rect 10140 13812 10192 13864
rect 10784 13812 10836 13864
rect 10048 13744 10100 13796
rect 11060 13744 11112 13796
rect 12164 13744 12216 13796
rect 12624 13744 12676 13796
rect 9588 13676 9640 13728
rect 9680 13676 9732 13728
rect 10232 13676 10284 13728
rect 10600 13676 10652 13728
rect 11336 13676 11388 13728
rect 11888 13676 11940 13728
rect 12808 13719 12860 13728
rect 12808 13685 12817 13719
rect 12817 13685 12851 13719
rect 12851 13685 12860 13719
rect 12808 13676 12860 13685
rect 13452 13676 13504 13728
rect 14004 13676 14056 13728
rect 5912 13574 5964 13626
rect 5976 13574 6028 13626
rect 6040 13574 6092 13626
rect 6104 13574 6156 13626
rect 10843 13574 10895 13626
rect 10907 13574 10959 13626
rect 10971 13574 11023 13626
rect 11035 13574 11087 13626
rect 2780 13515 2832 13524
rect 2780 13481 2789 13515
rect 2789 13481 2823 13515
rect 2823 13481 2832 13515
rect 2780 13472 2832 13481
rect 2596 13404 2648 13456
rect 6368 13472 6420 13524
rect 7196 13515 7248 13524
rect 7196 13481 7205 13515
rect 7205 13481 7239 13515
rect 7239 13481 7248 13515
rect 7196 13472 7248 13481
rect 7656 13515 7708 13524
rect 7656 13481 7665 13515
rect 7665 13481 7699 13515
rect 7699 13481 7708 13515
rect 7656 13472 7708 13481
rect 3792 13404 3844 13456
rect 1584 13243 1636 13252
rect 1584 13209 1593 13243
rect 1593 13209 1627 13243
rect 1627 13209 1636 13243
rect 1584 13200 1636 13209
rect 2964 13336 3016 13388
rect 2596 13200 2648 13252
rect 6276 13404 6328 13456
rect 7564 13404 7616 13456
rect 8576 13404 8628 13456
rect 9312 13404 9364 13456
rect 10048 13404 10100 13456
rect 10232 13472 10284 13524
rect 12808 13472 12860 13524
rect 5448 13336 5500 13388
rect 6368 13336 6420 13388
rect 6644 13336 6696 13388
rect 7288 13336 7340 13388
rect 8116 13336 8168 13388
rect 9496 13336 9548 13388
rect 12716 13404 12768 13456
rect 13268 13404 13320 13456
rect 13544 13404 13596 13456
rect 14004 13404 14056 13456
rect 10876 13336 10928 13388
rect 11888 13379 11940 13388
rect 4252 13311 4304 13320
rect 4252 13277 4261 13311
rect 4261 13277 4295 13311
rect 4295 13277 4304 13311
rect 4252 13268 4304 13277
rect 5080 13268 5132 13320
rect 4528 13200 4580 13252
rect 4804 13200 4856 13252
rect 4988 13200 5040 13252
rect 7748 13268 7800 13320
rect 8760 13268 8812 13320
rect 9036 13268 9088 13320
rect 2228 13132 2280 13184
rect 8116 13200 8168 13252
rect 8392 13200 8444 13252
rect 11244 13268 11296 13320
rect 10784 13200 10836 13252
rect 7012 13132 7064 13184
rect 7656 13132 7708 13184
rect 10876 13132 10928 13184
rect 11244 13132 11296 13184
rect 11888 13345 11897 13379
rect 11897 13345 11931 13379
rect 11931 13345 11940 13379
rect 11888 13336 11940 13345
rect 12992 13336 13044 13388
rect 11980 13311 12032 13320
rect 11980 13277 11989 13311
rect 11989 13277 12023 13311
rect 12023 13277 12032 13311
rect 11980 13268 12032 13277
rect 12164 13268 12216 13320
rect 13084 13268 13136 13320
rect 13912 13336 13964 13388
rect 12992 13200 13044 13252
rect 13084 13132 13136 13184
rect 3447 13030 3499 13082
rect 3511 13030 3563 13082
rect 3575 13030 3627 13082
rect 3639 13030 3691 13082
rect 8378 13030 8430 13082
rect 8442 13030 8494 13082
rect 8506 13030 8558 13082
rect 8570 13030 8622 13082
rect 13308 13030 13360 13082
rect 13372 13030 13424 13082
rect 13436 13030 13488 13082
rect 13500 13030 13552 13082
rect 3056 12928 3108 12980
rect 4436 12971 4488 12980
rect 4436 12937 4445 12971
rect 4445 12937 4479 12971
rect 4479 12937 4488 12971
rect 4436 12928 4488 12937
rect 4528 12928 4580 12980
rect 1492 12656 1544 12708
rect 4804 12724 4856 12776
rect 7104 12928 7156 12980
rect 8116 12928 8168 12980
rect 8668 12928 8720 12980
rect 10232 12928 10284 12980
rect 10876 12928 10928 12980
rect 11980 12928 12032 12980
rect 12716 12928 12768 12980
rect 13820 12928 13872 12980
rect 6828 12792 6880 12844
rect 8300 12792 8352 12844
rect 10232 12724 10284 12776
rect 10876 12792 10928 12844
rect 11428 12792 11480 12844
rect 11796 12903 11848 12912
rect 11796 12869 11805 12903
rect 11805 12869 11839 12903
rect 11839 12869 11848 12903
rect 11796 12860 11848 12869
rect 13268 12860 13320 12912
rect 14740 12860 14792 12912
rect 12992 12835 13044 12844
rect 12992 12801 13001 12835
rect 13001 12801 13035 12835
rect 13035 12801 13044 12835
rect 12992 12792 13044 12801
rect 13636 12792 13688 12844
rect 10784 12724 10836 12776
rect 11796 12724 11848 12776
rect 7012 12656 7064 12708
rect 4344 12588 4396 12640
rect 5632 12588 5684 12640
rect 8760 12656 8812 12708
rect 9220 12699 9272 12708
rect 9220 12665 9229 12699
rect 9229 12665 9263 12699
rect 9263 12665 9272 12699
rect 9220 12656 9272 12665
rect 7380 12588 7432 12640
rect 8852 12588 8904 12640
rect 10416 12656 10468 12708
rect 10600 12656 10652 12708
rect 10140 12588 10192 12640
rect 10232 12588 10284 12640
rect 11612 12656 11664 12708
rect 12164 12656 12216 12708
rect 12716 12588 12768 12640
rect 13084 12588 13136 12640
rect 14004 12631 14056 12640
rect 14004 12597 14013 12631
rect 14013 12597 14047 12631
rect 14047 12597 14056 12631
rect 14004 12588 14056 12597
rect 5912 12486 5964 12538
rect 5976 12486 6028 12538
rect 6040 12486 6092 12538
rect 6104 12486 6156 12538
rect 10843 12486 10895 12538
rect 10907 12486 10959 12538
rect 10971 12486 11023 12538
rect 11035 12486 11087 12538
rect 1584 12384 1636 12436
rect 4896 12384 4948 12436
rect 5632 12384 5684 12436
rect 6460 12384 6512 12436
rect 6644 12384 6696 12436
rect 7104 12384 7156 12436
rect 2688 12316 2740 12368
rect 4160 12316 4212 12368
rect 5356 12316 5408 12368
rect 6552 12316 6604 12368
rect 7472 12359 7524 12368
rect 7472 12325 7481 12359
rect 7481 12325 7515 12359
rect 7515 12325 7524 12359
rect 7472 12316 7524 12325
rect 8760 12384 8812 12436
rect 9312 12384 9364 12436
rect 9588 12384 9640 12436
rect 2780 12248 2832 12300
rect 7196 12248 7248 12300
rect 8024 12248 8076 12300
rect 8668 12316 8720 12368
rect 9864 12316 9916 12368
rect 10692 12384 10744 12436
rect 11612 12316 11664 12368
rect 12348 12384 12400 12436
rect 13176 12384 13228 12436
rect 14464 12384 14516 12436
rect 14740 12384 14792 12436
rect 15108 12384 15160 12436
rect 15292 12316 15344 12368
rect 10416 12248 10468 12300
rect 11152 12248 11204 12300
rect 12164 12248 12216 12300
rect 12440 12291 12492 12300
rect 12440 12257 12449 12291
rect 12449 12257 12483 12291
rect 12483 12257 12492 12291
rect 12440 12248 12492 12257
rect 2136 12223 2188 12232
rect 2136 12189 2145 12223
rect 2145 12189 2179 12223
rect 2179 12189 2188 12223
rect 2136 12180 2188 12189
rect 4896 12180 4948 12232
rect 5356 12223 5408 12232
rect 5356 12189 5365 12223
rect 5365 12189 5399 12223
rect 5399 12189 5408 12223
rect 5356 12180 5408 12189
rect 5724 12180 5776 12232
rect 6460 12180 6512 12232
rect 6644 12180 6696 12232
rect 6920 12180 6972 12232
rect 8852 12180 8904 12232
rect 9496 12180 9548 12232
rect 9680 12180 9732 12232
rect 10140 12180 10192 12232
rect 4344 12112 4396 12164
rect 6736 12112 6788 12164
rect 7840 12112 7892 12164
rect 3792 12044 3844 12096
rect 9036 12112 9088 12164
rect 9312 12112 9364 12164
rect 13268 12248 13320 12300
rect 13728 12291 13780 12300
rect 13728 12257 13737 12291
rect 13737 12257 13771 12291
rect 13771 12257 13780 12291
rect 13728 12248 13780 12257
rect 14740 12248 14792 12300
rect 14924 12248 14976 12300
rect 10508 12112 10560 12164
rect 8024 12044 8076 12096
rect 13820 12223 13872 12232
rect 12440 12112 12492 12164
rect 13820 12189 13829 12223
rect 13829 12189 13863 12223
rect 13863 12189 13872 12223
rect 13820 12180 13872 12189
rect 13728 12112 13780 12164
rect 13912 12112 13964 12164
rect 12348 12044 12400 12096
rect 12532 12044 12584 12096
rect 14004 12044 14056 12096
rect 3447 11942 3499 11994
rect 3511 11942 3563 11994
rect 3575 11942 3627 11994
rect 3639 11942 3691 11994
rect 8378 11942 8430 11994
rect 8442 11942 8494 11994
rect 8506 11942 8558 11994
rect 8570 11942 8622 11994
rect 13308 11942 13360 11994
rect 13372 11942 13424 11994
rect 13436 11942 13488 11994
rect 13500 11942 13552 11994
rect 2780 11772 2832 11824
rect 3332 11840 3384 11892
rect 7564 11840 7616 11892
rect 7840 11840 7892 11892
rect 10048 11883 10100 11892
rect 2964 11704 3016 11756
rect 6368 11772 6420 11824
rect 2320 11679 2372 11688
rect 2320 11645 2329 11679
rect 2329 11645 2363 11679
rect 2363 11645 2372 11679
rect 2320 11636 2372 11645
rect 4068 11636 4120 11688
rect 2412 11568 2464 11620
rect 4528 11704 4580 11756
rect 4804 11704 4856 11756
rect 6644 11704 6696 11756
rect 6828 11747 6880 11756
rect 6828 11713 6837 11747
rect 6837 11713 6871 11747
rect 6871 11713 6880 11747
rect 6828 11704 6880 11713
rect 8484 11772 8536 11824
rect 10048 11849 10057 11883
rect 10057 11849 10091 11883
rect 10091 11849 10100 11883
rect 10048 11840 10100 11849
rect 11152 11840 11204 11892
rect 11244 11840 11296 11892
rect 11980 11840 12032 11892
rect 13084 11840 13136 11892
rect 10508 11815 10560 11824
rect 10508 11781 10517 11815
rect 10517 11781 10551 11815
rect 10551 11781 10560 11815
rect 10508 11772 10560 11781
rect 10968 11772 11020 11824
rect 1584 11500 1636 11552
rect 6276 11636 6328 11688
rect 8116 11636 8168 11688
rect 8484 11636 8536 11688
rect 9680 11704 9732 11756
rect 11152 11704 11204 11756
rect 12992 11747 13044 11756
rect 12992 11713 13001 11747
rect 13001 11713 13035 11747
rect 13035 11713 13044 11747
rect 12992 11704 13044 11713
rect 8944 11679 8996 11688
rect 8944 11645 8967 11679
rect 8967 11645 8996 11679
rect 4804 11568 4856 11620
rect 5172 11611 5224 11620
rect 5172 11577 5184 11611
rect 5184 11577 5224 11611
rect 5172 11568 5224 11577
rect 7932 11568 7984 11620
rect 8944 11636 8996 11645
rect 10232 11636 10284 11688
rect 9588 11568 9640 11620
rect 10324 11568 10376 11620
rect 10876 11611 10928 11620
rect 10876 11577 10885 11611
rect 10885 11577 10919 11611
rect 10919 11577 10928 11611
rect 10876 11568 10928 11577
rect 11428 11636 11480 11688
rect 14004 11679 14056 11688
rect 14004 11645 14013 11679
rect 14013 11645 14047 11679
rect 14047 11645 14056 11679
rect 14004 11636 14056 11645
rect 14832 11679 14884 11688
rect 14832 11645 14841 11679
rect 14841 11645 14875 11679
rect 14875 11645 14884 11679
rect 14832 11636 14884 11645
rect 14372 11568 14424 11620
rect 8116 11500 8168 11552
rect 9680 11500 9732 11552
rect 11244 11500 11296 11552
rect 12624 11500 12676 11552
rect 13176 11500 13228 11552
rect 13636 11543 13688 11552
rect 13636 11509 13645 11543
rect 13645 11509 13679 11543
rect 13679 11509 13688 11543
rect 13636 11500 13688 11509
rect 14096 11543 14148 11552
rect 14096 11509 14105 11543
rect 14105 11509 14139 11543
rect 14139 11509 14148 11543
rect 14096 11500 14148 11509
rect 14464 11500 14516 11552
rect 5912 11398 5964 11450
rect 5976 11398 6028 11450
rect 6040 11398 6092 11450
rect 6104 11398 6156 11450
rect 10843 11398 10895 11450
rect 10907 11398 10959 11450
rect 10971 11398 11023 11450
rect 11035 11398 11087 11450
rect 1860 11271 1912 11280
rect 1860 11237 1869 11271
rect 1869 11237 1903 11271
rect 1903 11237 1912 11271
rect 1860 11228 1912 11237
rect 2780 11228 2832 11280
rect 2412 11203 2464 11212
rect 2412 11169 2446 11203
rect 2446 11169 2464 11203
rect 2412 11160 2464 11169
rect 2964 11160 3016 11212
rect 4436 11228 4488 11280
rect 5264 11296 5316 11348
rect 5448 11339 5500 11348
rect 5448 11305 5457 11339
rect 5457 11305 5491 11339
rect 5491 11305 5500 11339
rect 5448 11296 5500 11305
rect 5816 11296 5868 11348
rect 7656 11296 7708 11348
rect 8024 11296 8076 11348
rect 8760 11296 8812 11348
rect 6000 11228 6052 11280
rect 3700 11160 3752 11212
rect 4620 11160 4672 11212
rect 6736 11228 6788 11280
rect 8300 11228 8352 11280
rect 11796 11296 11848 11348
rect 12348 11296 12400 11348
rect 12900 11296 12952 11348
rect 14096 11296 14148 11348
rect 14372 11339 14424 11348
rect 14372 11305 14381 11339
rect 14381 11305 14415 11339
rect 14415 11305 14424 11339
rect 14372 11296 14424 11305
rect 9220 11228 9272 11280
rect 9680 11228 9732 11280
rect 8668 11160 8720 11212
rect 10048 11228 10100 11280
rect 10968 11228 11020 11280
rect 11060 11228 11112 11280
rect 15200 11228 15252 11280
rect 4068 11135 4120 11144
rect 4068 11101 4077 11135
rect 4077 11101 4111 11135
rect 4111 11101 4120 11135
rect 4068 11092 4120 11101
rect 6368 11135 6420 11144
rect 6368 11101 6377 11135
rect 6377 11101 6411 11135
rect 6411 11101 6420 11135
rect 6368 11092 6420 11101
rect 7472 11092 7524 11144
rect 10416 11160 10468 11212
rect 12440 11160 12492 11212
rect 13084 11160 13136 11212
rect 14280 11203 14332 11212
rect 14280 11169 14289 11203
rect 14289 11169 14323 11203
rect 14323 11169 14332 11203
rect 14280 11160 14332 11169
rect 14372 11160 14424 11212
rect 9588 11092 9640 11144
rect 10968 11092 11020 11144
rect 12348 11092 12400 11144
rect 3332 11024 3384 11076
rect 5080 11024 5132 11076
rect 5356 11024 5408 11076
rect 3976 10956 4028 11008
rect 5172 10956 5224 11008
rect 5448 10956 5500 11008
rect 8024 10956 8076 11008
rect 9220 10956 9272 11008
rect 13820 11024 13872 11076
rect 10968 10956 11020 11008
rect 11152 10956 11204 11008
rect 11796 10956 11848 11008
rect 13728 10956 13780 11008
rect 14556 10956 14608 11008
rect 3447 10854 3499 10906
rect 3511 10854 3563 10906
rect 3575 10854 3627 10906
rect 3639 10854 3691 10906
rect 8378 10854 8430 10906
rect 8442 10854 8494 10906
rect 8506 10854 8558 10906
rect 8570 10854 8622 10906
rect 13308 10854 13360 10906
rect 13372 10854 13424 10906
rect 13436 10854 13488 10906
rect 13500 10854 13552 10906
rect 1676 10752 1728 10804
rect 2136 10752 2188 10804
rect 2964 10752 3016 10804
rect 5172 10752 5224 10804
rect 5540 10752 5592 10804
rect 6276 10795 6328 10804
rect 6276 10761 6285 10795
rect 6285 10761 6319 10795
rect 6319 10761 6328 10795
rect 6276 10752 6328 10761
rect 6368 10752 6420 10804
rect 12992 10752 13044 10804
rect 4528 10684 4580 10736
rect 7840 10684 7892 10736
rect 9680 10684 9732 10736
rect 10508 10684 10560 10736
rect 12072 10684 12124 10736
rect 2504 10659 2556 10668
rect 2504 10625 2513 10659
rect 2513 10625 2547 10659
rect 2547 10625 2556 10659
rect 2504 10616 2556 10625
rect 2780 10616 2832 10668
rect 4068 10616 4120 10668
rect 6828 10659 6880 10668
rect 6828 10625 6837 10659
rect 6837 10625 6871 10659
rect 6871 10625 6880 10659
rect 6828 10616 6880 10625
rect 7932 10616 7984 10668
rect 11612 10616 11664 10668
rect 11980 10616 12032 10668
rect 1676 10548 1728 10600
rect 8208 10548 8260 10600
rect 10324 10548 10376 10600
rect 12992 10659 13044 10668
rect 12992 10625 13001 10659
rect 13001 10625 13035 10659
rect 13035 10625 13044 10659
rect 12992 10616 13044 10625
rect 13084 10616 13136 10668
rect 13360 10616 13412 10668
rect 13820 10616 13872 10668
rect 5264 10480 5316 10532
rect 5356 10480 5408 10532
rect 2320 10455 2372 10464
rect 2320 10421 2329 10455
rect 2329 10421 2363 10455
rect 2363 10421 2372 10455
rect 2320 10412 2372 10421
rect 4436 10412 4488 10464
rect 6368 10412 6420 10464
rect 7380 10480 7432 10532
rect 9772 10480 9824 10532
rect 10600 10480 10652 10532
rect 9220 10412 9272 10464
rect 12900 10548 12952 10600
rect 14280 10548 14332 10600
rect 15936 10548 15988 10600
rect 10784 10523 10836 10532
rect 10784 10489 10818 10523
rect 10818 10489 10836 10523
rect 10784 10480 10836 10489
rect 12348 10480 12400 10532
rect 13268 10480 13320 10532
rect 13360 10480 13412 10532
rect 12440 10455 12492 10464
rect 12440 10421 12449 10455
rect 12449 10421 12483 10455
rect 12483 10421 12492 10455
rect 12900 10455 12952 10464
rect 12440 10412 12492 10421
rect 12900 10421 12909 10455
rect 12909 10421 12943 10455
rect 12943 10421 12952 10455
rect 12900 10412 12952 10421
rect 13912 10412 13964 10464
rect 5912 10310 5964 10362
rect 5976 10310 6028 10362
rect 6040 10310 6092 10362
rect 6104 10310 6156 10362
rect 10843 10310 10895 10362
rect 10907 10310 10959 10362
rect 10971 10310 11023 10362
rect 11035 10310 11087 10362
rect 4528 10208 4580 10260
rect 5448 10251 5500 10260
rect 5448 10217 5457 10251
rect 5457 10217 5491 10251
rect 5491 10217 5500 10251
rect 5448 10208 5500 10217
rect 2504 10140 2556 10192
rect 2688 10140 2740 10192
rect 10508 10208 10560 10260
rect 10692 10208 10744 10260
rect 6276 10140 6328 10192
rect 8116 10140 8168 10192
rect 8668 10140 8720 10192
rect 12164 10208 12216 10260
rect 12348 10208 12400 10260
rect 12440 10208 12492 10260
rect 14004 10208 14056 10260
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 2780 10072 2832 10124
rect 5080 10072 5132 10124
rect 4068 10047 4120 10056
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 3792 9868 3844 9920
rect 10508 10072 10560 10124
rect 5908 10047 5960 10056
rect 5908 10013 5917 10047
rect 5917 10013 5951 10047
rect 5951 10013 5960 10047
rect 5908 10004 5960 10013
rect 7748 10047 7800 10056
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 9588 10004 9640 10056
rect 7104 9936 7156 9988
rect 5908 9868 5960 9920
rect 9312 9936 9364 9988
rect 10784 10072 10836 10124
rect 14372 10140 14424 10192
rect 12256 10072 12308 10124
rect 12440 10072 12492 10124
rect 13084 10115 13136 10124
rect 13084 10081 13093 10115
rect 13093 10081 13127 10115
rect 13127 10081 13136 10115
rect 13084 10072 13136 10081
rect 14004 10072 14056 10124
rect 12164 10047 12216 10056
rect 12164 10013 12173 10047
rect 12173 10013 12207 10047
rect 12207 10013 12216 10047
rect 12164 10004 12216 10013
rect 14372 10047 14424 10056
rect 10600 9868 10652 9920
rect 10784 9868 10836 9920
rect 11244 9868 11296 9920
rect 14372 10013 14381 10047
rect 14381 10013 14415 10047
rect 14415 10013 14424 10047
rect 14372 10004 14424 10013
rect 14188 9936 14240 9988
rect 3447 9766 3499 9818
rect 3511 9766 3563 9818
rect 3575 9766 3627 9818
rect 3639 9766 3691 9818
rect 8378 9766 8430 9818
rect 8442 9766 8494 9818
rect 8506 9766 8558 9818
rect 8570 9766 8622 9818
rect 13308 9766 13360 9818
rect 13372 9766 13424 9818
rect 13436 9766 13488 9818
rect 13500 9766 13552 9818
rect 2320 9664 2372 9716
rect 2596 9664 2648 9716
rect 2964 9664 3016 9716
rect 2504 9571 2556 9580
rect 2504 9537 2513 9571
rect 2513 9537 2547 9571
rect 2547 9537 2556 9571
rect 2504 9528 2556 9537
rect 4068 9664 4120 9716
rect 4436 9639 4488 9648
rect 4436 9605 4445 9639
rect 4445 9605 4479 9639
rect 4479 9605 4488 9639
rect 4436 9596 4488 9605
rect 5908 9664 5960 9716
rect 6000 9664 6052 9716
rect 8116 9664 8168 9716
rect 6276 9596 6328 9648
rect 8668 9596 8720 9648
rect 8208 9528 8260 9580
rect 10232 9596 10284 9648
rect 13084 9664 13136 9716
rect 14004 9596 14056 9648
rect 12992 9571 13044 9580
rect 3608 9460 3660 9512
rect 2964 9392 3016 9444
rect 8576 9460 8628 9512
rect 9128 9460 9180 9512
rect 9588 9460 9640 9512
rect 5540 9435 5592 9444
rect 5540 9401 5574 9435
rect 5574 9401 5592 9435
rect 5540 9392 5592 9401
rect 5816 9392 5868 9444
rect 6276 9392 6328 9444
rect 7196 9435 7248 9444
rect 4896 9367 4948 9376
rect 4896 9333 4905 9367
rect 4905 9333 4939 9367
rect 4939 9333 4948 9367
rect 4896 9324 4948 9333
rect 6920 9324 6972 9376
rect 7196 9401 7205 9435
rect 7205 9401 7239 9435
rect 7239 9401 7248 9435
rect 7196 9392 7248 9401
rect 8760 9435 8812 9444
rect 8760 9401 8769 9435
rect 8769 9401 8803 9435
rect 8803 9401 8812 9435
rect 8760 9392 8812 9401
rect 12072 9460 12124 9512
rect 12992 9537 13001 9571
rect 13001 9537 13035 9571
rect 13035 9537 13044 9571
rect 12992 9528 13044 9537
rect 11152 9392 11204 9444
rect 12164 9392 12216 9444
rect 9128 9324 9180 9376
rect 9588 9324 9640 9376
rect 11612 9324 11664 9376
rect 11888 9367 11940 9376
rect 11888 9333 11897 9367
rect 11897 9333 11931 9367
rect 11931 9333 11940 9367
rect 12624 9460 12676 9512
rect 13452 9460 13504 9512
rect 14280 9392 14332 9444
rect 14096 9367 14148 9376
rect 11888 9324 11940 9333
rect 14096 9333 14105 9367
rect 14105 9333 14139 9367
rect 14139 9333 14148 9367
rect 14096 9324 14148 9333
rect 15016 9367 15068 9376
rect 15016 9333 15025 9367
rect 15025 9333 15059 9367
rect 15059 9333 15068 9367
rect 15016 9324 15068 9333
rect 5912 9222 5964 9274
rect 5976 9222 6028 9274
rect 6040 9222 6092 9274
rect 6104 9222 6156 9274
rect 10843 9222 10895 9274
rect 10907 9222 10959 9274
rect 10971 9222 11023 9274
rect 11035 9222 11087 9274
rect 2964 9120 3016 9172
rect 2504 9052 2556 9104
rect 5816 9052 5868 9104
rect 6000 9095 6052 9104
rect 6000 9061 6034 9095
rect 6034 9061 6052 9095
rect 6000 9052 6052 9061
rect 6276 9052 6328 9104
rect 11888 9052 11940 9104
rect 2044 8984 2096 9036
rect 4160 8984 4212 9036
rect 5448 8984 5500 9036
rect 2136 8959 2188 8968
rect 2136 8925 2145 8959
rect 2145 8925 2179 8959
rect 2179 8925 2188 8959
rect 2136 8916 2188 8925
rect 4068 8916 4120 8968
rect 7288 8984 7340 9036
rect 8852 8984 8904 9036
rect 9036 8984 9088 9036
rect 9220 8984 9272 9036
rect 5724 8848 5776 8900
rect 3792 8780 3844 8832
rect 4896 8780 4948 8832
rect 6460 8780 6512 8832
rect 7288 8780 7340 8832
rect 8576 8916 8628 8968
rect 9588 8916 9640 8968
rect 10232 8984 10284 9036
rect 10508 8984 10560 9036
rect 12256 8984 12308 9036
rect 13544 8984 13596 9036
rect 13636 8984 13688 9036
rect 10968 8916 11020 8968
rect 12532 8916 12584 8968
rect 14464 8916 14516 8968
rect 15568 8916 15620 8968
rect 11244 8848 11296 8900
rect 12716 8848 12768 8900
rect 7840 8780 7892 8832
rect 8208 8780 8260 8832
rect 10324 8780 10376 8832
rect 10600 8780 10652 8832
rect 12440 8780 12492 8832
rect 13084 8780 13136 8832
rect 14004 8780 14056 8832
rect 3447 8678 3499 8730
rect 3511 8678 3563 8730
rect 3575 8678 3627 8730
rect 3639 8678 3691 8730
rect 8378 8678 8430 8730
rect 8442 8678 8494 8730
rect 8506 8678 8558 8730
rect 8570 8678 8622 8730
rect 13308 8678 13360 8730
rect 13372 8678 13424 8730
rect 13436 8678 13488 8730
rect 13500 8678 13552 8730
rect 2964 8576 3016 8628
rect 2136 8508 2188 8560
rect 4068 8576 4120 8628
rect 11152 8576 11204 8628
rect 6000 8508 6052 8560
rect 6276 8551 6328 8560
rect 6276 8517 6285 8551
rect 6285 8517 6319 8551
rect 6319 8517 6328 8551
rect 6276 8508 6328 8517
rect 9680 8508 9732 8560
rect 9864 8508 9916 8560
rect 2688 8415 2740 8424
rect 2688 8381 2697 8415
rect 2697 8381 2731 8415
rect 2731 8381 2740 8415
rect 2688 8372 2740 8381
rect 1768 8347 1820 8356
rect 1768 8313 1777 8347
rect 1777 8313 1811 8347
rect 1811 8313 1820 8347
rect 1768 8304 1820 8313
rect 2320 8304 2372 8356
rect 1032 8236 1084 8288
rect 2228 8236 2280 8288
rect 4068 8440 4120 8492
rect 4896 8483 4948 8492
rect 4896 8449 4905 8483
rect 4905 8449 4939 8483
rect 4939 8449 4948 8483
rect 4896 8440 4948 8449
rect 7840 8440 7892 8492
rect 10048 8440 10100 8492
rect 11888 8619 11940 8628
rect 11888 8585 11897 8619
rect 11897 8585 11931 8619
rect 11931 8585 11940 8619
rect 11888 8576 11940 8585
rect 14096 8576 14148 8628
rect 12348 8508 12400 8560
rect 12624 8508 12676 8560
rect 13820 8508 13872 8560
rect 3332 8415 3384 8424
rect 3332 8381 3366 8415
rect 3366 8381 3384 8415
rect 3332 8372 3384 8381
rect 5540 8372 5592 8424
rect 6736 8372 6788 8424
rect 6920 8372 6972 8424
rect 7932 8372 7984 8424
rect 8668 8415 8720 8424
rect 5172 8347 5224 8356
rect 5172 8313 5206 8347
rect 5206 8313 5224 8347
rect 5172 8304 5224 8313
rect 5816 8304 5868 8356
rect 7288 8304 7340 8356
rect 8668 8381 8677 8415
rect 8677 8381 8711 8415
rect 8711 8381 8720 8415
rect 8668 8372 8720 8381
rect 9220 8372 9272 8424
rect 14464 8508 14516 8560
rect 14188 8483 14240 8492
rect 14188 8449 14197 8483
rect 14197 8449 14231 8483
rect 14231 8449 14240 8483
rect 14188 8440 14240 8449
rect 3332 8236 3384 8288
rect 3792 8236 3844 8288
rect 4160 8236 4212 8288
rect 8208 8279 8260 8288
rect 8208 8245 8217 8279
rect 8217 8245 8251 8279
rect 8251 8245 8260 8279
rect 8208 8236 8260 8245
rect 8392 8236 8444 8288
rect 9864 8236 9916 8288
rect 15108 8372 15160 8424
rect 10692 8304 10744 8356
rect 10968 8304 11020 8356
rect 11336 8304 11388 8356
rect 11152 8236 11204 8288
rect 11612 8236 11664 8288
rect 12072 8304 12124 8356
rect 12716 8304 12768 8356
rect 14464 8304 14516 8356
rect 14004 8279 14056 8288
rect 14004 8245 14013 8279
rect 14013 8245 14047 8279
rect 14047 8245 14056 8279
rect 14004 8236 14056 8245
rect 15016 8279 15068 8288
rect 15016 8245 15025 8279
rect 15025 8245 15059 8279
rect 15059 8245 15068 8279
rect 15016 8236 15068 8245
rect 5912 8134 5964 8186
rect 5976 8134 6028 8186
rect 6040 8134 6092 8186
rect 6104 8134 6156 8186
rect 10843 8134 10895 8186
rect 10907 8134 10959 8186
rect 10971 8134 11023 8186
rect 11035 8134 11087 8186
rect 4160 8032 4212 8084
rect 11612 8032 11664 8084
rect 12532 8032 12584 8084
rect 12716 8075 12768 8084
rect 12716 8041 12725 8075
rect 12725 8041 12759 8075
rect 12759 8041 12768 8075
rect 12716 8032 12768 8041
rect 14004 8032 14056 8084
rect 2688 7964 2740 8016
rect 3056 7964 3108 8016
rect 4068 7964 4120 8016
rect 5172 7964 5224 8016
rect 1952 7896 2004 7948
rect 2136 7939 2188 7948
rect 2136 7905 2145 7939
rect 2145 7905 2179 7939
rect 2179 7905 2188 7939
rect 2136 7896 2188 7905
rect 5540 7896 5592 7948
rect 6828 7896 6880 7948
rect 7380 7896 7432 7948
rect 4252 7828 4304 7880
rect 5264 7760 5316 7812
rect 1492 7692 1544 7744
rect 4528 7735 4580 7744
rect 4528 7701 4537 7735
rect 4537 7701 4571 7735
rect 4571 7701 4580 7735
rect 4528 7692 4580 7701
rect 4620 7692 4672 7744
rect 5448 7871 5500 7880
rect 5448 7837 5457 7871
rect 5457 7837 5491 7871
rect 5491 7837 5500 7871
rect 5448 7828 5500 7837
rect 6736 7828 6788 7880
rect 8392 7964 8444 8016
rect 10416 7964 10468 8016
rect 12348 7964 12400 8016
rect 8760 7896 8812 7948
rect 10324 7896 10376 7948
rect 6092 7692 6144 7744
rect 6184 7692 6236 7744
rect 7564 7692 7616 7744
rect 9220 7828 9272 7880
rect 11060 7828 11112 7880
rect 12532 7828 12584 7880
rect 13728 7896 13780 7948
rect 13820 7828 13872 7880
rect 14832 7896 14884 7948
rect 10784 7760 10836 7812
rect 12348 7760 12400 7812
rect 13084 7760 13136 7812
rect 14188 7760 14240 7812
rect 9128 7735 9180 7744
rect 9128 7701 9137 7735
rect 9137 7701 9171 7735
rect 9171 7701 9180 7735
rect 9128 7692 9180 7701
rect 9220 7692 9272 7744
rect 9496 7692 9548 7744
rect 9864 7692 9916 7744
rect 10692 7692 10744 7744
rect 11612 7692 11664 7744
rect 14004 7692 14056 7744
rect 3447 7590 3499 7642
rect 3511 7590 3563 7642
rect 3575 7590 3627 7642
rect 3639 7590 3691 7642
rect 8378 7590 8430 7642
rect 8442 7590 8494 7642
rect 8506 7590 8558 7642
rect 8570 7590 8622 7642
rect 13308 7590 13360 7642
rect 13372 7590 13424 7642
rect 13436 7590 13488 7642
rect 13500 7590 13552 7642
rect 2964 7420 3016 7472
rect 4620 7488 4672 7540
rect 5172 7488 5224 7540
rect 5264 7488 5316 7540
rect 11612 7488 11664 7540
rect 11796 7488 11848 7540
rect 12256 7488 12308 7540
rect 2136 7284 2188 7336
rect 2504 7216 2556 7268
rect 6828 7420 6880 7472
rect 4252 7352 4304 7404
rect 4620 7352 4672 7404
rect 6092 7352 6144 7404
rect 4988 7284 5040 7336
rect 6000 7284 6052 7336
rect 6736 7284 6788 7336
rect 6184 7216 6236 7268
rect 7012 7216 7064 7268
rect 7656 7284 7708 7336
rect 9772 7420 9824 7472
rect 10232 7420 10284 7472
rect 10876 7420 10928 7472
rect 10968 7420 11020 7472
rect 14372 7488 14424 7540
rect 8300 7352 8352 7404
rect 8668 7327 8720 7336
rect 8668 7293 8677 7327
rect 8677 7293 8711 7327
rect 8711 7293 8720 7327
rect 8668 7284 8720 7293
rect 10784 7352 10836 7404
rect 11060 7395 11112 7404
rect 11060 7361 11069 7395
rect 11069 7361 11103 7395
rect 11103 7361 11112 7395
rect 11060 7352 11112 7361
rect 12256 7352 12308 7404
rect 10140 7284 10192 7336
rect 10876 7327 10928 7336
rect 9312 7216 9364 7268
rect 10876 7293 10885 7327
rect 10885 7293 10919 7327
rect 10919 7293 10928 7327
rect 10876 7284 10928 7293
rect 11336 7284 11388 7336
rect 11612 7284 11664 7336
rect 13912 7352 13964 7404
rect 14188 7352 14240 7404
rect 5264 7148 5316 7200
rect 5816 7148 5868 7200
rect 7196 7148 7248 7200
rect 11704 7216 11756 7268
rect 12900 7284 12952 7336
rect 14648 7284 14700 7336
rect 12256 7148 12308 7200
rect 12624 7148 12676 7200
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 14004 7148 14056 7200
rect 14372 7148 14424 7200
rect 15016 7191 15068 7200
rect 15016 7157 15025 7191
rect 15025 7157 15059 7191
rect 15059 7157 15068 7191
rect 15016 7148 15068 7157
rect 5912 7046 5964 7098
rect 5976 7046 6028 7098
rect 6040 7046 6092 7098
rect 6104 7046 6156 7098
rect 10843 7046 10895 7098
rect 10907 7046 10959 7098
rect 10971 7046 11023 7098
rect 11035 7046 11087 7098
rect 4988 6944 5040 6996
rect 5448 6944 5500 6996
rect 7012 6944 7064 6996
rect 9496 6944 9548 6996
rect 11520 6944 11572 6996
rect 11704 6944 11756 6996
rect 2780 6876 2832 6928
rect 10508 6876 10560 6928
rect 10692 6876 10744 6928
rect 13176 6944 13228 6996
rect 13636 6944 13688 6996
rect 14832 6944 14884 6996
rect 14096 6876 14148 6928
rect 1584 6851 1636 6860
rect 1584 6817 1593 6851
rect 1593 6817 1627 6851
rect 1627 6817 1636 6851
rect 1584 6808 1636 6817
rect 4436 6808 4488 6860
rect 5448 6808 5500 6860
rect 6552 6808 6604 6860
rect 6736 6808 6788 6860
rect 7564 6851 7616 6860
rect 7564 6817 7573 6851
rect 7573 6817 7607 6851
rect 7607 6817 7616 6851
rect 7564 6808 7616 6817
rect 7840 6851 7892 6860
rect 7840 6817 7874 6851
rect 7874 6817 7892 6851
rect 7840 6808 7892 6817
rect 8116 6808 8168 6860
rect 2136 6783 2188 6792
rect 2136 6749 2145 6783
rect 2145 6749 2179 6783
rect 2179 6749 2188 6783
rect 2136 6740 2188 6749
rect 3792 6672 3844 6724
rect 4896 6604 4948 6656
rect 5632 6740 5684 6792
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 10324 6783 10376 6792
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 11152 6808 11204 6860
rect 11336 6851 11388 6860
rect 11336 6817 11345 6851
rect 11345 6817 11379 6851
rect 11379 6817 11388 6851
rect 11336 6808 11388 6817
rect 11704 6808 11756 6860
rect 11888 6808 11940 6860
rect 13636 6851 13688 6860
rect 10324 6740 10376 6749
rect 12532 6783 12584 6792
rect 12532 6749 12541 6783
rect 12541 6749 12575 6783
rect 12575 6749 12584 6783
rect 12532 6740 12584 6749
rect 13636 6817 13645 6851
rect 13645 6817 13679 6851
rect 13679 6817 13688 6851
rect 13636 6808 13688 6817
rect 13728 6851 13780 6860
rect 13728 6817 13737 6851
rect 13737 6817 13771 6851
rect 13771 6817 13780 6851
rect 13728 6808 13780 6817
rect 14188 6808 14240 6860
rect 6920 6604 6972 6656
rect 8668 6672 8720 6724
rect 8852 6604 8904 6656
rect 9680 6647 9732 6656
rect 9680 6613 9689 6647
rect 9689 6613 9723 6647
rect 9723 6613 9732 6647
rect 9680 6604 9732 6613
rect 10324 6604 10376 6656
rect 10600 6604 10652 6656
rect 10692 6604 10744 6656
rect 11336 6604 11388 6656
rect 12532 6604 12584 6656
rect 14740 6672 14792 6724
rect 13176 6604 13228 6656
rect 3447 6502 3499 6554
rect 3511 6502 3563 6554
rect 3575 6502 3627 6554
rect 3639 6502 3691 6554
rect 8378 6502 8430 6554
rect 8442 6502 8494 6554
rect 8506 6502 8558 6554
rect 8570 6502 8622 6554
rect 13308 6502 13360 6554
rect 13372 6502 13424 6554
rect 13436 6502 13488 6554
rect 13500 6502 13552 6554
rect 1952 6332 2004 6384
rect 2320 6332 2372 6384
rect 1308 6264 1360 6316
rect 2136 6264 2188 6316
rect 5264 6400 5316 6452
rect 5632 6400 5684 6452
rect 6460 6400 6512 6452
rect 10508 6443 10560 6452
rect 10508 6409 10517 6443
rect 10517 6409 10551 6443
rect 10551 6409 10560 6443
rect 10508 6400 10560 6409
rect 10600 6400 10652 6452
rect 10784 6400 10836 6452
rect 13636 6400 13688 6452
rect 9772 6332 9824 6384
rect 12716 6332 12768 6384
rect 13084 6332 13136 6384
rect 5448 6196 5500 6248
rect 5724 6196 5776 6248
rect 6828 6239 6880 6248
rect 6828 6205 6837 6239
rect 6837 6205 6871 6239
rect 6871 6205 6880 6239
rect 6828 6196 6880 6205
rect 8116 6196 8168 6248
rect 2504 6128 2556 6180
rect 3332 6171 3384 6180
rect 3332 6137 3366 6171
rect 3366 6137 3384 6171
rect 3332 6128 3384 6137
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 1860 6103 1912 6112
rect 1860 6069 1869 6103
rect 1869 6069 1903 6103
rect 1903 6069 1912 6103
rect 1860 6060 1912 6069
rect 2228 6103 2280 6112
rect 2228 6069 2237 6103
rect 2237 6069 2271 6103
rect 2271 6069 2280 6103
rect 2228 6060 2280 6069
rect 2320 6103 2372 6112
rect 2320 6069 2329 6103
rect 2329 6069 2363 6103
rect 2363 6069 2372 6103
rect 4436 6103 4488 6112
rect 2320 6060 2372 6069
rect 4436 6069 4445 6103
rect 4445 6069 4479 6103
rect 4479 6069 4488 6103
rect 4436 6060 4488 6069
rect 5724 6060 5776 6112
rect 6920 6128 6972 6180
rect 7564 6128 7616 6180
rect 9220 6196 9272 6248
rect 9496 6196 9548 6248
rect 10140 6196 10192 6248
rect 10508 6264 10560 6316
rect 12164 6264 12216 6316
rect 13268 6264 13320 6316
rect 10692 6196 10744 6248
rect 10968 6239 11020 6248
rect 10968 6205 10977 6239
rect 10977 6205 11011 6239
rect 11011 6205 11020 6239
rect 10968 6196 11020 6205
rect 7380 6060 7432 6112
rect 8208 6103 8260 6112
rect 8208 6069 8217 6103
rect 8217 6069 8251 6103
rect 8251 6069 8260 6103
rect 8208 6060 8260 6069
rect 8760 6060 8812 6112
rect 9404 6128 9456 6180
rect 9956 6060 10008 6112
rect 10692 6060 10744 6112
rect 11980 6128 12032 6180
rect 12348 6060 12400 6112
rect 13728 6128 13780 6180
rect 14188 6128 14240 6180
rect 13636 6103 13688 6112
rect 13636 6069 13645 6103
rect 13645 6069 13679 6103
rect 13679 6069 13688 6103
rect 13636 6060 13688 6069
rect 13820 6060 13872 6112
rect 5912 5958 5964 6010
rect 5976 5958 6028 6010
rect 6040 5958 6092 6010
rect 6104 5958 6156 6010
rect 10843 5958 10895 6010
rect 10907 5958 10959 6010
rect 10971 5958 11023 6010
rect 11035 5958 11087 6010
rect 1860 5856 1912 5908
rect 4896 5899 4948 5908
rect 4436 5788 4488 5840
rect 4896 5865 4905 5899
rect 4905 5865 4939 5899
rect 4939 5865 4948 5899
rect 4896 5856 4948 5865
rect 5448 5856 5500 5908
rect 5724 5856 5776 5908
rect 6092 5788 6144 5840
rect 6552 5856 6604 5908
rect 9680 5788 9732 5840
rect 10232 5856 10284 5908
rect 11980 5856 12032 5908
rect 12348 5856 12400 5908
rect 13452 5856 13504 5908
rect 11336 5831 11388 5840
rect 11336 5797 11345 5831
rect 11345 5797 11379 5831
rect 11379 5797 11388 5831
rect 11336 5788 11388 5797
rect 12532 5788 12584 5840
rect 12716 5788 12768 5840
rect 12992 5788 13044 5840
rect 13544 5788 13596 5840
rect 2780 5652 2832 5704
rect 6828 5720 6880 5772
rect 7564 5720 7616 5772
rect 9772 5720 9824 5772
rect 9956 5720 10008 5772
rect 13268 5720 13320 5772
rect 4068 5652 4120 5704
rect 4988 5695 5040 5704
rect 4988 5661 4997 5695
rect 4997 5661 5031 5695
rect 5031 5661 5040 5695
rect 4988 5652 5040 5661
rect 5540 5652 5592 5704
rect 5724 5695 5776 5704
rect 5724 5661 5733 5695
rect 5733 5661 5767 5695
rect 5767 5661 5776 5695
rect 5724 5652 5776 5661
rect 4436 5516 4488 5568
rect 4896 5516 4948 5568
rect 6736 5584 6788 5636
rect 7012 5516 7064 5568
rect 8852 5584 8904 5636
rect 10232 5652 10284 5704
rect 10508 5652 10560 5704
rect 11612 5652 11664 5704
rect 12532 5695 12584 5704
rect 12532 5661 12541 5695
rect 12541 5661 12575 5695
rect 12575 5661 12584 5695
rect 12532 5652 12584 5661
rect 11336 5584 11388 5636
rect 11888 5584 11940 5636
rect 12164 5584 12216 5636
rect 12808 5652 12860 5704
rect 13176 5584 13228 5636
rect 14556 5720 14608 5772
rect 9128 5516 9180 5568
rect 9404 5516 9456 5568
rect 13728 5516 13780 5568
rect 3447 5414 3499 5466
rect 3511 5414 3563 5466
rect 3575 5414 3627 5466
rect 3639 5414 3691 5466
rect 8378 5414 8430 5466
rect 8442 5414 8494 5466
rect 8506 5414 8558 5466
rect 8570 5414 8622 5466
rect 13308 5414 13360 5466
rect 13372 5414 13424 5466
rect 13436 5414 13488 5466
rect 13500 5414 13552 5466
rect 1400 5355 1452 5364
rect 1400 5321 1409 5355
rect 1409 5321 1443 5355
rect 1443 5321 1452 5355
rect 1400 5312 1452 5321
rect 2596 5244 2648 5296
rect 2688 5176 2740 5228
rect 2964 5219 3016 5228
rect 2964 5185 2973 5219
rect 2973 5185 3007 5219
rect 3007 5185 3016 5219
rect 2964 5176 3016 5185
rect 5264 5312 5316 5364
rect 5540 5312 5592 5364
rect 7012 5312 7064 5364
rect 3424 5244 3476 5296
rect 4804 5244 4856 5296
rect 9680 5312 9732 5364
rect 12256 5312 12308 5364
rect 12348 5312 12400 5364
rect 9128 5244 9180 5296
rect 9588 5244 9640 5296
rect 9772 5244 9824 5296
rect 10232 5244 10284 5296
rect 10324 5244 10376 5296
rect 4068 5176 4120 5228
rect 6644 5176 6696 5228
rect 1676 5108 1728 5160
rect 4528 5108 4580 5160
rect 4804 5108 4856 5160
rect 5632 5108 5684 5160
rect 6092 5108 6144 5160
rect 6368 5108 6420 5160
rect 7012 5108 7064 5160
rect 8576 5176 8628 5228
rect 9956 5176 10008 5228
rect 10876 5176 10928 5228
rect 8392 5108 8444 5160
rect 10784 5151 10836 5160
rect 7472 5040 7524 5092
rect 7840 5040 7892 5092
rect 3516 4972 3568 5024
rect 3700 5015 3752 5024
rect 3700 4981 3709 5015
rect 3709 4981 3743 5015
rect 3743 4981 3752 5015
rect 3700 4972 3752 4981
rect 5540 4972 5592 5024
rect 5724 4972 5776 5024
rect 7932 4972 7984 5024
rect 9128 5040 9180 5092
rect 9220 5040 9272 5092
rect 10784 5117 10793 5151
rect 10793 5117 10827 5151
rect 10827 5117 10836 5151
rect 10784 5108 10836 5117
rect 8760 5015 8812 5024
rect 8760 4981 8769 5015
rect 8769 4981 8803 5015
rect 8803 4981 8812 5015
rect 8760 4972 8812 4981
rect 9496 4972 9548 5024
rect 9772 4972 9824 5024
rect 11520 5108 11572 5160
rect 11796 5176 11848 5228
rect 12348 5176 12400 5228
rect 12440 5176 12492 5228
rect 12624 5176 12676 5228
rect 12716 5176 12768 5228
rect 12992 5219 13044 5228
rect 12992 5185 13001 5219
rect 13001 5185 13035 5219
rect 13035 5185 13044 5219
rect 12992 5176 13044 5185
rect 13360 5176 13412 5228
rect 11888 5108 11940 5160
rect 12256 5108 12308 5160
rect 13084 5108 13136 5160
rect 13636 5108 13688 5160
rect 13544 5040 13596 5092
rect 11796 5015 11848 5024
rect 11796 4981 11805 5015
rect 11805 4981 11839 5015
rect 11839 4981 11848 5015
rect 11796 4972 11848 4981
rect 12992 4972 13044 5024
rect 13728 4972 13780 5024
rect 14832 4972 14884 5024
rect 15016 5015 15068 5024
rect 15016 4981 15025 5015
rect 15025 4981 15059 5015
rect 15059 4981 15068 5015
rect 15016 4972 15068 4981
rect 5912 4870 5964 4922
rect 5976 4870 6028 4922
rect 6040 4870 6092 4922
rect 6104 4870 6156 4922
rect 10843 4870 10895 4922
rect 10907 4870 10959 4922
rect 10971 4870 11023 4922
rect 11035 4870 11087 4922
rect 3424 4768 3476 4820
rect 3700 4768 3752 4820
rect 4988 4768 5040 4820
rect 5356 4768 5408 4820
rect 7196 4768 7248 4820
rect 7472 4768 7524 4820
rect 8392 4768 8444 4820
rect 9128 4768 9180 4820
rect 9312 4768 9364 4820
rect 9496 4768 9548 4820
rect 9956 4768 10008 4820
rect 10416 4768 10468 4820
rect 3976 4700 4028 4752
rect 4436 4743 4488 4752
rect 4436 4709 4445 4743
rect 4445 4709 4479 4743
rect 4479 4709 4488 4743
rect 4436 4700 4488 4709
rect 2136 4632 2188 4684
rect 4068 4632 4120 4684
rect 3056 4564 3108 4616
rect 3332 4607 3384 4616
rect 3332 4573 3341 4607
rect 3341 4573 3375 4607
rect 3375 4573 3384 4607
rect 3332 4564 3384 4573
rect 3516 4607 3568 4616
rect 3516 4573 3525 4607
rect 3525 4573 3559 4607
rect 3559 4573 3568 4607
rect 3516 4564 3568 4573
rect 6276 4700 6328 4752
rect 4804 4632 4856 4684
rect 5264 4632 5316 4684
rect 5632 4675 5684 4684
rect 5632 4641 5641 4675
rect 5641 4641 5675 4675
rect 5675 4641 5684 4675
rect 5632 4632 5684 4641
rect 6184 4632 6236 4684
rect 7564 4700 7616 4752
rect 7932 4700 7984 4752
rect 8576 4700 8628 4752
rect 11336 4768 11388 4820
rect 13084 4768 13136 4820
rect 13268 4811 13320 4820
rect 13268 4777 13277 4811
rect 13277 4777 13311 4811
rect 13311 4777 13320 4811
rect 13268 4768 13320 4777
rect 13544 4768 13596 4820
rect 14648 4811 14700 4820
rect 14648 4777 14657 4811
rect 14657 4777 14691 4811
rect 14691 4777 14700 4811
rect 14648 4768 14700 4777
rect 7012 4632 7064 4684
rect 10140 4675 10192 4684
rect 10140 4641 10149 4675
rect 10149 4641 10183 4675
rect 10183 4641 10192 4675
rect 10140 4632 10192 4641
rect 5724 4607 5776 4616
rect 5724 4573 5733 4607
rect 5733 4573 5767 4607
rect 5767 4573 5776 4607
rect 5724 4564 5776 4573
rect 5816 4607 5868 4616
rect 5816 4573 5825 4607
rect 5825 4573 5859 4607
rect 5859 4573 5868 4607
rect 5816 4564 5868 4573
rect 7472 4564 7524 4616
rect 8116 4564 8168 4616
rect 8576 4564 8628 4616
rect 10048 4564 10100 4616
rect 10692 4632 10744 4684
rect 10784 4632 10836 4684
rect 10324 4564 10376 4616
rect 10968 4564 11020 4616
rect 12808 4700 12860 4752
rect 13452 4700 13504 4752
rect 2964 4496 3016 4548
rect 3608 4496 3660 4548
rect 5356 4496 5408 4548
rect 5448 4496 5500 4548
rect 6276 4496 6328 4548
rect 8484 4496 8536 4548
rect 11152 4496 11204 4548
rect 14464 4675 14516 4684
rect 14464 4641 14473 4675
rect 14473 4641 14507 4675
rect 14507 4641 14516 4675
rect 14464 4632 14516 4641
rect 12256 4564 12308 4616
rect 12716 4607 12768 4616
rect 12716 4573 12725 4607
rect 12725 4573 12759 4607
rect 12759 4573 12768 4607
rect 12716 4564 12768 4573
rect 13360 4564 13412 4616
rect 4068 4471 4120 4480
rect 4068 4437 4077 4471
rect 4077 4437 4111 4471
rect 4111 4437 4120 4471
rect 4068 4428 4120 4437
rect 4804 4428 4856 4480
rect 6368 4428 6420 4480
rect 6828 4428 6880 4480
rect 7472 4428 7524 4480
rect 7840 4471 7892 4480
rect 7840 4437 7849 4471
rect 7849 4437 7883 4471
rect 7883 4437 7892 4471
rect 7840 4428 7892 4437
rect 8760 4428 8812 4480
rect 9312 4428 9364 4480
rect 9588 4428 9640 4480
rect 10140 4428 10192 4480
rect 10600 4428 10652 4480
rect 11060 4428 11112 4480
rect 11520 4428 11572 4480
rect 12716 4428 12768 4480
rect 3447 4326 3499 4378
rect 3511 4326 3563 4378
rect 3575 4326 3627 4378
rect 3639 4326 3691 4378
rect 8378 4326 8430 4378
rect 8442 4326 8494 4378
rect 8506 4326 8558 4378
rect 8570 4326 8622 4378
rect 13308 4326 13360 4378
rect 13372 4326 13424 4378
rect 13436 4326 13488 4378
rect 13500 4326 13552 4378
rect 5356 4224 5408 4276
rect 5540 4267 5592 4276
rect 5540 4233 5549 4267
rect 5549 4233 5583 4267
rect 5583 4233 5592 4267
rect 5540 4224 5592 4233
rect 5632 4224 5684 4276
rect 7472 4224 7524 4276
rect 9036 4224 9088 4276
rect 9312 4224 9364 4276
rect 10324 4224 10376 4276
rect 10968 4224 11020 4276
rect 11428 4224 11480 4276
rect 11520 4224 11572 4276
rect 11888 4224 11940 4276
rect 12716 4224 12768 4276
rect 4252 4156 4304 4208
rect 4528 4088 4580 4140
rect 6460 4156 6512 4208
rect 1308 4020 1360 4072
rect 3332 4020 3384 4072
rect 4804 4020 4856 4072
rect 5540 4020 5592 4072
rect 5908 4020 5960 4072
rect 6828 4088 6880 4140
rect 7380 4131 7432 4140
rect 7380 4097 7389 4131
rect 7389 4097 7423 4131
rect 7423 4097 7432 4131
rect 7380 4088 7432 4097
rect 7932 4088 7984 4140
rect 9680 4156 9732 4208
rect 9864 4156 9916 4208
rect 10876 4156 10928 4208
rect 6368 4020 6420 4072
rect 7196 4020 7248 4072
rect 7840 4020 7892 4072
rect 9036 4020 9088 4072
rect 9128 4020 9180 4072
rect 9312 4063 9364 4072
rect 9312 4029 9321 4063
rect 9321 4029 9355 4063
rect 9355 4029 9364 4063
rect 9312 4020 9364 4029
rect 9496 4020 9548 4072
rect 11336 4088 11388 4140
rect 2136 3952 2188 4004
rect 2780 3952 2832 4004
rect 3056 3952 3108 4004
rect 5632 3952 5684 4004
rect 6184 3952 6236 4004
rect 6276 3952 6328 4004
rect 6460 3952 6512 4004
rect 1676 3884 1728 3936
rect 2964 3884 3016 3936
rect 4252 3884 4304 3936
rect 4436 3927 4488 3936
rect 4436 3893 4445 3927
rect 4445 3893 4479 3927
rect 4479 3893 4488 3927
rect 4436 3884 4488 3893
rect 4528 3927 4580 3936
rect 4528 3893 4537 3927
rect 4537 3893 4571 3927
rect 4571 3893 4580 3927
rect 4528 3884 4580 3893
rect 4804 3884 4856 3936
rect 6828 3952 6880 4004
rect 7012 3952 7064 4004
rect 8116 3952 8168 4004
rect 9864 3952 9916 4004
rect 11428 4020 11480 4072
rect 12256 4156 12308 4208
rect 11704 4088 11756 4140
rect 13084 4224 13136 4276
rect 13268 4156 13320 4208
rect 13084 4088 13136 4140
rect 12072 4020 12124 4072
rect 12532 4020 12584 4072
rect 13360 4020 13412 4072
rect 7288 3884 7340 3936
rect 9036 3884 9088 3936
rect 10232 3884 10284 3936
rect 10416 3927 10468 3936
rect 10416 3893 10425 3927
rect 10425 3893 10459 3927
rect 10459 3893 10468 3927
rect 10416 3884 10468 3893
rect 10692 3884 10744 3936
rect 11888 3952 11940 4004
rect 12808 3995 12860 4004
rect 12808 3961 12817 3995
rect 12817 3961 12851 3995
rect 12851 3961 12860 3995
rect 12808 3952 12860 3961
rect 14004 3995 14056 4004
rect 11336 3884 11388 3936
rect 11796 3884 11848 3936
rect 12256 3884 12308 3936
rect 13636 3927 13688 3936
rect 13636 3893 13645 3927
rect 13645 3893 13679 3927
rect 13679 3893 13688 3927
rect 13636 3884 13688 3893
rect 14004 3961 14013 3995
rect 14013 3961 14047 3995
rect 14047 3961 14056 3995
rect 14004 3952 14056 3961
rect 15108 3952 15160 4004
rect 14280 3884 14332 3936
rect 15016 3927 15068 3936
rect 15016 3893 15025 3927
rect 15025 3893 15059 3927
rect 15059 3893 15068 3927
rect 15016 3884 15068 3893
rect 5912 3782 5964 3834
rect 5976 3782 6028 3834
rect 6040 3782 6092 3834
rect 6104 3782 6156 3834
rect 10843 3782 10895 3834
rect 10907 3782 10959 3834
rect 10971 3782 11023 3834
rect 11035 3782 11087 3834
rect 2412 3612 2464 3664
rect 2872 3723 2924 3732
rect 2872 3689 2881 3723
rect 2881 3689 2915 3723
rect 2915 3689 2924 3723
rect 2872 3680 2924 3689
rect 3240 3680 3292 3732
rect 4528 3680 4580 3732
rect 3976 3612 4028 3664
rect 4160 3612 4212 3664
rect 572 3544 624 3596
rect 1492 3544 1544 3596
rect 2136 3544 2188 3596
rect 3240 3587 3292 3596
rect 1308 3476 1360 3528
rect 3240 3553 3249 3587
rect 3249 3553 3283 3587
rect 3283 3553 3292 3587
rect 3240 3544 3292 3553
rect 3608 3544 3660 3596
rect 5356 3587 5408 3596
rect 5356 3553 5365 3587
rect 5365 3553 5399 3587
rect 5399 3553 5408 3587
rect 5356 3544 5408 3553
rect 7748 3680 7800 3732
rect 8300 3723 8352 3732
rect 8300 3689 8309 3723
rect 8309 3689 8343 3723
rect 8343 3689 8352 3723
rect 8300 3680 8352 3689
rect 8484 3680 8536 3732
rect 10692 3680 10744 3732
rect 11796 3680 11848 3732
rect 12072 3680 12124 3732
rect 12624 3680 12676 3732
rect 13268 3723 13320 3732
rect 13268 3689 13277 3723
rect 13277 3689 13311 3723
rect 13311 3689 13320 3723
rect 13268 3680 13320 3689
rect 13912 3680 13964 3732
rect 14648 3723 14700 3732
rect 14648 3689 14657 3723
rect 14657 3689 14691 3723
rect 14691 3689 14700 3723
rect 14648 3680 14700 3689
rect 6184 3655 6236 3664
rect 6184 3621 6193 3655
rect 6193 3621 6227 3655
rect 6227 3621 6236 3655
rect 6184 3612 6236 3621
rect 8392 3612 8444 3664
rect 6276 3587 6328 3596
rect 6276 3553 6285 3587
rect 6285 3553 6319 3587
rect 6319 3553 6328 3587
rect 6276 3544 6328 3553
rect 7196 3544 7248 3596
rect 7840 3587 7892 3596
rect 7840 3553 7849 3587
rect 7849 3553 7883 3587
rect 7883 3553 7892 3587
rect 7840 3544 7892 3553
rect 4528 3519 4580 3528
rect 4528 3485 4537 3519
rect 4537 3485 4571 3519
rect 4571 3485 4580 3519
rect 4528 3476 4580 3485
rect 4988 3476 5040 3528
rect 5448 3519 5500 3528
rect 5448 3485 5457 3519
rect 5457 3485 5491 3519
rect 5491 3485 5500 3519
rect 5448 3476 5500 3485
rect 4804 3408 4856 3460
rect 5816 3476 5868 3528
rect 6184 3476 6236 3528
rect 6920 3476 6972 3528
rect 7380 3476 7432 3528
rect 8576 3544 8628 3596
rect 8208 3476 8260 3528
rect 5724 3408 5776 3460
rect 8668 3408 8720 3460
rect 9312 3612 9364 3664
rect 9680 3544 9732 3596
rect 11520 3612 11572 3664
rect 10232 3544 10284 3596
rect 10508 3544 10560 3596
rect 10968 3544 11020 3596
rect 11244 3587 11296 3596
rect 11244 3553 11253 3587
rect 11253 3553 11287 3587
rect 11287 3553 11296 3587
rect 11244 3544 11296 3553
rect 9128 3476 9180 3528
rect 9588 3476 9640 3528
rect 9864 3476 9916 3528
rect 10140 3476 10192 3528
rect 15200 3612 15252 3664
rect 15936 3612 15988 3664
rect 13176 3544 13228 3596
rect 13268 3544 13320 3596
rect 14464 3587 14516 3596
rect 14464 3553 14473 3587
rect 14473 3553 14507 3587
rect 14507 3553 14516 3587
rect 14464 3544 14516 3553
rect 11612 3476 11664 3528
rect 12072 3476 12124 3528
rect 12624 3519 12676 3528
rect 12624 3485 12633 3519
rect 12633 3485 12667 3519
rect 12667 3485 12676 3519
rect 12624 3476 12676 3485
rect 9036 3408 9088 3460
rect 10692 3408 10744 3460
rect 10876 3451 10928 3460
rect 10876 3417 10885 3451
rect 10885 3417 10919 3451
rect 10919 3417 10928 3451
rect 10876 3408 10928 3417
rect 2320 3340 2372 3392
rect 4988 3383 5040 3392
rect 4988 3349 4997 3383
rect 4997 3349 5031 3383
rect 5031 3349 5040 3383
rect 4988 3340 5040 3349
rect 5632 3340 5684 3392
rect 11244 3340 11296 3392
rect 11704 3340 11756 3392
rect 11888 3383 11940 3392
rect 11888 3349 11897 3383
rect 11897 3349 11931 3383
rect 11931 3349 11940 3383
rect 11888 3340 11940 3349
rect 11980 3340 12032 3392
rect 13820 3340 13872 3392
rect 14556 3340 14608 3392
rect 3447 3238 3499 3290
rect 3511 3238 3563 3290
rect 3575 3238 3627 3290
rect 3639 3238 3691 3290
rect 8378 3238 8430 3290
rect 8442 3238 8494 3290
rect 8506 3238 8558 3290
rect 8570 3238 8622 3290
rect 13308 3238 13360 3290
rect 13372 3238 13424 3290
rect 13436 3238 13488 3290
rect 13500 3238 13552 3290
rect 1032 3136 1084 3188
rect 1584 3136 1636 3188
rect 4344 3136 4396 3188
rect 4528 3136 4580 3188
rect 2872 3068 2924 3120
rect 5448 3068 5500 3120
rect 6368 3068 6420 3120
rect 1308 3000 1360 3052
rect 4252 3000 4304 3052
rect 4620 3000 4672 3052
rect 5632 3000 5684 3052
rect 3700 2932 3752 2984
rect 6184 3043 6236 3052
rect 6184 3009 6193 3043
rect 6193 3009 6227 3043
rect 6227 3009 6236 3043
rect 6184 3000 6236 3009
rect 6460 2932 6512 2984
rect 1768 2864 1820 2916
rect 2504 2864 2556 2916
rect 4712 2907 4764 2916
rect 4712 2873 4721 2907
rect 4721 2873 4755 2907
rect 4755 2873 4764 2907
rect 4712 2864 4764 2873
rect 6092 2864 6144 2916
rect 7380 3136 7432 3188
rect 8668 3136 8720 3188
rect 9220 3179 9272 3188
rect 9220 3145 9229 3179
rect 9229 3145 9263 3179
rect 9263 3145 9272 3179
rect 9220 3136 9272 3145
rect 12440 3136 12492 3188
rect 12532 3136 12584 3188
rect 10508 3068 10560 3120
rect 11612 3068 11664 3120
rect 13268 3068 13320 3120
rect 13912 3068 13964 3120
rect 14004 3068 14056 3120
rect 14924 3068 14976 3120
rect 7196 3000 7248 3052
rect 7380 3043 7432 3052
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 7472 3000 7524 3052
rect 8852 3000 8904 3052
rect 10324 3000 10376 3052
rect 11152 3000 11204 3052
rect 13084 3043 13136 3052
rect 13084 3009 13093 3043
rect 13093 3009 13127 3043
rect 13127 3009 13136 3043
rect 13084 3000 13136 3009
rect 14740 3000 14792 3052
rect 8484 2932 8536 2984
rect 8576 2975 8628 2984
rect 8576 2941 8585 2975
rect 8585 2941 8619 2975
rect 8619 2941 8628 2975
rect 8576 2932 8628 2941
rect 7104 2864 7156 2916
rect 7656 2864 7708 2916
rect 9220 2932 9272 2984
rect 10416 2932 10468 2984
rect 10600 2932 10652 2984
rect 12348 2932 12400 2984
rect 12440 2932 12492 2984
rect 9128 2864 9180 2916
rect 2872 2796 2924 2848
rect 3884 2796 3936 2848
rect 4344 2839 4396 2848
rect 4344 2805 4353 2839
rect 4353 2805 4387 2839
rect 4387 2805 4396 2839
rect 4344 2796 4396 2805
rect 4804 2839 4856 2848
rect 4804 2805 4813 2839
rect 4813 2805 4847 2839
rect 4847 2805 4856 2839
rect 4804 2796 4856 2805
rect 5356 2796 5408 2848
rect 5448 2796 5500 2848
rect 7840 2796 7892 2848
rect 9496 2796 9548 2848
rect 9772 2796 9824 2848
rect 11244 2864 11296 2916
rect 11888 2864 11940 2916
rect 12992 2932 13044 2984
rect 14096 2932 14148 2984
rect 14556 2975 14608 2984
rect 14556 2941 14565 2975
rect 14565 2941 14599 2975
rect 14599 2941 14608 2975
rect 14556 2932 14608 2941
rect 14832 2932 14884 2984
rect 12164 2796 12216 2848
rect 12348 2796 12400 2848
rect 14648 2864 14700 2916
rect 14004 2796 14056 2848
rect 14740 2839 14792 2848
rect 14740 2805 14749 2839
rect 14749 2805 14783 2839
rect 14783 2805 14792 2839
rect 14740 2796 14792 2805
rect 15108 2864 15160 2916
rect 16764 2864 16816 2916
rect 15292 2796 15344 2848
rect 5912 2694 5964 2746
rect 5976 2694 6028 2746
rect 6040 2694 6092 2746
rect 6104 2694 6156 2746
rect 10843 2694 10895 2746
rect 10907 2694 10959 2746
rect 10971 2694 11023 2746
rect 11035 2694 11087 2746
rect 2320 2592 2372 2644
rect 2872 2635 2924 2644
rect 2872 2601 2881 2635
rect 2881 2601 2915 2635
rect 2915 2601 2924 2635
rect 2872 2592 2924 2601
rect 3332 2592 3384 2644
rect 2228 2524 2280 2576
rect 3976 2592 4028 2644
rect 5540 2635 5592 2644
rect 5540 2601 5549 2635
rect 5549 2601 5583 2635
rect 5583 2601 5592 2635
rect 5540 2592 5592 2601
rect 5816 2592 5868 2644
rect 6736 2592 6788 2644
rect 2228 2431 2280 2440
rect 2228 2397 2237 2431
rect 2237 2397 2271 2431
rect 2271 2397 2280 2431
rect 2228 2388 2280 2397
rect 3240 2388 3292 2440
rect 3424 2431 3476 2440
rect 3424 2397 3433 2431
rect 3433 2397 3467 2431
rect 3467 2397 3476 2431
rect 3700 2431 3752 2440
rect 3424 2388 3476 2397
rect 3700 2397 3709 2431
rect 3709 2397 3743 2431
rect 3743 2397 3752 2431
rect 3700 2388 3752 2397
rect 7840 2592 7892 2644
rect 9588 2592 9640 2644
rect 12256 2592 12308 2644
rect 12348 2592 12400 2644
rect 13268 2592 13320 2644
rect 5540 2456 5592 2508
rect 7012 2456 7064 2508
rect 7104 2456 7156 2508
rect 8208 2456 8260 2508
rect 8944 2456 8996 2508
rect 10048 2524 10100 2576
rect 10600 2456 10652 2508
rect 6552 2388 6604 2440
rect 7472 2431 7524 2440
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 7472 2388 7524 2397
rect 8760 2431 8812 2440
rect 8760 2397 8769 2431
rect 8769 2397 8803 2431
rect 8803 2397 8812 2431
rect 8760 2388 8812 2397
rect 9220 2388 9272 2440
rect 10048 2388 10100 2440
rect 10324 2388 10376 2440
rect 10416 2431 10468 2440
rect 10416 2397 10425 2431
rect 10425 2397 10459 2431
rect 10459 2397 10468 2431
rect 13636 2524 13688 2576
rect 15108 2524 15160 2576
rect 11612 2456 11664 2508
rect 12348 2456 12400 2508
rect 12624 2499 12676 2508
rect 12624 2465 12633 2499
rect 12633 2465 12667 2499
rect 12667 2465 12676 2499
rect 12624 2456 12676 2465
rect 12716 2456 12768 2508
rect 14464 2499 14516 2508
rect 14464 2465 14473 2499
rect 14473 2465 14507 2499
rect 14507 2465 14516 2499
rect 14464 2456 14516 2465
rect 10416 2388 10468 2397
rect 11704 2388 11756 2440
rect 11980 2388 12032 2440
rect 12808 2431 12860 2440
rect 12808 2397 12817 2431
rect 12817 2397 12851 2431
rect 12851 2397 12860 2431
rect 12808 2388 12860 2397
rect 13728 2431 13780 2440
rect 13728 2397 13737 2431
rect 13737 2397 13771 2431
rect 13771 2397 13780 2431
rect 13728 2388 13780 2397
rect 5356 2320 5408 2372
rect 5816 2320 5868 2372
rect 14188 2320 14240 2372
rect 3792 2252 3844 2304
rect 4068 2252 4120 2304
rect 4252 2252 4304 2304
rect 6920 2295 6972 2304
rect 6920 2261 6929 2295
rect 6929 2261 6963 2295
rect 6963 2261 6972 2295
rect 6920 2252 6972 2261
rect 7932 2252 7984 2304
rect 9128 2252 9180 2304
rect 9404 2295 9456 2304
rect 9404 2261 9413 2295
rect 9413 2261 9447 2295
rect 9447 2261 9456 2295
rect 9404 2252 9456 2261
rect 9772 2295 9824 2304
rect 9772 2261 9781 2295
rect 9781 2261 9815 2295
rect 9815 2261 9824 2295
rect 9772 2252 9824 2261
rect 10048 2252 10100 2304
rect 11704 2252 11756 2304
rect 11980 2295 12032 2304
rect 11980 2261 11989 2295
rect 11989 2261 12023 2295
rect 12023 2261 12032 2295
rect 11980 2252 12032 2261
rect 3447 2150 3499 2202
rect 3511 2150 3563 2202
rect 3575 2150 3627 2202
rect 3639 2150 3691 2202
rect 8378 2150 8430 2202
rect 8442 2150 8494 2202
rect 8506 2150 8558 2202
rect 8570 2150 8622 2202
rect 13308 2150 13360 2202
rect 13372 2150 13424 2202
rect 13436 2150 13488 2202
rect 13500 2150 13552 2202
rect 5264 2048 5316 2100
rect 9404 2048 9456 2100
rect 10692 2048 10744 2100
rect 13176 2048 13228 2100
rect 14464 2091 14516 2100
rect 14464 2057 14473 2091
rect 14473 2057 14507 2091
rect 14507 2057 14516 2091
rect 14464 2048 14516 2057
rect 2044 1980 2096 2032
rect 12808 1980 12860 2032
rect 204 1912 256 1964
rect 11980 1912 12032 1964
rect 4160 1844 4212 1896
rect 7012 1844 7064 1896
rect 11612 1844 11664 1896
rect 13728 1844 13780 1896
rect 4896 1776 4948 1828
rect 7288 1776 7340 1828
rect 10968 1776 11020 1828
rect 12624 1776 12676 1828
rect 2964 1708 3016 1760
rect 9772 1708 9824 1760
rect 10600 1708 10652 1760
rect 15476 1708 15528 1760
rect 1952 1640 2004 1692
rect 6920 1640 6972 1692
rect 12716 1640 12768 1692
rect 2228 1572 2280 1624
rect 10232 1572 10284 1624
rect 11152 1572 11204 1624
rect 16304 1572 16356 1624
rect 6276 1504 6328 1556
rect 8484 1504 8536 1556
rect 8852 1504 8904 1556
rect 9864 1504 9916 1556
rect 11428 1504 11480 1556
rect 15108 1504 15160 1556
rect 1400 1436 1452 1488
rect 6644 1436 6696 1488
rect 1124 1368 1176 1420
rect 2228 1300 2280 1352
rect 9496 1300 9548 1352
rect 6000 1232 6052 1284
rect 6736 1232 6788 1284
rect 1860 1164 1912 1216
rect 7564 1164 7616 1216
rect 4712 1096 4764 1148
rect 9312 1096 9364 1148
rect 7380 1028 7432 1080
rect 13084 1028 13136 1080
rect 8208 960 8260 1012
rect 9312 960 9364 1012
rect 4436 892 4488 944
rect 9588 892 9640 944
rect 8944 620 8996 672
rect 12624 620 12676 672
<< metal2 >>
rect 202 19520 258 20000
rect 570 19520 626 20000
rect 938 19520 994 20000
rect 1398 19520 1454 20000
rect 1766 19520 1822 20000
rect 2226 19520 2282 20000
rect 2594 19520 2650 20000
rect 2870 19544 2926 19553
rect 216 16182 244 19520
rect 584 17610 612 19520
rect 572 17604 624 17610
rect 572 17546 624 17552
rect 204 16176 256 16182
rect 204 16118 256 16124
rect 952 15638 980 19520
rect 1412 16522 1440 19520
rect 1780 17746 1808 19520
rect 1768 17740 1820 17746
rect 1768 17682 1820 17688
rect 2136 17060 2188 17066
rect 2136 17002 2188 17008
rect 2148 16697 2176 17002
rect 2134 16688 2190 16697
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1860 16652 1912 16658
rect 2134 16623 2190 16632
rect 1860 16594 1912 16600
rect 1400 16516 1452 16522
rect 1400 16458 1452 16464
rect 940 15632 992 15638
rect 940 15574 992 15580
rect 1596 14618 1624 16594
rect 1676 16040 1728 16046
rect 1676 15982 1728 15988
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 1492 13864 1544 13870
rect 1492 13806 1544 13812
rect 572 13796 624 13802
rect 572 13738 624 13744
rect 584 10033 612 13738
rect 1504 13138 1532 13806
rect 1582 13288 1638 13297
rect 1582 13223 1584 13232
rect 1636 13223 1638 13232
rect 1584 13194 1636 13200
rect 1504 13110 1624 13138
rect 1492 12708 1544 12714
rect 1492 12650 1544 12656
rect 1398 10160 1454 10169
rect 1398 10095 1400 10104
rect 1452 10095 1454 10104
rect 1400 10066 1452 10072
rect 570 10024 626 10033
rect 570 9959 626 9968
rect 1504 9738 1532 12650
rect 1596 12442 1624 13110
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1412 9710 1532 9738
rect 1032 8288 1084 8294
rect 1032 8230 1084 8236
rect 572 3596 624 3602
rect 572 3538 624 3544
rect 204 1964 256 1970
rect 204 1906 256 1912
rect 216 480 244 1906
rect 584 480 612 3538
rect 1044 3505 1072 8230
rect 1308 6316 1360 6322
rect 1308 6258 1360 6264
rect 1214 6216 1270 6225
rect 1214 6151 1270 6160
rect 1122 4312 1178 4321
rect 1122 4247 1178 4256
rect 1030 3496 1086 3505
rect 1030 3431 1086 3440
rect 1032 3188 1084 3194
rect 1032 3130 1084 3136
rect 1044 480 1072 3130
rect 1136 1426 1164 4247
rect 1228 2009 1256 6151
rect 1320 4078 1348 6258
rect 1412 5370 1440 9710
rect 1492 7744 1544 7750
rect 1492 7686 1544 7692
rect 1400 5364 1452 5370
rect 1400 5306 1452 5312
rect 1308 4072 1360 4078
rect 1308 4014 1360 4020
rect 1320 3534 1348 4014
rect 1504 3602 1532 7686
rect 1596 6866 1624 11494
rect 1688 10810 1716 15982
rect 1872 15745 1900 16594
rect 2240 16590 2268 19520
rect 2412 16652 2464 16658
rect 2412 16594 2464 16600
rect 2228 16584 2280 16590
rect 2228 16526 2280 16532
rect 2228 16448 2280 16454
rect 2228 16390 2280 16396
rect 1858 15736 1914 15745
rect 1858 15671 1914 15680
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1858 11928 1914 11937
rect 1858 11863 1914 11872
rect 1872 11286 1900 11863
rect 1860 11280 1912 11286
rect 1964 11257 1992 14758
rect 2240 13870 2268 16390
rect 2318 16144 2374 16153
rect 2318 16079 2374 16088
rect 2332 15570 2360 16079
rect 2320 15564 2372 15570
rect 2320 15506 2372 15512
rect 2320 14816 2372 14822
rect 2320 14758 2372 14764
rect 2228 13864 2280 13870
rect 2228 13806 2280 13812
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 1860 11222 1912 11228
rect 1950 11248 2006 11257
rect 1950 11183 2006 11192
rect 2148 10810 2176 12174
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1858 10568 1914 10577
rect 1688 9489 1716 10542
rect 1858 10503 1914 10512
rect 1674 9480 1730 9489
rect 1674 9415 1730 9424
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1492 3596 1544 3602
rect 1492 3538 1544 3544
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1320 3058 1348 3470
rect 1596 3194 1624 6054
rect 1688 5166 1716 9415
rect 1768 8356 1820 8362
rect 1768 8298 1820 8304
rect 1780 7857 1808 8298
rect 1766 7848 1822 7857
rect 1766 7783 1822 7792
rect 1872 7698 1900 10503
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 2056 8945 2084 8978
rect 2136 8968 2188 8974
rect 2042 8936 2098 8945
rect 2136 8910 2188 8916
rect 2042 8871 2098 8880
rect 2148 8566 2176 8910
rect 2136 8560 2188 8566
rect 2136 8502 2188 8508
rect 2148 7954 2176 8502
rect 2240 8294 2268 13126
rect 2332 12481 2360 14758
rect 2424 14074 2452 16594
rect 2502 15056 2558 15065
rect 2502 14991 2558 15000
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 2516 13734 2544 14991
rect 2608 14929 2636 19520
rect 2962 19520 3018 20000
rect 3422 19520 3478 20000
rect 3790 19520 3846 20000
rect 4250 19520 4306 20000
rect 4618 19520 4674 20000
rect 4986 19520 5042 20000
rect 5446 19520 5502 20000
rect 5814 19520 5870 20000
rect 6274 19520 6330 20000
rect 6642 19520 6698 20000
rect 7010 19520 7066 20000
rect 7470 19520 7526 20000
rect 7838 19520 7894 20000
rect 8298 19520 8354 20000
rect 8666 19520 8722 20000
rect 9034 19520 9090 20000
rect 9494 19520 9550 20000
rect 9862 19520 9918 20000
rect 10322 19520 10378 20000
rect 10690 19520 10746 20000
rect 11058 19520 11114 20000
rect 11518 19520 11574 20000
rect 11886 19520 11942 20000
rect 12346 19520 12402 20000
rect 12714 19520 12770 20000
rect 13082 19530 13138 20000
rect 12912 19520 13138 19530
rect 13542 19520 13598 20000
rect 13910 19520 13966 20000
rect 14370 19520 14426 20000
rect 14738 19520 14794 20000
rect 15106 19520 15162 20000
rect 15566 19520 15622 20000
rect 15934 19520 15990 20000
rect 16394 19520 16450 20000
rect 16762 19520 16818 20000
rect 2870 19479 2926 19488
rect 2778 17640 2834 17649
rect 2778 17575 2834 17584
rect 2792 16114 2820 17575
rect 2884 16250 2912 19479
rect 2976 17626 3004 19520
rect 3436 18154 3464 19520
rect 3514 18592 3570 18601
rect 3514 18527 3570 18536
rect 3424 18148 3476 18154
rect 3424 18090 3476 18096
rect 3528 18018 3556 18527
rect 3516 18012 3568 18018
rect 3516 17954 3568 17960
rect 2976 17598 3188 17626
rect 3056 17060 3108 17066
rect 3056 17002 3108 17008
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2792 15609 2820 15642
rect 2778 15600 2834 15609
rect 2778 15535 2834 15544
rect 2780 15428 2832 15434
rect 2780 15370 2832 15376
rect 2792 15094 2820 15370
rect 2780 15088 2832 15094
rect 2976 15042 3004 16594
rect 2780 15030 2832 15036
rect 2884 15014 3004 15042
rect 2594 14920 2650 14929
rect 2594 14855 2650 14864
rect 2780 14884 2832 14890
rect 2780 14826 2832 14832
rect 2688 14544 2740 14550
rect 2688 14486 2740 14492
rect 2596 14408 2648 14414
rect 2596 14350 2648 14356
rect 2504 13728 2556 13734
rect 2504 13670 2556 13676
rect 2608 13462 2636 14350
rect 2596 13456 2648 13462
rect 2596 13398 2648 13404
rect 2596 13252 2648 13258
rect 2596 13194 2648 13200
rect 2502 12744 2558 12753
rect 2502 12679 2558 12688
rect 2318 12472 2374 12481
rect 2318 12407 2374 12416
rect 2320 11688 2372 11694
rect 2318 11656 2320 11665
rect 2372 11656 2374 11665
rect 2318 11591 2374 11600
rect 2412 11620 2464 11626
rect 2412 11562 2464 11568
rect 2424 11218 2452 11562
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2516 10826 2544 12679
rect 2424 10798 2544 10826
rect 2320 10464 2372 10470
rect 2320 10406 2372 10412
rect 2332 9722 2360 10406
rect 2320 9716 2372 9722
rect 2320 9658 2372 9664
rect 2320 8356 2372 8362
rect 2320 8298 2372 8304
rect 2228 8288 2280 8294
rect 2228 8230 2280 8236
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 2136 7948 2188 7954
rect 2136 7890 2188 7896
rect 1780 7670 1900 7698
rect 1676 5160 1728 5166
rect 1676 5102 1728 5108
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1584 3188 1636 3194
rect 1584 3130 1636 3136
rect 1308 3052 1360 3058
rect 1308 2994 1360 3000
rect 1688 2553 1716 3878
rect 1780 2922 1808 7670
rect 1964 7313 1992 7890
rect 2136 7336 2188 7342
rect 1950 7304 2006 7313
rect 2136 7278 2188 7284
rect 1950 7239 2006 7248
rect 2148 6798 2176 7278
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 1952 6384 2004 6390
rect 1952 6326 2004 6332
rect 1858 6216 1914 6225
rect 1858 6151 1914 6160
rect 1872 6118 1900 6151
rect 1860 6112 1912 6118
rect 1860 6054 1912 6060
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 1872 5817 1900 5850
rect 1858 5808 1914 5817
rect 1858 5743 1914 5752
rect 1768 2916 1820 2922
rect 1768 2858 1820 2864
rect 1674 2544 1730 2553
rect 1674 2479 1730 2488
rect 1214 2000 1270 2009
rect 1214 1935 1270 1944
rect 1964 1698 1992 6326
rect 2148 6322 2176 6734
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2240 6202 2268 8230
rect 2332 6390 2360 8298
rect 2320 6384 2372 6390
rect 2320 6326 2372 6332
rect 2148 6174 2268 6202
rect 2042 5128 2098 5137
rect 2042 5063 2098 5072
rect 2056 2038 2084 5063
rect 2148 4690 2176 6174
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 2136 4684 2188 4690
rect 2136 4626 2188 4632
rect 2136 4004 2188 4010
rect 2136 3946 2188 3952
rect 2148 3602 2176 3946
rect 2136 3596 2188 3602
rect 2136 3538 2188 3544
rect 2240 2582 2268 6054
rect 2332 3398 2360 6054
rect 2424 3670 2452 10798
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 2516 10305 2544 10610
rect 2502 10296 2558 10305
rect 2502 10231 2558 10240
rect 2516 10198 2544 10231
rect 2504 10192 2556 10198
rect 2504 10134 2556 10140
rect 2608 10010 2636 13194
rect 2700 12458 2728 14486
rect 2792 13530 2820 14826
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2884 12889 2912 15014
rect 2964 14952 3016 14958
rect 2964 14894 3016 14900
rect 2976 14482 3004 14894
rect 3068 14793 3096 17002
rect 3160 16561 3188 17598
rect 3421 17436 3717 17456
rect 3477 17434 3501 17436
rect 3557 17434 3581 17436
rect 3637 17434 3661 17436
rect 3499 17382 3501 17434
rect 3563 17382 3575 17434
rect 3637 17382 3639 17434
rect 3477 17380 3501 17382
rect 3557 17380 3581 17382
rect 3637 17380 3661 17382
rect 3421 17360 3717 17380
rect 3804 16946 3832 19520
rect 4264 17490 4292 19520
rect 4264 17462 4476 17490
rect 4252 17332 4304 17338
rect 4252 17274 4304 17280
rect 3804 16918 4108 16946
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 3146 16552 3202 16561
rect 3146 16487 3202 16496
rect 3238 16008 3294 16017
rect 3238 15943 3294 15952
rect 3148 15904 3200 15910
rect 3148 15846 3200 15852
rect 3160 15473 3188 15846
rect 3146 15464 3202 15473
rect 3146 15399 3202 15408
rect 3148 15360 3200 15366
rect 3148 15302 3200 15308
rect 3054 14784 3110 14793
rect 3054 14719 3110 14728
rect 2964 14476 3016 14482
rect 2964 14418 3016 14424
rect 3056 14408 3108 14414
rect 2962 14376 3018 14385
rect 3056 14350 3108 14356
rect 2962 14311 3018 14320
rect 2976 13394 3004 14311
rect 2964 13388 3016 13394
rect 2964 13330 3016 13336
rect 3068 12986 3096 14350
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 2870 12880 2926 12889
rect 2870 12815 2926 12824
rect 3160 12594 3188 15302
rect 3252 15026 3280 15943
rect 3240 15020 3292 15026
rect 3240 14962 3292 14968
rect 3240 14816 3292 14822
rect 3240 14758 3292 14764
rect 3068 12566 3188 12594
rect 2700 12430 2820 12458
rect 2792 12424 2820 12430
rect 2792 12396 2912 12424
rect 2688 12368 2740 12374
rect 2688 12310 2740 12316
rect 2700 10198 2728 12310
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2792 12209 2820 12242
rect 2778 12200 2834 12209
rect 2778 12135 2834 12144
rect 2780 11824 2832 11830
rect 2780 11766 2832 11772
rect 2792 11286 2820 11766
rect 2780 11280 2832 11286
rect 2780 11222 2832 11228
rect 2792 10674 2820 11222
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 2688 10192 2740 10198
rect 2688 10134 2740 10140
rect 2792 10130 2820 10610
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 2686 10024 2742 10033
rect 2608 9982 2686 10010
rect 2686 9959 2742 9968
rect 2596 9716 2648 9722
rect 2596 9658 2648 9664
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 2516 9110 2544 9522
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2608 7528 2636 9658
rect 2700 8430 2728 9959
rect 2778 9072 2834 9081
rect 2778 9007 2834 9016
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2700 8022 2728 8366
rect 2688 8016 2740 8022
rect 2688 7958 2740 7964
rect 2608 7500 2728 7528
rect 2504 7268 2556 7274
rect 2504 7210 2556 7216
rect 2516 6769 2544 7210
rect 2594 6896 2650 6905
rect 2594 6831 2650 6840
rect 2502 6760 2558 6769
rect 2502 6695 2558 6704
rect 2504 6180 2556 6186
rect 2504 6122 2556 6128
rect 2412 3664 2464 3670
rect 2412 3606 2464 3612
rect 2320 3392 2372 3398
rect 2320 3334 2372 3340
rect 2332 2650 2360 3334
rect 2516 2922 2544 6122
rect 2608 5302 2636 6831
rect 2596 5296 2648 5302
rect 2596 5238 2648 5244
rect 2700 5234 2728 7500
rect 2792 6934 2820 9007
rect 2780 6928 2832 6934
rect 2780 6870 2832 6876
rect 2780 5704 2832 5710
rect 2778 5672 2780 5681
rect 2832 5672 2834 5681
rect 2778 5607 2834 5616
rect 2688 5228 2740 5234
rect 2688 5170 2740 5176
rect 2686 4040 2742 4049
rect 2686 3975 2742 3984
rect 2780 4004 2832 4010
rect 2504 2916 2556 2922
rect 2504 2858 2556 2864
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 2228 2576 2280 2582
rect 2228 2518 2280 2524
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 2044 2032 2096 2038
rect 2044 1974 2096 1980
rect 1952 1692 2004 1698
rect 1952 1634 2004 1640
rect 2240 1630 2268 2382
rect 2228 1624 2280 1630
rect 2228 1566 2280 1572
rect 1400 1488 1452 1494
rect 1400 1430 1452 1436
rect 1124 1420 1176 1426
rect 1124 1362 1176 1368
rect 1412 480 1440 1430
rect 2228 1352 2280 1358
rect 2228 1294 2280 1300
rect 1860 1216 1912 1222
rect 1860 1158 1912 1164
rect 1872 480 1900 1158
rect 2240 480 2268 1294
rect 2700 480 2728 3975
rect 2780 3946 2832 3952
rect 2792 1465 2820 3946
rect 2884 3738 2912 12396
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2976 11218 3004 11698
rect 2964 11212 3016 11218
rect 2964 11154 3016 11160
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 2976 9722 3004 10746
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2976 9178 3004 9386
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 2976 8537 3004 8570
rect 2962 8528 3018 8537
rect 2962 8463 3018 8472
rect 3068 8129 3096 12566
rect 3146 12336 3202 12345
rect 3146 12271 3202 12280
rect 3054 8120 3110 8129
rect 3054 8055 3110 8064
rect 3056 8016 3108 8022
rect 3056 7958 3108 7964
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 2976 5234 3004 7414
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 3068 4622 3096 7958
rect 3056 4616 3108 4622
rect 2962 4584 3018 4593
rect 3056 4558 3108 4564
rect 2962 4519 2964 4528
rect 3016 4519 3018 4528
rect 2964 4490 3016 4496
rect 3056 4004 3108 4010
rect 3056 3946 3108 3952
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 2872 3120 2924 3126
rect 2872 3062 2924 3068
rect 2884 2854 2912 3062
rect 2872 2848 2924 2854
rect 2872 2790 2924 2796
rect 2870 2680 2926 2689
rect 2870 2615 2872 2624
rect 2924 2615 2926 2624
rect 2872 2586 2924 2592
rect 2976 1766 3004 3878
rect 3068 3369 3096 3946
rect 3054 3360 3110 3369
rect 3054 3295 3110 3304
rect 3054 3088 3110 3097
rect 3054 3023 3110 3032
rect 2964 1760 3016 1766
rect 2964 1702 3016 1708
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 3068 480 3096 3023
rect 3160 513 3188 12271
rect 3252 3738 3280 14758
rect 3344 11898 3372 16730
rect 3790 16688 3846 16697
rect 3790 16623 3846 16632
rect 3421 16348 3717 16368
rect 3477 16346 3501 16348
rect 3557 16346 3581 16348
rect 3637 16346 3661 16348
rect 3499 16294 3501 16346
rect 3563 16294 3575 16346
rect 3637 16294 3639 16346
rect 3477 16292 3501 16294
rect 3557 16292 3581 16294
rect 3637 16292 3661 16294
rect 3421 16272 3717 16292
rect 3516 15904 3568 15910
rect 3514 15872 3516 15881
rect 3804 15892 3832 16623
rect 4080 16266 4108 16918
rect 4264 16522 4292 17274
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 4252 16516 4304 16522
rect 4252 16458 4304 16464
rect 4356 16425 4384 16526
rect 4342 16416 4398 16425
rect 4342 16351 4398 16360
rect 4080 16238 4292 16266
rect 4068 16176 4120 16182
rect 4066 16144 4068 16153
rect 4120 16144 4122 16153
rect 3976 16108 4028 16114
rect 4066 16079 4122 16088
rect 4160 16108 4212 16114
rect 3976 16050 4028 16056
rect 4160 16050 4212 16056
rect 3568 15872 3832 15892
rect 3570 15864 3832 15872
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3514 15807 3570 15816
rect 3424 15564 3476 15570
rect 3424 15506 3476 15512
rect 3436 15473 3464 15506
rect 3792 15496 3844 15502
rect 3422 15464 3478 15473
rect 3792 15438 3844 15444
rect 3422 15399 3478 15408
rect 3421 15260 3717 15280
rect 3477 15258 3501 15260
rect 3557 15258 3581 15260
rect 3637 15258 3661 15260
rect 3499 15206 3501 15258
rect 3563 15206 3575 15258
rect 3637 15206 3639 15258
rect 3477 15204 3501 15206
rect 3557 15204 3581 15206
rect 3637 15204 3661 15206
rect 3421 15184 3717 15204
rect 3804 15162 3832 15438
rect 3792 15156 3844 15162
rect 3792 15098 3844 15104
rect 3896 15008 3924 15846
rect 3804 14980 3924 15008
rect 3804 14385 3832 14980
rect 3790 14376 3846 14385
rect 3790 14311 3846 14320
rect 3421 14172 3717 14192
rect 3477 14170 3501 14172
rect 3557 14170 3581 14172
rect 3637 14170 3661 14172
rect 3499 14118 3501 14170
rect 3563 14118 3575 14170
rect 3637 14118 3639 14170
rect 3477 14116 3501 14118
rect 3557 14116 3581 14118
rect 3637 14116 3661 14118
rect 3421 14096 3717 14116
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 3436 13705 3464 13874
rect 3422 13696 3478 13705
rect 3422 13631 3478 13640
rect 3804 13462 3832 14311
rect 3882 14240 3938 14249
rect 3882 14175 3938 14184
rect 3896 13841 3924 14175
rect 3882 13832 3938 13841
rect 3882 13767 3938 13776
rect 3884 13728 3936 13734
rect 3884 13670 3936 13676
rect 3792 13456 3844 13462
rect 3792 13398 3844 13404
rect 3421 13084 3717 13104
rect 3477 13082 3501 13084
rect 3557 13082 3581 13084
rect 3637 13082 3661 13084
rect 3499 13030 3501 13082
rect 3563 13030 3575 13082
rect 3637 13030 3639 13082
rect 3477 13028 3501 13030
rect 3557 13028 3581 13030
rect 3637 13028 3661 13030
rect 3421 13008 3717 13028
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3421 11996 3717 12016
rect 3477 11994 3501 11996
rect 3557 11994 3581 11996
rect 3637 11994 3661 11996
rect 3499 11942 3501 11994
rect 3563 11942 3575 11994
rect 3637 11942 3639 11994
rect 3477 11940 3501 11942
rect 3557 11940 3581 11942
rect 3637 11940 3661 11942
rect 3421 11920 3717 11940
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 3700 11212 3752 11218
rect 3700 11154 3752 11160
rect 3712 11121 3740 11154
rect 3698 11112 3754 11121
rect 3332 11076 3384 11082
rect 3698 11047 3754 11056
rect 3332 11018 3384 11024
rect 3344 8430 3372 11018
rect 3421 10908 3717 10928
rect 3477 10906 3501 10908
rect 3557 10906 3581 10908
rect 3637 10906 3661 10908
rect 3499 10854 3501 10906
rect 3563 10854 3575 10906
rect 3637 10854 3639 10906
rect 3477 10852 3501 10854
rect 3557 10852 3581 10854
rect 3637 10852 3661 10854
rect 3421 10832 3717 10852
rect 3606 10704 3662 10713
rect 3606 10639 3662 10648
rect 3620 10169 3648 10639
rect 3606 10160 3662 10169
rect 3606 10095 3662 10104
rect 3804 9926 3832 12038
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3421 9820 3717 9840
rect 3477 9818 3501 9820
rect 3557 9818 3581 9820
rect 3637 9818 3661 9820
rect 3499 9766 3501 9818
rect 3563 9766 3575 9818
rect 3637 9766 3639 9818
rect 3477 9764 3501 9766
rect 3557 9764 3581 9766
rect 3637 9764 3661 9766
rect 3421 9744 3717 9764
rect 3606 9616 3662 9625
rect 3606 9551 3662 9560
rect 3620 9518 3648 9551
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3421 8732 3717 8752
rect 3477 8730 3501 8732
rect 3557 8730 3581 8732
rect 3637 8730 3661 8732
rect 3499 8678 3501 8730
rect 3563 8678 3575 8730
rect 3637 8678 3639 8730
rect 3477 8676 3501 8678
rect 3557 8676 3581 8678
rect 3637 8676 3661 8678
rect 3421 8656 3717 8676
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3804 8294 3832 8774
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3344 6186 3372 8230
rect 3790 7984 3846 7993
rect 3790 7919 3846 7928
rect 3421 7644 3717 7664
rect 3477 7642 3501 7644
rect 3557 7642 3581 7644
rect 3637 7642 3661 7644
rect 3499 7590 3501 7642
rect 3563 7590 3575 7642
rect 3637 7590 3639 7642
rect 3477 7588 3501 7590
rect 3557 7588 3581 7590
rect 3637 7588 3661 7590
rect 3421 7568 3717 7588
rect 3804 6730 3832 7919
rect 3792 6724 3844 6730
rect 3792 6666 3844 6672
rect 3421 6556 3717 6576
rect 3477 6554 3501 6556
rect 3557 6554 3581 6556
rect 3637 6554 3661 6556
rect 3499 6502 3501 6554
rect 3563 6502 3575 6554
rect 3637 6502 3639 6554
rect 3477 6500 3501 6502
rect 3557 6500 3581 6502
rect 3637 6500 3661 6502
rect 3421 6480 3717 6500
rect 3790 6352 3846 6361
rect 3790 6287 3846 6296
rect 3332 6180 3384 6186
rect 3332 6122 3384 6128
rect 3344 6089 3372 6122
rect 3330 6080 3386 6089
rect 3330 6015 3386 6024
rect 3421 5468 3717 5488
rect 3477 5466 3501 5468
rect 3557 5466 3581 5468
rect 3637 5466 3661 5468
rect 3499 5414 3501 5466
rect 3563 5414 3575 5466
rect 3637 5414 3639 5466
rect 3477 5412 3501 5414
rect 3557 5412 3581 5414
rect 3637 5412 3661 5414
rect 3421 5392 3717 5412
rect 3424 5296 3476 5302
rect 3424 5238 3476 5244
rect 3436 4826 3464 5238
rect 3516 5024 3568 5030
rect 3700 5024 3752 5030
rect 3568 4984 3648 5012
rect 3516 4966 3568 4972
rect 3514 4856 3570 4865
rect 3424 4820 3476 4826
rect 3514 4791 3570 4800
rect 3424 4762 3476 4768
rect 3528 4622 3556 4791
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 3516 4616 3568 4622
rect 3516 4558 3568 4564
rect 3344 4078 3372 4558
rect 3620 4554 3648 4984
rect 3700 4966 3752 4972
rect 3712 4826 3740 4966
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3608 4548 3660 4554
rect 3608 4490 3660 4496
rect 3421 4380 3717 4400
rect 3477 4378 3501 4380
rect 3557 4378 3581 4380
rect 3637 4378 3661 4380
rect 3499 4326 3501 4378
rect 3563 4326 3575 4378
rect 3637 4326 3639 4378
rect 3477 4324 3501 4326
rect 3557 4324 3581 4326
rect 3637 4324 3661 4326
rect 3421 4304 3717 4324
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3238 3632 3294 3641
rect 3238 3567 3240 3576
rect 3292 3567 3294 3576
rect 3240 3538 3292 3544
rect 3344 2650 3372 4014
rect 3606 3768 3662 3777
rect 3606 3703 3662 3712
rect 3620 3602 3648 3703
rect 3608 3596 3660 3602
rect 3608 3538 3660 3544
rect 3421 3292 3717 3312
rect 3477 3290 3501 3292
rect 3557 3290 3581 3292
rect 3637 3290 3661 3292
rect 3499 3238 3501 3290
rect 3563 3238 3575 3290
rect 3637 3238 3639 3290
rect 3477 3236 3501 3238
rect 3557 3236 3581 3238
rect 3637 3236 3661 3238
rect 3421 3216 3717 3236
rect 3700 2984 3752 2990
rect 3422 2952 3478 2961
rect 3804 2972 3832 6287
rect 3752 2944 3832 2972
rect 3700 2926 3752 2932
rect 3422 2887 3478 2896
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3436 2446 3464 2887
rect 3896 2854 3924 13670
rect 3988 11014 4016 16050
rect 4172 15688 4200 16050
rect 4080 15660 4200 15688
rect 4080 15502 4108 15660
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 4080 13818 4108 15302
rect 4264 14657 4292 16238
rect 4344 15904 4396 15910
rect 4344 15846 4396 15852
rect 4356 15337 4384 15846
rect 4342 15328 4398 15337
rect 4342 15263 4398 15272
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 4356 14906 4384 15098
rect 4448 15065 4476 17462
rect 4528 17060 4580 17066
rect 4528 17002 4580 17008
rect 4434 15056 4490 15065
rect 4434 14991 4490 15000
rect 4356 14890 4476 14906
rect 4356 14884 4488 14890
rect 4356 14878 4436 14884
rect 4436 14826 4488 14832
rect 4344 14816 4396 14822
rect 4344 14758 4396 14764
rect 4250 14648 4306 14657
rect 4250 14583 4306 14592
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 4264 14074 4292 14418
rect 4252 14068 4304 14074
rect 4252 14010 4304 14016
rect 4252 13932 4304 13938
rect 4252 13874 4304 13880
rect 4080 13802 4200 13818
rect 4080 13796 4212 13802
rect 4080 13790 4160 13796
rect 4160 13738 4212 13744
rect 4264 13705 4292 13874
rect 4066 13696 4122 13705
rect 4066 13631 4122 13640
rect 4250 13696 4306 13705
rect 4250 13631 4306 13640
rect 4080 12220 4108 13631
rect 4158 13560 4214 13569
rect 4158 13495 4214 13504
rect 4172 12374 4200 13495
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 4160 12368 4212 12374
rect 4160 12310 4212 12316
rect 4080 12192 4200 12220
rect 4066 11928 4122 11937
rect 4066 11863 4122 11872
rect 4080 11694 4108 11863
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 4080 10674 4108 11086
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 4172 10554 4200 12192
rect 3988 10526 4200 10554
rect 3988 4758 4016 10526
rect 4066 10432 4122 10441
rect 4264 10418 4292 13262
rect 4356 12646 4384 14758
rect 4436 14544 4488 14550
rect 4434 14512 4436 14521
rect 4488 14512 4490 14521
rect 4434 14447 4490 14456
rect 4436 14408 4488 14414
rect 4436 14350 4488 14356
rect 4448 12986 4476 14350
rect 4540 14006 4568 17002
rect 4632 16250 4660 19520
rect 5000 17542 5028 19520
rect 4988 17536 5040 17542
rect 4988 17478 5040 17484
rect 5172 17196 5224 17202
rect 5172 17138 5224 17144
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 4988 17060 5040 17066
rect 4988 17002 5040 17008
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 4712 16176 4764 16182
rect 4712 16118 4764 16124
rect 4724 15881 4752 16118
rect 4710 15872 4766 15881
rect 4710 15807 4766 15816
rect 4710 15736 4766 15745
rect 4710 15671 4766 15680
rect 4724 15502 4752 15671
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4632 14793 4660 15438
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 4618 14784 4674 14793
rect 4618 14719 4674 14728
rect 4620 14544 4672 14550
rect 4620 14486 4672 14492
rect 4528 14000 4580 14006
rect 4528 13942 4580 13948
rect 4632 13841 4660 14486
rect 4618 13832 4674 13841
rect 4618 13767 4674 13776
rect 4724 13716 4752 14962
rect 4816 14618 4844 16934
rect 4894 16824 4950 16833
rect 4894 16759 4950 16768
rect 4908 16658 4936 16759
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 4894 16416 4950 16425
rect 4894 16351 4950 16360
rect 4908 16114 4936 16351
rect 5000 16182 5028 17002
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 4988 16176 5040 16182
rect 4988 16118 5040 16124
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 4908 16017 4936 16050
rect 4894 16008 4950 16017
rect 4894 15943 4950 15952
rect 4986 15872 5042 15881
rect 4986 15807 5042 15816
rect 4896 15496 4948 15502
rect 4896 15438 4948 15444
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 4908 14498 4936 15438
rect 4816 14470 4936 14498
rect 4816 13870 4844 14470
rect 5000 14056 5028 15807
rect 5092 14890 5120 16934
rect 5080 14884 5132 14890
rect 5080 14826 5132 14832
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 5092 14278 5120 14418
rect 5080 14272 5132 14278
rect 5080 14214 5132 14220
rect 4908 14028 5028 14056
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 4632 13688 4752 13716
rect 4528 13252 4580 13258
rect 4528 13194 4580 13200
rect 4540 12986 4568 13194
rect 4436 12980 4488 12986
rect 4436 12922 4488 12928
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4344 12640 4396 12646
rect 4344 12582 4396 12588
rect 4344 12164 4396 12170
rect 4344 12106 4396 12112
rect 4122 10390 4292 10418
rect 4066 10367 4122 10376
rect 4068 10056 4120 10062
rect 4066 10024 4068 10033
rect 4120 10024 4122 10033
rect 4066 9959 4122 9968
rect 4080 9722 4108 9959
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 4080 8974 4108 9658
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4080 8634 4108 8910
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4080 8498 4108 8570
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 4172 8401 4200 8978
rect 4158 8392 4214 8401
rect 4158 8327 4214 8336
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 4172 8090 4200 8230
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4068 8016 4120 8022
rect 4068 7958 4120 7964
rect 4080 5710 4108 7958
rect 4172 5930 4200 8026
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4264 7410 4292 7822
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 4172 5902 4292 5930
rect 4158 5808 4214 5817
rect 4158 5743 4214 5752
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4080 5234 4108 5646
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 4066 5128 4122 5137
rect 4066 5063 4122 5072
rect 3976 4752 4028 4758
rect 3976 4694 4028 4700
rect 4080 4690 4108 5063
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 3974 4312 4030 4321
rect 3974 4247 4030 4256
rect 3988 3670 4016 4247
rect 3976 3664 4028 3670
rect 3976 3606 4028 3612
rect 3974 3360 4030 3369
rect 3974 3295 4030 3304
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3988 2650 4016 3295
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 3700 2440 3752 2446
rect 4080 2394 4108 4422
rect 4172 3670 4200 5743
rect 4264 4214 4292 5902
rect 4252 4208 4304 4214
rect 4252 4150 4304 4156
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4160 3664 4212 3670
rect 4160 3606 4212 3612
rect 4264 3058 4292 3878
rect 4356 3194 4384 12106
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4436 11280 4488 11286
rect 4436 11222 4488 11228
rect 4448 10724 4476 11222
rect 4540 11098 4568 11698
rect 4632 11218 4660 13688
rect 4710 13424 4766 13433
rect 4710 13359 4766 13368
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4540 11070 4660 11098
rect 4528 10736 4580 10742
rect 4448 10696 4528 10724
rect 4528 10678 4580 10684
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4448 9654 4476 10406
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4540 10033 4568 10202
rect 4526 10024 4582 10033
rect 4526 9959 4582 9968
rect 4632 9897 4660 11070
rect 4618 9888 4674 9897
rect 4618 9823 4674 9832
rect 4436 9648 4488 9654
rect 4436 9590 4488 9596
rect 4528 7744 4580 7750
rect 4528 7686 4580 7692
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4436 6860 4488 6866
rect 4436 6802 4488 6808
rect 4448 6118 4476 6802
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4436 5840 4488 5846
rect 4434 5808 4436 5817
rect 4488 5808 4490 5817
rect 4434 5743 4490 5752
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4448 4758 4476 5510
rect 4540 5166 4568 7686
rect 4632 7546 4660 7686
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 4436 4752 4488 4758
rect 4632 4729 4660 7346
rect 4436 4694 4488 4700
rect 4618 4720 4674 4729
rect 4618 4655 4674 4664
rect 4724 4321 4752 13359
rect 4804 13252 4856 13258
rect 4804 13194 4856 13200
rect 4816 12782 4844 13194
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4816 11762 4844 12718
rect 4908 12442 4936 14028
rect 4986 13968 5042 13977
rect 4986 13903 5042 13912
rect 5000 13870 5028 13903
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 5000 13258 5028 13806
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 4988 13252 5040 13258
rect 4988 13194 5040 13200
rect 4896 12436 4948 12442
rect 4896 12378 4948 12384
rect 4896 12232 4948 12238
rect 4894 12200 4896 12209
rect 4948 12200 4950 12209
rect 4894 12135 4950 12144
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 4804 11620 4856 11626
rect 4804 11562 4856 11568
rect 4816 5302 4844 11562
rect 5092 11200 5120 13262
rect 5184 11626 5212 17138
rect 5276 15162 5304 17138
rect 5356 17128 5408 17134
rect 5356 17070 5408 17076
rect 5368 15366 5396 17070
rect 5460 15978 5488 19520
rect 5632 16788 5684 16794
rect 5632 16730 5684 16736
rect 5448 15972 5500 15978
rect 5448 15914 5500 15920
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5460 15434 5488 15506
rect 5552 15473 5580 15642
rect 5538 15464 5594 15473
rect 5448 15428 5500 15434
rect 5538 15399 5594 15408
rect 5448 15370 5500 15376
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5264 15156 5316 15162
rect 5264 15098 5316 15104
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 5356 15088 5408 15094
rect 5356 15030 5408 15036
rect 5264 14884 5316 14890
rect 5264 14826 5316 14832
rect 5276 14521 5304 14826
rect 5262 14512 5318 14521
rect 5262 14447 5318 14456
rect 5368 14396 5396 15030
rect 5276 14368 5396 14396
rect 5276 12220 5304 14368
rect 5460 13569 5488 15098
rect 5552 14958 5580 15302
rect 5644 15162 5672 16730
rect 5724 16516 5776 16522
rect 5724 16458 5776 16464
rect 5632 15156 5684 15162
rect 5632 15098 5684 15104
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 5644 14346 5672 14894
rect 5736 14618 5764 16458
rect 5828 16017 5856 19520
rect 6092 17944 6144 17950
rect 6092 17886 6144 17892
rect 6104 17202 6132 17886
rect 6288 17626 6316 19520
rect 6288 17598 6500 17626
rect 6276 17536 6328 17542
rect 6276 17478 6328 17484
rect 6368 17536 6420 17542
rect 6368 17478 6420 17484
rect 6092 17196 6144 17202
rect 6092 17138 6144 17144
rect 5886 16892 6182 16912
rect 5942 16890 5966 16892
rect 6022 16890 6046 16892
rect 6102 16890 6126 16892
rect 5964 16838 5966 16890
rect 6028 16838 6040 16890
rect 6102 16838 6104 16890
rect 5942 16836 5966 16838
rect 6022 16836 6046 16838
rect 6102 16836 6126 16838
rect 5886 16816 6182 16836
rect 6288 16794 6316 17478
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 6380 16658 6408 17478
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 5814 16008 5870 16017
rect 5814 15943 5870 15952
rect 6276 15904 6328 15910
rect 6274 15872 6276 15881
rect 6328 15872 6330 15881
rect 5886 15804 6182 15824
rect 6274 15807 6330 15816
rect 5942 15802 5966 15804
rect 6022 15802 6046 15804
rect 6102 15802 6126 15804
rect 5964 15750 5966 15802
rect 6028 15750 6040 15802
rect 6102 15750 6104 15802
rect 5942 15748 5966 15750
rect 6022 15748 6046 15750
rect 6102 15748 6126 15750
rect 5886 15728 6182 15748
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 6276 14816 6328 14822
rect 6276 14758 6328 14764
rect 6368 14816 6420 14822
rect 6472 14793 6500 17598
rect 6656 17202 6684 19520
rect 7024 17678 7052 19520
rect 7484 18086 7512 19520
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6736 16992 6788 16998
rect 6734 16960 6736 16969
rect 6788 16960 6790 16969
rect 6734 16895 6790 16904
rect 7116 16794 7144 17818
rect 7852 17270 7880 19520
rect 8312 18222 8340 19520
rect 8300 18216 8352 18222
rect 8300 18158 8352 18164
rect 7932 17808 7984 17814
rect 7932 17750 7984 17756
rect 7840 17264 7892 17270
rect 7286 17232 7342 17241
rect 7840 17206 7892 17212
rect 7286 17167 7342 17176
rect 7380 17196 7432 17202
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 7104 16788 7156 16794
rect 7104 16730 7156 16736
rect 6748 16454 6776 16730
rect 6736 16448 6788 16454
rect 6736 16390 6788 16396
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 6736 16108 6788 16114
rect 6736 16050 6788 16056
rect 6642 15464 6698 15473
rect 6642 15399 6698 15408
rect 6368 14758 6420 14764
rect 6458 14784 6514 14793
rect 5828 14618 5856 14758
rect 5886 14716 6182 14736
rect 5942 14714 5966 14716
rect 6022 14714 6046 14716
rect 6102 14714 6126 14716
rect 5964 14662 5966 14714
rect 6028 14662 6040 14714
rect 6102 14662 6104 14714
rect 5942 14660 5966 14662
rect 6022 14660 6046 14662
rect 6102 14660 6126 14662
rect 5886 14640 6182 14660
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5908 14544 5960 14550
rect 5908 14486 5960 14492
rect 5724 14476 5776 14482
rect 5724 14418 5776 14424
rect 5632 14340 5684 14346
rect 5632 14282 5684 14288
rect 5538 13696 5594 13705
rect 5538 13631 5594 13640
rect 5446 13560 5502 13569
rect 5446 13495 5502 13504
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5354 12472 5410 12481
rect 5354 12407 5410 12416
rect 5368 12374 5396 12407
rect 5356 12368 5408 12374
rect 5356 12310 5408 12316
rect 5356 12232 5408 12238
rect 5276 12192 5356 12220
rect 5356 12174 5408 12180
rect 5172 11620 5224 11626
rect 5172 11562 5224 11568
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5000 11172 5120 11200
rect 4894 10296 4950 10305
rect 4894 10231 4950 10240
rect 4908 9761 4936 10231
rect 5000 10010 5028 11172
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 5092 10130 5120 11018
rect 5172 11008 5224 11014
rect 5172 10950 5224 10956
rect 5184 10810 5212 10950
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5184 10418 5212 10746
rect 5276 10538 5304 11290
rect 5368 11121 5396 12174
rect 5460 11801 5488 13330
rect 5446 11792 5502 11801
rect 5446 11727 5502 11736
rect 5446 11384 5502 11393
rect 5446 11319 5448 11328
rect 5500 11319 5502 11328
rect 5448 11290 5500 11296
rect 5354 11112 5410 11121
rect 5354 11047 5356 11056
rect 5408 11047 5410 11056
rect 5356 11018 5408 11024
rect 5368 10987 5396 11018
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 5368 10418 5396 10474
rect 5184 10390 5396 10418
rect 5460 10266 5488 10950
rect 5552 10810 5580 13631
rect 5632 12640 5684 12646
rect 5630 12608 5632 12617
rect 5684 12608 5686 12617
rect 5630 12543 5686 12552
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 5000 9982 5120 10010
rect 4894 9752 4950 9761
rect 4894 9687 4950 9696
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4908 8838 4936 9318
rect 5092 8945 5120 9982
rect 5354 9888 5410 9897
rect 5354 9823 5410 9832
rect 5078 8936 5134 8945
rect 5078 8871 5134 8880
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4896 8492 4948 8498
rect 4948 8452 5028 8480
rect 4896 8434 4948 8440
rect 5000 7342 5028 8452
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 5184 8022 5212 8298
rect 5172 8016 5224 8022
rect 5172 7958 5224 7964
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 5170 7576 5226 7585
rect 5276 7546 5304 7754
rect 5170 7511 5172 7520
rect 5224 7511 5226 7520
rect 5264 7540 5316 7546
rect 5172 7482 5224 7488
rect 5264 7482 5316 7488
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 5000 7002 5028 7278
rect 5264 7200 5316 7206
rect 5078 7168 5134 7177
rect 5264 7142 5316 7148
rect 5078 7103 5134 7112
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4908 5914 4936 6598
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4804 5296 4856 5302
rect 4804 5238 4856 5244
rect 4804 5160 4856 5166
rect 4804 5102 4856 5108
rect 4816 4690 4844 5102
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4710 4312 4766 4321
rect 4710 4247 4766 4256
rect 4816 4196 4844 4422
rect 4724 4168 4844 4196
rect 4528 4140 4580 4146
rect 4580 4100 4660 4128
rect 4528 4082 4580 4088
rect 4436 3936 4488 3942
rect 4436 3878 4488 3884
rect 4528 3936 4580 3942
rect 4528 3878 4580 3884
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4250 2952 4306 2961
rect 4250 2887 4306 2896
rect 3752 2388 3832 2394
rect 3700 2382 3832 2388
rect 3252 1465 3280 2382
rect 3712 2366 3832 2382
rect 4080 2366 4200 2394
rect 3804 2310 3832 2366
rect 3792 2304 3844 2310
rect 3792 2246 3844 2252
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 3421 2204 3717 2224
rect 3477 2202 3501 2204
rect 3557 2202 3581 2204
rect 3637 2202 3661 2204
rect 3499 2150 3501 2202
rect 3563 2150 3575 2202
rect 3637 2150 3639 2202
rect 3477 2148 3501 2150
rect 3557 2148 3581 2150
rect 3637 2148 3661 2150
rect 3421 2128 3717 2148
rect 4080 1873 4108 2246
rect 4172 1902 4200 2366
rect 4264 2310 4292 2887
rect 4344 2848 4396 2854
rect 4342 2816 4344 2825
rect 4396 2816 4398 2825
rect 4342 2751 4398 2760
rect 4252 2304 4304 2310
rect 4252 2246 4304 2252
rect 4160 1896 4212 1902
rect 4066 1864 4122 1873
rect 4160 1838 4212 1844
rect 4066 1799 4122 1808
rect 3882 1728 3938 1737
rect 3882 1663 3938 1672
rect 3514 1592 3570 1601
rect 3514 1527 3570 1536
rect 3238 1456 3294 1465
rect 3238 1391 3294 1400
rect 3146 504 3202 513
rect 202 0 258 480
rect 570 0 626 480
rect 1030 0 1086 480
rect 1398 0 1454 480
rect 1858 0 1914 480
rect 2226 0 2282 480
rect 2686 0 2742 480
rect 3054 0 3110 480
rect 3528 480 3556 1527
rect 3896 480 3924 1663
rect 4342 1184 4398 1193
rect 4342 1119 4398 1128
rect 4356 480 4384 1119
rect 4448 950 4476 3878
rect 4540 3738 4568 3878
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4540 3194 4568 3470
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4632 3058 4660 4100
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4724 2922 4752 4168
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4816 3942 4844 4014
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4802 3632 4858 3641
rect 4802 3567 4858 3576
rect 4816 3466 4844 3567
rect 4804 3460 4856 3466
rect 4804 3402 4856 3408
rect 4712 2916 4764 2922
rect 4712 2858 4764 2864
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 4816 2417 4844 2790
rect 4802 2408 4858 2417
rect 4802 2343 4858 2352
rect 4908 1834 4936 5510
rect 5000 4826 5028 5646
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4986 4720 5042 4729
rect 4986 4655 5042 4664
rect 5000 3534 5028 4655
rect 5092 4321 5120 7103
rect 5276 6458 5304 7142
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 5170 5672 5226 5681
rect 5170 5607 5226 5616
rect 5078 4312 5134 4321
rect 5078 4247 5134 4256
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 5000 2145 5028 3334
rect 4986 2136 5042 2145
rect 4986 2071 5042 2080
rect 4896 1828 4948 1834
rect 4896 1770 4948 1776
rect 4712 1148 4764 1154
rect 4712 1090 4764 1096
rect 4436 944 4488 950
rect 4436 886 4488 892
rect 4724 480 4752 1090
rect 5184 480 5212 5607
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 5276 4842 5304 5306
rect 5368 5001 5396 9823
rect 5460 9042 5488 10202
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5552 8809 5580 9386
rect 5538 8800 5594 8809
rect 5538 8735 5594 8744
rect 5552 8430 5580 8735
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5460 7002 5488 7822
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5460 6866 5488 6938
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5460 5914 5488 6190
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5354 4992 5410 5001
rect 5354 4927 5410 4936
rect 5276 4826 5396 4842
rect 5276 4820 5408 4826
rect 5276 4814 5356 4820
rect 5356 4762 5408 4768
rect 5460 4706 5488 5850
rect 5552 5710 5580 7890
rect 5644 6905 5672 12378
rect 5736 12238 5764 14418
rect 5816 14272 5868 14278
rect 5920 14249 5948 14486
rect 5816 14214 5868 14220
rect 5906 14240 5962 14249
rect 5828 13025 5856 14214
rect 5906 14175 5962 14184
rect 6288 13870 6316 14758
rect 6276 13864 6328 13870
rect 6276 13806 6328 13812
rect 6276 13728 6328 13734
rect 6276 13670 6328 13676
rect 5886 13628 6182 13648
rect 5942 13626 5966 13628
rect 6022 13626 6046 13628
rect 6102 13626 6126 13628
rect 5964 13574 5966 13626
rect 6028 13574 6040 13626
rect 6102 13574 6104 13626
rect 5942 13572 5966 13574
rect 6022 13572 6046 13574
rect 6102 13572 6126 13574
rect 5886 13552 6182 13572
rect 6288 13462 6316 13670
rect 6380 13530 6408 14758
rect 6458 14719 6514 14728
rect 6460 14340 6512 14346
rect 6460 14282 6512 14288
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 6276 13456 6328 13462
rect 6276 13398 6328 13404
rect 5814 13016 5870 13025
rect 5814 12951 5870 12960
rect 5814 12744 5870 12753
rect 5814 12679 5870 12688
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5722 11928 5778 11937
rect 5722 11863 5778 11872
rect 5736 8906 5764 11863
rect 5828 11354 5856 12679
rect 5886 12540 6182 12560
rect 5942 12538 5966 12540
rect 6022 12538 6046 12540
rect 6102 12538 6126 12540
rect 5964 12486 5966 12538
rect 6028 12486 6040 12538
rect 6102 12486 6104 12538
rect 5942 12484 5966 12486
rect 6022 12484 6046 12486
rect 6102 12484 6126 12486
rect 5886 12464 6182 12484
rect 6288 11694 6316 13398
rect 6380 13394 6408 13466
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6472 12753 6500 14282
rect 6550 13968 6606 13977
rect 6550 13903 6606 13912
rect 6458 12744 6514 12753
rect 6458 12679 6514 12688
rect 6458 12472 6514 12481
rect 6458 12407 6460 12416
rect 6512 12407 6514 12416
rect 6460 12378 6512 12384
rect 6564 12374 6592 13903
rect 6656 13705 6684 15399
rect 6642 13696 6698 13705
rect 6642 13631 6698 13640
rect 6748 13569 6776 16050
rect 6826 15736 6882 15745
rect 6826 15671 6882 15680
rect 6840 15638 6868 15671
rect 6828 15632 6880 15638
rect 6828 15574 6880 15580
rect 6828 15428 6880 15434
rect 6828 15370 6880 15376
rect 6840 15042 6868 15370
rect 6932 15201 6960 16390
rect 7024 15638 7052 16390
rect 7104 16108 7156 16114
rect 7208 16096 7236 17070
rect 7300 16658 7328 17167
rect 7656 17196 7708 17202
rect 7380 17138 7432 17144
rect 7576 17156 7656 17184
rect 7288 16652 7340 16658
rect 7288 16594 7340 16600
rect 7208 16068 7328 16096
rect 7104 16050 7156 16056
rect 7012 15632 7064 15638
rect 7012 15574 7064 15580
rect 6918 15192 6974 15201
rect 6918 15127 6974 15136
rect 6840 15014 6960 15042
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6840 14414 6868 14894
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 6840 13802 6868 14350
rect 6828 13796 6880 13802
rect 6828 13738 6880 13744
rect 6734 13560 6790 13569
rect 6734 13495 6790 13504
rect 6644 13388 6696 13394
rect 6644 13330 6696 13336
rect 6656 12442 6684 13330
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6552 12368 6604 12374
rect 6552 12310 6604 12316
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6368 11824 6420 11830
rect 6368 11766 6420 11772
rect 6276 11688 6328 11694
rect 6276 11630 6328 11636
rect 6274 11520 6330 11529
rect 5886 11452 6182 11472
rect 6274 11455 6330 11464
rect 5942 11450 5966 11452
rect 6022 11450 6046 11452
rect 6102 11450 6126 11452
rect 5964 11398 5966 11450
rect 6028 11398 6040 11450
rect 6102 11398 6104 11450
rect 5942 11396 5966 11398
rect 6022 11396 6046 11398
rect 6102 11396 6126 11398
rect 5886 11376 6182 11396
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 6000 11280 6052 11286
rect 6288 11268 6316 11455
rect 6052 11240 6316 11268
rect 6000 11222 6052 11228
rect 6380 11150 6408 11766
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 5886 10364 6182 10384
rect 5942 10362 5966 10364
rect 6022 10362 6046 10364
rect 6102 10362 6126 10364
rect 5964 10310 5966 10362
rect 6028 10310 6040 10362
rect 6102 10310 6104 10362
rect 5942 10308 5966 10310
rect 6022 10308 6046 10310
rect 6102 10308 6126 10310
rect 5886 10288 6182 10308
rect 6288 10198 6316 10746
rect 6380 10470 6408 10746
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6276 10192 6328 10198
rect 6276 10134 6328 10140
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 5920 9926 5948 9998
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 5920 9722 5948 9862
rect 5998 9752 6054 9761
rect 5908 9716 5960 9722
rect 5998 9687 6000 9696
rect 5908 9658 5960 9664
rect 6052 9687 6054 9696
rect 6000 9658 6052 9664
rect 6276 9648 6328 9654
rect 6274 9616 6276 9625
rect 6328 9616 6330 9625
rect 6274 9551 6330 9560
rect 5816 9444 5868 9450
rect 5816 9386 5868 9392
rect 6276 9444 6328 9450
rect 6276 9386 6328 9392
rect 5828 9110 5856 9386
rect 5886 9276 6182 9296
rect 5942 9274 5966 9276
rect 6022 9274 6046 9276
rect 6102 9274 6126 9276
rect 5964 9222 5966 9274
rect 6028 9222 6040 9274
rect 6102 9222 6104 9274
rect 5942 9220 5966 9222
rect 6022 9220 6046 9222
rect 6102 9220 6126 9222
rect 5886 9200 6182 9220
rect 6288 9110 6316 9386
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 6000 9104 6052 9110
rect 6000 9046 6052 9052
rect 6276 9104 6328 9110
rect 6276 9046 6328 9052
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 6012 8566 6040 9046
rect 6472 8838 6500 12174
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5828 7206 5856 8298
rect 5886 8188 6182 8208
rect 5942 8186 5966 8188
rect 6022 8186 6046 8188
rect 6102 8186 6126 8188
rect 5964 8134 5966 8186
rect 6028 8134 6040 8186
rect 6102 8134 6104 8186
rect 5942 8132 5966 8134
rect 6022 8132 6046 8134
rect 6102 8132 6126 8134
rect 5886 8112 6182 8132
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 5998 7440 6054 7449
rect 6104 7410 6132 7686
rect 5998 7375 6054 7384
rect 6092 7404 6144 7410
rect 6012 7342 6040 7375
rect 6092 7346 6144 7352
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 6196 7274 6224 7686
rect 6184 7268 6236 7274
rect 6184 7210 6236 7216
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5886 7100 6182 7120
rect 5942 7098 5966 7100
rect 6022 7098 6046 7100
rect 6102 7098 6126 7100
rect 5964 7046 5966 7098
rect 6028 7046 6040 7098
rect 6102 7046 6104 7098
rect 5942 7044 5966 7046
rect 6022 7044 6046 7046
rect 6102 7044 6126 7046
rect 5886 7024 6182 7044
rect 5630 6896 5686 6905
rect 5630 6831 5686 6840
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5644 6458 5672 6734
rect 5814 6488 5870 6497
rect 5632 6452 5684 6458
rect 5814 6423 5870 6432
rect 5632 6394 5684 6400
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5552 5370 5580 5646
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5644 5166 5672 6394
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 5736 6118 5764 6190
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 5736 5710 5764 5850
rect 5828 5794 5856 6423
rect 5886 6012 6182 6032
rect 5942 6010 5966 6012
rect 6022 6010 6046 6012
rect 6102 6010 6126 6012
rect 5964 5958 5966 6010
rect 6028 5958 6040 6010
rect 6102 5958 6104 6010
rect 5942 5956 5966 5958
rect 6022 5956 6046 5958
rect 6102 5956 6126 5958
rect 5886 5936 6182 5956
rect 6092 5840 6144 5846
rect 5828 5788 6092 5794
rect 5828 5782 6144 5788
rect 5828 5766 6132 5782
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 6104 5166 6132 5766
rect 5632 5160 5684 5166
rect 6092 5160 6144 5166
rect 5684 5108 5856 5114
rect 5632 5102 5856 5108
rect 6092 5102 6144 5108
rect 5644 5086 5856 5102
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5276 4690 5488 4706
rect 5264 4684 5488 4690
rect 5316 4678 5488 4684
rect 5264 4626 5316 4632
rect 5276 2106 5304 4626
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5448 4548 5500 4554
rect 5448 4490 5500 4496
rect 5368 4457 5396 4490
rect 5354 4448 5410 4457
rect 5354 4383 5410 4392
rect 5356 4276 5408 4282
rect 5460 4264 5488 4490
rect 5552 4282 5580 4966
rect 5736 4865 5764 4966
rect 5722 4856 5778 4865
rect 5722 4791 5778 4800
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5644 4282 5672 4626
rect 5828 4622 5856 5086
rect 5886 4924 6182 4944
rect 5942 4922 5966 4924
rect 6022 4922 6046 4924
rect 6102 4922 6126 4924
rect 5964 4870 5966 4922
rect 6028 4870 6040 4922
rect 6102 4870 6104 4922
rect 5942 4868 5966 4870
rect 6022 4868 6046 4870
rect 6102 4868 6126 4870
rect 5886 4848 6182 4868
rect 6288 4758 6316 8502
rect 6472 7188 6500 8774
rect 6564 7721 6592 12310
rect 6656 12238 6684 12378
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6748 12170 6776 13495
rect 6840 12850 6868 13738
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6736 12164 6788 12170
rect 6736 12106 6788 12112
rect 6840 11762 6868 12786
rect 6932 12345 6960 15014
rect 7010 14784 7066 14793
rect 7010 14719 7066 14728
rect 7024 13841 7052 14719
rect 7116 14482 7144 16050
rect 7196 15972 7248 15978
rect 7196 15914 7248 15920
rect 7208 15706 7236 15914
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7196 15496 7248 15502
rect 7196 15438 7248 15444
rect 7208 14890 7236 15438
rect 7196 14884 7248 14890
rect 7196 14826 7248 14832
rect 7208 14793 7236 14826
rect 7194 14784 7250 14793
rect 7194 14719 7250 14728
rect 7194 14648 7250 14657
rect 7194 14583 7250 14592
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 7116 13870 7144 14418
rect 7208 14113 7236 14583
rect 7194 14104 7250 14113
rect 7194 14039 7250 14048
rect 7104 13864 7156 13870
rect 7010 13832 7066 13841
rect 7104 13806 7156 13812
rect 7010 13767 7066 13776
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 7024 12714 7052 13126
rect 7116 12986 7144 13670
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 7208 13433 7236 13466
rect 7194 13424 7250 13433
rect 7300 13394 7328 16068
rect 7392 15366 7420 17138
rect 7472 16992 7524 16998
rect 7472 16934 7524 16940
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 7484 13938 7512 16934
rect 7576 14890 7604 17156
rect 7656 17138 7708 17144
rect 7748 16992 7800 16998
rect 7748 16934 7800 16940
rect 7760 16046 7788 16934
rect 7944 16726 7972 17750
rect 8206 17640 8262 17649
rect 8206 17575 8262 17584
rect 8220 17252 8248 17575
rect 8352 17436 8648 17456
rect 8408 17434 8432 17436
rect 8488 17434 8512 17436
rect 8568 17434 8592 17436
rect 8430 17382 8432 17434
rect 8494 17382 8506 17434
rect 8568 17382 8570 17434
rect 8408 17380 8432 17382
rect 8488 17380 8512 17382
rect 8568 17380 8592 17382
rect 8352 17360 8648 17380
rect 8220 17224 8340 17252
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 7932 16720 7984 16726
rect 7932 16662 7984 16668
rect 7932 16584 7984 16590
rect 7932 16526 7984 16532
rect 7944 16425 7972 16526
rect 7930 16416 7986 16425
rect 7930 16351 7986 16360
rect 7748 16040 7800 16046
rect 7748 15982 7800 15988
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7852 15892 7880 15982
rect 7760 15881 7880 15892
rect 7746 15872 7880 15881
rect 7802 15864 7880 15872
rect 7746 15807 7802 15816
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7564 14272 7616 14278
rect 7564 14214 7616 14220
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7576 13818 7604 14214
rect 7392 13790 7604 13818
rect 7194 13359 7250 13368
rect 7288 13388 7340 13394
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7208 12889 7236 13359
rect 7288 13330 7340 13336
rect 7392 13138 7420 13790
rect 7668 13530 7696 15506
rect 7760 13734 7788 15807
rect 8036 15434 8064 17138
rect 8114 16824 8170 16833
rect 8114 16759 8170 16768
rect 8128 16658 8156 16759
rect 8312 16726 8340 17224
rect 8680 17184 8708 19520
rect 8852 18148 8904 18154
rect 9048 18136 9076 19520
rect 9048 18108 9168 18136
rect 8852 18090 8904 18096
rect 8588 17156 8708 17184
rect 8482 17096 8538 17105
rect 8482 17031 8484 17040
rect 8536 17031 8538 17040
rect 8484 17002 8536 17008
rect 8300 16720 8352 16726
rect 8588 16697 8616 17156
rect 8668 17060 8720 17066
rect 8668 17002 8720 17008
rect 8680 16810 8708 17002
rect 8680 16782 8800 16810
rect 8300 16662 8352 16668
rect 8574 16688 8630 16697
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8208 16652 8260 16658
rect 8574 16623 8630 16632
rect 8208 16594 8260 16600
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 7840 15428 7892 15434
rect 7840 15370 7892 15376
rect 8024 15428 8076 15434
rect 8024 15370 8076 15376
rect 7748 13728 7800 13734
rect 7748 13670 7800 13676
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 7564 13456 7616 13462
rect 7564 13398 7616 13404
rect 7300 13110 7420 13138
rect 7194 12880 7250 12889
rect 7194 12815 7250 12824
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 7300 12594 7328 13110
rect 7024 12566 7328 12594
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 6918 12336 6974 12345
rect 6918 12271 6974 12280
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6656 9625 6684 11698
rect 6734 11384 6790 11393
rect 6734 11319 6790 11328
rect 6748 11286 6776 11319
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6840 10674 6868 11698
rect 6932 10985 6960 12174
rect 6918 10976 6974 10985
rect 6918 10911 6974 10920
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 6642 9616 6698 9625
rect 6642 9551 6698 9560
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6932 8430 6960 9318
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6748 7886 6776 8366
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6550 7712 6606 7721
rect 6550 7647 6606 7656
rect 6748 7342 6776 7822
rect 6840 7478 6868 7890
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 7024 7392 7052 12566
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7116 9994 7144 12378
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 7208 9450 7236 12242
rect 7286 12200 7342 12209
rect 7286 12135 7342 12144
rect 7300 9874 7328 12135
rect 7392 10538 7420 12582
rect 7472 12368 7524 12374
rect 7472 12310 7524 12316
rect 7484 12209 7512 12310
rect 7470 12200 7526 12209
rect 7470 12135 7526 12144
rect 7576 11898 7604 13398
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7668 11354 7696 13126
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7484 10849 7512 11086
rect 7470 10840 7526 10849
rect 7470 10775 7526 10784
rect 7760 10724 7788 13262
rect 7852 12889 7880 15370
rect 7932 15360 7984 15366
rect 7932 15302 7984 15308
rect 7944 15162 7972 15302
rect 7932 15156 7984 15162
rect 7932 15098 7984 15104
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 7944 14482 7972 14554
rect 7932 14476 7984 14482
rect 7932 14418 7984 14424
rect 8036 14278 8064 15370
rect 8128 14618 8156 15438
rect 8116 14612 8168 14618
rect 8116 14554 8168 14560
rect 8116 14340 8168 14346
rect 8116 14282 8168 14288
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 7932 13728 7984 13734
rect 7932 13670 7984 13676
rect 7944 13161 7972 13670
rect 8128 13394 8156 14282
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 8116 13252 8168 13258
rect 8116 13194 8168 13200
rect 7930 13152 7986 13161
rect 7930 13087 7986 13096
rect 8128 12986 8156 13194
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 7838 12880 7894 12889
rect 7838 12815 7894 12824
rect 7838 12472 7894 12481
rect 8220 12424 8248 16594
rect 8352 16348 8648 16368
rect 8408 16346 8432 16348
rect 8488 16346 8512 16348
rect 8568 16346 8592 16348
rect 8430 16294 8432 16346
rect 8494 16294 8506 16346
rect 8568 16294 8570 16346
rect 8408 16292 8432 16294
rect 8488 16292 8512 16294
rect 8568 16292 8592 16294
rect 8352 16272 8648 16292
rect 8668 15972 8720 15978
rect 8668 15914 8720 15920
rect 8352 15260 8648 15280
rect 8408 15258 8432 15260
rect 8488 15258 8512 15260
rect 8568 15258 8592 15260
rect 8430 15206 8432 15258
rect 8494 15206 8506 15258
rect 8568 15206 8570 15258
rect 8408 15204 8432 15206
rect 8488 15204 8512 15206
rect 8568 15204 8592 15206
rect 8352 15184 8648 15204
rect 8680 15094 8708 15914
rect 8772 15722 8800 16782
rect 8864 16522 8892 18090
rect 8944 17944 8996 17950
rect 8942 17912 8944 17921
rect 8996 17912 8998 17921
rect 8942 17847 8998 17856
rect 8944 16992 8996 16998
rect 8944 16934 8996 16940
rect 8852 16516 8904 16522
rect 8852 16458 8904 16464
rect 8956 16266 8984 16934
rect 8864 16238 8984 16266
rect 8864 16114 8892 16238
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 8944 16040 8996 16046
rect 8944 15982 8996 15988
rect 8772 15694 8892 15722
rect 8760 15564 8812 15570
rect 8760 15506 8812 15512
rect 8668 15088 8720 15094
rect 8668 15030 8720 15036
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8482 14784 8538 14793
rect 8482 14719 8538 14728
rect 8496 14414 8524 14719
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8588 14260 8616 14894
rect 8668 14884 8720 14890
rect 8668 14826 8720 14832
rect 8680 14385 8708 14826
rect 8666 14376 8722 14385
rect 8666 14311 8722 14320
rect 8588 14232 8708 14260
rect 8352 14172 8648 14192
rect 8408 14170 8432 14172
rect 8488 14170 8512 14172
rect 8568 14170 8592 14172
rect 8430 14118 8432 14170
rect 8494 14118 8506 14170
rect 8568 14118 8570 14170
rect 8408 14116 8432 14118
rect 8488 14116 8512 14118
rect 8568 14116 8592 14118
rect 8352 14096 8648 14116
rect 8680 14056 8708 14232
rect 8588 14028 8708 14056
rect 8390 13560 8446 13569
rect 8390 13495 8446 13504
rect 8404 13258 8432 13495
rect 8588 13462 8616 14028
rect 8772 13802 8800 15506
rect 8864 14074 8892 15694
rect 8956 15366 8984 15982
rect 9036 15904 9088 15910
rect 9036 15846 9088 15852
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8942 15192 8998 15201
rect 8942 15127 8998 15136
rect 8956 14822 8984 15127
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 8942 14240 8998 14249
rect 8942 14175 8998 14184
rect 8852 14068 8904 14074
rect 8852 14010 8904 14016
rect 8760 13796 8812 13802
rect 8760 13738 8812 13744
rect 8852 13796 8904 13802
rect 8852 13738 8904 13744
rect 8758 13560 8814 13569
rect 8758 13495 8814 13504
rect 8576 13456 8628 13462
rect 8576 13398 8628 13404
rect 8772 13326 8800 13495
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 8758 13152 8814 13161
rect 8352 13084 8648 13104
rect 8758 13087 8814 13096
rect 8408 13082 8432 13084
rect 8488 13082 8512 13084
rect 8568 13082 8592 13084
rect 8430 13030 8432 13082
rect 8494 13030 8506 13082
rect 8568 13030 8570 13082
rect 8408 13028 8432 13030
rect 8488 13028 8512 13030
rect 8568 13028 8592 13030
rect 8352 13008 8648 13028
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 7838 12407 7894 12416
rect 7852 12170 7880 12407
rect 7944 12396 8248 12424
rect 7840 12164 7892 12170
rect 7840 12106 7892 12112
rect 7838 12064 7894 12073
rect 7838 11999 7894 12008
rect 7852 11898 7880 11999
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7944 11744 7972 12396
rect 8312 12356 8340 12786
rect 8680 12374 8708 12922
rect 8772 12714 8800 13087
rect 8760 12708 8812 12714
rect 8760 12650 8812 12656
rect 8864 12646 8892 13738
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 8220 12328 8340 12356
rect 8668 12368 8720 12374
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 8036 12102 8064 12242
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8114 11928 8170 11937
rect 8114 11863 8170 11872
rect 7944 11716 8064 11744
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 7840 10736 7892 10742
rect 7760 10696 7840 10724
rect 7840 10678 7892 10684
rect 7852 10577 7880 10678
rect 7944 10674 7972 11562
rect 8036 11354 8064 11716
rect 8128 11694 8156 11863
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8024 11348 8076 11354
rect 8024 11290 8076 11296
rect 8024 11008 8076 11014
rect 8024 10950 8076 10956
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 7838 10568 7894 10577
rect 7380 10532 7432 10538
rect 7838 10503 7894 10512
rect 7380 10474 7432 10480
rect 7748 10056 7800 10062
rect 7944 10044 7972 10610
rect 7800 10016 7972 10044
rect 7748 9998 7800 10004
rect 7300 9846 7512 9874
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7288 9036 7340 9042
rect 7208 8996 7288 9024
rect 7102 8528 7158 8537
rect 7102 8463 7158 8472
rect 6932 7364 7052 7392
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6472 7160 6684 7188
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6276 4752 6328 4758
rect 6276 4694 6328 4700
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 5408 4236 5488 4264
rect 5540 4276 5592 4282
rect 5356 4218 5408 4224
rect 5540 4218 5592 4224
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5368 2961 5396 3538
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5460 3233 5488 3470
rect 5446 3224 5502 3233
rect 5446 3159 5502 3168
rect 5448 3120 5500 3126
rect 5448 3062 5500 3068
rect 5354 2952 5410 2961
rect 5354 2887 5410 2896
rect 5460 2854 5488 3062
rect 5356 2848 5408 2854
rect 5356 2790 5408 2796
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 5368 2378 5396 2790
rect 5552 2650 5580 4014
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5644 3398 5672 3946
rect 5736 3466 5764 4558
rect 5814 4312 5870 4321
rect 5998 4312 6054 4321
rect 5814 4247 5870 4256
rect 5920 4270 5998 4298
rect 5828 3534 5856 4247
rect 5920 4078 5948 4270
rect 5998 4247 6054 4256
rect 5908 4072 5960 4078
rect 5908 4014 5960 4020
rect 6196 4010 6224 4626
rect 6380 4570 6408 5102
rect 6288 4554 6408 4570
rect 6276 4548 6408 4554
rect 6328 4542 6408 4548
rect 6276 4490 6328 4496
rect 6288 4010 6316 4490
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 6380 4078 6408 4422
rect 6472 4214 6500 6394
rect 6564 5914 6592 6802
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 6184 4004 6236 4010
rect 6184 3946 6236 3952
rect 6276 4004 6328 4010
rect 6276 3946 6328 3952
rect 6460 4004 6512 4010
rect 6460 3946 6512 3952
rect 6366 3904 6422 3913
rect 5886 3836 6182 3856
rect 6366 3839 6422 3848
rect 5942 3834 5966 3836
rect 6022 3834 6046 3836
rect 6102 3834 6126 3836
rect 5964 3782 5966 3834
rect 6028 3782 6040 3834
rect 6102 3782 6104 3834
rect 5942 3780 5966 3782
rect 6022 3780 6046 3782
rect 6102 3780 6126 3782
rect 5886 3760 6182 3780
rect 6184 3664 6236 3670
rect 6104 3624 6184 3652
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5632 3392 5684 3398
rect 6104 3369 6132 3624
rect 6184 3606 6236 3612
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 5632 3334 5684 3340
rect 6090 3360 6146 3369
rect 5644 3058 5672 3334
rect 6090 3295 6146 3304
rect 6196 3058 6224 3470
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 6092 2916 6144 2922
rect 5828 2876 6092 2904
rect 5722 2816 5778 2825
rect 5828 2802 5856 2876
rect 6092 2858 6144 2864
rect 5778 2774 5856 2802
rect 5722 2751 5778 2760
rect 5886 2748 6182 2768
rect 5942 2746 5966 2748
rect 6022 2746 6046 2748
rect 6102 2746 6126 2748
rect 5964 2694 5966 2746
rect 6028 2694 6040 2746
rect 6102 2694 6104 2746
rect 5942 2692 5966 2694
rect 6022 2692 6046 2694
rect 6102 2692 6126 2694
rect 5886 2672 6182 2692
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 5446 2544 5502 2553
rect 5630 2544 5686 2553
rect 5540 2508 5592 2514
rect 5502 2488 5540 2496
rect 5446 2479 5540 2488
rect 5460 2468 5540 2479
rect 5630 2479 5686 2488
rect 5540 2450 5592 2456
rect 5356 2372 5408 2378
rect 5356 2314 5408 2320
rect 5264 2100 5316 2106
rect 5264 2042 5316 2048
rect 5644 1442 5672 2479
rect 5828 2378 5856 2586
rect 5816 2372 5868 2378
rect 5816 2314 5868 2320
rect 6288 1562 6316 3538
rect 6380 3126 6408 3839
rect 6368 3120 6420 3126
rect 6368 3062 6420 3068
rect 6472 2990 6500 3946
rect 6460 2984 6512 2990
rect 6460 2926 6512 2932
rect 6458 2544 6514 2553
rect 6458 2479 6514 2488
rect 6276 1556 6328 1562
rect 6276 1498 6328 1504
rect 6472 1442 6500 2479
rect 6564 2446 6592 5850
rect 6656 5522 6684 7160
rect 6748 6866 6776 7278
rect 6932 6882 6960 7364
rect 7012 7268 7064 7274
rect 7012 7210 7064 7216
rect 7024 7002 7052 7210
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 6736 6860 6788 6866
rect 6932 6854 7052 6882
rect 6788 6820 6868 6848
rect 6736 6802 6788 6808
rect 6734 6760 6790 6769
rect 6734 6695 6790 6704
rect 6748 5642 6776 6695
rect 6840 6254 6868 6820
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6932 6186 6960 6598
rect 7024 6361 7052 6854
rect 7010 6352 7066 6361
rect 7010 6287 7066 6296
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 6656 5494 6776 5522
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6656 5137 6684 5170
rect 6642 5128 6698 5137
rect 6642 5063 6698 5072
rect 6642 4992 6698 5001
rect 6642 4927 6698 4936
rect 6656 3913 6684 4927
rect 6642 3904 6698 3913
rect 6642 3839 6698 3848
rect 6642 3768 6698 3777
rect 6642 3703 6698 3712
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 6656 1494 6684 3703
rect 6748 2650 6776 5494
rect 6840 4486 6868 5714
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6840 4010 6868 4082
rect 6828 4004 6880 4010
rect 6828 3946 6880 3952
rect 6826 3904 6882 3913
rect 6826 3839 6882 3848
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 6734 2272 6790 2281
rect 6734 2207 6790 2216
rect 5552 1414 5672 1442
rect 6380 1414 6500 1442
rect 6644 1488 6696 1494
rect 6644 1430 6696 1436
rect 5552 480 5580 1414
rect 6000 1284 6052 1290
rect 6000 1226 6052 1232
rect 6012 480 6040 1226
rect 6380 480 6408 1414
rect 6748 1290 6776 2207
rect 6736 1284 6788 1290
rect 6736 1226 6788 1232
rect 6840 480 6868 3839
rect 6932 3534 6960 6122
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 7024 5370 7052 5510
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 7010 5264 7066 5273
rect 7010 5199 7066 5208
rect 7024 5166 7052 5199
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 7024 4690 7052 5102
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 7010 4448 7066 4457
rect 7010 4383 7066 4392
rect 7024 4010 7052 4383
rect 7012 4004 7064 4010
rect 7012 3946 7064 3952
rect 7010 3904 7066 3913
rect 7010 3839 7066 3848
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6918 3360 6974 3369
rect 6918 3295 6974 3304
rect 6932 2394 6960 3295
rect 7024 2514 7052 3839
rect 7116 2922 7144 8463
rect 7208 7206 7236 8996
rect 7288 8978 7340 8984
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7300 8362 7328 8774
rect 7288 8356 7340 8362
rect 7288 8298 7340 8304
rect 7300 8129 7328 8298
rect 7286 8120 7342 8129
rect 7286 8055 7342 8064
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7286 7712 7342 7721
rect 7286 7647 7342 7656
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7208 4826 7236 7142
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 7208 3602 7236 4014
rect 7300 3942 7328 7647
rect 7392 6202 7420 7890
rect 7484 6769 7512 9846
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7852 8498 7880 8774
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7564 7744 7616 7750
rect 7562 7712 7564 7721
rect 7616 7712 7618 7721
rect 7562 7647 7618 7656
rect 7746 7440 7802 7449
rect 7746 7375 7802 7384
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 7470 6760 7526 6769
rect 7470 6695 7526 6704
rect 7392 6174 7512 6202
rect 7576 6186 7604 6802
rect 7668 6497 7696 7278
rect 7654 6488 7710 6497
rect 7654 6423 7710 6432
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7392 4146 7420 6054
rect 7484 5216 7512 6174
rect 7564 6180 7616 6186
rect 7564 6122 7616 6128
rect 7576 5778 7604 6122
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7576 5409 7604 5714
rect 7562 5400 7618 5409
rect 7562 5335 7618 5344
rect 7484 5188 7584 5216
rect 7556 5148 7584 5188
rect 7556 5120 7604 5148
rect 7472 5092 7524 5098
rect 7472 5034 7524 5040
rect 7484 4826 7512 5034
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7576 4758 7604 5120
rect 7654 5128 7710 5137
rect 7654 5063 7710 5072
rect 7564 4752 7616 4758
rect 7564 4694 7616 4700
rect 7472 4616 7524 4622
rect 7524 4564 7604 4570
rect 7472 4558 7604 4564
rect 7484 4542 7604 4558
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7484 4282 7512 4422
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7470 4176 7526 4185
rect 7380 4140 7432 4146
rect 7470 4111 7526 4120
rect 7380 4082 7432 4088
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 7194 3224 7250 3233
rect 7194 3159 7250 3168
rect 7208 3058 7236 3159
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7104 2916 7156 2922
rect 7104 2858 7156 2864
rect 7194 2816 7250 2825
rect 7194 2751 7250 2760
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7116 2417 7144 2450
rect 7102 2408 7158 2417
rect 6932 2366 7052 2394
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 6932 1698 6960 2246
rect 7024 1902 7052 2366
rect 7102 2343 7158 2352
rect 7012 1896 7064 1902
rect 7012 1838 7064 1844
rect 6920 1692 6972 1698
rect 6920 1634 6972 1640
rect 7208 480 7236 2751
rect 7300 1834 7328 3878
rect 7392 3534 7420 4082
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7378 3224 7434 3233
rect 7378 3159 7380 3168
rect 7432 3159 7434 3168
rect 7380 3130 7432 3136
rect 7484 3058 7512 4111
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7392 2938 7420 2994
rect 7576 2938 7604 4542
rect 7392 2910 7604 2938
rect 7668 2922 7696 5063
rect 7760 3738 7788 7375
rect 7840 6860 7892 6866
rect 7840 6802 7892 6808
rect 7852 5386 7880 6802
rect 7944 5545 7972 8366
rect 7930 5536 7986 5545
rect 7930 5471 7986 5480
rect 7852 5358 7972 5386
rect 7840 5092 7892 5098
rect 7840 5034 7892 5040
rect 7852 4486 7880 5034
rect 7944 5030 7972 5358
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7932 4752 7984 4758
rect 7932 4694 7984 4700
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7944 4321 7972 4694
rect 7930 4312 7986 4321
rect 7930 4247 7986 4256
rect 7944 4146 7972 4247
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7852 3602 7880 4014
rect 7840 3596 7892 3602
rect 7840 3538 7892 3544
rect 8036 3482 8064 10950
rect 8128 10198 8156 11494
rect 8220 11393 8248 12328
rect 8668 12310 8720 12316
rect 8352 11996 8648 12016
rect 8408 11994 8432 11996
rect 8488 11994 8512 11996
rect 8568 11994 8592 11996
rect 8430 11942 8432 11994
rect 8494 11942 8506 11994
rect 8568 11942 8570 11994
rect 8408 11940 8432 11942
rect 8488 11940 8512 11942
rect 8568 11940 8592 11942
rect 8352 11920 8648 11940
rect 8484 11824 8536 11830
rect 8484 11766 8536 11772
rect 8496 11694 8524 11766
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8206 11384 8262 11393
rect 8772 11354 8800 12378
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 8864 12073 8892 12174
rect 8850 12064 8906 12073
rect 8850 11999 8906 12008
rect 8956 11694 8984 14175
rect 9048 13870 9076 15846
rect 9140 15434 9168 18108
rect 9402 17368 9458 17377
rect 9402 17303 9458 17312
rect 9310 16824 9366 16833
rect 9310 16759 9366 16768
rect 9324 16590 9352 16759
rect 9312 16584 9364 16590
rect 9312 16526 9364 16532
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9220 15904 9272 15910
rect 9220 15846 9272 15852
rect 9128 15428 9180 15434
rect 9128 15370 9180 15376
rect 9126 14648 9182 14657
rect 9126 14583 9182 14592
rect 9140 14385 9168 14583
rect 9126 14376 9182 14385
rect 9232 14346 9260 15846
rect 9324 15026 9352 16050
rect 9416 15881 9444 17303
rect 9508 16969 9536 19520
rect 9588 18216 9640 18222
rect 9588 18158 9640 18164
rect 9494 16960 9550 16969
rect 9494 16895 9550 16904
rect 9508 16425 9536 16895
rect 9600 16640 9628 18158
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9692 16794 9720 17818
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9784 16697 9812 16934
rect 9770 16688 9826 16697
rect 9600 16612 9720 16640
rect 9876 16658 9904 19520
rect 10232 17808 10284 17814
rect 10232 17750 10284 17756
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 10152 16794 10180 17478
rect 10244 16794 10272 17750
rect 10336 17134 10364 19520
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 10414 17232 10470 17241
rect 10414 17167 10416 17176
rect 10468 17167 10470 17176
rect 10416 17138 10468 17144
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 10232 16788 10284 16794
rect 10232 16730 10284 16736
rect 9770 16623 9826 16632
rect 9864 16652 9916 16658
rect 9494 16416 9550 16425
rect 9494 16351 9550 16360
rect 9692 16289 9720 16612
rect 9864 16594 9916 16600
rect 9678 16280 9734 16289
rect 9588 16244 9640 16250
rect 9678 16215 9734 16224
rect 9588 16186 9640 16192
rect 9496 16040 9548 16046
rect 9496 15982 9548 15988
rect 9402 15872 9458 15881
rect 9402 15807 9458 15816
rect 9508 15722 9536 15982
rect 9600 15910 9628 16186
rect 9680 16176 9732 16182
rect 9680 16118 9732 16124
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 9692 15745 9720 16118
rect 9678 15736 9734 15745
rect 9508 15694 9628 15722
rect 9600 15620 9628 15694
rect 9678 15671 9734 15680
rect 9600 15592 9812 15620
rect 9404 15496 9456 15502
rect 9680 15496 9732 15502
rect 9404 15438 9456 15444
rect 9494 15464 9550 15473
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9310 14784 9366 14793
rect 9310 14719 9366 14728
rect 9324 14550 9352 14719
rect 9312 14544 9364 14550
rect 9312 14486 9364 14492
rect 9126 14311 9182 14320
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 9140 14113 9168 14214
rect 9126 14104 9182 14113
rect 9126 14039 9182 14048
rect 9036 13864 9088 13870
rect 9036 13806 9088 13812
rect 9048 13326 9076 13806
rect 9416 13546 9444 15438
rect 9680 15438 9732 15444
rect 9494 15399 9550 15408
rect 9508 15201 9536 15399
rect 9692 15366 9720 15438
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9494 15192 9550 15201
rect 9494 15127 9550 15136
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9496 14952 9548 14958
rect 9496 14894 9548 14900
rect 9508 14346 9536 14894
rect 9496 14340 9548 14346
rect 9496 14282 9548 14288
rect 9600 13734 9628 14962
rect 9692 14657 9720 15302
rect 9784 14958 9812 15592
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 9876 14770 9904 16594
rect 9956 16108 10008 16114
rect 9956 16050 10008 16056
rect 9968 14770 9996 16050
rect 10048 15972 10100 15978
rect 10048 15914 10100 15920
rect 10060 15881 10088 15914
rect 10046 15872 10102 15881
rect 10046 15807 10102 15816
rect 10152 15473 10180 16730
rect 10232 16584 10284 16590
rect 10232 16526 10284 16532
rect 10244 15994 10272 16526
rect 10336 16114 10364 17070
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10428 16454 10456 16526
rect 10416 16448 10468 16454
rect 10416 16390 10468 16396
rect 10428 16114 10456 16390
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10416 16108 10468 16114
rect 10416 16050 10468 16056
rect 10244 15966 10364 15994
rect 10232 15904 10284 15910
rect 10232 15846 10284 15852
rect 10138 15464 10194 15473
rect 10138 15399 10194 15408
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 9784 14742 9904 14770
rect 9959 14742 9996 14770
rect 10060 14770 10088 15302
rect 10060 14742 10180 14770
rect 9678 14648 9734 14657
rect 9678 14583 9734 14592
rect 9784 14498 9812 14742
rect 9862 14648 9918 14657
rect 9862 14583 9918 14592
rect 9876 14550 9904 14583
rect 9692 14470 9812 14498
rect 9864 14544 9916 14550
rect 9959 14532 9987 14742
rect 9959 14504 9996 14532
rect 9864 14486 9916 14492
rect 9692 14260 9720 14470
rect 9692 14232 9904 14260
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9680 13728 9732 13734
rect 9680 13670 9732 13676
rect 9140 13518 9444 13546
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 8944 11688 8996 11694
rect 8944 11630 8996 11636
rect 9048 11393 9076 12106
rect 9034 11384 9090 11393
rect 8206 11319 8262 11328
rect 8760 11348 8812 11354
rect 8220 11268 8248 11319
rect 9034 11319 9090 11328
rect 8760 11290 8812 11296
rect 8300 11280 8352 11286
rect 8220 11240 8300 11268
rect 8300 11222 8352 11228
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 8352 10908 8648 10928
rect 8408 10906 8432 10908
rect 8488 10906 8512 10908
rect 8568 10906 8592 10908
rect 8430 10854 8432 10906
rect 8494 10854 8506 10906
rect 8568 10854 8570 10906
rect 8408 10852 8432 10854
rect 8488 10852 8512 10854
rect 8568 10852 8592 10854
rect 8352 10832 8648 10852
rect 8680 10724 8708 11154
rect 9140 11064 9168 13518
rect 9312 13456 9364 13462
rect 9312 13398 9364 13404
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 9232 12617 9260 12650
rect 9218 12608 9274 12617
rect 9218 12543 9274 12552
rect 9324 12442 9352 13398
rect 9496 13388 9548 13394
rect 9692 13376 9720 13670
rect 9548 13348 9720 13376
rect 9496 13330 9548 13336
rect 9678 13016 9734 13025
rect 9678 12951 9734 12960
rect 9692 12900 9720 12951
rect 9692 12872 9812 12900
rect 9678 12472 9734 12481
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9588 12436 9640 12442
rect 9678 12407 9734 12416
rect 9588 12378 9640 12384
rect 9600 12345 9628 12378
rect 9586 12336 9642 12345
rect 9586 12271 9642 12280
rect 9692 12238 9720 12407
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9218 12064 9274 12073
rect 9218 11999 9274 12008
rect 9232 11286 9260 11999
rect 9220 11280 9272 11286
rect 9220 11222 9272 11228
rect 8864 11036 9168 11064
rect 8680 10696 8800 10724
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8128 9353 8156 9658
rect 8220 9586 8248 10542
rect 8668 10192 8720 10198
rect 8668 10134 8720 10140
rect 8352 9820 8648 9840
rect 8408 9818 8432 9820
rect 8488 9818 8512 9820
rect 8568 9818 8592 9820
rect 8430 9766 8432 9818
rect 8494 9766 8506 9818
rect 8568 9766 8570 9818
rect 8408 9764 8432 9766
rect 8488 9764 8512 9766
rect 8568 9764 8592 9766
rect 8352 9744 8648 9764
rect 8680 9654 8708 10134
rect 8668 9648 8720 9654
rect 8668 9590 8720 9596
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8114 9344 8170 9353
rect 8114 9279 8170 9288
rect 8588 8974 8616 9454
rect 8772 9450 8800 10696
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8208 8832 8260 8838
rect 8206 8800 8208 8809
rect 8260 8800 8262 8809
rect 8206 8735 8262 8744
rect 8352 8732 8648 8752
rect 8408 8730 8432 8732
rect 8488 8730 8512 8732
rect 8568 8730 8592 8732
rect 8430 8678 8432 8730
rect 8494 8678 8506 8730
rect 8568 8678 8570 8730
rect 8408 8676 8432 8678
rect 8488 8676 8512 8678
rect 8568 8676 8592 8678
rect 8352 8656 8648 8676
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8114 7712 8170 7721
rect 8114 7647 8170 7656
rect 8128 6866 8156 7647
rect 8220 7585 8248 8230
rect 8404 8022 8432 8230
rect 8392 8016 8444 8022
rect 8392 7958 8444 7964
rect 8352 7644 8648 7664
rect 8408 7642 8432 7644
rect 8488 7642 8512 7644
rect 8568 7642 8592 7644
rect 8430 7590 8432 7642
rect 8494 7590 8506 7642
rect 8568 7590 8570 7642
rect 8408 7588 8432 7590
rect 8488 7588 8512 7590
rect 8568 7588 8592 7590
rect 8206 7576 8262 7585
rect 8352 7568 8648 7588
rect 8206 7511 8262 7520
rect 8220 7392 8248 7511
rect 8300 7404 8352 7410
rect 8220 7364 8300 7392
rect 8300 7346 8352 7352
rect 8680 7342 8708 8366
rect 8772 7954 8800 9386
rect 8864 9042 8892 11036
rect 9220 11008 9272 11014
rect 9034 10976 9090 10985
rect 9220 10950 9272 10956
rect 9034 10911 9090 10920
rect 8942 10432 8998 10441
rect 8942 10367 8998 10376
rect 8852 9036 8904 9042
rect 8852 8978 8904 8984
rect 8850 8664 8906 8673
rect 8850 8599 8906 8608
rect 8864 8265 8892 8599
rect 8850 8256 8906 8265
rect 8850 8191 8906 8200
rect 8850 8120 8906 8129
rect 8850 8055 8906 8064
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8864 7154 8892 8055
rect 8680 7126 8892 7154
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 8680 6730 8708 7126
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8352 6556 8648 6576
rect 8408 6554 8432 6556
rect 8488 6554 8512 6556
rect 8568 6554 8592 6556
rect 8430 6502 8432 6554
rect 8494 6502 8506 6554
rect 8568 6502 8570 6554
rect 8408 6500 8432 6502
rect 8488 6500 8512 6502
rect 8568 6500 8592 6502
rect 8352 6480 8648 6500
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 8128 5794 8156 6190
rect 8208 6112 8260 6118
rect 8206 6080 8208 6089
rect 8260 6080 8262 6089
rect 8206 6015 8262 6024
rect 8128 5766 8248 5794
rect 8114 5536 8170 5545
rect 8114 5471 8170 5480
rect 8128 4622 8156 5471
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8116 4004 8168 4010
rect 8116 3946 8168 3952
rect 7760 3454 8064 3482
rect 7656 2916 7708 2922
rect 7288 1828 7340 1834
rect 7288 1770 7340 1776
rect 7392 1086 7420 2910
rect 7656 2858 7708 2864
rect 7562 2816 7618 2825
rect 7760 2802 7788 3454
rect 7930 3224 7986 3233
rect 7930 3159 7986 3168
rect 7838 2952 7894 2961
rect 7838 2887 7894 2896
rect 7852 2854 7880 2887
rect 7562 2751 7618 2760
rect 7668 2774 7788 2802
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 7470 2544 7526 2553
rect 7470 2479 7526 2488
rect 7484 2446 7512 2479
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7576 1222 7604 2751
rect 7564 1216 7616 1222
rect 7564 1158 7616 1164
rect 7380 1080 7432 1086
rect 7380 1022 7432 1028
rect 7668 480 7696 2774
rect 7944 2689 7972 3159
rect 8022 2952 8078 2961
rect 8128 2938 8156 3946
rect 8220 3534 8248 5766
rect 8352 5468 8648 5488
rect 8408 5466 8432 5468
rect 8488 5466 8512 5468
rect 8568 5466 8592 5468
rect 8430 5414 8432 5466
rect 8494 5414 8506 5466
rect 8568 5414 8570 5466
rect 8408 5412 8432 5414
rect 8488 5412 8512 5414
rect 8568 5412 8592 5414
rect 8352 5392 8648 5412
rect 8482 5264 8538 5273
rect 8482 5199 8538 5208
rect 8576 5228 8628 5234
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8404 4826 8432 5102
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8496 4554 8524 5199
rect 8576 5170 8628 5176
rect 8588 4758 8616 5170
rect 8576 4752 8628 4758
rect 8576 4694 8628 4700
rect 8588 4622 8616 4694
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8484 4548 8536 4554
rect 8484 4490 8536 4496
rect 8352 4380 8648 4400
rect 8408 4378 8432 4380
rect 8488 4378 8512 4380
rect 8568 4378 8592 4380
rect 8430 4326 8432 4378
rect 8494 4326 8506 4378
rect 8568 4326 8570 4378
rect 8408 4324 8432 4326
rect 8488 4324 8512 4326
rect 8568 4324 8592 4326
rect 8352 4304 8648 4324
rect 8298 4176 8354 4185
rect 8298 4111 8354 4120
rect 8312 3738 8340 4111
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8404 3380 8432 3606
rect 8496 3505 8524 3674
rect 8576 3596 8628 3602
rect 8680 3584 8708 6666
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 8772 5030 8800 6054
rect 8864 5642 8892 6598
rect 8852 5636 8904 5642
rect 8852 5578 8904 5584
rect 8760 5024 8812 5030
rect 8812 4984 8892 5012
rect 8760 4966 8812 4972
rect 8760 4480 8812 4486
rect 8760 4422 8812 4428
rect 8628 3556 8708 3584
rect 8576 3538 8628 3544
rect 8482 3496 8538 3505
rect 8482 3431 8538 3440
rect 8668 3460 8720 3466
rect 8668 3402 8720 3408
rect 8078 2910 8156 2938
rect 8220 3352 8432 3380
rect 8022 2887 8078 2896
rect 7930 2680 7986 2689
rect 7840 2644 7892 2650
rect 7930 2615 7986 2624
rect 7840 2586 7892 2592
rect 7852 2145 7880 2586
rect 8022 2544 8078 2553
rect 8220 2514 8248 3352
rect 8352 3292 8648 3312
rect 8408 3290 8432 3292
rect 8488 3290 8512 3292
rect 8568 3290 8592 3292
rect 8430 3238 8432 3290
rect 8494 3238 8506 3290
rect 8568 3238 8570 3290
rect 8408 3236 8432 3238
rect 8488 3236 8512 3238
rect 8568 3236 8592 3238
rect 8352 3216 8648 3236
rect 8680 3194 8708 3402
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 8484 2984 8536 2990
rect 8576 2984 8628 2990
rect 8484 2926 8536 2932
rect 8574 2952 8576 2961
rect 8628 2952 8630 2961
rect 8496 2553 8524 2926
rect 8574 2887 8630 2896
rect 8482 2544 8538 2553
rect 8022 2479 8078 2488
rect 8208 2508 8260 2514
rect 7932 2304 7984 2310
rect 7932 2246 7984 2252
rect 7838 2136 7894 2145
rect 7838 2071 7894 2080
rect 7944 2009 7972 2246
rect 7930 2000 7986 2009
rect 7930 1935 7986 1944
rect 8036 480 8064 2479
rect 8482 2479 8538 2488
rect 8208 2450 8260 2456
rect 8220 1018 8248 2450
rect 8772 2446 8800 4422
rect 8864 3058 8892 4984
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 8956 2514 8984 10367
rect 9048 10305 9076 10911
rect 9232 10470 9260 10950
rect 9324 10713 9352 12106
rect 9310 10704 9366 10713
rect 9310 10639 9366 10648
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9034 10296 9090 10305
rect 9034 10231 9090 10240
rect 9324 9994 9352 10639
rect 9312 9988 9364 9994
rect 9312 9930 9364 9936
rect 9218 9888 9274 9897
rect 9218 9823 9274 9832
rect 9126 9752 9182 9761
rect 9126 9687 9182 9696
rect 9140 9518 9168 9687
rect 9232 9602 9260 9823
rect 9232 9574 9352 9602
rect 9128 9512 9180 9518
rect 9180 9472 9260 9500
rect 9128 9454 9180 9460
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 9048 6633 9076 8978
rect 9140 7750 9168 9318
rect 9232 9042 9260 9472
rect 9220 9036 9272 9042
rect 9220 8978 9272 8984
rect 9232 8430 9260 8978
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 9232 7886 9260 8366
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 9034 6624 9090 6633
rect 9034 6559 9090 6568
rect 9034 6352 9090 6361
rect 9034 6287 9090 6296
rect 9048 5953 9076 6287
rect 9034 5944 9090 5953
rect 9034 5879 9090 5888
rect 9140 5828 9168 7686
rect 9232 6610 9260 7686
rect 9324 7274 9352 9574
rect 9508 7750 9536 12174
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9600 11150 9628 11562
rect 9692 11558 9720 11698
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9784 11370 9812 12872
rect 9876 12374 9904 14232
rect 9968 13138 9996 14504
rect 10152 14482 10180 14742
rect 10140 14476 10192 14482
rect 10140 14418 10192 14424
rect 10140 14340 10192 14346
rect 10140 14282 10192 14288
rect 10152 13870 10180 14282
rect 10244 14074 10272 15846
rect 10336 15706 10364 15966
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10324 15700 10376 15706
rect 10324 15642 10376 15648
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10336 15201 10364 15438
rect 10322 15192 10378 15201
rect 10322 15127 10378 15136
rect 10324 14816 10376 14822
rect 10428 14793 10456 15846
rect 10520 15570 10548 18158
rect 10508 15564 10560 15570
rect 10508 15506 10560 15512
rect 10508 15428 10560 15434
rect 10508 15370 10560 15376
rect 10324 14758 10376 14764
rect 10414 14784 10470 14793
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 10060 13462 10088 13738
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 10244 13530 10272 13670
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 10048 13456 10100 13462
rect 10048 13398 10100 13404
rect 9968 13110 10088 13138
rect 9954 13016 10010 13025
rect 9954 12951 10010 12960
rect 9864 12368 9916 12374
rect 9864 12310 9916 12316
rect 9784 11342 9904 11370
rect 9680 11280 9732 11286
rect 9732 11240 9812 11268
rect 9680 11222 9732 11228
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9678 11112 9734 11121
rect 9600 10062 9628 11086
rect 9678 11047 9734 11056
rect 9692 10742 9720 11047
rect 9784 10849 9812 11240
rect 9770 10840 9826 10849
rect 9770 10775 9826 10784
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9772 10532 9824 10538
rect 9772 10474 9824 10480
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9600 9518 9628 9998
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9600 9217 9628 9318
rect 9586 9208 9642 9217
rect 9586 9143 9642 9152
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9312 7268 9364 7274
rect 9312 7210 9364 7216
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9402 6624 9458 6633
rect 9232 6582 9352 6610
rect 9218 6488 9274 6497
rect 9218 6423 9274 6432
rect 9232 6254 9260 6423
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9324 5896 9352 6582
rect 9402 6559 9458 6568
rect 9416 6186 9444 6559
rect 9508 6254 9536 6938
rect 9600 6905 9628 8910
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 9586 6896 9642 6905
rect 9586 6831 9642 6840
rect 9692 6746 9720 8502
rect 9784 7478 9812 10474
rect 9876 8566 9904 11342
rect 9968 10305 9996 12951
rect 10060 12050 10088 13110
rect 10232 12980 10284 12986
rect 10232 12922 10284 12928
rect 10244 12782 10272 12922
rect 10232 12776 10284 12782
rect 10232 12718 10284 12724
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 10152 12481 10180 12582
rect 10138 12472 10194 12481
rect 10138 12407 10194 12416
rect 10140 12232 10192 12238
rect 10244 12220 10272 12582
rect 10192 12192 10272 12220
rect 10140 12174 10192 12180
rect 10060 12022 10180 12050
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 10060 11286 10088 11834
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 10046 11112 10102 11121
rect 10046 11047 10102 11056
rect 9954 10296 10010 10305
rect 9954 10231 10010 10240
rect 10060 10180 10088 11047
rect 9968 10152 10088 10180
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 9864 8288 9916 8294
rect 9862 8256 9864 8265
rect 9916 8256 9918 8265
rect 9862 8191 9918 8200
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9772 7472 9824 7478
rect 9772 7414 9824 7420
rect 9600 6718 9720 6746
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 9324 5868 9536 5896
rect 9140 5800 9352 5828
rect 9034 5672 9090 5681
rect 9034 5607 9090 5616
rect 9048 4282 9076 5607
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 9140 5302 9168 5510
rect 9128 5296 9180 5302
rect 9128 5238 9180 5244
rect 9140 5098 9168 5238
rect 9128 5092 9180 5098
rect 9128 5034 9180 5040
rect 9220 5092 9272 5098
rect 9220 5034 9272 5040
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 9036 4276 9088 4282
rect 9036 4218 9088 4224
rect 9034 4176 9090 4185
rect 9034 4111 9090 4120
rect 9048 4078 9076 4111
rect 9140 4078 9168 4762
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 9048 3466 9076 3878
rect 9128 3528 9180 3534
rect 9126 3496 9128 3505
rect 9180 3496 9182 3505
rect 9036 3460 9088 3466
rect 9126 3431 9182 3440
rect 9036 3402 9088 3408
rect 9232 3194 9260 5034
rect 9324 4826 9352 5800
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9324 4282 9352 4422
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9324 3670 9352 4014
rect 9312 3664 9364 3670
rect 9312 3606 9364 3612
rect 9416 3584 9444 5510
rect 9508 5030 9536 5868
rect 9600 5692 9628 6718
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9692 5846 9720 6598
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9784 5778 9812 6326
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9600 5664 9720 5692
rect 9692 5522 9720 5664
rect 9770 5536 9826 5545
rect 9692 5494 9770 5522
rect 9770 5471 9826 5480
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9588 5296 9640 5302
rect 9588 5238 9640 5244
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9508 4078 9536 4762
rect 9600 4486 9628 5238
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9692 4298 9720 5306
rect 9772 5296 9824 5302
rect 9772 5238 9824 5244
rect 9784 5030 9812 5238
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9770 4856 9826 4865
rect 9770 4791 9826 4800
rect 9784 4604 9812 4791
rect 9876 4706 9904 7686
rect 9968 6633 9996 10152
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 9954 6624 10010 6633
rect 9954 6559 10010 6568
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 9968 5778 9996 6054
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 9968 5137 9996 5170
rect 9954 5128 10010 5137
rect 9954 5063 10010 5072
rect 10060 4978 10088 8434
rect 10152 7342 10180 12022
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 10244 11393 10272 11630
rect 10336 11626 10364 14758
rect 10414 14719 10470 14728
rect 10520 14657 10548 15370
rect 10612 15337 10640 18226
rect 10704 18154 10732 19520
rect 11072 18290 11100 19520
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 10692 18148 10744 18154
rect 10692 18090 10744 18096
rect 11428 18148 11480 18154
rect 11428 18090 11480 18096
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 11164 16998 11192 18022
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 10704 16640 10732 16934
rect 10817 16892 11113 16912
rect 10873 16890 10897 16892
rect 10953 16890 10977 16892
rect 11033 16890 11057 16892
rect 10895 16838 10897 16890
rect 10959 16838 10971 16890
rect 11033 16838 11035 16890
rect 10873 16836 10897 16838
rect 10953 16836 10977 16838
rect 11033 16836 11057 16838
rect 10817 16816 11113 16836
rect 11060 16720 11112 16726
rect 11060 16662 11112 16668
rect 10784 16652 10836 16658
rect 10704 16612 10784 16640
rect 10784 16594 10836 16600
rect 10796 15978 10824 16594
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10888 16289 10916 16390
rect 10874 16280 10930 16289
rect 10874 16215 10930 16224
rect 11072 15978 11100 16662
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 10784 15972 10836 15978
rect 10784 15914 10836 15920
rect 11060 15972 11112 15978
rect 11060 15914 11112 15920
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10704 15502 10732 15846
rect 10817 15804 11113 15824
rect 10873 15802 10897 15804
rect 10953 15802 10977 15804
rect 11033 15802 11057 15804
rect 10895 15750 10897 15802
rect 10959 15750 10971 15802
rect 11033 15750 11035 15802
rect 10873 15748 10897 15750
rect 10953 15748 10977 15750
rect 11033 15748 11057 15750
rect 10817 15728 11113 15748
rect 11164 15688 11192 16594
rect 11334 16552 11390 16561
rect 11334 16487 11390 16496
rect 11348 16250 11376 16487
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 11072 15660 11192 15688
rect 10784 15632 10836 15638
rect 10968 15632 11020 15638
rect 10784 15574 10836 15580
rect 10888 15592 10968 15620
rect 10692 15496 10744 15502
rect 10692 15438 10744 15444
rect 10796 15348 10824 15574
rect 10888 15473 10916 15592
rect 10968 15574 11020 15580
rect 10874 15464 10930 15473
rect 10874 15399 10930 15408
rect 10598 15328 10654 15337
rect 10598 15263 10654 15272
rect 10704 15320 10824 15348
rect 10506 14648 10562 14657
rect 10506 14583 10562 14592
rect 10508 14544 10560 14550
rect 10704 14532 10732 15320
rect 11072 15201 11100 15660
rect 11058 15192 11114 15201
rect 11058 15127 11114 15136
rect 10876 14884 10928 14890
rect 11072 14872 11100 15127
rect 10928 14844 11100 14872
rect 10876 14826 10928 14832
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 10817 14716 11113 14736
rect 10873 14714 10897 14716
rect 10953 14714 10977 14716
rect 11033 14714 11057 14716
rect 10895 14662 10897 14714
rect 10959 14662 10971 14714
rect 11033 14662 11035 14714
rect 10873 14660 10897 14662
rect 10953 14660 10977 14662
rect 11033 14660 11057 14662
rect 10817 14640 11113 14660
rect 11164 14618 11192 14758
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 10704 14504 11008 14532
rect 10508 14486 10560 14492
rect 10520 14362 10548 14486
rect 10600 14476 10652 14482
rect 10652 14436 10824 14464
rect 10600 14418 10652 14424
rect 10416 14340 10468 14346
rect 10520 14334 10640 14362
rect 10416 14282 10468 14288
rect 10612 14328 10640 14334
rect 10692 14340 10744 14346
rect 10612 14300 10692 14328
rect 10428 13569 10456 14282
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10414 13560 10470 13569
rect 10414 13495 10470 13504
rect 10414 13016 10470 13025
rect 10414 12951 10470 12960
rect 10428 12714 10456 12951
rect 10416 12708 10468 12714
rect 10416 12650 10468 12656
rect 10416 12300 10468 12306
rect 10416 12242 10468 12248
rect 10324 11620 10376 11626
rect 10324 11562 10376 11568
rect 10230 11384 10286 11393
rect 10230 11319 10286 11328
rect 10336 10606 10364 11562
rect 10428 11218 10456 12242
rect 10520 12170 10548 14214
rect 10612 13734 10640 14300
rect 10692 14282 10744 14288
rect 10692 14000 10744 14006
rect 10692 13942 10744 13948
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 10598 13560 10654 13569
rect 10598 13495 10654 13504
rect 10612 12714 10640 13495
rect 10704 13240 10732 13942
rect 10796 13870 10824 14436
rect 10980 14278 11008 14504
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 11072 13802 11100 14418
rect 11060 13796 11112 13802
rect 11060 13738 11112 13744
rect 10817 13628 11113 13648
rect 10873 13626 10897 13628
rect 10953 13626 10977 13628
rect 11033 13626 11057 13628
rect 10895 13574 10897 13626
rect 10959 13574 10971 13626
rect 11033 13574 11035 13626
rect 10873 13572 10897 13574
rect 10953 13572 10977 13574
rect 11033 13572 11057 13574
rect 10817 13552 11113 13572
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10784 13252 10836 13258
rect 10704 13212 10784 13240
rect 10784 13194 10836 13200
rect 10888 13190 10916 13330
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 11164 13025 11192 14418
rect 11256 13326 11284 16186
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11348 13818 11376 15438
rect 11440 14770 11468 18090
rect 11532 15745 11560 19520
rect 11900 18306 11928 19520
rect 12256 18828 12308 18834
rect 12256 18770 12308 18776
rect 11624 18278 11928 18306
rect 11518 15736 11574 15745
rect 11518 15671 11574 15680
rect 11440 14742 11560 14770
rect 11426 14648 11482 14657
rect 11426 14583 11482 14592
rect 11440 14113 11468 14583
rect 11426 14104 11482 14113
rect 11426 14039 11482 14048
rect 11348 13790 11468 13818
rect 11336 13728 11388 13734
rect 11334 13696 11336 13705
rect 11388 13696 11390 13705
rect 11334 13631 11390 13640
rect 11334 13560 11390 13569
rect 11334 13495 11390 13504
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11244 13184 11296 13190
rect 11244 13126 11296 13132
rect 11150 13016 11206 13025
rect 10876 12980 10928 12986
rect 11150 12951 11206 12960
rect 10876 12922 10928 12928
rect 10888 12850 10916 12922
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10784 12776 10836 12782
rect 10704 12736 10784 12764
rect 10600 12708 10652 12714
rect 10600 12650 10652 12656
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10508 11824 10560 11830
rect 10508 11766 10560 11772
rect 10520 11393 10548 11766
rect 10506 11384 10562 11393
rect 10506 11319 10562 11328
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10508 10736 10560 10742
rect 10506 10704 10508 10713
rect 10560 10704 10562 10713
rect 10506 10639 10562 10648
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10612 10538 10640 12650
rect 10704 12442 10732 12736
rect 10784 12718 10836 12724
rect 10817 12540 11113 12560
rect 10873 12538 10897 12540
rect 10953 12538 10977 12540
rect 11033 12538 11057 12540
rect 10895 12486 10897 12538
rect 10959 12486 10971 12538
rect 11033 12486 11035 12538
rect 10873 12484 10897 12486
rect 10953 12484 10977 12486
rect 11033 12484 11057 12486
rect 10817 12464 11113 12484
rect 10692 12436 10744 12442
rect 11164 12424 11192 12951
rect 11256 12617 11284 13126
rect 11242 12608 11298 12617
rect 11242 12543 11298 12552
rect 10692 12378 10744 12384
rect 11072 12396 11192 12424
rect 10874 12064 10930 12073
rect 10874 11999 10930 12008
rect 10888 11626 10916 11999
rect 10968 11824 11020 11830
rect 10966 11792 10968 11801
rect 11020 11792 11022 11801
rect 10966 11727 11022 11736
rect 10876 11620 10928 11626
rect 10876 11562 10928 11568
rect 11072 11540 11100 12396
rect 11152 12300 11204 12306
rect 11348 12288 11376 13495
rect 11440 13433 11468 13790
rect 11426 13424 11482 13433
rect 11426 13359 11482 13368
rect 11426 13152 11482 13161
rect 11426 13087 11482 13096
rect 11440 12850 11468 13087
rect 11428 12844 11480 12850
rect 11428 12786 11480 12792
rect 11204 12260 11376 12288
rect 11152 12242 11204 12248
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11164 11762 11192 11834
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11256 11558 11284 11834
rect 11348 11801 11376 12260
rect 11334 11792 11390 11801
rect 11334 11727 11390 11736
rect 11428 11688 11480 11694
rect 11428 11630 11480 11636
rect 11244 11552 11296 11558
rect 11072 11512 11192 11540
rect 10817 11452 11113 11472
rect 10873 11450 10897 11452
rect 10953 11450 10977 11452
rect 11033 11450 11057 11452
rect 10895 11398 10897 11450
rect 10959 11398 10971 11450
rect 11033 11398 11035 11450
rect 10873 11396 10897 11398
rect 10953 11396 10977 11398
rect 11033 11396 11057 11398
rect 10817 11376 11113 11396
rect 10968 11280 11020 11286
rect 10968 11222 11020 11228
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 10980 11150 11008 11222
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10980 11014 11008 11086
rect 10968 11008 11020 11014
rect 10968 10950 11020 10956
rect 11072 10849 11100 11222
rect 11164 11014 11192 11512
rect 11244 11494 11296 11500
rect 11334 11520 11390 11529
rect 11334 11455 11390 11464
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 11058 10840 11114 10849
rect 11058 10775 11114 10784
rect 10600 10532 10652 10538
rect 10784 10532 10836 10538
rect 10600 10474 10652 10480
rect 10704 10492 10784 10520
rect 10414 10432 10470 10441
rect 10414 10367 10470 10376
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 10244 9042 10272 9590
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 10336 7954 10364 8774
rect 10428 8022 10456 10367
rect 10704 10266 10732 10492
rect 10784 10474 10836 10480
rect 10817 10364 11113 10384
rect 10873 10362 10897 10364
rect 10953 10362 10977 10364
rect 11033 10362 11057 10364
rect 10895 10310 10897 10362
rect 10959 10310 10971 10362
rect 11033 10310 11035 10362
rect 10873 10308 10897 10310
rect 10953 10308 10977 10310
rect 11033 10308 11057 10310
rect 10817 10288 11113 10308
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10520 10130 10548 10202
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 10506 9344 10562 9353
rect 10506 9279 10562 9288
rect 10520 9042 10548 9279
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10612 8922 10640 9862
rect 10704 9058 10732 10202
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 10796 9926 10824 10066
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 10817 9276 11113 9296
rect 10873 9274 10897 9276
rect 10953 9274 10977 9276
rect 11033 9274 11057 9276
rect 10895 9222 10897 9274
rect 10959 9222 10971 9274
rect 11033 9222 11035 9274
rect 10873 9220 10897 9222
rect 10953 9220 10977 9222
rect 11033 9220 11057 9222
rect 10817 9200 11113 9220
rect 10704 9030 11100 9058
rect 10968 8968 11020 8974
rect 10612 8894 10732 8922
rect 10968 8910 11020 8916
rect 10600 8832 10652 8838
rect 10520 8792 10600 8820
rect 10416 8016 10468 8022
rect 10416 7958 10468 7964
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10232 7472 10284 7478
rect 10232 7414 10284 7420
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 10138 7032 10194 7041
rect 10138 6967 10194 6976
rect 10152 6798 10180 6967
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10140 6248 10192 6254
rect 10140 6190 10192 6196
rect 9968 4950 10088 4978
rect 10152 4978 10180 6190
rect 10244 5914 10272 7414
rect 10336 6798 10364 7890
rect 10520 7041 10548 8792
rect 10600 8774 10652 8780
rect 10704 8514 10732 8894
rect 10612 8486 10732 8514
rect 10506 7032 10562 7041
rect 10506 6967 10562 6976
rect 10508 6928 10560 6934
rect 10508 6870 10560 6876
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 10232 5908 10284 5914
rect 10232 5850 10284 5856
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10244 5545 10272 5646
rect 10230 5536 10286 5545
rect 10230 5471 10286 5480
rect 10336 5302 10364 6598
rect 10520 6458 10548 6870
rect 10612 6662 10640 8486
rect 10980 8362 11008 8910
rect 11072 8378 11100 9030
rect 11164 8634 11192 9386
rect 11256 8906 11284 9862
rect 11244 8900 11296 8906
rect 11244 8842 11296 8848
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10968 8356 11020 8362
rect 11072 8350 11284 8378
rect 11348 8362 11376 11455
rect 10968 8298 11020 8304
rect 10704 7750 10732 8298
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 10817 8188 11113 8208
rect 10873 8186 10897 8188
rect 10953 8186 10977 8188
rect 11033 8186 11057 8188
rect 10895 8134 10897 8186
rect 10959 8134 10971 8186
rect 11033 8134 11035 8186
rect 10873 8132 10897 8134
rect 10953 8132 10977 8134
rect 11033 8132 11057 8134
rect 10817 8112 11113 8132
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10784 7812 10836 7818
rect 10784 7754 10836 7760
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10690 7576 10746 7585
rect 10796 7562 10824 7754
rect 10746 7534 10824 7562
rect 10690 7511 10746 7520
rect 10704 6934 10732 7511
rect 10876 7472 10928 7478
rect 10876 7414 10928 7420
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10796 7188 10824 7346
rect 10888 7342 10916 7414
rect 10876 7336 10928 7342
rect 10980 7313 11008 7414
rect 11072 7410 11100 7822
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 10876 7278 10928 7284
rect 10966 7304 11022 7313
rect 10966 7239 11022 7248
rect 11072 7188 11100 7346
rect 10796 7160 11100 7188
rect 10817 7100 11113 7120
rect 10873 7098 10897 7100
rect 10953 7098 10977 7100
rect 11033 7098 11057 7100
rect 10895 7046 10897 7098
rect 10959 7046 10971 7098
rect 11033 7046 11035 7098
rect 10873 7044 10897 7046
rect 10953 7044 10977 7046
rect 11033 7044 11057 7046
rect 10817 7024 11113 7044
rect 11164 6984 11192 8230
rect 10980 6956 11192 6984
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10782 6624 10838 6633
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10414 6080 10470 6089
rect 10414 6015 10470 6024
rect 10232 5296 10284 5302
rect 10232 5238 10284 5244
rect 10324 5296 10376 5302
rect 10324 5238 10376 5244
rect 10244 5148 10272 5238
rect 10244 5120 10364 5148
rect 10152 4950 10272 4978
rect 9968 4826 9996 4950
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 10138 4822 10194 4831
rect 10138 4757 10194 4766
rect 9876 4678 9996 4706
rect 10152 4690 10180 4757
rect 9784 4576 9904 4604
rect 9600 4270 9720 4298
rect 9600 4185 9628 4270
rect 9876 4214 9904 4576
rect 9680 4208 9732 4214
rect 9586 4176 9642 4185
rect 9680 4150 9732 4156
rect 9864 4208 9916 4214
rect 9864 4150 9916 4156
rect 9586 4111 9642 4120
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9692 3992 9720 4150
rect 9600 3964 9720 3992
rect 9864 4004 9916 4010
rect 9416 3556 9536 3584
rect 9402 3496 9458 3505
rect 9402 3431 9458 3440
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 9128 2916 9180 2922
rect 9128 2858 9180 2864
rect 8944 2508 8996 2514
rect 8944 2450 8996 2456
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 8352 2204 8648 2224
rect 8408 2202 8432 2204
rect 8488 2202 8512 2204
rect 8568 2202 8592 2204
rect 8430 2150 8432 2202
rect 8494 2150 8506 2202
rect 8568 2150 8570 2202
rect 8408 2148 8432 2150
rect 8488 2148 8512 2150
rect 8568 2148 8592 2150
rect 8352 2128 8648 2148
rect 8484 1556 8536 1562
rect 8484 1498 8536 1504
rect 8852 1556 8904 1562
rect 8852 1498 8904 1504
rect 8496 1329 8524 1498
rect 8482 1320 8538 1329
rect 8482 1255 8538 1264
rect 8208 1012 8260 1018
rect 8208 954 8260 960
rect 8496 480 8524 1255
rect 8864 480 8892 1498
rect 8956 678 8984 2450
rect 9140 2310 9168 2858
rect 9232 2446 9260 2926
rect 9220 2440 9272 2446
rect 9416 2394 9444 3431
rect 9508 2854 9536 3556
rect 9600 3534 9628 3964
rect 9864 3946 9916 3952
rect 9876 3652 9904 3946
rect 9968 3754 9996 4678
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 10060 3913 10088 4558
rect 10140 4480 10192 4486
rect 10140 4422 10192 4428
rect 10046 3904 10102 3913
rect 10046 3839 10102 3848
rect 9968 3726 10088 3754
rect 9770 3632 9826 3641
rect 9680 3596 9732 3602
rect 9876 3624 9996 3652
rect 9770 3567 9826 3576
rect 9680 3538 9732 3544
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9220 2382 9272 2388
rect 9324 2366 9444 2394
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 9324 1154 9352 2366
rect 9404 2304 9456 2310
rect 9404 2246 9456 2252
rect 9416 2106 9444 2246
rect 9494 2136 9550 2145
rect 9404 2100 9456 2106
rect 9494 2071 9550 2080
rect 9404 2042 9456 2048
rect 9508 1358 9536 2071
rect 9496 1352 9548 1358
rect 9496 1294 9548 1300
rect 9312 1148 9364 1154
rect 9312 1090 9364 1096
rect 9312 1012 9364 1018
rect 9312 954 9364 960
rect 8944 672 8996 678
rect 8944 614 8996 620
rect 9324 480 9352 954
rect 9600 950 9628 2586
rect 9588 944 9640 950
rect 9588 886 9640 892
rect 9692 480 9720 3538
rect 9784 2854 9812 3567
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 9784 1766 9812 2246
rect 9772 1760 9824 1766
rect 9772 1702 9824 1708
rect 9876 1562 9904 3470
rect 9968 2417 9996 3624
rect 10060 2972 10088 3726
rect 10152 3534 10180 4422
rect 10244 4026 10272 4950
rect 10336 4729 10364 5120
rect 10428 4826 10456 6015
rect 10520 5953 10548 6258
rect 10506 5944 10562 5953
rect 10506 5879 10562 5888
rect 10520 5710 10548 5879
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10612 5545 10640 6394
rect 10704 6254 10732 6598
rect 10782 6559 10838 6568
rect 10796 6458 10824 6559
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 10980 6254 11008 6956
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10598 5536 10654 5545
rect 10598 5471 10654 5480
rect 10704 5080 10732 6054
rect 10817 6012 11113 6032
rect 10873 6010 10897 6012
rect 10953 6010 10977 6012
rect 11033 6010 11057 6012
rect 10895 5958 10897 6010
rect 10959 5958 10971 6010
rect 11033 5958 11035 6010
rect 10873 5956 10897 5958
rect 10953 5956 10977 5958
rect 11033 5956 11057 5958
rect 10817 5936 11113 5956
rect 10874 5808 10930 5817
rect 10874 5743 10930 5752
rect 10782 5536 10838 5545
rect 10782 5471 10838 5480
rect 10796 5166 10824 5471
rect 10888 5234 10916 5743
rect 11164 5273 11192 6802
rect 11150 5264 11206 5273
rect 10876 5228 10928 5234
rect 11150 5199 11206 5208
rect 10876 5170 10928 5176
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10612 5052 10732 5080
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10322 4720 10378 4729
rect 10322 4655 10378 4664
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 10336 4282 10364 4558
rect 10324 4276 10376 4282
rect 10324 4218 10376 4224
rect 10428 4196 10456 4762
rect 10612 4486 10640 5052
rect 10888 5012 10916 5170
rect 10704 4984 10916 5012
rect 10704 4690 10732 4984
rect 10817 4924 11113 4944
rect 10873 4922 10897 4924
rect 10953 4922 10977 4924
rect 11033 4922 11057 4924
rect 10895 4870 10897 4922
rect 10959 4870 10971 4922
rect 11033 4870 11035 4922
rect 10873 4868 10897 4870
rect 10953 4868 10977 4870
rect 11033 4868 11057 4870
rect 10817 4848 11113 4868
rect 11256 4706 11284 8350
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11348 7342 11376 8298
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11334 7168 11390 7177
rect 11334 7103 11390 7112
rect 11348 6866 11376 7103
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 11348 5846 11376 6598
rect 11336 5840 11388 5846
rect 11336 5782 11388 5788
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 11348 4826 11376 5578
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10888 4678 11284 4706
rect 10600 4480 10652 4486
rect 10600 4422 10652 4428
rect 10428 4168 10548 4196
rect 10244 3998 10364 4026
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10244 3777 10272 3878
rect 10230 3768 10286 3777
rect 10230 3703 10286 3712
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10244 3097 10272 3538
rect 10230 3088 10286 3097
rect 10336 3058 10364 3998
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 10230 3023 10286 3032
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10060 2944 10272 2972
rect 10046 2680 10102 2689
rect 10046 2615 10102 2624
rect 10060 2582 10088 2615
rect 10048 2576 10100 2582
rect 10048 2518 10100 2524
rect 10138 2544 10194 2553
rect 10138 2479 10194 2488
rect 10048 2440 10100 2446
rect 9954 2408 10010 2417
rect 10048 2382 10100 2388
rect 9954 2343 10010 2352
rect 10060 2310 10088 2382
rect 10048 2304 10100 2310
rect 10048 2246 10100 2252
rect 9864 1556 9916 1562
rect 9864 1498 9916 1504
rect 10152 480 10180 2479
rect 10244 1630 10272 2944
rect 10336 2836 10364 2994
rect 10428 2990 10456 3878
rect 10520 3602 10548 4168
rect 10796 4026 10824 4626
rect 10888 4214 10916 4678
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 11058 4584 11114 4593
rect 10980 4282 11008 4558
rect 11242 4584 11298 4593
rect 11164 4554 11242 4570
rect 11058 4519 11114 4528
rect 11152 4548 11242 4554
rect 11072 4486 11100 4519
rect 11204 4542 11242 4548
rect 11242 4519 11298 4528
rect 11152 4490 11204 4496
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11348 4298 11376 4762
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 11256 4270 11376 4298
rect 11440 4282 11468 11630
rect 11532 7002 11560 14742
rect 11624 13025 11652 18278
rect 11794 17912 11850 17921
rect 11794 17847 11850 17856
rect 11704 17808 11756 17814
rect 11704 17750 11756 17756
rect 11610 13016 11666 13025
rect 11610 12951 11666 12960
rect 11612 12708 11664 12714
rect 11612 12650 11664 12656
rect 11624 12374 11652 12650
rect 11612 12368 11664 12374
rect 11612 12310 11664 12316
rect 11624 10674 11652 12310
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11624 8294 11652 9318
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11624 8090 11652 8230
rect 11612 8084 11664 8090
rect 11612 8026 11664 8032
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 11624 7546 11652 7686
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 11716 7392 11744 17750
rect 11808 17134 11836 17847
rect 11980 17604 12032 17610
rect 11980 17546 12032 17552
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11808 16969 11836 17070
rect 11794 16960 11850 16969
rect 11794 16895 11850 16904
rect 11992 16522 12020 17546
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 11980 16516 12032 16522
rect 11980 16458 12032 16464
rect 12070 16144 12126 16153
rect 12070 16079 12072 16088
rect 12124 16079 12126 16088
rect 12072 16050 12124 16056
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11900 15706 11928 15982
rect 11980 15972 12032 15978
rect 11980 15914 12032 15920
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 11796 15428 11848 15434
rect 11796 15370 11848 15376
rect 11808 15065 11836 15370
rect 11794 15056 11850 15065
rect 11794 14991 11850 15000
rect 11796 14952 11848 14958
rect 11796 14894 11848 14900
rect 11808 12918 11836 14894
rect 11900 14362 11928 15642
rect 11992 15502 12020 15914
rect 12072 15632 12124 15638
rect 12072 15574 12124 15580
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 11980 15360 12032 15366
rect 11978 15328 11980 15337
rect 12032 15328 12034 15337
rect 11978 15263 12034 15272
rect 11980 14884 12032 14890
rect 11980 14826 12032 14832
rect 11992 14793 12020 14826
rect 11978 14784 12034 14793
rect 11978 14719 12034 14728
rect 12084 14482 12112 15574
rect 12176 14822 12204 17138
rect 12268 17066 12296 18770
rect 12360 17814 12388 19520
rect 12348 17808 12400 17814
rect 12348 17750 12400 17756
rect 12532 17740 12584 17746
rect 12532 17682 12584 17688
rect 12346 17368 12402 17377
rect 12346 17303 12402 17312
rect 12256 17060 12308 17066
rect 12256 17002 12308 17008
rect 12268 14890 12296 17002
rect 12360 16658 12388 17303
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12544 16522 12572 17682
rect 12532 16516 12584 16522
rect 12532 16458 12584 16464
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 12544 15609 12572 15982
rect 12728 15638 12756 19520
rect 12912 19502 13124 19520
rect 12808 18012 12860 18018
rect 12808 17954 12860 17960
rect 12820 17066 12848 17954
rect 12808 17060 12860 17066
rect 12808 17002 12860 17008
rect 12912 16726 12940 19502
rect 13556 17610 13584 19520
rect 13924 18834 13952 19520
rect 13912 18828 13964 18834
rect 13912 18770 13964 18776
rect 14004 17672 14056 17678
rect 14004 17614 14056 17620
rect 13544 17604 13596 17610
rect 13544 17546 13596 17552
rect 13282 17436 13578 17456
rect 13338 17434 13362 17436
rect 13418 17434 13442 17436
rect 13498 17434 13522 17436
rect 13360 17382 13362 17434
rect 13424 17382 13436 17434
rect 13498 17382 13500 17434
rect 13338 17380 13362 17382
rect 13418 17380 13442 17382
rect 13498 17380 13522 17382
rect 13282 17360 13578 17380
rect 13174 17232 13230 17241
rect 13174 17167 13230 17176
rect 13636 17196 13688 17202
rect 12900 16720 12952 16726
rect 12900 16662 12952 16668
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 12808 16584 12860 16590
rect 13096 16561 13124 16594
rect 12808 16526 12860 16532
rect 13082 16552 13138 16561
rect 12820 15706 12848 16526
rect 13082 16487 13138 16496
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12992 16040 13044 16046
rect 12992 15982 13044 15988
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 12716 15632 12768 15638
rect 12530 15600 12586 15609
rect 12716 15574 12768 15580
rect 12806 15600 12862 15609
rect 12530 15535 12586 15544
rect 12806 15535 12862 15544
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12624 15496 12676 15502
rect 12624 15438 12676 15444
rect 12256 14884 12308 14890
rect 12256 14826 12308 14832
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 11900 14334 12112 14362
rect 11888 13728 11940 13734
rect 11940 13676 12020 13682
rect 11888 13670 12020 13676
rect 11900 13654 12020 13670
rect 11992 13433 12020 13654
rect 11978 13424 12034 13433
rect 11888 13388 11940 13394
rect 11978 13359 12034 13368
rect 11888 13330 11940 13336
rect 11796 12912 11848 12918
rect 11796 12854 11848 12860
rect 11796 12776 11848 12782
rect 11794 12744 11796 12753
rect 11848 12744 11850 12753
rect 11794 12679 11850 12688
rect 11796 11348 11848 11354
rect 11900 11336 11928 13330
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 11992 12986 12020 13262
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 12084 12866 12112 14334
rect 12268 13841 12296 14418
rect 12254 13832 12310 13841
rect 12164 13796 12216 13802
rect 12254 13767 12310 13776
rect 12164 13738 12216 13744
rect 12176 13433 12204 13738
rect 12360 13682 12388 15438
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12452 14074 12480 14418
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12438 13968 12494 13977
rect 12636 13920 12664 15438
rect 12820 15026 12848 15535
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12808 15020 12860 15026
rect 12808 14962 12860 14968
rect 12728 13938 12756 14962
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12820 14006 12848 14758
rect 12808 14000 12860 14006
rect 12808 13942 12860 13948
rect 12438 13903 12494 13912
rect 12268 13654 12388 13682
rect 12162 13424 12218 13433
rect 12162 13359 12218 13368
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 11992 12838 12112 12866
rect 11992 11898 12020 12838
rect 12176 12714 12204 13262
rect 12164 12708 12216 12714
rect 12164 12650 12216 12656
rect 12268 12594 12296 13654
rect 12346 13152 12402 13161
rect 12346 13087 12402 13096
rect 12084 12566 12296 12594
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 11848 11308 11928 11336
rect 11796 11290 11848 11296
rect 11796 11008 11848 11014
rect 11796 10950 11848 10956
rect 11808 7546 11836 10950
rect 12084 10742 12112 12566
rect 12360 12442 12388 13087
rect 12348 12436 12400 12442
rect 12268 12396 12348 12424
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11900 9110 11928 9318
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 11886 8664 11942 8673
rect 11886 8599 11888 8608
rect 11940 8599 11942 8608
rect 11888 8570 11940 8576
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 11886 7440 11942 7449
rect 11716 7364 11836 7392
rect 11886 7375 11942 7384
rect 11612 7336 11664 7342
rect 11612 7278 11664 7284
rect 11520 6996 11572 7002
rect 11520 6938 11572 6944
rect 11532 5166 11560 6938
rect 11624 5710 11652 7278
rect 11704 7268 11756 7274
rect 11704 7210 11756 7216
rect 11716 7002 11744 7210
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11520 5160 11572 5166
rect 11572 5120 11652 5148
rect 11520 5102 11572 5108
rect 11518 4584 11574 4593
rect 11518 4519 11574 4528
rect 11532 4486 11560 4519
rect 11520 4480 11572 4486
rect 11520 4422 11572 4428
rect 11428 4276 11480 4282
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 10612 3998 10824 4026
rect 10612 3913 10640 3998
rect 10692 3936 10744 3942
rect 10598 3904 10654 3913
rect 10888 3924 10916 4150
rect 10888 3896 11192 3924
rect 10692 3878 10744 3884
rect 10598 3839 10654 3848
rect 10598 3768 10654 3777
rect 10704 3738 10732 3878
rect 10817 3836 11113 3856
rect 10873 3834 10897 3836
rect 10953 3834 10977 3836
rect 11033 3834 11057 3836
rect 10895 3782 10897 3834
rect 10959 3782 10971 3834
rect 11033 3782 11035 3834
rect 10873 3780 10897 3782
rect 10953 3780 10977 3782
rect 11033 3780 11057 3782
rect 10817 3760 11113 3780
rect 10598 3703 10654 3712
rect 10692 3732 10744 3738
rect 10508 3596 10560 3602
rect 10508 3538 10560 3544
rect 10612 3369 10640 3703
rect 10692 3674 10744 3680
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10692 3460 10744 3466
rect 10692 3402 10744 3408
rect 10876 3460 10928 3466
rect 10876 3402 10928 3408
rect 10598 3360 10654 3369
rect 10598 3295 10654 3304
rect 10508 3120 10560 3126
rect 10508 3062 10560 3068
rect 10416 2984 10468 2990
rect 10416 2926 10468 2932
rect 10336 2808 10456 2836
rect 10322 2680 10378 2689
rect 10322 2615 10378 2624
rect 10336 2446 10364 2615
rect 10428 2446 10456 2808
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 10428 2281 10456 2382
rect 10414 2272 10470 2281
rect 10414 2207 10470 2216
rect 10232 1624 10284 1630
rect 10232 1566 10284 1572
rect 10520 480 10548 3062
rect 10600 2984 10652 2990
rect 10600 2926 10652 2932
rect 10612 2825 10640 2926
rect 10598 2816 10654 2825
rect 10598 2751 10654 2760
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 10612 1766 10640 2450
rect 10704 2106 10732 3402
rect 10888 3097 10916 3402
rect 10874 3088 10930 3097
rect 10874 3023 10930 3032
rect 10980 2938 11008 3538
rect 11164 3058 11192 3896
rect 11256 3754 11284 4270
rect 11428 4218 11480 4224
rect 11520 4276 11572 4282
rect 11520 4218 11572 4224
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11348 3942 11376 4082
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11440 3777 11468 4014
rect 11426 3768 11482 3777
rect 11256 3726 11376 3754
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11256 3398 11284 3538
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 10980 2910 11192 2938
rect 10817 2748 11113 2768
rect 10873 2746 10897 2748
rect 10953 2746 10977 2748
rect 11033 2746 11057 2748
rect 10895 2694 10897 2746
rect 10959 2694 10971 2746
rect 11033 2694 11035 2746
rect 10873 2692 10897 2694
rect 10953 2692 10977 2694
rect 11033 2692 11057 2694
rect 10817 2672 11113 2692
rect 10692 2100 10744 2106
rect 10692 2042 10744 2048
rect 10968 1828 11020 1834
rect 10968 1770 11020 1776
rect 10600 1760 10652 1766
rect 10600 1702 10652 1708
rect 10980 480 11008 1770
rect 11164 1630 11192 2910
rect 11244 2916 11296 2922
rect 11244 2858 11296 2864
rect 11256 2689 11284 2858
rect 11242 2680 11298 2689
rect 11242 2615 11298 2624
rect 11152 1624 11204 1630
rect 11152 1566 11204 1572
rect 11348 480 11376 3726
rect 11426 3703 11482 3712
rect 11440 1562 11468 3703
rect 11532 3670 11560 4218
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 11624 3618 11652 5120
rect 11716 4146 11744 6802
rect 11808 5234 11836 7364
rect 11900 7041 11928 7375
rect 11886 7032 11942 7041
rect 11886 6967 11942 6976
rect 11886 6896 11942 6905
rect 11886 6831 11888 6840
rect 11940 6831 11942 6840
rect 11888 6802 11940 6808
rect 11992 6712 12020 10610
rect 12084 9518 12112 10678
rect 12176 10266 12204 12242
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12268 10130 12296 12396
rect 12348 12378 12400 12384
rect 12452 12306 12480 13903
rect 12544 13892 12664 13920
rect 12716 13932 12768 13938
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12360 11354 12388 12038
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12452 11218 12480 12106
rect 12544 12102 12572 13892
rect 12716 13874 12768 13880
rect 12624 13796 12676 13802
rect 12624 13738 12676 13744
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12636 11676 12664 13738
rect 12808 13728 12860 13734
rect 12808 13670 12860 13676
rect 12820 13530 12848 13670
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12716 13456 12768 13462
rect 12716 13398 12768 13404
rect 12728 12986 12756 13398
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12806 12608 12862 12617
rect 12728 12073 12756 12582
rect 12912 12594 12940 15982
rect 13004 14657 13032 15982
rect 13084 15564 13136 15570
rect 13084 15506 13136 15512
rect 12990 14648 13046 14657
rect 12990 14583 13046 14592
rect 12990 14512 13046 14521
rect 12990 14447 13046 14456
rect 13004 14414 13032 14447
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 12990 14240 13046 14249
rect 12990 14175 13046 14184
rect 13004 13394 13032 14175
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 13096 13326 13124 15506
rect 13188 15502 13216 17167
rect 13636 17138 13688 17144
rect 13282 16348 13578 16368
rect 13338 16346 13362 16348
rect 13418 16346 13442 16348
rect 13498 16346 13522 16348
rect 13360 16294 13362 16346
rect 13424 16294 13436 16346
rect 13498 16294 13500 16346
rect 13338 16292 13362 16294
rect 13418 16292 13442 16294
rect 13498 16292 13522 16294
rect 13282 16272 13578 16292
rect 13176 15496 13228 15502
rect 13176 15438 13228 15444
rect 13282 15260 13578 15280
rect 13338 15258 13362 15260
rect 13418 15258 13442 15260
rect 13498 15258 13522 15260
rect 13360 15206 13362 15258
rect 13424 15206 13436 15258
rect 13498 15206 13500 15258
rect 13338 15204 13362 15206
rect 13418 15204 13442 15206
rect 13498 15204 13522 15206
rect 13282 15184 13578 15204
rect 13176 15156 13228 15162
rect 13176 15098 13228 15104
rect 13188 14618 13216 15098
rect 13268 15088 13320 15094
rect 13268 15030 13320 15036
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 13280 14550 13308 15030
rect 13648 14634 13676 17138
rect 13728 17060 13780 17066
rect 13728 17002 13780 17008
rect 13740 15978 13768 17002
rect 14016 16794 14044 17614
rect 14188 17604 14240 17610
rect 14188 17546 14240 17552
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13728 15972 13780 15978
rect 13728 15914 13780 15920
rect 13740 15502 13768 15914
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13728 15360 13780 15366
rect 13728 15302 13780 15308
rect 13556 14606 13676 14634
rect 13268 14544 13320 14550
rect 13268 14486 13320 14492
rect 13176 14272 13228 14278
rect 13556 14260 13584 14606
rect 13740 14550 13768 15302
rect 13924 15162 13952 16594
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 13820 15088 13872 15094
rect 13818 15056 13820 15065
rect 13872 15056 13874 15065
rect 13818 14991 13874 15000
rect 14004 14952 14056 14958
rect 13818 14920 13874 14929
rect 14004 14894 14056 14900
rect 13818 14855 13874 14864
rect 13832 14822 13860 14855
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13728 14544 13780 14550
rect 13728 14486 13780 14492
rect 13636 14476 13688 14482
rect 13636 14418 13688 14424
rect 13648 14385 13676 14418
rect 13634 14376 13690 14385
rect 13634 14311 13690 14320
rect 13556 14232 13676 14260
rect 13176 14214 13228 14220
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 12992 13252 13044 13258
rect 12992 13194 13044 13200
rect 13004 12850 13032 13194
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 13096 12889 13124 13126
rect 13082 12880 13138 12889
rect 12992 12844 13044 12850
rect 13082 12815 13138 12824
rect 12992 12786 13044 12792
rect 12862 12566 12940 12594
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 12806 12543 12862 12552
rect 12714 12064 12770 12073
rect 12714 11999 12770 12008
rect 12544 11648 12664 11676
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12360 10538 12388 11086
rect 12348 10532 12400 10538
rect 12348 10474 12400 10480
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 10266 12480 10406
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 12072 9512 12124 9518
rect 12072 9454 12124 9460
rect 12084 8480 12112 9454
rect 12176 9450 12204 9998
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 12084 8452 12204 8480
rect 12072 8356 12124 8362
rect 12072 8298 12124 8304
rect 11900 6684 12020 6712
rect 11900 5642 11928 6684
rect 11978 6624 12034 6633
rect 11978 6559 12034 6568
rect 11992 6186 12020 6559
rect 11980 6180 12032 6186
rect 11980 6122 12032 6128
rect 11980 5908 12032 5914
rect 12084 5896 12112 8298
rect 12176 6322 12204 8452
rect 12268 7993 12296 8978
rect 12360 8566 12388 10202
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12452 9353 12480 10066
rect 12438 9344 12494 9353
rect 12438 9279 12494 9288
rect 12544 9058 12572 11648
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12714 11520 12770 11529
rect 12636 9518 12664 11494
rect 12714 11455 12770 11464
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 12728 9160 12756 11455
rect 12452 9030 12572 9058
rect 12636 9132 12756 9160
rect 12452 8838 12480 9030
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12440 8832 12492 8838
rect 12544 8809 12572 8910
rect 12440 8774 12492 8780
rect 12530 8800 12586 8809
rect 12348 8560 12400 8566
rect 12348 8502 12400 8508
rect 12346 8256 12402 8265
rect 12346 8191 12402 8200
rect 12360 8022 12388 8191
rect 12348 8016 12400 8022
rect 12254 7984 12310 7993
rect 12348 7958 12400 7964
rect 12254 7919 12310 7928
rect 12360 7818 12388 7958
rect 12348 7812 12400 7818
rect 12348 7754 12400 7760
rect 12256 7540 12308 7546
rect 12308 7500 12388 7528
rect 12256 7482 12308 7488
rect 12254 7440 12310 7449
rect 12254 7375 12256 7384
rect 12308 7375 12310 7384
rect 12256 7346 12308 7352
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12268 6905 12296 7142
rect 12254 6896 12310 6905
rect 12254 6831 12310 6840
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 12032 5868 12112 5896
rect 11980 5850 12032 5856
rect 11888 5636 11940 5642
rect 11888 5578 11940 5584
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11888 5160 11940 5166
rect 11888 5102 11940 5108
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11808 4457 11836 4966
rect 11794 4448 11850 4457
rect 11794 4383 11850 4392
rect 11900 4282 11928 5102
rect 11888 4276 11940 4282
rect 11888 4218 11940 4224
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11886 4040 11942 4049
rect 11886 3975 11888 3984
rect 11940 3975 11942 3984
rect 11888 3946 11940 3952
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11808 3738 11836 3878
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11624 3590 11744 3618
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11518 3360 11574 3369
rect 11518 3295 11574 3304
rect 11532 2825 11560 3295
rect 11624 3126 11652 3470
rect 11716 3398 11744 3590
rect 11992 3584 12020 5850
rect 12070 5672 12126 5681
rect 12176 5642 12204 6258
rect 12360 6202 12388 7500
rect 12268 6174 12388 6202
rect 12070 5607 12126 5616
rect 12164 5636 12216 5642
rect 12084 4078 12112 5607
rect 12164 5578 12216 5584
rect 12268 5522 12296 6174
rect 12348 6112 12400 6118
rect 12346 6080 12348 6089
rect 12400 6080 12402 6089
rect 12346 6015 12402 6024
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12360 5681 12388 5850
rect 12346 5672 12402 5681
rect 12346 5607 12402 5616
rect 12176 5494 12296 5522
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 12176 3777 12204 5494
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12268 5166 12296 5306
rect 12360 5234 12388 5306
rect 12452 5234 12480 8774
rect 12530 8735 12586 8744
rect 12636 8650 12664 9132
rect 12716 8900 12768 8906
rect 12716 8842 12768 8848
rect 12544 8622 12664 8650
rect 12544 8090 12572 8622
rect 12624 8560 12676 8566
rect 12624 8502 12676 8508
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12530 7984 12586 7993
rect 12530 7919 12586 7928
rect 12544 7886 12572 7919
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12544 7177 12572 7822
rect 12636 7313 12664 8502
rect 12728 8362 12756 8842
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12622 7304 12678 7313
rect 12622 7239 12678 7248
rect 12624 7200 12676 7206
rect 12530 7168 12586 7177
rect 12624 7142 12676 7148
rect 12530 7103 12586 7112
rect 12636 7041 12664 7142
rect 12622 7032 12678 7041
rect 12622 6967 12678 6976
rect 12532 6792 12584 6798
rect 12530 6760 12532 6769
rect 12584 6760 12586 6769
rect 12530 6695 12586 6704
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12544 5846 12572 6598
rect 12728 6474 12756 8026
rect 12636 6446 12756 6474
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12532 5704 12584 5710
rect 12532 5646 12584 5652
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 12256 5160 12308 5166
rect 12256 5102 12308 5108
rect 12256 4616 12308 4622
rect 12256 4558 12308 4564
rect 12268 4214 12296 4558
rect 12256 4208 12308 4214
rect 12256 4150 12308 4156
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 12162 3768 12218 3777
rect 12072 3732 12124 3738
rect 12162 3703 12218 3712
rect 12072 3674 12124 3680
rect 11808 3556 12020 3584
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11612 3120 11664 3126
rect 11612 3062 11664 3068
rect 11702 3088 11758 3097
rect 11702 3023 11758 3032
rect 11518 2816 11574 2825
rect 11518 2751 11574 2760
rect 11716 2553 11744 3023
rect 11702 2544 11758 2553
rect 11612 2508 11664 2514
rect 11702 2479 11758 2488
rect 11612 2450 11664 2456
rect 11624 1902 11652 2450
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 11716 2310 11744 2382
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 11612 1896 11664 1902
rect 11612 1838 11664 1844
rect 11428 1556 11480 1562
rect 11428 1498 11480 1504
rect 11808 480 11836 3556
rect 12084 3534 12112 3674
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 11888 3392 11940 3398
rect 11886 3360 11888 3369
rect 11980 3392 12032 3398
rect 11940 3360 11942 3369
rect 11980 3334 12032 3340
rect 11886 3295 11942 3304
rect 11888 2916 11940 2922
rect 11888 2858 11940 2864
rect 11900 2009 11928 2858
rect 11992 2446 12020 3334
rect 12268 2938 12296 3878
rect 12360 2990 12388 5170
rect 12544 4672 12572 5646
rect 12636 5409 12664 6446
rect 12716 6384 12768 6390
rect 12716 6326 12768 6332
rect 12728 5846 12756 6326
rect 12820 6066 12848 12543
rect 12898 12064 12954 12073
rect 12898 11999 12954 12008
rect 12912 11354 12940 11999
rect 13096 11898 13124 12582
rect 13188 12442 13216 14214
rect 13282 14172 13578 14192
rect 13338 14170 13362 14172
rect 13418 14170 13442 14172
rect 13498 14170 13522 14172
rect 13360 14118 13362 14170
rect 13424 14118 13436 14170
rect 13498 14118 13500 14170
rect 13338 14116 13362 14118
rect 13418 14116 13442 14118
rect 13498 14116 13522 14118
rect 13282 14096 13578 14116
rect 13648 14056 13676 14232
rect 13556 14028 13676 14056
rect 13452 14000 13504 14006
rect 13452 13942 13504 13948
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13266 13560 13322 13569
rect 13266 13495 13322 13504
rect 13280 13462 13308 13495
rect 13268 13456 13320 13462
rect 13268 13398 13320 13404
rect 13372 13308 13400 13874
rect 13464 13734 13492 13942
rect 13452 13728 13504 13734
rect 13452 13670 13504 13676
rect 13464 13433 13492 13670
rect 13556 13462 13584 14028
rect 13634 13968 13690 13977
rect 13634 13903 13636 13912
rect 13688 13903 13690 13912
rect 13636 13874 13688 13880
rect 13544 13456 13596 13462
rect 13450 13424 13506 13433
rect 13544 13398 13596 13404
rect 13450 13359 13506 13368
rect 13372 13280 13676 13308
rect 13282 13084 13578 13104
rect 13338 13082 13362 13084
rect 13418 13082 13442 13084
rect 13498 13082 13522 13084
rect 13360 13030 13362 13082
rect 13424 13030 13436 13082
rect 13498 13030 13500 13082
rect 13338 13028 13362 13030
rect 13418 13028 13442 13030
rect 13498 13028 13522 13030
rect 13282 13008 13578 13028
rect 13268 12912 13320 12918
rect 13268 12854 13320 12860
rect 13176 12436 13228 12442
rect 13176 12378 13228 12384
rect 13280 12306 13308 12854
rect 13648 12850 13676 13280
rect 13740 13025 13768 14486
rect 13910 13832 13966 13841
rect 13910 13767 13966 13776
rect 13818 13696 13874 13705
rect 13818 13631 13874 13640
rect 13726 13016 13782 13025
rect 13832 12986 13860 13631
rect 13924 13394 13952 13767
rect 14016 13734 14044 14894
rect 14094 14512 14150 14521
rect 14094 14447 14150 14456
rect 14108 13938 14136 14447
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 14004 13728 14056 13734
rect 14004 13670 14056 13676
rect 14004 13456 14056 13462
rect 14002 13424 14004 13433
rect 14056 13424 14058 13433
rect 13912 13388 13964 13394
rect 14002 13359 14058 13368
rect 13912 13330 13964 13336
rect 13726 12951 13782 12960
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13726 12336 13782 12345
rect 13268 12300 13320 12306
rect 13726 12271 13728 12280
rect 13268 12242 13320 12248
rect 13780 12271 13782 12280
rect 13728 12242 13780 12248
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13282 11996 13578 12016
rect 13338 11994 13362 11996
rect 13418 11994 13442 11996
rect 13498 11994 13522 11996
rect 13360 11942 13362 11994
rect 13424 11942 13436 11994
rect 13498 11942 13500 11994
rect 13338 11940 13362 11942
rect 13418 11940 13442 11942
rect 13498 11940 13522 11942
rect 13282 11920 13578 11940
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12912 10985 12940 11290
rect 12898 10976 12954 10985
rect 12898 10911 12954 10920
rect 12912 10606 12940 10911
rect 13004 10810 13032 11698
rect 13096 11218 13124 11834
rect 13634 11656 13690 11665
rect 13634 11591 13690 11600
rect 13648 11558 13676 11591
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 13096 10674 13124 11154
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12900 10464 12952 10470
rect 12898 10432 12900 10441
rect 12952 10432 12954 10441
rect 12898 10367 12954 10376
rect 12898 10160 12954 10169
rect 12898 10095 12954 10104
rect 12912 7342 12940 10095
rect 13004 9586 13032 10610
rect 13096 10577 13124 10610
rect 13082 10568 13138 10577
rect 13082 10503 13138 10512
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 13096 9722 13124 10066
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 13084 8832 13136 8838
rect 13084 8774 13136 8780
rect 13096 7818 13124 8774
rect 13084 7812 13136 7818
rect 13004 7772 13084 7800
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12912 6225 12940 7142
rect 12898 6216 12954 6225
rect 12898 6151 12954 6160
rect 12820 6038 12940 6066
rect 12716 5840 12768 5846
rect 12716 5782 12768 5788
rect 12808 5704 12860 5710
rect 12714 5672 12770 5681
rect 12808 5646 12860 5652
rect 12714 5607 12770 5616
rect 12622 5400 12678 5409
rect 12622 5335 12678 5344
rect 12728 5234 12756 5607
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12452 4644 12572 4672
rect 12452 3194 12480 4644
rect 12530 4584 12586 4593
rect 12530 4519 12586 4528
rect 12544 4078 12572 4519
rect 12532 4072 12584 4078
rect 12532 4014 12584 4020
rect 12636 3738 12664 5170
rect 12820 4758 12848 5646
rect 12808 4752 12860 4758
rect 12808 4694 12860 4700
rect 12716 4616 12768 4622
rect 12714 4584 12716 4593
rect 12768 4584 12770 4593
rect 12714 4519 12770 4528
rect 12716 4480 12768 4486
rect 12714 4448 12716 4457
rect 12768 4448 12770 4457
rect 12714 4383 12770 4392
rect 12728 4282 12756 4383
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 12714 4176 12770 4185
rect 12770 4134 12848 4162
rect 12714 4111 12770 4120
rect 12820 4010 12848 4134
rect 12808 4004 12860 4010
rect 12808 3946 12860 3952
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12622 3632 12678 3641
rect 12622 3567 12678 3576
rect 12636 3534 12664 3567
rect 12624 3528 12676 3534
rect 12624 3470 12676 3476
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12544 3097 12572 3130
rect 12530 3088 12586 3097
rect 12530 3023 12586 3032
rect 12176 2910 12296 2938
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12176 2854 12204 2910
rect 12164 2848 12216 2854
rect 12348 2848 12400 2854
rect 12164 2790 12216 2796
rect 12268 2808 12348 2836
rect 12268 2650 12296 2808
rect 12348 2790 12400 2796
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 12360 2514 12388 2586
rect 12348 2508 12400 2514
rect 12348 2450 12400 2456
rect 11980 2440 12032 2446
rect 12452 2417 12480 2926
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 12716 2508 12768 2514
rect 12716 2450 12768 2456
rect 11980 2382 12032 2388
rect 12438 2408 12494 2417
rect 12438 2343 12494 2352
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 11886 2000 11942 2009
rect 11992 1970 12020 2246
rect 11886 1935 11942 1944
rect 11980 1964 12032 1970
rect 11900 1850 11928 1935
rect 11980 1906 12032 1912
rect 11900 1822 12204 1850
rect 12636 1834 12664 2450
rect 12176 480 12204 1822
rect 12624 1828 12676 1834
rect 12624 1770 12676 1776
rect 12728 1698 12756 2450
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 12820 2038 12848 2382
rect 12808 2032 12860 2038
rect 12912 2009 12940 6038
rect 13004 5953 13032 7772
rect 13084 7754 13136 7760
rect 13082 7712 13138 7721
rect 13082 7647 13138 7656
rect 13096 6390 13124 7647
rect 13188 7002 13216 11494
rect 13740 11014 13768 12106
rect 13832 11082 13860 12174
rect 13924 12170 13952 13330
rect 14002 13288 14058 13297
rect 14002 13223 14058 13232
rect 14016 12646 14044 13223
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 14200 12481 14228 17546
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 14186 12472 14242 12481
rect 14186 12407 14242 12416
rect 13912 12164 13964 12170
rect 13912 12106 13964 12112
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 13910 11792 13966 11801
rect 13910 11727 13966 11736
rect 13924 11506 13952 11727
rect 14016 11694 14044 12038
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 14096 11552 14148 11558
rect 13924 11478 14044 11506
rect 14200 11529 14228 12407
rect 14292 12209 14320 16594
rect 14384 15366 14412 19520
rect 14554 17912 14610 17921
rect 14554 17847 14610 17856
rect 14568 17202 14596 17847
rect 14556 17196 14608 17202
rect 14556 17138 14608 17144
rect 14556 16040 14608 16046
rect 14462 16008 14518 16017
rect 14556 15982 14608 15988
rect 14462 15943 14518 15952
rect 14372 15360 14424 15366
rect 14372 15302 14424 15308
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14278 12200 14334 12209
rect 14278 12135 14334 12144
rect 14384 11778 14412 14894
rect 14476 12442 14504 15943
rect 14464 12436 14516 12442
rect 14464 12378 14516 12384
rect 14292 11750 14412 11778
rect 14096 11494 14148 11500
rect 14186 11520 14242 11529
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 13728 11008 13780 11014
rect 13728 10950 13780 10956
rect 13282 10908 13578 10928
rect 13338 10906 13362 10908
rect 13418 10906 13442 10908
rect 13498 10906 13522 10908
rect 13360 10854 13362 10906
rect 13424 10854 13436 10906
rect 13498 10854 13500 10906
rect 13338 10852 13362 10854
rect 13418 10852 13442 10854
rect 13498 10852 13522 10854
rect 13282 10832 13578 10852
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13266 10568 13322 10577
rect 13372 10538 13400 10610
rect 13266 10503 13268 10512
rect 13320 10503 13322 10512
rect 13360 10532 13412 10538
rect 13268 10474 13320 10480
rect 13360 10474 13412 10480
rect 13282 9820 13578 9840
rect 13338 9818 13362 9820
rect 13418 9818 13442 9820
rect 13498 9818 13522 9820
rect 13360 9766 13362 9818
rect 13424 9766 13436 9818
rect 13498 9766 13500 9818
rect 13338 9764 13362 9766
rect 13418 9764 13442 9766
rect 13498 9764 13522 9766
rect 13282 9744 13578 9764
rect 13832 9704 13860 10610
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 13556 9676 13860 9704
rect 13452 9512 13504 9518
rect 13450 9480 13452 9489
rect 13504 9480 13506 9489
rect 13450 9415 13506 9424
rect 13556 9042 13584 9676
rect 13818 9616 13874 9625
rect 13818 9551 13874 9560
rect 13634 9208 13690 9217
rect 13634 9143 13690 9152
rect 13648 9042 13676 9143
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13282 8732 13578 8752
rect 13338 8730 13362 8732
rect 13418 8730 13442 8732
rect 13498 8730 13522 8732
rect 13360 8678 13362 8730
rect 13424 8678 13436 8730
rect 13498 8678 13500 8730
rect 13338 8676 13362 8678
rect 13418 8676 13442 8678
rect 13498 8676 13522 8678
rect 13282 8656 13578 8676
rect 13282 7644 13578 7664
rect 13338 7642 13362 7644
rect 13418 7642 13442 7644
rect 13498 7642 13522 7644
rect 13360 7590 13362 7642
rect 13424 7590 13436 7642
rect 13498 7590 13500 7642
rect 13338 7588 13362 7590
rect 13418 7588 13442 7590
rect 13498 7588 13522 7590
rect 13282 7568 13578 7588
rect 13648 7002 13676 8978
rect 13832 8566 13860 9551
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13740 7449 13768 7890
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 13726 7440 13782 7449
rect 13726 7375 13782 7384
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13726 6896 13782 6905
rect 13636 6860 13688 6866
rect 13726 6831 13728 6840
rect 13636 6802 13688 6808
rect 13780 6831 13782 6840
rect 13728 6802 13780 6808
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 13084 6384 13136 6390
rect 13084 6326 13136 6332
rect 12990 5944 13046 5953
rect 12990 5879 13046 5888
rect 12992 5840 13044 5846
rect 13188 5817 13216 6598
rect 13282 6556 13578 6576
rect 13338 6554 13362 6556
rect 13418 6554 13442 6556
rect 13498 6554 13522 6556
rect 13360 6502 13362 6554
rect 13424 6502 13436 6554
rect 13498 6502 13500 6554
rect 13338 6500 13362 6502
rect 13418 6500 13442 6502
rect 13498 6500 13522 6502
rect 13282 6480 13578 6500
rect 13648 6458 13676 6802
rect 13832 6746 13860 7822
rect 13924 7410 13952 10406
rect 14016 10266 14044 11478
rect 14108 11354 14136 11494
rect 14186 11455 14242 11464
rect 14096 11348 14148 11354
rect 14292 11336 14320 11750
rect 14372 11620 14424 11626
rect 14372 11562 14424 11568
rect 14384 11354 14412 11562
rect 14464 11552 14516 11558
rect 14464 11494 14516 11500
rect 14096 11290 14148 11296
rect 14200 11308 14320 11336
rect 14372 11348 14424 11354
rect 14004 10260 14056 10266
rect 14200 10248 14228 11308
rect 14372 11290 14424 11296
rect 14278 11248 14334 11257
rect 14278 11183 14280 11192
rect 14332 11183 14334 11192
rect 14372 11212 14424 11218
rect 14280 11154 14332 11160
rect 14372 11154 14424 11160
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14004 10202 14056 10208
rect 14108 10220 14228 10248
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 14016 9654 14044 10066
rect 14004 9648 14056 9654
rect 14002 9616 14004 9625
rect 14056 9616 14058 9625
rect 14002 9551 14058 9560
rect 14016 9525 14044 9551
rect 14108 9466 14136 10220
rect 14186 10024 14242 10033
rect 14186 9959 14188 9968
rect 14240 9959 14242 9968
rect 14188 9930 14240 9936
rect 14016 9438 14136 9466
rect 14016 8838 14044 9438
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14004 8832 14056 8838
rect 14004 8774 14056 8780
rect 14108 8634 14136 9318
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 14200 8498 14228 9930
rect 14292 9450 14320 10542
rect 14384 10198 14412 11154
rect 14372 10192 14424 10198
rect 14372 10134 14424 10140
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14280 9444 14332 9450
rect 14280 9386 14332 9392
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14004 8288 14056 8294
rect 14004 8230 14056 8236
rect 14016 8090 14044 8230
rect 14004 8084 14056 8090
rect 14004 8026 14056 8032
rect 14188 7812 14240 7818
rect 14188 7754 14240 7760
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 13910 7304 13966 7313
rect 13910 7239 13966 7248
rect 13740 6718 13860 6746
rect 13636 6452 13688 6458
rect 13636 6394 13688 6400
rect 13268 6316 13320 6322
rect 13268 6258 13320 6264
rect 12992 5782 13044 5788
rect 13174 5808 13230 5817
rect 13004 5234 13032 5782
rect 13280 5778 13308 6258
rect 13740 6186 13768 6718
rect 13728 6180 13780 6186
rect 13728 6122 13780 6128
rect 13636 6112 13688 6118
rect 13450 6080 13506 6089
rect 13636 6054 13688 6060
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13450 6015 13506 6024
rect 13464 5914 13492 6015
rect 13542 5944 13598 5953
rect 13452 5908 13504 5914
rect 13542 5879 13598 5888
rect 13452 5850 13504 5856
rect 13556 5846 13584 5879
rect 13544 5840 13596 5846
rect 13544 5782 13596 5788
rect 13174 5743 13230 5752
rect 13268 5772 13320 5778
rect 13268 5714 13320 5720
rect 13648 5681 13676 6054
rect 13634 5672 13690 5681
rect 13176 5636 13228 5642
rect 13634 5607 13690 5616
rect 13176 5578 13228 5584
rect 13082 5536 13138 5545
rect 13082 5471 13138 5480
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 13096 5166 13124 5471
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 13004 2990 13032 4966
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 13096 4282 13124 4762
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 13096 3058 13124 4082
rect 13188 3602 13216 5578
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13282 5468 13578 5488
rect 13338 5466 13362 5468
rect 13418 5466 13442 5468
rect 13498 5466 13522 5468
rect 13360 5414 13362 5466
rect 13424 5414 13436 5466
rect 13498 5414 13500 5466
rect 13338 5412 13362 5414
rect 13418 5412 13442 5414
rect 13498 5412 13522 5414
rect 13282 5392 13578 5412
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13266 4992 13322 5001
rect 13266 4927 13322 4936
rect 13280 4826 13308 4927
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 13372 4622 13400 5170
rect 13636 5160 13688 5166
rect 13740 5137 13768 5510
rect 13636 5102 13688 5108
rect 13726 5128 13782 5137
rect 13544 5092 13596 5098
rect 13544 5034 13596 5040
rect 13450 4856 13506 4865
rect 13556 4826 13584 5034
rect 13450 4791 13506 4800
rect 13544 4820 13596 4826
rect 13464 4758 13492 4791
rect 13544 4762 13596 4768
rect 13452 4752 13504 4758
rect 13452 4694 13504 4700
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13282 4380 13578 4400
rect 13338 4378 13362 4380
rect 13418 4378 13442 4380
rect 13498 4378 13522 4380
rect 13360 4326 13362 4378
rect 13424 4326 13436 4378
rect 13498 4326 13500 4378
rect 13338 4324 13362 4326
rect 13418 4324 13442 4326
rect 13498 4324 13522 4326
rect 13282 4304 13578 4324
rect 13268 4208 13320 4214
rect 13648 4185 13676 5102
rect 13726 5063 13782 5072
rect 13728 5024 13780 5030
rect 13728 4966 13780 4972
rect 13268 4150 13320 4156
rect 13634 4176 13690 4185
rect 13280 3738 13308 4150
rect 13634 4111 13690 4120
rect 13360 4072 13412 4078
rect 13360 4014 13412 4020
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13266 3632 13322 3641
rect 13176 3596 13228 3602
rect 13266 3567 13268 3576
rect 13176 3538 13228 3544
rect 13320 3567 13322 3576
rect 13268 3538 13320 3544
rect 13372 3482 13400 4014
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13188 3454 13400 3482
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 12992 2984 13044 2990
rect 12992 2926 13044 2932
rect 12990 2408 13046 2417
rect 12990 2343 13046 2352
rect 12808 1974 12860 1980
rect 12898 2000 12954 2009
rect 12898 1935 12954 1944
rect 12716 1692 12768 1698
rect 12716 1634 12768 1640
rect 12622 1456 12678 1465
rect 12622 1391 12678 1400
rect 12636 678 12664 1391
rect 12624 672 12676 678
rect 12624 614 12676 620
rect 12636 480 12664 614
rect 13004 480 13032 2343
rect 13096 1086 13124 2994
rect 13188 2106 13216 3454
rect 13282 3292 13578 3312
rect 13338 3290 13362 3292
rect 13418 3290 13442 3292
rect 13498 3290 13522 3292
rect 13360 3238 13362 3290
rect 13424 3238 13436 3290
rect 13498 3238 13500 3290
rect 13338 3236 13362 3238
rect 13418 3236 13442 3238
rect 13498 3236 13522 3238
rect 13282 3216 13578 3236
rect 13268 3120 13320 3126
rect 13268 3062 13320 3068
rect 13280 2650 13308 3062
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 13648 2582 13676 3878
rect 13636 2576 13688 2582
rect 13740 2553 13768 4966
rect 13832 3505 13860 6054
rect 13924 3738 13952 7239
rect 14016 7206 14044 7686
rect 14200 7410 14228 7754
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14186 7304 14242 7313
rect 14186 7239 14242 7248
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 14096 6928 14148 6934
rect 14096 6870 14148 6876
rect 14002 6760 14058 6769
rect 14002 6695 14058 6704
rect 14016 4010 14044 6695
rect 14004 4004 14056 4010
rect 14004 3946 14056 3952
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 13818 3496 13874 3505
rect 13818 3431 13874 3440
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13636 2518 13688 2524
rect 13726 2544 13782 2553
rect 13726 2479 13782 2488
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 13282 2204 13578 2224
rect 13338 2202 13362 2204
rect 13418 2202 13442 2204
rect 13498 2202 13522 2204
rect 13360 2150 13362 2202
rect 13424 2150 13436 2202
rect 13498 2150 13500 2202
rect 13338 2148 13362 2150
rect 13418 2148 13442 2150
rect 13498 2148 13522 2150
rect 13282 2128 13578 2148
rect 13176 2100 13228 2106
rect 13176 2042 13228 2048
rect 13740 1902 13768 2382
rect 13728 1896 13780 1902
rect 13728 1838 13780 1844
rect 13450 1320 13506 1329
rect 13450 1255 13506 1264
rect 13084 1080 13136 1086
rect 13084 1022 13136 1028
rect 13464 480 13492 1255
rect 13832 480 13860 3334
rect 13924 3126 13952 3674
rect 13912 3120 13964 3126
rect 13912 3062 13964 3068
rect 14004 3120 14056 3126
rect 14004 3062 14056 3068
rect 14016 2854 14044 3062
rect 14108 2990 14136 6870
rect 14200 6866 14228 7239
rect 14188 6860 14240 6866
rect 14188 6802 14240 6808
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 14096 2984 14148 2990
rect 14096 2926 14148 2932
rect 14004 2848 14056 2854
rect 14004 2790 14056 2796
rect 14200 2378 14228 6122
rect 14292 3942 14320 9386
rect 14384 7546 14412 9998
rect 14476 9081 14504 11494
rect 14568 11121 14596 15982
rect 14646 14784 14702 14793
rect 14646 14719 14702 14728
rect 14554 11112 14610 11121
rect 14554 11047 14610 11056
rect 14556 11008 14608 11014
rect 14556 10950 14608 10956
rect 14462 9072 14518 9081
rect 14462 9007 14518 9016
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14476 8566 14504 8910
rect 14464 8560 14516 8566
rect 14464 8502 14516 8508
rect 14464 8356 14516 8362
rect 14464 8298 14516 8304
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 14384 2972 14412 7142
rect 14476 4690 14504 8298
rect 14568 5778 14596 10950
rect 14660 7342 14688 14719
rect 14752 12918 14780 19520
rect 15120 18222 15148 19520
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 15120 15858 15148 18158
rect 14832 14884 14884 14890
rect 14832 14826 14884 14832
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 14752 12442 14780 12854
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14752 6730 14780 12242
rect 14844 11694 14872 14826
rect 14936 12306 14964 15846
rect 15120 15830 15240 15858
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 14924 12300 14976 12306
rect 14924 12242 14976 12248
rect 15028 11914 15056 15506
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 14936 11886 15056 11914
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14844 7954 14872 11630
rect 14832 7948 14884 7954
rect 14832 7890 14884 7896
rect 14832 6996 14884 7002
rect 14832 6938 14884 6944
rect 14740 6724 14792 6730
rect 14660 6684 14740 6712
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 14660 5352 14688 6684
rect 14740 6666 14792 6672
rect 14738 5944 14794 5953
rect 14738 5879 14794 5888
rect 14568 5324 14688 5352
rect 14464 4684 14516 4690
rect 14464 4626 14516 4632
rect 14462 4040 14518 4049
rect 14462 3975 14518 3984
rect 14476 3602 14504 3975
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14568 3398 14596 5324
rect 14646 5264 14702 5273
rect 14646 5199 14702 5208
rect 14660 4826 14688 5199
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14646 3904 14702 3913
rect 14646 3839 14702 3848
rect 14660 3738 14688 3839
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 14752 3058 14780 5879
rect 14844 5030 14872 6938
rect 14832 5024 14884 5030
rect 14832 4966 14884 4972
rect 14936 3126 14964 11886
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 15028 8537 15056 9318
rect 15014 8528 15070 8537
rect 15014 8463 15070 8472
rect 15120 8430 15148 12378
rect 15212 11286 15240 15830
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15292 14476 15344 14482
rect 15292 14418 15344 14424
rect 15304 12374 15332 14418
rect 15292 12368 15344 12374
rect 15292 12310 15344 12316
rect 15200 11280 15252 11286
rect 15200 11222 15252 11228
rect 15198 10568 15254 10577
rect 15198 10503 15254 10512
rect 15108 8424 15160 8430
rect 15014 8392 15070 8401
rect 15108 8366 15160 8372
rect 15014 8327 15070 8336
rect 15028 8294 15056 8327
rect 15016 8288 15068 8294
rect 15016 8230 15068 8236
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 15028 6361 15056 7142
rect 15014 6352 15070 6361
rect 15014 6287 15070 6296
rect 15016 5024 15068 5030
rect 15016 4966 15068 4972
rect 15028 4593 15056 4966
rect 15120 4729 15148 8366
rect 15106 4720 15162 4729
rect 15106 4655 15162 4664
rect 15014 4584 15070 4593
rect 15014 4519 15070 4528
rect 15120 4010 15148 4655
rect 15108 4004 15160 4010
rect 15108 3946 15160 3952
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 14924 3120 14976 3126
rect 15028 3097 15056 3878
rect 15212 3670 15240 10503
rect 15200 3664 15252 3670
rect 15200 3606 15252 3612
rect 14924 3062 14976 3068
rect 15014 3088 15070 3097
rect 14740 3052 14792 3058
rect 15014 3023 15070 3032
rect 14740 2994 14792 3000
rect 14292 2944 14412 2972
rect 14556 2984 14608 2990
rect 14188 2372 14240 2378
rect 14188 2314 14240 2320
rect 14292 480 14320 2944
rect 14832 2984 14884 2990
rect 14556 2926 14608 2932
rect 14738 2952 14794 2961
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 14476 2106 14504 2450
rect 14464 2100 14516 2106
rect 14464 2042 14516 2048
rect 14568 1601 14596 2926
rect 14648 2916 14700 2922
rect 14832 2926 14884 2932
rect 14738 2887 14794 2896
rect 14648 2858 14700 2864
rect 14554 1592 14610 1601
rect 14554 1527 14610 1536
rect 14660 480 14688 2858
rect 14752 2854 14780 2887
rect 14740 2848 14792 2854
rect 14844 2825 14872 2926
rect 15108 2916 15160 2922
rect 15108 2858 15160 2864
rect 14740 2790 14792 2796
rect 14830 2816 14886 2825
rect 14830 2751 14886 2760
rect 15120 2582 15148 2858
rect 15304 2854 15332 12310
rect 15396 9738 15424 14962
rect 15488 9897 15516 15438
rect 15580 14006 15608 19520
rect 15948 17649 15976 19520
rect 15934 17640 15990 17649
rect 15934 17575 15990 17584
rect 15568 14000 15620 14006
rect 15568 13942 15620 13948
rect 15948 10606 15976 17575
rect 16408 14890 16436 19520
rect 16776 16114 16804 19520
rect 16764 16108 16816 16114
rect 16764 16050 16816 16056
rect 16396 14884 16448 14890
rect 16396 14826 16448 14832
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 15474 9888 15530 9897
rect 15474 9823 15530 9832
rect 15396 9710 15516 9738
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 15108 2576 15160 2582
rect 15108 2518 15160 2524
rect 15488 1766 15516 9710
rect 15568 8968 15620 8974
rect 15568 8910 15620 8916
rect 15580 2689 15608 8910
rect 15936 3664 15988 3670
rect 15936 3606 15988 3612
rect 15566 2680 15622 2689
rect 15566 2615 15622 2624
rect 15476 1760 15528 1766
rect 15476 1702 15528 1708
rect 15108 1556 15160 1562
rect 15108 1498 15160 1504
rect 15120 480 15148 1498
rect 15488 480 15516 1702
rect 15948 480 15976 3606
rect 16764 2916 16816 2922
rect 16764 2858 16816 2864
rect 16304 1624 16356 1630
rect 16304 1566 16356 1572
rect 16316 480 16344 1566
rect 16776 480 16804 2858
rect 3146 439 3202 448
rect 3514 0 3570 480
rect 3882 0 3938 480
rect 4342 0 4398 480
rect 4710 0 4766 480
rect 5170 0 5226 480
rect 5538 0 5594 480
rect 5998 0 6054 480
rect 6366 0 6422 480
rect 6826 0 6882 480
rect 7194 0 7250 480
rect 7654 0 7710 480
rect 8022 0 8078 480
rect 8482 0 8538 480
rect 8850 0 8906 480
rect 9310 0 9366 480
rect 9678 0 9734 480
rect 10138 0 10194 480
rect 10506 0 10562 480
rect 10966 0 11022 480
rect 11334 0 11390 480
rect 11794 0 11850 480
rect 12162 0 12218 480
rect 12622 0 12678 480
rect 12990 0 13046 480
rect 13450 0 13506 480
rect 13818 0 13874 480
rect 14278 0 14334 480
rect 14646 0 14702 480
rect 15106 0 15162 480
rect 15474 0 15530 480
rect 15934 0 15990 480
rect 16302 0 16358 480
rect 16762 0 16818 480
<< via2 >>
rect 2134 16632 2190 16688
rect 1582 13252 1638 13288
rect 1582 13232 1584 13252
rect 1584 13232 1636 13252
rect 1636 13232 1638 13252
rect 1398 10124 1454 10160
rect 1398 10104 1400 10124
rect 1400 10104 1452 10124
rect 1452 10104 1454 10124
rect 570 9968 626 10024
rect 1214 6160 1270 6216
rect 1122 4256 1178 4312
rect 1030 3440 1086 3496
rect 1858 15680 1914 15736
rect 1858 11872 1914 11928
rect 2318 16088 2374 16144
rect 1950 11192 2006 11248
rect 1858 10512 1914 10568
rect 1674 9424 1730 9480
rect 1766 7792 1822 7848
rect 2042 8880 2098 8936
rect 2502 15000 2558 15056
rect 2870 19488 2926 19544
rect 2778 17584 2834 17640
rect 3514 18536 3570 18592
rect 2778 15544 2834 15600
rect 2594 14864 2650 14920
rect 2502 12688 2558 12744
rect 2318 12416 2374 12472
rect 2318 11636 2320 11656
rect 2320 11636 2372 11656
rect 2372 11636 2374 11656
rect 2318 11600 2374 11636
rect 1950 7248 2006 7304
rect 1858 6160 1914 6216
rect 1858 5752 1914 5808
rect 1674 2488 1730 2544
rect 1214 1944 1270 2000
rect 2042 5072 2098 5128
rect 2502 10240 2558 10296
rect 3421 17434 3477 17436
rect 3501 17434 3557 17436
rect 3581 17434 3637 17436
rect 3661 17434 3717 17436
rect 3421 17382 3447 17434
rect 3447 17382 3477 17434
rect 3501 17382 3511 17434
rect 3511 17382 3557 17434
rect 3581 17382 3627 17434
rect 3627 17382 3637 17434
rect 3661 17382 3691 17434
rect 3691 17382 3717 17434
rect 3421 17380 3477 17382
rect 3501 17380 3557 17382
rect 3581 17380 3637 17382
rect 3661 17380 3717 17382
rect 3146 16496 3202 16552
rect 3238 15952 3294 16008
rect 3146 15408 3202 15464
rect 3054 14728 3110 14784
rect 2962 14320 3018 14376
rect 2870 12824 2926 12880
rect 2778 12144 2834 12200
rect 2686 9968 2742 10024
rect 2778 9016 2834 9072
rect 2594 6840 2650 6896
rect 2502 6704 2558 6760
rect 2778 5652 2780 5672
rect 2780 5652 2832 5672
rect 2832 5652 2834 5672
rect 2778 5616 2834 5652
rect 2686 3984 2742 4040
rect 2962 8472 3018 8528
rect 3146 12280 3202 12336
rect 3054 8064 3110 8120
rect 2962 4548 3018 4584
rect 2962 4528 2964 4548
rect 2964 4528 3016 4548
rect 3016 4528 3018 4548
rect 2870 2644 2926 2680
rect 2870 2624 2872 2644
rect 2872 2624 2924 2644
rect 2924 2624 2926 2644
rect 3054 3304 3110 3360
rect 3054 3032 3110 3088
rect 2778 1400 2834 1456
rect 3790 16632 3846 16688
rect 3421 16346 3477 16348
rect 3501 16346 3557 16348
rect 3581 16346 3637 16348
rect 3661 16346 3717 16348
rect 3421 16294 3447 16346
rect 3447 16294 3477 16346
rect 3501 16294 3511 16346
rect 3511 16294 3557 16346
rect 3581 16294 3627 16346
rect 3627 16294 3637 16346
rect 3661 16294 3691 16346
rect 3691 16294 3717 16346
rect 3421 16292 3477 16294
rect 3501 16292 3557 16294
rect 3581 16292 3637 16294
rect 3661 16292 3717 16294
rect 4342 16360 4398 16416
rect 4066 16124 4068 16144
rect 4068 16124 4120 16144
rect 4120 16124 4122 16144
rect 4066 16088 4122 16124
rect 3514 15852 3516 15872
rect 3516 15852 3568 15872
rect 3568 15852 3570 15872
rect 3514 15816 3570 15852
rect 3422 15408 3478 15464
rect 3421 15258 3477 15260
rect 3501 15258 3557 15260
rect 3581 15258 3637 15260
rect 3661 15258 3717 15260
rect 3421 15206 3447 15258
rect 3447 15206 3477 15258
rect 3501 15206 3511 15258
rect 3511 15206 3557 15258
rect 3581 15206 3627 15258
rect 3627 15206 3637 15258
rect 3661 15206 3691 15258
rect 3691 15206 3717 15258
rect 3421 15204 3477 15206
rect 3501 15204 3557 15206
rect 3581 15204 3637 15206
rect 3661 15204 3717 15206
rect 3790 14320 3846 14376
rect 3421 14170 3477 14172
rect 3501 14170 3557 14172
rect 3581 14170 3637 14172
rect 3661 14170 3717 14172
rect 3421 14118 3447 14170
rect 3447 14118 3477 14170
rect 3501 14118 3511 14170
rect 3511 14118 3557 14170
rect 3581 14118 3627 14170
rect 3627 14118 3637 14170
rect 3661 14118 3691 14170
rect 3691 14118 3717 14170
rect 3421 14116 3477 14118
rect 3501 14116 3557 14118
rect 3581 14116 3637 14118
rect 3661 14116 3717 14118
rect 3422 13640 3478 13696
rect 3882 14184 3938 14240
rect 3882 13776 3938 13832
rect 3421 13082 3477 13084
rect 3501 13082 3557 13084
rect 3581 13082 3637 13084
rect 3661 13082 3717 13084
rect 3421 13030 3447 13082
rect 3447 13030 3477 13082
rect 3501 13030 3511 13082
rect 3511 13030 3557 13082
rect 3581 13030 3627 13082
rect 3627 13030 3637 13082
rect 3661 13030 3691 13082
rect 3691 13030 3717 13082
rect 3421 13028 3477 13030
rect 3501 13028 3557 13030
rect 3581 13028 3637 13030
rect 3661 13028 3717 13030
rect 3421 11994 3477 11996
rect 3501 11994 3557 11996
rect 3581 11994 3637 11996
rect 3661 11994 3717 11996
rect 3421 11942 3447 11994
rect 3447 11942 3477 11994
rect 3501 11942 3511 11994
rect 3511 11942 3557 11994
rect 3581 11942 3627 11994
rect 3627 11942 3637 11994
rect 3661 11942 3691 11994
rect 3691 11942 3717 11994
rect 3421 11940 3477 11942
rect 3501 11940 3557 11942
rect 3581 11940 3637 11942
rect 3661 11940 3717 11942
rect 3698 11056 3754 11112
rect 3421 10906 3477 10908
rect 3501 10906 3557 10908
rect 3581 10906 3637 10908
rect 3661 10906 3717 10908
rect 3421 10854 3447 10906
rect 3447 10854 3477 10906
rect 3501 10854 3511 10906
rect 3511 10854 3557 10906
rect 3581 10854 3627 10906
rect 3627 10854 3637 10906
rect 3661 10854 3691 10906
rect 3691 10854 3717 10906
rect 3421 10852 3477 10854
rect 3501 10852 3557 10854
rect 3581 10852 3637 10854
rect 3661 10852 3717 10854
rect 3606 10648 3662 10704
rect 3606 10104 3662 10160
rect 3421 9818 3477 9820
rect 3501 9818 3557 9820
rect 3581 9818 3637 9820
rect 3661 9818 3717 9820
rect 3421 9766 3447 9818
rect 3447 9766 3477 9818
rect 3501 9766 3511 9818
rect 3511 9766 3557 9818
rect 3581 9766 3627 9818
rect 3627 9766 3637 9818
rect 3661 9766 3691 9818
rect 3691 9766 3717 9818
rect 3421 9764 3477 9766
rect 3501 9764 3557 9766
rect 3581 9764 3637 9766
rect 3661 9764 3717 9766
rect 3606 9560 3662 9616
rect 3421 8730 3477 8732
rect 3501 8730 3557 8732
rect 3581 8730 3637 8732
rect 3661 8730 3717 8732
rect 3421 8678 3447 8730
rect 3447 8678 3477 8730
rect 3501 8678 3511 8730
rect 3511 8678 3557 8730
rect 3581 8678 3627 8730
rect 3627 8678 3637 8730
rect 3661 8678 3691 8730
rect 3691 8678 3717 8730
rect 3421 8676 3477 8678
rect 3501 8676 3557 8678
rect 3581 8676 3637 8678
rect 3661 8676 3717 8678
rect 3790 7928 3846 7984
rect 3421 7642 3477 7644
rect 3501 7642 3557 7644
rect 3581 7642 3637 7644
rect 3661 7642 3717 7644
rect 3421 7590 3447 7642
rect 3447 7590 3477 7642
rect 3501 7590 3511 7642
rect 3511 7590 3557 7642
rect 3581 7590 3627 7642
rect 3627 7590 3637 7642
rect 3661 7590 3691 7642
rect 3691 7590 3717 7642
rect 3421 7588 3477 7590
rect 3501 7588 3557 7590
rect 3581 7588 3637 7590
rect 3661 7588 3717 7590
rect 3421 6554 3477 6556
rect 3501 6554 3557 6556
rect 3581 6554 3637 6556
rect 3661 6554 3717 6556
rect 3421 6502 3447 6554
rect 3447 6502 3477 6554
rect 3501 6502 3511 6554
rect 3511 6502 3557 6554
rect 3581 6502 3627 6554
rect 3627 6502 3637 6554
rect 3661 6502 3691 6554
rect 3691 6502 3717 6554
rect 3421 6500 3477 6502
rect 3501 6500 3557 6502
rect 3581 6500 3637 6502
rect 3661 6500 3717 6502
rect 3790 6296 3846 6352
rect 3330 6024 3386 6080
rect 3421 5466 3477 5468
rect 3501 5466 3557 5468
rect 3581 5466 3637 5468
rect 3661 5466 3717 5468
rect 3421 5414 3447 5466
rect 3447 5414 3477 5466
rect 3501 5414 3511 5466
rect 3511 5414 3557 5466
rect 3581 5414 3627 5466
rect 3627 5414 3637 5466
rect 3661 5414 3691 5466
rect 3691 5414 3717 5466
rect 3421 5412 3477 5414
rect 3501 5412 3557 5414
rect 3581 5412 3637 5414
rect 3661 5412 3717 5414
rect 3514 4800 3570 4856
rect 3421 4378 3477 4380
rect 3501 4378 3557 4380
rect 3581 4378 3637 4380
rect 3661 4378 3717 4380
rect 3421 4326 3447 4378
rect 3447 4326 3477 4378
rect 3501 4326 3511 4378
rect 3511 4326 3557 4378
rect 3581 4326 3627 4378
rect 3627 4326 3637 4378
rect 3661 4326 3691 4378
rect 3691 4326 3717 4378
rect 3421 4324 3477 4326
rect 3501 4324 3557 4326
rect 3581 4324 3637 4326
rect 3661 4324 3717 4326
rect 3238 3596 3294 3632
rect 3238 3576 3240 3596
rect 3240 3576 3292 3596
rect 3292 3576 3294 3596
rect 3606 3712 3662 3768
rect 3421 3290 3477 3292
rect 3501 3290 3557 3292
rect 3581 3290 3637 3292
rect 3661 3290 3717 3292
rect 3421 3238 3447 3290
rect 3447 3238 3477 3290
rect 3501 3238 3511 3290
rect 3511 3238 3557 3290
rect 3581 3238 3627 3290
rect 3627 3238 3637 3290
rect 3661 3238 3691 3290
rect 3691 3238 3717 3290
rect 3421 3236 3477 3238
rect 3501 3236 3557 3238
rect 3581 3236 3637 3238
rect 3661 3236 3717 3238
rect 3422 2896 3478 2952
rect 4342 15272 4398 15328
rect 4434 15000 4490 15056
rect 4250 14592 4306 14648
rect 4066 13640 4122 13696
rect 4250 13640 4306 13696
rect 4158 13504 4214 13560
rect 4066 11872 4122 11928
rect 4066 10376 4122 10432
rect 4434 14492 4436 14512
rect 4436 14492 4488 14512
rect 4488 14492 4490 14512
rect 4434 14456 4490 14492
rect 4710 15816 4766 15872
rect 4710 15680 4766 15736
rect 4618 14728 4674 14784
rect 4618 13776 4674 13832
rect 4894 16768 4950 16824
rect 4894 16360 4950 16416
rect 4894 15952 4950 16008
rect 4986 15816 5042 15872
rect 4066 10004 4068 10024
rect 4068 10004 4120 10024
rect 4120 10004 4122 10024
rect 4066 9968 4122 10004
rect 4158 8336 4214 8392
rect 4158 5752 4214 5808
rect 4066 5072 4122 5128
rect 3974 4256 4030 4312
rect 3974 3304 4030 3360
rect 4710 13368 4766 13424
rect 4526 9968 4582 10024
rect 4618 9832 4674 9888
rect 4434 5788 4436 5808
rect 4436 5788 4488 5808
rect 4488 5788 4490 5808
rect 4434 5752 4490 5788
rect 4618 4664 4674 4720
rect 4986 13912 5042 13968
rect 4894 12180 4896 12200
rect 4896 12180 4948 12200
rect 4948 12180 4950 12200
rect 4894 12144 4950 12180
rect 5538 15408 5594 15464
rect 5262 14456 5318 14512
rect 5886 16890 5942 16892
rect 5966 16890 6022 16892
rect 6046 16890 6102 16892
rect 6126 16890 6182 16892
rect 5886 16838 5912 16890
rect 5912 16838 5942 16890
rect 5966 16838 5976 16890
rect 5976 16838 6022 16890
rect 6046 16838 6092 16890
rect 6092 16838 6102 16890
rect 6126 16838 6156 16890
rect 6156 16838 6182 16890
rect 5886 16836 5942 16838
rect 5966 16836 6022 16838
rect 6046 16836 6102 16838
rect 6126 16836 6182 16838
rect 5814 15952 5870 16008
rect 6274 15852 6276 15872
rect 6276 15852 6328 15872
rect 6328 15852 6330 15872
rect 6274 15816 6330 15852
rect 5886 15802 5942 15804
rect 5966 15802 6022 15804
rect 6046 15802 6102 15804
rect 6126 15802 6182 15804
rect 5886 15750 5912 15802
rect 5912 15750 5942 15802
rect 5966 15750 5976 15802
rect 5976 15750 6022 15802
rect 6046 15750 6092 15802
rect 6092 15750 6102 15802
rect 6126 15750 6156 15802
rect 6156 15750 6182 15802
rect 5886 15748 5942 15750
rect 5966 15748 6022 15750
rect 6046 15748 6102 15750
rect 6126 15748 6182 15750
rect 6734 16940 6736 16960
rect 6736 16940 6788 16960
rect 6788 16940 6790 16960
rect 6734 16904 6790 16940
rect 7286 17176 7342 17232
rect 6642 15408 6698 15464
rect 5886 14714 5942 14716
rect 5966 14714 6022 14716
rect 6046 14714 6102 14716
rect 6126 14714 6182 14716
rect 5886 14662 5912 14714
rect 5912 14662 5942 14714
rect 5966 14662 5976 14714
rect 5976 14662 6022 14714
rect 6046 14662 6092 14714
rect 6092 14662 6102 14714
rect 6126 14662 6156 14714
rect 6156 14662 6182 14714
rect 5886 14660 5942 14662
rect 5966 14660 6022 14662
rect 6046 14660 6102 14662
rect 6126 14660 6182 14662
rect 5538 13640 5594 13696
rect 5446 13504 5502 13560
rect 5354 12416 5410 12472
rect 4894 10240 4950 10296
rect 5446 11736 5502 11792
rect 5446 11348 5502 11384
rect 5446 11328 5448 11348
rect 5448 11328 5500 11348
rect 5500 11328 5502 11348
rect 5354 11076 5410 11112
rect 5354 11056 5356 11076
rect 5356 11056 5408 11076
rect 5408 11056 5410 11076
rect 5630 12588 5632 12608
rect 5632 12588 5684 12608
rect 5684 12588 5686 12608
rect 5630 12552 5686 12588
rect 4894 9696 4950 9752
rect 5354 9832 5410 9888
rect 5078 8880 5134 8936
rect 5170 7540 5226 7576
rect 5170 7520 5172 7540
rect 5172 7520 5224 7540
rect 5224 7520 5226 7540
rect 5078 7112 5134 7168
rect 4710 4256 4766 4312
rect 4250 2896 4306 2952
rect 3421 2202 3477 2204
rect 3501 2202 3557 2204
rect 3581 2202 3637 2204
rect 3661 2202 3717 2204
rect 3421 2150 3447 2202
rect 3447 2150 3477 2202
rect 3501 2150 3511 2202
rect 3511 2150 3557 2202
rect 3581 2150 3627 2202
rect 3627 2150 3637 2202
rect 3661 2150 3691 2202
rect 3691 2150 3717 2202
rect 3421 2148 3477 2150
rect 3501 2148 3557 2150
rect 3581 2148 3637 2150
rect 3661 2148 3717 2150
rect 4342 2796 4344 2816
rect 4344 2796 4396 2816
rect 4396 2796 4398 2816
rect 4342 2760 4398 2796
rect 4066 1808 4122 1864
rect 3882 1672 3938 1728
rect 3514 1536 3570 1592
rect 3238 1400 3294 1456
rect 3146 448 3202 504
rect 4342 1128 4398 1184
rect 4802 3576 4858 3632
rect 4802 2352 4858 2408
rect 4986 4664 5042 4720
rect 5170 5616 5226 5672
rect 5078 4256 5134 4312
rect 4986 2080 5042 2136
rect 5538 8744 5594 8800
rect 5354 4936 5410 4992
rect 5906 14184 5962 14240
rect 5886 13626 5942 13628
rect 5966 13626 6022 13628
rect 6046 13626 6102 13628
rect 6126 13626 6182 13628
rect 5886 13574 5912 13626
rect 5912 13574 5942 13626
rect 5966 13574 5976 13626
rect 5976 13574 6022 13626
rect 6046 13574 6092 13626
rect 6092 13574 6102 13626
rect 6126 13574 6156 13626
rect 6156 13574 6182 13626
rect 5886 13572 5942 13574
rect 5966 13572 6022 13574
rect 6046 13572 6102 13574
rect 6126 13572 6182 13574
rect 6458 14728 6514 14784
rect 5814 12960 5870 13016
rect 5814 12688 5870 12744
rect 5722 11872 5778 11928
rect 5886 12538 5942 12540
rect 5966 12538 6022 12540
rect 6046 12538 6102 12540
rect 6126 12538 6182 12540
rect 5886 12486 5912 12538
rect 5912 12486 5942 12538
rect 5966 12486 5976 12538
rect 5976 12486 6022 12538
rect 6046 12486 6092 12538
rect 6092 12486 6102 12538
rect 6126 12486 6156 12538
rect 6156 12486 6182 12538
rect 5886 12484 5942 12486
rect 5966 12484 6022 12486
rect 6046 12484 6102 12486
rect 6126 12484 6182 12486
rect 6550 13912 6606 13968
rect 6458 12688 6514 12744
rect 6458 12436 6514 12472
rect 6458 12416 6460 12436
rect 6460 12416 6512 12436
rect 6512 12416 6514 12436
rect 6642 13640 6698 13696
rect 6826 15680 6882 15736
rect 6918 15136 6974 15192
rect 6734 13504 6790 13560
rect 6274 11464 6330 11520
rect 5886 11450 5942 11452
rect 5966 11450 6022 11452
rect 6046 11450 6102 11452
rect 6126 11450 6182 11452
rect 5886 11398 5912 11450
rect 5912 11398 5942 11450
rect 5966 11398 5976 11450
rect 5976 11398 6022 11450
rect 6046 11398 6092 11450
rect 6092 11398 6102 11450
rect 6126 11398 6156 11450
rect 6156 11398 6182 11450
rect 5886 11396 5942 11398
rect 5966 11396 6022 11398
rect 6046 11396 6102 11398
rect 6126 11396 6182 11398
rect 5886 10362 5942 10364
rect 5966 10362 6022 10364
rect 6046 10362 6102 10364
rect 6126 10362 6182 10364
rect 5886 10310 5912 10362
rect 5912 10310 5942 10362
rect 5966 10310 5976 10362
rect 5976 10310 6022 10362
rect 6046 10310 6092 10362
rect 6092 10310 6102 10362
rect 6126 10310 6156 10362
rect 6156 10310 6182 10362
rect 5886 10308 5942 10310
rect 5966 10308 6022 10310
rect 6046 10308 6102 10310
rect 6126 10308 6182 10310
rect 5998 9716 6054 9752
rect 5998 9696 6000 9716
rect 6000 9696 6052 9716
rect 6052 9696 6054 9716
rect 6274 9596 6276 9616
rect 6276 9596 6328 9616
rect 6328 9596 6330 9616
rect 6274 9560 6330 9596
rect 5886 9274 5942 9276
rect 5966 9274 6022 9276
rect 6046 9274 6102 9276
rect 6126 9274 6182 9276
rect 5886 9222 5912 9274
rect 5912 9222 5942 9274
rect 5966 9222 5976 9274
rect 5976 9222 6022 9274
rect 6046 9222 6092 9274
rect 6092 9222 6102 9274
rect 6126 9222 6156 9274
rect 6156 9222 6182 9274
rect 5886 9220 5942 9222
rect 5966 9220 6022 9222
rect 6046 9220 6102 9222
rect 6126 9220 6182 9222
rect 5886 8186 5942 8188
rect 5966 8186 6022 8188
rect 6046 8186 6102 8188
rect 6126 8186 6182 8188
rect 5886 8134 5912 8186
rect 5912 8134 5942 8186
rect 5966 8134 5976 8186
rect 5976 8134 6022 8186
rect 6046 8134 6092 8186
rect 6092 8134 6102 8186
rect 6126 8134 6156 8186
rect 6156 8134 6182 8186
rect 5886 8132 5942 8134
rect 5966 8132 6022 8134
rect 6046 8132 6102 8134
rect 6126 8132 6182 8134
rect 5998 7384 6054 7440
rect 5886 7098 5942 7100
rect 5966 7098 6022 7100
rect 6046 7098 6102 7100
rect 6126 7098 6182 7100
rect 5886 7046 5912 7098
rect 5912 7046 5942 7098
rect 5966 7046 5976 7098
rect 5976 7046 6022 7098
rect 6046 7046 6092 7098
rect 6092 7046 6102 7098
rect 6126 7046 6156 7098
rect 6156 7046 6182 7098
rect 5886 7044 5942 7046
rect 5966 7044 6022 7046
rect 6046 7044 6102 7046
rect 6126 7044 6182 7046
rect 5630 6840 5686 6896
rect 5814 6432 5870 6488
rect 5886 6010 5942 6012
rect 5966 6010 6022 6012
rect 6046 6010 6102 6012
rect 6126 6010 6182 6012
rect 5886 5958 5912 6010
rect 5912 5958 5942 6010
rect 5966 5958 5976 6010
rect 5976 5958 6022 6010
rect 6046 5958 6092 6010
rect 6092 5958 6102 6010
rect 6126 5958 6156 6010
rect 6156 5958 6182 6010
rect 5886 5956 5942 5958
rect 5966 5956 6022 5958
rect 6046 5956 6102 5958
rect 6126 5956 6182 5958
rect 5354 4392 5410 4448
rect 5722 4800 5778 4856
rect 5886 4922 5942 4924
rect 5966 4922 6022 4924
rect 6046 4922 6102 4924
rect 6126 4922 6182 4924
rect 5886 4870 5912 4922
rect 5912 4870 5942 4922
rect 5966 4870 5976 4922
rect 5976 4870 6022 4922
rect 6046 4870 6092 4922
rect 6092 4870 6102 4922
rect 6126 4870 6156 4922
rect 6156 4870 6182 4922
rect 5886 4868 5942 4870
rect 5966 4868 6022 4870
rect 6046 4868 6102 4870
rect 6126 4868 6182 4870
rect 7010 14728 7066 14784
rect 7194 14728 7250 14784
rect 7194 14592 7250 14648
rect 7194 14048 7250 14104
rect 7010 13776 7066 13832
rect 7194 13368 7250 13424
rect 8206 17584 8262 17640
rect 8352 17434 8408 17436
rect 8432 17434 8488 17436
rect 8512 17434 8568 17436
rect 8592 17434 8648 17436
rect 8352 17382 8378 17434
rect 8378 17382 8408 17434
rect 8432 17382 8442 17434
rect 8442 17382 8488 17434
rect 8512 17382 8558 17434
rect 8558 17382 8568 17434
rect 8592 17382 8622 17434
rect 8622 17382 8648 17434
rect 8352 17380 8408 17382
rect 8432 17380 8488 17382
rect 8512 17380 8568 17382
rect 8592 17380 8648 17382
rect 7930 16360 7986 16416
rect 7746 15816 7802 15872
rect 8114 16768 8170 16824
rect 8482 17060 8538 17096
rect 8482 17040 8484 17060
rect 8484 17040 8536 17060
rect 8536 17040 8538 17060
rect 8574 16632 8630 16688
rect 7194 12824 7250 12880
rect 6918 12280 6974 12336
rect 6734 11328 6790 11384
rect 6918 10920 6974 10976
rect 6642 9560 6698 9616
rect 6550 7656 6606 7712
rect 7286 12144 7342 12200
rect 7470 12144 7526 12200
rect 7470 10784 7526 10840
rect 7930 13096 7986 13152
rect 7838 12824 7894 12880
rect 7838 12416 7894 12472
rect 8352 16346 8408 16348
rect 8432 16346 8488 16348
rect 8512 16346 8568 16348
rect 8592 16346 8648 16348
rect 8352 16294 8378 16346
rect 8378 16294 8408 16346
rect 8432 16294 8442 16346
rect 8442 16294 8488 16346
rect 8512 16294 8558 16346
rect 8558 16294 8568 16346
rect 8592 16294 8622 16346
rect 8622 16294 8648 16346
rect 8352 16292 8408 16294
rect 8432 16292 8488 16294
rect 8512 16292 8568 16294
rect 8592 16292 8648 16294
rect 8352 15258 8408 15260
rect 8432 15258 8488 15260
rect 8512 15258 8568 15260
rect 8592 15258 8648 15260
rect 8352 15206 8378 15258
rect 8378 15206 8408 15258
rect 8432 15206 8442 15258
rect 8442 15206 8488 15258
rect 8512 15206 8558 15258
rect 8558 15206 8568 15258
rect 8592 15206 8622 15258
rect 8622 15206 8648 15258
rect 8352 15204 8408 15206
rect 8432 15204 8488 15206
rect 8512 15204 8568 15206
rect 8592 15204 8648 15206
rect 8942 17892 8944 17912
rect 8944 17892 8996 17912
rect 8996 17892 8998 17912
rect 8942 17856 8998 17892
rect 8482 14728 8538 14784
rect 8666 14320 8722 14376
rect 8352 14170 8408 14172
rect 8432 14170 8488 14172
rect 8512 14170 8568 14172
rect 8592 14170 8648 14172
rect 8352 14118 8378 14170
rect 8378 14118 8408 14170
rect 8432 14118 8442 14170
rect 8442 14118 8488 14170
rect 8512 14118 8558 14170
rect 8558 14118 8568 14170
rect 8592 14118 8622 14170
rect 8622 14118 8648 14170
rect 8352 14116 8408 14118
rect 8432 14116 8488 14118
rect 8512 14116 8568 14118
rect 8592 14116 8648 14118
rect 8390 13504 8446 13560
rect 8942 15136 8998 15192
rect 8942 14184 8998 14240
rect 8758 13504 8814 13560
rect 8758 13096 8814 13152
rect 8352 13082 8408 13084
rect 8432 13082 8488 13084
rect 8512 13082 8568 13084
rect 8592 13082 8648 13084
rect 8352 13030 8378 13082
rect 8378 13030 8408 13082
rect 8432 13030 8442 13082
rect 8442 13030 8488 13082
rect 8512 13030 8558 13082
rect 8558 13030 8568 13082
rect 8592 13030 8622 13082
rect 8622 13030 8648 13082
rect 8352 13028 8408 13030
rect 8432 13028 8488 13030
rect 8512 13028 8568 13030
rect 8592 13028 8648 13030
rect 7838 12008 7894 12064
rect 8114 11872 8170 11928
rect 7838 10512 7894 10568
rect 7102 8472 7158 8528
rect 5446 3168 5502 3224
rect 5354 2896 5410 2952
rect 5814 4256 5870 4312
rect 5998 4256 6054 4312
rect 6366 3848 6422 3904
rect 5886 3834 5942 3836
rect 5966 3834 6022 3836
rect 6046 3834 6102 3836
rect 6126 3834 6182 3836
rect 5886 3782 5912 3834
rect 5912 3782 5942 3834
rect 5966 3782 5976 3834
rect 5976 3782 6022 3834
rect 6046 3782 6092 3834
rect 6092 3782 6102 3834
rect 6126 3782 6156 3834
rect 6156 3782 6182 3834
rect 5886 3780 5942 3782
rect 5966 3780 6022 3782
rect 6046 3780 6102 3782
rect 6126 3780 6182 3782
rect 6090 3304 6146 3360
rect 5722 2760 5778 2816
rect 5886 2746 5942 2748
rect 5966 2746 6022 2748
rect 6046 2746 6102 2748
rect 6126 2746 6182 2748
rect 5886 2694 5912 2746
rect 5912 2694 5942 2746
rect 5966 2694 5976 2746
rect 5976 2694 6022 2746
rect 6046 2694 6092 2746
rect 6092 2694 6102 2746
rect 6126 2694 6156 2746
rect 6156 2694 6182 2746
rect 5886 2692 5942 2694
rect 5966 2692 6022 2694
rect 6046 2692 6102 2694
rect 6126 2692 6182 2694
rect 5446 2488 5502 2544
rect 5630 2488 5686 2544
rect 6458 2488 6514 2544
rect 6734 6704 6790 6760
rect 7010 6296 7066 6352
rect 6642 5072 6698 5128
rect 6642 4936 6698 4992
rect 6642 3848 6698 3904
rect 6642 3712 6698 3768
rect 6826 3848 6882 3904
rect 6734 2216 6790 2272
rect 7010 5208 7066 5264
rect 7010 4392 7066 4448
rect 7010 3848 7066 3904
rect 6918 3304 6974 3360
rect 7286 8064 7342 8120
rect 7286 7656 7342 7712
rect 7562 7692 7564 7712
rect 7564 7692 7616 7712
rect 7616 7692 7618 7712
rect 7562 7656 7618 7692
rect 7746 7384 7802 7440
rect 7470 6704 7526 6760
rect 7654 6432 7710 6488
rect 7562 5344 7618 5400
rect 7654 5072 7710 5128
rect 7470 4120 7526 4176
rect 7194 3168 7250 3224
rect 7194 2760 7250 2816
rect 7102 2352 7158 2408
rect 7378 3188 7434 3224
rect 7378 3168 7380 3188
rect 7380 3168 7432 3188
rect 7432 3168 7434 3188
rect 7930 5480 7986 5536
rect 7930 4256 7986 4312
rect 8352 11994 8408 11996
rect 8432 11994 8488 11996
rect 8512 11994 8568 11996
rect 8592 11994 8648 11996
rect 8352 11942 8378 11994
rect 8378 11942 8408 11994
rect 8432 11942 8442 11994
rect 8442 11942 8488 11994
rect 8512 11942 8558 11994
rect 8558 11942 8568 11994
rect 8592 11942 8622 11994
rect 8622 11942 8648 11994
rect 8352 11940 8408 11942
rect 8432 11940 8488 11942
rect 8512 11940 8568 11942
rect 8592 11940 8648 11942
rect 8206 11328 8262 11384
rect 8850 12008 8906 12064
rect 9402 17312 9458 17368
rect 9310 16768 9366 16824
rect 9126 14592 9182 14648
rect 9126 14320 9182 14376
rect 9494 16904 9550 16960
rect 9770 16632 9826 16688
rect 10414 17196 10470 17232
rect 10414 17176 10416 17196
rect 10416 17176 10468 17196
rect 10468 17176 10470 17196
rect 9494 16360 9550 16416
rect 9678 16224 9734 16280
rect 9402 15816 9458 15872
rect 9678 15680 9734 15736
rect 9310 14728 9366 14784
rect 9126 14048 9182 14104
rect 9494 15408 9550 15464
rect 9494 15136 9550 15192
rect 10046 15816 10102 15872
rect 10138 15408 10194 15464
rect 9678 14592 9734 14648
rect 9862 14592 9918 14648
rect 9034 11328 9090 11384
rect 8352 10906 8408 10908
rect 8432 10906 8488 10908
rect 8512 10906 8568 10908
rect 8592 10906 8648 10908
rect 8352 10854 8378 10906
rect 8378 10854 8408 10906
rect 8432 10854 8442 10906
rect 8442 10854 8488 10906
rect 8512 10854 8558 10906
rect 8558 10854 8568 10906
rect 8592 10854 8622 10906
rect 8622 10854 8648 10906
rect 8352 10852 8408 10854
rect 8432 10852 8488 10854
rect 8512 10852 8568 10854
rect 8592 10852 8648 10854
rect 9218 12552 9274 12608
rect 9678 12960 9734 13016
rect 9678 12416 9734 12472
rect 9586 12280 9642 12336
rect 9218 12008 9274 12064
rect 8352 9818 8408 9820
rect 8432 9818 8488 9820
rect 8512 9818 8568 9820
rect 8592 9818 8648 9820
rect 8352 9766 8378 9818
rect 8378 9766 8408 9818
rect 8432 9766 8442 9818
rect 8442 9766 8488 9818
rect 8512 9766 8558 9818
rect 8558 9766 8568 9818
rect 8592 9766 8622 9818
rect 8622 9766 8648 9818
rect 8352 9764 8408 9766
rect 8432 9764 8488 9766
rect 8512 9764 8568 9766
rect 8592 9764 8648 9766
rect 8114 9288 8170 9344
rect 8206 8780 8208 8800
rect 8208 8780 8260 8800
rect 8260 8780 8262 8800
rect 8206 8744 8262 8780
rect 8352 8730 8408 8732
rect 8432 8730 8488 8732
rect 8512 8730 8568 8732
rect 8592 8730 8648 8732
rect 8352 8678 8378 8730
rect 8378 8678 8408 8730
rect 8432 8678 8442 8730
rect 8442 8678 8488 8730
rect 8512 8678 8558 8730
rect 8558 8678 8568 8730
rect 8592 8678 8622 8730
rect 8622 8678 8648 8730
rect 8352 8676 8408 8678
rect 8432 8676 8488 8678
rect 8512 8676 8568 8678
rect 8592 8676 8648 8678
rect 8114 7656 8170 7712
rect 8352 7642 8408 7644
rect 8432 7642 8488 7644
rect 8512 7642 8568 7644
rect 8592 7642 8648 7644
rect 8352 7590 8378 7642
rect 8378 7590 8408 7642
rect 8432 7590 8442 7642
rect 8442 7590 8488 7642
rect 8512 7590 8558 7642
rect 8558 7590 8568 7642
rect 8592 7590 8622 7642
rect 8622 7590 8648 7642
rect 8352 7588 8408 7590
rect 8432 7588 8488 7590
rect 8512 7588 8568 7590
rect 8592 7588 8648 7590
rect 8206 7520 8262 7576
rect 9034 10920 9090 10976
rect 8942 10376 8998 10432
rect 8850 8608 8906 8664
rect 8850 8200 8906 8256
rect 8850 8064 8906 8120
rect 8352 6554 8408 6556
rect 8432 6554 8488 6556
rect 8512 6554 8568 6556
rect 8592 6554 8648 6556
rect 8352 6502 8378 6554
rect 8378 6502 8408 6554
rect 8432 6502 8442 6554
rect 8442 6502 8488 6554
rect 8512 6502 8558 6554
rect 8558 6502 8568 6554
rect 8592 6502 8622 6554
rect 8622 6502 8648 6554
rect 8352 6500 8408 6502
rect 8432 6500 8488 6502
rect 8512 6500 8568 6502
rect 8592 6500 8648 6502
rect 8206 6060 8208 6080
rect 8208 6060 8260 6080
rect 8260 6060 8262 6080
rect 8206 6024 8262 6060
rect 8114 5480 8170 5536
rect 7562 2760 7618 2816
rect 7930 3168 7986 3224
rect 7838 2896 7894 2952
rect 7470 2488 7526 2544
rect 8022 2896 8078 2952
rect 8352 5466 8408 5468
rect 8432 5466 8488 5468
rect 8512 5466 8568 5468
rect 8592 5466 8648 5468
rect 8352 5414 8378 5466
rect 8378 5414 8408 5466
rect 8432 5414 8442 5466
rect 8442 5414 8488 5466
rect 8512 5414 8558 5466
rect 8558 5414 8568 5466
rect 8592 5414 8622 5466
rect 8622 5414 8648 5466
rect 8352 5412 8408 5414
rect 8432 5412 8488 5414
rect 8512 5412 8568 5414
rect 8592 5412 8648 5414
rect 8482 5208 8538 5264
rect 8352 4378 8408 4380
rect 8432 4378 8488 4380
rect 8512 4378 8568 4380
rect 8592 4378 8648 4380
rect 8352 4326 8378 4378
rect 8378 4326 8408 4378
rect 8432 4326 8442 4378
rect 8442 4326 8488 4378
rect 8512 4326 8558 4378
rect 8558 4326 8568 4378
rect 8592 4326 8622 4378
rect 8622 4326 8648 4378
rect 8352 4324 8408 4326
rect 8432 4324 8488 4326
rect 8512 4324 8568 4326
rect 8592 4324 8648 4326
rect 8298 4120 8354 4176
rect 8482 3440 8538 3496
rect 7930 2624 7986 2680
rect 8022 2488 8078 2544
rect 8352 3290 8408 3292
rect 8432 3290 8488 3292
rect 8512 3290 8568 3292
rect 8592 3290 8648 3292
rect 8352 3238 8378 3290
rect 8378 3238 8408 3290
rect 8432 3238 8442 3290
rect 8442 3238 8488 3290
rect 8512 3238 8558 3290
rect 8558 3238 8568 3290
rect 8592 3238 8622 3290
rect 8622 3238 8648 3290
rect 8352 3236 8408 3238
rect 8432 3236 8488 3238
rect 8512 3236 8568 3238
rect 8592 3236 8648 3238
rect 8574 2932 8576 2952
rect 8576 2932 8628 2952
rect 8628 2932 8630 2952
rect 8574 2896 8630 2932
rect 7838 2080 7894 2136
rect 7930 1944 7986 2000
rect 8482 2488 8538 2544
rect 9310 10648 9366 10704
rect 9034 10240 9090 10296
rect 9218 9832 9274 9888
rect 9126 9696 9182 9752
rect 9034 6568 9090 6624
rect 9034 6296 9090 6352
rect 9034 5888 9090 5944
rect 10322 15136 10378 15192
rect 9954 12960 10010 13016
rect 9678 11056 9734 11112
rect 9770 10784 9826 10840
rect 9586 9152 9642 9208
rect 9218 6432 9274 6488
rect 9402 6568 9458 6624
rect 9586 6840 9642 6896
rect 10138 12416 10194 12472
rect 10046 11056 10102 11112
rect 9954 10240 10010 10296
rect 9862 8236 9864 8256
rect 9864 8236 9916 8256
rect 9916 8236 9918 8256
rect 9862 8200 9918 8236
rect 9034 5616 9090 5672
rect 9034 4120 9090 4176
rect 9126 3476 9128 3496
rect 9128 3476 9180 3496
rect 9180 3476 9182 3496
rect 9126 3440 9182 3476
rect 9770 5480 9826 5536
rect 9770 4800 9826 4856
rect 9954 6568 10010 6624
rect 9954 5072 10010 5128
rect 10414 14728 10470 14784
rect 10817 16890 10873 16892
rect 10897 16890 10953 16892
rect 10977 16890 11033 16892
rect 11057 16890 11113 16892
rect 10817 16838 10843 16890
rect 10843 16838 10873 16890
rect 10897 16838 10907 16890
rect 10907 16838 10953 16890
rect 10977 16838 11023 16890
rect 11023 16838 11033 16890
rect 11057 16838 11087 16890
rect 11087 16838 11113 16890
rect 10817 16836 10873 16838
rect 10897 16836 10953 16838
rect 10977 16836 11033 16838
rect 11057 16836 11113 16838
rect 10874 16224 10930 16280
rect 10817 15802 10873 15804
rect 10897 15802 10953 15804
rect 10977 15802 11033 15804
rect 11057 15802 11113 15804
rect 10817 15750 10843 15802
rect 10843 15750 10873 15802
rect 10897 15750 10907 15802
rect 10907 15750 10953 15802
rect 10977 15750 11023 15802
rect 11023 15750 11033 15802
rect 11057 15750 11087 15802
rect 11087 15750 11113 15802
rect 10817 15748 10873 15750
rect 10897 15748 10953 15750
rect 10977 15748 11033 15750
rect 11057 15748 11113 15750
rect 11334 16496 11390 16552
rect 10874 15408 10930 15464
rect 10598 15272 10654 15328
rect 10506 14592 10562 14648
rect 11058 15136 11114 15192
rect 10817 14714 10873 14716
rect 10897 14714 10953 14716
rect 10977 14714 11033 14716
rect 11057 14714 11113 14716
rect 10817 14662 10843 14714
rect 10843 14662 10873 14714
rect 10897 14662 10907 14714
rect 10907 14662 10953 14714
rect 10977 14662 11023 14714
rect 11023 14662 11033 14714
rect 11057 14662 11087 14714
rect 11087 14662 11113 14714
rect 10817 14660 10873 14662
rect 10897 14660 10953 14662
rect 10977 14660 11033 14662
rect 11057 14660 11113 14662
rect 10414 13504 10470 13560
rect 10414 12960 10470 13016
rect 10230 11328 10286 11384
rect 10598 13504 10654 13560
rect 10817 13626 10873 13628
rect 10897 13626 10953 13628
rect 10977 13626 11033 13628
rect 11057 13626 11113 13628
rect 10817 13574 10843 13626
rect 10843 13574 10873 13626
rect 10897 13574 10907 13626
rect 10907 13574 10953 13626
rect 10977 13574 11023 13626
rect 11023 13574 11033 13626
rect 11057 13574 11087 13626
rect 11087 13574 11113 13626
rect 10817 13572 10873 13574
rect 10897 13572 10953 13574
rect 10977 13572 11033 13574
rect 11057 13572 11113 13574
rect 11518 15680 11574 15736
rect 11426 14592 11482 14648
rect 11426 14048 11482 14104
rect 11334 13676 11336 13696
rect 11336 13676 11388 13696
rect 11388 13676 11390 13696
rect 11334 13640 11390 13676
rect 11334 13504 11390 13560
rect 11150 12960 11206 13016
rect 10506 11328 10562 11384
rect 10506 10684 10508 10704
rect 10508 10684 10560 10704
rect 10560 10684 10562 10704
rect 10506 10648 10562 10684
rect 10817 12538 10873 12540
rect 10897 12538 10953 12540
rect 10977 12538 11033 12540
rect 11057 12538 11113 12540
rect 10817 12486 10843 12538
rect 10843 12486 10873 12538
rect 10897 12486 10907 12538
rect 10907 12486 10953 12538
rect 10977 12486 11023 12538
rect 11023 12486 11033 12538
rect 11057 12486 11087 12538
rect 11087 12486 11113 12538
rect 10817 12484 10873 12486
rect 10897 12484 10953 12486
rect 10977 12484 11033 12486
rect 11057 12484 11113 12486
rect 11242 12552 11298 12608
rect 10874 12008 10930 12064
rect 10966 11772 10968 11792
rect 10968 11772 11020 11792
rect 11020 11772 11022 11792
rect 10966 11736 11022 11772
rect 11426 13368 11482 13424
rect 11426 13096 11482 13152
rect 11334 11736 11390 11792
rect 10817 11450 10873 11452
rect 10897 11450 10953 11452
rect 10977 11450 11033 11452
rect 11057 11450 11113 11452
rect 10817 11398 10843 11450
rect 10843 11398 10873 11450
rect 10897 11398 10907 11450
rect 10907 11398 10953 11450
rect 10977 11398 11023 11450
rect 11023 11398 11033 11450
rect 11057 11398 11087 11450
rect 11087 11398 11113 11450
rect 10817 11396 10873 11398
rect 10897 11396 10953 11398
rect 10977 11396 11033 11398
rect 11057 11396 11113 11398
rect 11334 11464 11390 11520
rect 11058 10784 11114 10840
rect 10414 10376 10470 10432
rect 10817 10362 10873 10364
rect 10897 10362 10953 10364
rect 10977 10362 11033 10364
rect 11057 10362 11113 10364
rect 10817 10310 10843 10362
rect 10843 10310 10873 10362
rect 10897 10310 10907 10362
rect 10907 10310 10953 10362
rect 10977 10310 11023 10362
rect 11023 10310 11033 10362
rect 11057 10310 11087 10362
rect 11087 10310 11113 10362
rect 10817 10308 10873 10310
rect 10897 10308 10953 10310
rect 10977 10308 11033 10310
rect 11057 10308 11113 10310
rect 10506 9288 10562 9344
rect 10817 9274 10873 9276
rect 10897 9274 10953 9276
rect 10977 9274 11033 9276
rect 11057 9274 11113 9276
rect 10817 9222 10843 9274
rect 10843 9222 10873 9274
rect 10897 9222 10907 9274
rect 10907 9222 10953 9274
rect 10977 9222 11023 9274
rect 11023 9222 11033 9274
rect 11057 9222 11087 9274
rect 11087 9222 11113 9274
rect 10817 9220 10873 9222
rect 10897 9220 10953 9222
rect 10977 9220 11033 9222
rect 11057 9220 11113 9222
rect 10138 6976 10194 7032
rect 10506 6976 10562 7032
rect 10230 5480 10286 5536
rect 10817 8186 10873 8188
rect 10897 8186 10953 8188
rect 10977 8186 11033 8188
rect 11057 8186 11113 8188
rect 10817 8134 10843 8186
rect 10843 8134 10873 8186
rect 10897 8134 10907 8186
rect 10907 8134 10953 8186
rect 10977 8134 11023 8186
rect 11023 8134 11033 8186
rect 11057 8134 11087 8186
rect 11087 8134 11113 8186
rect 10817 8132 10873 8134
rect 10897 8132 10953 8134
rect 10977 8132 11033 8134
rect 11057 8132 11113 8134
rect 10690 7520 10746 7576
rect 10966 7248 11022 7304
rect 10817 7098 10873 7100
rect 10897 7098 10953 7100
rect 10977 7098 11033 7100
rect 11057 7098 11113 7100
rect 10817 7046 10843 7098
rect 10843 7046 10873 7098
rect 10897 7046 10907 7098
rect 10907 7046 10953 7098
rect 10977 7046 11023 7098
rect 11023 7046 11033 7098
rect 11057 7046 11087 7098
rect 11087 7046 11113 7098
rect 10817 7044 10873 7046
rect 10897 7044 10953 7046
rect 10977 7044 11033 7046
rect 11057 7044 11113 7046
rect 10414 6024 10470 6080
rect 10138 4766 10194 4822
rect 9586 4120 9642 4176
rect 9402 3440 9458 3496
rect 8352 2202 8408 2204
rect 8432 2202 8488 2204
rect 8512 2202 8568 2204
rect 8592 2202 8648 2204
rect 8352 2150 8378 2202
rect 8378 2150 8408 2202
rect 8432 2150 8442 2202
rect 8442 2150 8488 2202
rect 8512 2150 8558 2202
rect 8558 2150 8568 2202
rect 8592 2150 8622 2202
rect 8622 2150 8648 2202
rect 8352 2148 8408 2150
rect 8432 2148 8488 2150
rect 8512 2148 8568 2150
rect 8592 2148 8648 2150
rect 8482 1264 8538 1320
rect 10046 3848 10102 3904
rect 9770 3576 9826 3632
rect 9494 2080 9550 2136
rect 10506 5888 10562 5944
rect 10782 6568 10838 6624
rect 10598 5480 10654 5536
rect 10817 6010 10873 6012
rect 10897 6010 10953 6012
rect 10977 6010 11033 6012
rect 11057 6010 11113 6012
rect 10817 5958 10843 6010
rect 10843 5958 10873 6010
rect 10897 5958 10907 6010
rect 10907 5958 10953 6010
rect 10977 5958 11023 6010
rect 11023 5958 11033 6010
rect 11057 5958 11087 6010
rect 11087 5958 11113 6010
rect 10817 5956 10873 5958
rect 10897 5956 10953 5958
rect 10977 5956 11033 5958
rect 11057 5956 11113 5958
rect 10874 5752 10930 5808
rect 10782 5480 10838 5536
rect 11150 5208 11206 5264
rect 10322 4664 10378 4720
rect 10817 4922 10873 4924
rect 10897 4922 10953 4924
rect 10977 4922 11033 4924
rect 11057 4922 11113 4924
rect 10817 4870 10843 4922
rect 10843 4870 10873 4922
rect 10897 4870 10907 4922
rect 10907 4870 10953 4922
rect 10977 4870 11023 4922
rect 11023 4870 11033 4922
rect 11057 4870 11087 4922
rect 11087 4870 11113 4922
rect 10817 4868 10873 4870
rect 10897 4868 10953 4870
rect 10977 4868 11033 4870
rect 11057 4868 11113 4870
rect 11334 7112 11390 7168
rect 10230 3712 10286 3768
rect 10230 3032 10286 3088
rect 10046 2624 10102 2680
rect 10138 2488 10194 2544
rect 9954 2352 10010 2408
rect 11058 4528 11114 4584
rect 11242 4528 11298 4584
rect 11794 17856 11850 17912
rect 11610 12960 11666 13016
rect 11794 16904 11850 16960
rect 12070 16108 12126 16144
rect 12070 16088 12072 16108
rect 12072 16088 12124 16108
rect 12124 16088 12126 16108
rect 11794 15000 11850 15056
rect 11978 15308 11980 15328
rect 11980 15308 12032 15328
rect 12032 15308 12034 15328
rect 11978 15272 12034 15308
rect 11978 14728 12034 14784
rect 12346 17312 12402 17368
rect 13282 17434 13338 17436
rect 13362 17434 13418 17436
rect 13442 17434 13498 17436
rect 13522 17434 13578 17436
rect 13282 17382 13308 17434
rect 13308 17382 13338 17434
rect 13362 17382 13372 17434
rect 13372 17382 13418 17434
rect 13442 17382 13488 17434
rect 13488 17382 13498 17434
rect 13522 17382 13552 17434
rect 13552 17382 13578 17434
rect 13282 17380 13338 17382
rect 13362 17380 13418 17382
rect 13442 17380 13498 17382
rect 13522 17380 13578 17382
rect 13174 17176 13230 17232
rect 13082 16496 13138 16552
rect 12530 15544 12586 15600
rect 12806 15544 12862 15600
rect 11978 13368 12034 13424
rect 11794 12724 11796 12744
rect 11796 12724 11848 12744
rect 11848 12724 11850 12744
rect 11794 12688 11850 12724
rect 12254 13776 12310 13832
rect 12438 13912 12494 13968
rect 12162 13368 12218 13424
rect 12346 13096 12402 13152
rect 11886 8628 11942 8664
rect 11886 8608 11888 8628
rect 11888 8608 11940 8628
rect 11940 8608 11942 8628
rect 11886 7384 11942 7440
rect 11518 4528 11574 4584
rect 10598 3848 10654 3904
rect 10598 3712 10654 3768
rect 10817 3834 10873 3836
rect 10897 3834 10953 3836
rect 10977 3834 11033 3836
rect 11057 3834 11113 3836
rect 10817 3782 10843 3834
rect 10843 3782 10873 3834
rect 10897 3782 10907 3834
rect 10907 3782 10953 3834
rect 10977 3782 11023 3834
rect 11023 3782 11033 3834
rect 11057 3782 11087 3834
rect 11087 3782 11113 3834
rect 10817 3780 10873 3782
rect 10897 3780 10953 3782
rect 10977 3780 11033 3782
rect 11057 3780 11113 3782
rect 10598 3304 10654 3360
rect 10322 2624 10378 2680
rect 10414 2216 10470 2272
rect 10598 2760 10654 2816
rect 10874 3032 10930 3088
rect 10817 2746 10873 2748
rect 10897 2746 10953 2748
rect 10977 2746 11033 2748
rect 11057 2746 11113 2748
rect 10817 2694 10843 2746
rect 10843 2694 10873 2746
rect 10897 2694 10907 2746
rect 10907 2694 10953 2746
rect 10977 2694 11023 2746
rect 11023 2694 11033 2746
rect 11057 2694 11087 2746
rect 11087 2694 11113 2746
rect 10817 2692 10873 2694
rect 10897 2692 10953 2694
rect 10977 2692 11033 2694
rect 11057 2692 11113 2694
rect 11242 2624 11298 2680
rect 11426 3712 11482 3768
rect 11886 6976 11942 7032
rect 11886 6860 11942 6896
rect 11886 6840 11888 6860
rect 11888 6840 11940 6860
rect 11940 6840 11942 6860
rect 12806 12552 12862 12608
rect 12990 14592 13046 14648
rect 12990 14456 13046 14512
rect 12990 14184 13046 14240
rect 13282 16346 13338 16348
rect 13362 16346 13418 16348
rect 13442 16346 13498 16348
rect 13522 16346 13578 16348
rect 13282 16294 13308 16346
rect 13308 16294 13338 16346
rect 13362 16294 13372 16346
rect 13372 16294 13418 16346
rect 13442 16294 13488 16346
rect 13488 16294 13498 16346
rect 13522 16294 13552 16346
rect 13552 16294 13578 16346
rect 13282 16292 13338 16294
rect 13362 16292 13418 16294
rect 13442 16292 13498 16294
rect 13522 16292 13578 16294
rect 13282 15258 13338 15260
rect 13362 15258 13418 15260
rect 13442 15258 13498 15260
rect 13522 15258 13578 15260
rect 13282 15206 13308 15258
rect 13308 15206 13338 15258
rect 13362 15206 13372 15258
rect 13372 15206 13418 15258
rect 13442 15206 13488 15258
rect 13488 15206 13498 15258
rect 13522 15206 13552 15258
rect 13552 15206 13578 15258
rect 13282 15204 13338 15206
rect 13362 15204 13418 15206
rect 13442 15204 13498 15206
rect 13522 15204 13578 15206
rect 13818 15036 13820 15056
rect 13820 15036 13872 15056
rect 13872 15036 13874 15056
rect 13818 15000 13874 15036
rect 13818 14864 13874 14920
rect 13634 14320 13690 14376
rect 13082 12824 13138 12880
rect 12714 12008 12770 12064
rect 11978 6568 12034 6624
rect 12438 9288 12494 9344
rect 12714 11464 12770 11520
rect 12346 8200 12402 8256
rect 12254 7928 12310 7984
rect 12254 7404 12310 7440
rect 12254 7384 12256 7404
rect 12256 7384 12308 7404
rect 12308 7384 12310 7404
rect 12254 6840 12310 6896
rect 11794 4392 11850 4448
rect 11886 4004 11942 4040
rect 11886 3984 11888 4004
rect 11888 3984 11940 4004
rect 11940 3984 11942 4004
rect 11518 3304 11574 3360
rect 12070 5616 12126 5672
rect 12346 6060 12348 6080
rect 12348 6060 12400 6080
rect 12400 6060 12402 6080
rect 12346 6024 12402 6060
rect 12346 5616 12402 5672
rect 12530 8744 12586 8800
rect 12530 7928 12586 7984
rect 12622 7248 12678 7304
rect 12530 7112 12586 7168
rect 12622 6976 12678 7032
rect 12530 6740 12532 6760
rect 12532 6740 12584 6760
rect 12584 6740 12586 6760
rect 12530 6704 12586 6740
rect 12162 3712 12218 3768
rect 11702 3032 11758 3088
rect 11518 2760 11574 2816
rect 11702 2488 11758 2544
rect 11886 3340 11888 3360
rect 11888 3340 11940 3360
rect 11940 3340 11942 3360
rect 11886 3304 11942 3340
rect 12898 12008 12954 12064
rect 13282 14170 13338 14172
rect 13362 14170 13418 14172
rect 13442 14170 13498 14172
rect 13522 14170 13578 14172
rect 13282 14118 13308 14170
rect 13308 14118 13338 14170
rect 13362 14118 13372 14170
rect 13372 14118 13418 14170
rect 13442 14118 13488 14170
rect 13488 14118 13498 14170
rect 13522 14118 13552 14170
rect 13552 14118 13578 14170
rect 13282 14116 13338 14118
rect 13362 14116 13418 14118
rect 13442 14116 13498 14118
rect 13522 14116 13578 14118
rect 13266 13504 13322 13560
rect 13634 13932 13690 13968
rect 13634 13912 13636 13932
rect 13636 13912 13688 13932
rect 13688 13912 13690 13932
rect 13450 13368 13506 13424
rect 13282 13082 13338 13084
rect 13362 13082 13418 13084
rect 13442 13082 13498 13084
rect 13522 13082 13578 13084
rect 13282 13030 13308 13082
rect 13308 13030 13338 13082
rect 13362 13030 13372 13082
rect 13372 13030 13418 13082
rect 13442 13030 13488 13082
rect 13488 13030 13498 13082
rect 13522 13030 13552 13082
rect 13552 13030 13578 13082
rect 13282 13028 13338 13030
rect 13362 13028 13418 13030
rect 13442 13028 13498 13030
rect 13522 13028 13578 13030
rect 13910 13776 13966 13832
rect 13818 13640 13874 13696
rect 13726 12960 13782 13016
rect 14094 14456 14150 14512
rect 14002 13404 14004 13424
rect 14004 13404 14056 13424
rect 14056 13404 14058 13424
rect 14002 13368 14058 13404
rect 13726 12300 13782 12336
rect 13726 12280 13728 12300
rect 13728 12280 13780 12300
rect 13780 12280 13782 12300
rect 13282 11994 13338 11996
rect 13362 11994 13418 11996
rect 13442 11994 13498 11996
rect 13522 11994 13578 11996
rect 13282 11942 13308 11994
rect 13308 11942 13338 11994
rect 13362 11942 13372 11994
rect 13372 11942 13418 11994
rect 13442 11942 13488 11994
rect 13488 11942 13498 11994
rect 13522 11942 13552 11994
rect 13552 11942 13578 11994
rect 13282 11940 13338 11942
rect 13362 11940 13418 11942
rect 13442 11940 13498 11942
rect 13522 11940 13578 11942
rect 12898 10920 12954 10976
rect 13634 11600 13690 11656
rect 12898 10412 12900 10432
rect 12900 10412 12952 10432
rect 12952 10412 12954 10432
rect 12898 10376 12954 10412
rect 12898 10104 12954 10160
rect 13082 10512 13138 10568
rect 12898 6160 12954 6216
rect 12714 5616 12770 5672
rect 12622 5344 12678 5400
rect 12530 4528 12586 4584
rect 12714 4564 12716 4584
rect 12716 4564 12768 4584
rect 12768 4564 12770 4584
rect 12714 4528 12770 4564
rect 12714 4428 12716 4448
rect 12716 4428 12768 4448
rect 12768 4428 12770 4448
rect 12714 4392 12770 4428
rect 12714 4120 12770 4176
rect 12622 3576 12678 3632
rect 12530 3032 12586 3088
rect 12438 2352 12494 2408
rect 11886 1944 11942 2000
rect 13082 7656 13138 7712
rect 14002 13232 14058 13288
rect 14186 12416 14242 12472
rect 13910 11736 13966 11792
rect 14554 17856 14610 17912
rect 14462 15952 14518 16008
rect 14278 12144 14334 12200
rect 13282 10906 13338 10908
rect 13362 10906 13418 10908
rect 13442 10906 13498 10908
rect 13522 10906 13578 10908
rect 13282 10854 13308 10906
rect 13308 10854 13338 10906
rect 13362 10854 13372 10906
rect 13372 10854 13418 10906
rect 13442 10854 13488 10906
rect 13488 10854 13498 10906
rect 13522 10854 13552 10906
rect 13552 10854 13578 10906
rect 13282 10852 13338 10854
rect 13362 10852 13418 10854
rect 13442 10852 13498 10854
rect 13522 10852 13578 10854
rect 13266 10532 13322 10568
rect 13266 10512 13268 10532
rect 13268 10512 13320 10532
rect 13320 10512 13322 10532
rect 13282 9818 13338 9820
rect 13362 9818 13418 9820
rect 13442 9818 13498 9820
rect 13522 9818 13578 9820
rect 13282 9766 13308 9818
rect 13308 9766 13338 9818
rect 13362 9766 13372 9818
rect 13372 9766 13418 9818
rect 13442 9766 13488 9818
rect 13488 9766 13498 9818
rect 13522 9766 13552 9818
rect 13552 9766 13578 9818
rect 13282 9764 13338 9766
rect 13362 9764 13418 9766
rect 13442 9764 13498 9766
rect 13522 9764 13578 9766
rect 13450 9460 13452 9480
rect 13452 9460 13504 9480
rect 13504 9460 13506 9480
rect 13450 9424 13506 9460
rect 13818 9560 13874 9616
rect 13634 9152 13690 9208
rect 13282 8730 13338 8732
rect 13362 8730 13418 8732
rect 13442 8730 13498 8732
rect 13522 8730 13578 8732
rect 13282 8678 13308 8730
rect 13308 8678 13338 8730
rect 13362 8678 13372 8730
rect 13372 8678 13418 8730
rect 13442 8678 13488 8730
rect 13488 8678 13498 8730
rect 13522 8678 13552 8730
rect 13552 8678 13578 8730
rect 13282 8676 13338 8678
rect 13362 8676 13418 8678
rect 13442 8676 13498 8678
rect 13522 8676 13578 8678
rect 13282 7642 13338 7644
rect 13362 7642 13418 7644
rect 13442 7642 13498 7644
rect 13522 7642 13578 7644
rect 13282 7590 13308 7642
rect 13308 7590 13338 7642
rect 13362 7590 13372 7642
rect 13372 7590 13418 7642
rect 13442 7590 13488 7642
rect 13488 7590 13498 7642
rect 13522 7590 13552 7642
rect 13552 7590 13578 7642
rect 13282 7588 13338 7590
rect 13362 7588 13418 7590
rect 13442 7588 13498 7590
rect 13522 7588 13578 7590
rect 13726 7384 13782 7440
rect 13726 6860 13782 6896
rect 13726 6840 13728 6860
rect 13728 6840 13780 6860
rect 13780 6840 13782 6860
rect 12990 5888 13046 5944
rect 13282 6554 13338 6556
rect 13362 6554 13418 6556
rect 13442 6554 13498 6556
rect 13522 6554 13578 6556
rect 13282 6502 13308 6554
rect 13308 6502 13338 6554
rect 13362 6502 13372 6554
rect 13372 6502 13418 6554
rect 13442 6502 13488 6554
rect 13488 6502 13498 6554
rect 13522 6502 13552 6554
rect 13552 6502 13578 6554
rect 13282 6500 13338 6502
rect 13362 6500 13418 6502
rect 13442 6500 13498 6502
rect 13522 6500 13578 6502
rect 14186 11464 14242 11520
rect 14278 11212 14334 11248
rect 14278 11192 14280 11212
rect 14280 11192 14332 11212
rect 14332 11192 14334 11212
rect 14002 9596 14004 9616
rect 14004 9596 14056 9616
rect 14056 9596 14058 9616
rect 14002 9560 14058 9596
rect 14186 9988 14242 10024
rect 14186 9968 14188 9988
rect 14188 9968 14240 9988
rect 14240 9968 14242 9988
rect 13910 7248 13966 7304
rect 13174 5752 13230 5808
rect 13450 6024 13506 6080
rect 13542 5888 13598 5944
rect 13634 5616 13690 5672
rect 13082 5480 13138 5536
rect 13282 5466 13338 5468
rect 13362 5466 13418 5468
rect 13442 5466 13498 5468
rect 13522 5466 13578 5468
rect 13282 5414 13308 5466
rect 13308 5414 13338 5466
rect 13362 5414 13372 5466
rect 13372 5414 13418 5466
rect 13442 5414 13488 5466
rect 13488 5414 13498 5466
rect 13522 5414 13552 5466
rect 13552 5414 13578 5466
rect 13282 5412 13338 5414
rect 13362 5412 13418 5414
rect 13442 5412 13498 5414
rect 13522 5412 13578 5414
rect 13266 4936 13322 4992
rect 13450 4800 13506 4856
rect 13282 4378 13338 4380
rect 13362 4378 13418 4380
rect 13442 4378 13498 4380
rect 13522 4378 13578 4380
rect 13282 4326 13308 4378
rect 13308 4326 13338 4378
rect 13362 4326 13372 4378
rect 13372 4326 13418 4378
rect 13442 4326 13488 4378
rect 13488 4326 13498 4378
rect 13522 4326 13552 4378
rect 13552 4326 13578 4378
rect 13282 4324 13338 4326
rect 13362 4324 13418 4326
rect 13442 4324 13498 4326
rect 13522 4324 13578 4326
rect 13726 5072 13782 5128
rect 13634 4120 13690 4176
rect 13266 3596 13322 3632
rect 13266 3576 13268 3596
rect 13268 3576 13320 3596
rect 13320 3576 13322 3596
rect 12990 2352 13046 2408
rect 12898 1944 12954 2000
rect 12622 1400 12678 1456
rect 13282 3290 13338 3292
rect 13362 3290 13418 3292
rect 13442 3290 13498 3292
rect 13522 3290 13578 3292
rect 13282 3238 13308 3290
rect 13308 3238 13338 3290
rect 13362 3238 13372 3290
rect 13372 3238 13418 3290
rect 13442 3238 13488 3290
rect 13488 3238 13498 3290
rect 13522 3238 13552 3290
rect 13552 3238 13578 3290
rect 13282 3236 13338 3238
rect 13362 3236 13418 3238
rect 13442 3236 13498 3238
rect 13522 3236 13578 3238
rect 14186 7248 14242 7304
rect 14002 6704 14058 6760
rect 13818 3440 13874 3496
rect 13726 2488 13782 2544
rect 13282 2202 13338 2204
rect 13362 2202 13418 2204
rect 13442 2202 13498 2204
rect 13522 2202 13578 2204
rect 13282 2150 13308 2202
rect 13308 2150 13338 2202
rect 13362 2150 13372 2202
rect 13372 2150 13418 2202
rect 13442 2150 13488 2202
rect 13488 2150 13498 2202
rect 13522 2150 13552 2202
rect 13552 2150 13578 2202
rect 13282 2148 13338 2150
rect 13362 2148 13418 2150
rect 13442 2148 13498 2150
rect 13522 2148 13578 2150
rect 13450 1264 13506 1320
rect 14646 14728 14702 14784
rect 14554 11056 14610 11112
rect 14462 9016 14518 9072
rect 14738 5888 14794 5944
rect 14462 3984 14518 4040
rect 14646 5208 14702 5264
rect 14646 3848 14702 3904
rect 15014 8472 15070 8528
rect 15198 10512 15254 10568
rect 15014 8336 15070 8392
rect 15014 6296 15070 6352
rect 15106 4664 15162 4720
rect 15014 4528 15070 4584
rect 15014 3032 15070 3088
rect 14738 2896 14794 2952
rect 14554 1536 14610 1592
rect 14830 2760 14886 2816
rect 15934 17584 15990 17640
rect 15474 9832 15530 9888
rect 15566 2624 15622 2680
<< metal3 >>
rect 0 19546 480 19576
rect 2865 19546 2931 19549
rect 0 19544 2931 19546
rect 0 19488 2870 19544
rect 2926 19488 2931 19544
rect 0 19486 2931 19488
rect 0 19456 480 19486
rect 2865 19483 2931 19486
rect 0 18594 480 18624
rect 3509 18594 3575 18597
rect 0 18592 3575 18594
rect 0 18536 3514 18592
rect 3570 18536 3575 18592
rect 0 18534 3575 18536
rect 0 18504 480 18534
rect 3509 18531 3575 18534
rect 8937 17914 9003 17917
rect 11789 17914 11855 17917
rect 8937 17912 11855 17914
rect 8937 17856 8942 17912
rect 8998 17856 11794 17912
rect 11850 17856 11855 17912
rect 8937 17854 11855 17856
rect 8937 17851 9003 17854
rect 11789 17851 11855 17854
rect 14549 17914 14615 17917
rect 16520 17914 17000 17944
rect 14549 17912 17000 17914
rect 14549 17856 14554 17912
rect 14610 17856 17000 17912
rect 14549 17854 17000 17856
rect 14549 17851 14615 17854
rect 16520 17824 17000 17854
rect 0 17642 480 17672
rect 2773 17642 2839 17645
rect 0 17640 2839 17642
rect 0 17584 2778 17640
rect 2834 17584 2839 17640
rect 0 17582 2839 17584
rect 0 17552 480 17582
rect 2773 17579 2839 17582
rect 8201 17642 8267 17645
rect 15929 17642 15995 17645
rect 8201 17640 15995 17642
rect 8201 17584 8206 17640
rect 8262 17584 15934 17640
rect 15990 17584 15995 17640
rect 8201 17582 15995 17584
rect 8201 17579 8267 17582
rect 15929 17579 15995 17582
rect 3409 17440 3729 17441
rect 3409 17376 3417 17440
rect 3481 17376 3497 17440
rect 3561 17376 3577 17440
rect 3641 17376 3657 17440
rect 3721 17376 3729 17440
rect 3409 17375 3729 17376
rect 8340 17440 8660 17441
rect 8340 17376 8348 17440
rect 8412 17376 8428 17440
rect 8492 17376 8508 17440
rect 8572 17376 8588 17440
rect 8652 17376 8660 17440
rect 8340 17375 8660 17376
rect 13270 17440 13590 17441
rect 13270 17376 13278 17440
rect 13342 17376 13358 17440
rect 13422 17376 13438 17440
rect 13502 17376 13518 17440
rect 13582 17376 13590 17440
rect 13270 17375 13590 17376
rect 9397 17370 9463 17373
rect 12341 17370 12407 17373
rect 8894 17368 12407 17370
rect 8894 17312 9402 17368
rect 9458 17312 12346 17368
rect 12402 17312 12407 17368
rect 8894 17310 12407 17312
rect 7281 17234 7347 17237
rect 8894 17234 8954 17310
rect 9397 17307 9463 17310
rect 12341 17307 12407 17310
rect 7281 17232 8954 17234
rect 7281 17176 7286 17232
rect 7342 17176 8954 17232
rect 7281 17174 8954 17176
rect 10409 17234 10475 17237
rect 13169 17234 13235 17237
rect 10409 17232 13235 17234
rect 10409 17176 10414 17232
rect 10470 17176 13174 17232
rect 13230 17176 13235 17232
rect 10409 17174 13235 17176
rect 7281 17171 7347 17174
rect 10409 17171 10475 17174
rect 13169 17171 13235 17174
rect 8477 17098 8543 17101
rect 12750 17098 12756 17100
rect 8477 17096 12756 17098
rect 8477 17040 8482 17096
rect 8538 17040 12756 17096
rect 8477 17038 12756 17040
rect 8477 17035 8543 17038
rect 12750 17036 12756 17038
rect 12820 17036 12826 17100
rect 6729 16962 6795 16965
rect 9489 16962 9555 16965
rect 6729 16960 9555 16962
rect 6729 16904 6734 16960
rect 6790 16904 9494 16960
rect 9550 16904 9555 16960
rect 6729 16902 9555 16904
rect 6729 16899 6795 16902
rect 9489 16899 9555 16902
rect 11789 16962 11855 16965
rect 12198 16962 12204 16964
rect 11789 16960 12204 16962
rect 11789 16904 11794 16960
rect 11850 16904 12204 16960
rect 11789 16902 12204 16904
rect 11789 16899 11855 16902
rect 12198 16900 12204 16902
rect 12268 16900 12274 16964
rect 5874 16896 6194 16897
rect 5874 16832 5882 16896
rect 5946 16832 5962 16896
rect 6026 16832 6042 16896
rect 6106 16832 6122 16896
rect 6186 16832 6194 16896
rect 5874 16831 6194 16832
rect 10805 16896 11125 16897
rect 10805 16832 10813 16896
rect 10877 16832 10893 16896
rect 10957 16832 10973 16896
rect 11037 16832 11053 16896
rect 11117 16832 11125 16896
rect 10805 16831 11125 16832
rect 4889 16826 4955 16829
rect 5022 16826 5028 16828
rect 4889 16824 5028 16826
rect 4889 16768 4894 16824
rect 4950 16768 5028 16824
rect 4889 16766 5028 16768
rect 4889 16763 4955 16766
rect 5022 16764 5028 16766
rect 5092 16764 5098 16828
rect 8109 16826 8175 16829
rect 9305 16826 9371 16829
rect 8109 16824 9371 16826
rect 8109 16768 8114 16824
rect 8170 16768 9310 16824
rect 9366 16768 9371 16824
rect 8109 16766 9371 16768
rect 8109 16763 8175 16766
rect 9305 16763 9371 16766
rect 0 16690 480 16720
rect 2129 16690 2195 16693
rect 0 16688 2195 16690
rect 0 16632 2134 16688
rect 2190 16632 2195 16688
rect 0 16630 2195 16632
rect 0 16600 480 16630
rect 2129 16627 2195 16630
rect 3785 16690 3851 16693
rect 8569 16690 8635 16693
rect 9254 16690 9260 16692
rect 3785 16688 9260 16690
rect 3785 16632 3790 16688
rect 3846 16632 8574 16688
rect 8630 16632 9260 16688
rect 3785 16630 9260 16632
rect 3785 16627 3851 16630
rect 8569 16627 8635 16630
rect 9254 16628 9260 16630
rect 9324 16628 9330 16692
rect 9765 16690 9831 16693
rect 13118 16690 13124 16692
rect 9765 16688 13124 16690
rect 9765 16632 9770 16688
rect 9826 16632 13124 16688
rect 9765 16630 13124 16632
rect 9765 16627 9831 16630
rect 13118 16628 13124 16630
rect 13188 16628 13194 16692
rect 3141 16554 3207 16557
rect 11329 16554 11395 16557
rect 3141 16552 11395 16554
rect 3141 16496 3146 16552
rect 3202 16496 11334 16552
rect 11390 16496 11395 16552
rect 3141 16494 11395 16496
rect 3141 16491 3207 16494
rect 11329 16491 11395 16494
rect 12750 16492 12756 16556
rect 12820 16554 12826 16556
rect 13077 16554 13143 16557
rect 12820 16552 13143 16554
rect 12820 16496 13082 16552
rect 13138 16496 13143 16552
rect 12820 16494 13143 16496
rect 12820 16492 12826 16494
rect 13077 16491 13143 16494
rect 4337 16420 4403 16421
rect 4286 16418 4292 16420
rect 4246 16358 4292 16418
rect 4356 16416 4403 16420
rect 4398 16360 4403 16416
rect 4286 16356 4292 16358
rect 4356 16356 4403 16360
rect 4337 16355 4403 16356
rect 4889 16418 4955 16421
rect 7782 16418 7788 16420
rect 4889 16416 7788 16418
rect 4889 16360 4894 16416
rect 4950 16360 7788 16416
rect 4889 16358 7788 16360
rect 4889 16355 4955 16358
rect 7782 16356 7788 16358
rect 7852 16418 7858 16420
rect 7925 16418 7991 16421
rect 7852 16416 7991 16418
rect 7852 16360 7930 16416
rect 7986 16360 7991 16416
rect 7852 16358 7991 16360
rect 7852 16356 7858 16358
rect 7925 16355 7991 16358
rect 9489 16418 9555 16421
rect 11462 16418 11468 16420
rect 9489 16416 11468 16418
rect 9489 16360 9494 16416
rect 9550 16360 11468 16416
rect 9489 16358 11468 16360
rect 9489 16355 9555 16358
rect 11462 16356 11468 16358
rect 11532 16356 11538 16420
rect 3409 16352 3729 16353
rect 3409 16288 3417 16352
rect 3481 16288 3497 16352
rect 3561 16288 3577 16352
rect 3641 16288 3657 16352
rect 3721 16288 3729 16352
rect 3409 16287 3729 16288
rect 8340 16352 8660 16353
rect 8340 16288 8348 16352
rect 8412 16288 8428 16352
rect 8492 16288 8508 16352
rect 8572 16288 8588 16352
rect 8652 16288 8660 16352
rect 8340 16287 8660 16288
rect 13270 16352 13590 16353
rect 13270 16288 13278 16352
rect 13342 16288 13358 16352
rect 13422 16288 13438 16352
rect 13502 16288 13518 16352
rect 13582 16288 13590 16352
rect 13270 16287 13590 16288
rect 7598 16282 7604 16284
rect 3926 16222 7604 16282
rect 2313 16146 2379 16149
rect 3926 16146 3986 16222
rect 7598 16220 7604 16222
rect 7668 16220 7674 16284
rect 9673 16282 9739 16285
rect 10869 16282 10935 16285
rect 9673 16280 10935 16282
rect 9673 16224 9678 16280
rect 9734 16224 10874 16280
rect 10930 16224 10935 16280
rect 9673 16222 10935 16224
rect 9673 16219 9739 16222
rect 10869 16219 10935 16222
rect 2313 16144 3986 16146
rect 2313 16088 2318 16144
rect 2374 16088 3986 16144
rect 2313 16086 3986 16088
rect 4061 16146 4127 16149
rect 12065 16146 12131 16149
rect 4061 16144 12131 16146
rect 4061 16088 4066 16144
rect 4122 16088 12070 16144
rect 12126 16088 12131 16144
rect 4061 16086 12131 16088
rect 2313 16083 2379 16086
rect 4061 16083 4127 16086
rect 12065 16083 12131 16086
rect 3233 16010 3299 16013
rect 4889 16010 4955 16013
rect 3233 16008 4955 16010
rect 3233 15952 3238 16008
rect 3294 15952 4894 16008
rect 4950 15952 4955 16008
rect 3233 15950 4955 15952
rect 3233 15947 3299 15950
rect 4889 15947 4955 15950
rect 5809 16010 5875 16013
rect 14457 16010 14523 16013
rect 5809 16008 14523 16010
rect 5809 15952 5814 16008
rect 5870 15952 14462 16008
rect 14518 15952 14523 16008
rect 5809 15950 14523 15952
rect 5809 15947 5875 15950
rect 14457 15947 14523 15950
rect 2998 15812 3004 15876
rect 3068 15874 3074 15876
rect 3509 15874 3575 15877
rect 3068 15872 3575 15874
rect 3068 15816 3514 15872
rect 3570 15816 3575 15872
rect 3068 15814 3575 15816
rect 3068 15812 3074 15814
rect 3509 15811 3575 15814
rect 4705 15874 4771 15877
rect 4981 15874 5047 15877
rect 4705 15872 5047 15874
rect 4705 15816 4710 15872
rect 4766 15816 4986 15872
rect 5042 15816 5047 15872
rect 4705 15814 5047 15816
rect 4705 15811 4771 15814
rect 4981 15811 5047 15814
rect 6269 15874 6335 15877
rect 7741 15874 7807 15877
rect 6269 15872 7807 15874
rect 6269 15816 6274 15872
rect 6330 15816 7746 15872
rect 7802 15816 7807 15872
rect 6269 15814 7807 15816
rect 6269 15811 6335 15814
rect 7741 15811 7807 15814
rect 9397 15876 9463 15877
rect 9397 15872 9444 15876
rect 9508 15874 9514 15876
rect 10041 15874 10107 15877
rect 10174 15874 10180 15876
rect 9397 15816 9402 15872
rect 9397 15812 9444 15816
rect 9508 15814 9554 15874
rect 10041 15872 10180 15874
rect 10041 15816 10046 15872
rect 10102 15816 10180 15872
rect 10041 15814 10180 15816
rect 9508 15812 9514 15814
rect 9397 15811 9463 15812
rect 10041 15811 10107 15814
rect 10174 15812 10180 15814
rect 10244 15812 10250 15876
rect 5874 15808 6194 15809
rect 0 15738 480 15768
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6194 15808
rect 5874 15743 6194 15744
rect 10805 15808 11125 15809
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10805 15743 11125 15744
rect 1853 15738 1919 15741
rect 0 15736 1919 15738
rect 0 15680 1858 15736
rect 1914 15680 1919 15736
rect 0 15678 1919 15680
rect 0 15648 480 15678
rect 1853 15675 1919 15678
rect 4705 15738 4771 15741
rect 5390 15738 5396 15740
rect 4705 15736 5396 15738
rect 4705 15680 4710 15736
rect 4766 15680 5396 15736
rect 4705 15678 5396 15680
rect 4705 15675 4771 15678
rect 5390 15676 5396 15678
rect 5460 15676 5466 15740
rect 6821 15738 6887 15741
rect 9673 15738 9739 15741
rect 6821 15736 9739 15738
rect 6821 15680 6826 15736
rect 6882 15680 9678 15736
rect 9734 15680 9739 15736
rect 6821 15678 9739 15680
rect 6821 15675 6887 15678
rect 9673 15675 9739 15678
rect 11513 15738 11579 15741
rect 12566 15738 12572 15740
rect 11513 15736 12572 15738
rect 11513 15680 11518 15736
rect 11574 15680 12572 15736
rect 11513 15678 12572 15680
rect 11513 15675 11579 15678
rect 12566 15676 12572 15678
rect 12636 15676 12642 15740
rect 2773 15602 2839 15605
rect 12382 15602 12388 15604
rect 2773 15600 12388 15602
rect 2773 15544 2778 15600
rect 2834 15544 12388 15600
rect 2773 15542 12388 15544
rect 2773 15539 2839 15542
rect 12382 15540 12388 15542
rect 12452 15540 12458 15604
rect 12525 15602 12591 15605
rect 12801 15602 12867 15605
rect 12525 15600 12867 15602
rect 12525 15544 12530 15600
rect 12586 15544 12806 15600
rect 12862 15544 12867 15600
rect 12525 15542 12867 15544
rect 12525 15539 12591 15542
rect 12801 15539 12867 15542
rect 3141 15466 3207 15469
rect 3417 15466 3483 15469
rect 5533 15466 5599 15469
rect 6637 15466 6703 15469
rect 3141 15464 3250 15466
rect 3141 15408 3146 15464
rect 3202 15408 3250 15464
rect 3141 15403 3250 15408
rect 3417 15464 4676 15466
rect 3417 15408 3422 15464
rect 3478 15408 4676 15464
rect 3417 15406 4676 15408
rect 3417 15403 3483 15406
rect 3190 15196 3250 15403
rect 4337 15330 4403 15333
rect 4470 15330 4476 15332
rect 4337 15328 4476 15330
rect 4337 15272 4342 15328
rect 4398 15272 4476 15328
rect 4337 15270 4476 15272
rect 4337 15267 4403 15270
rect 4470 15268 4476 15270
rect 4540 15268 4546 15332
rect 4616 15330 4676 15406
rect 5533 15464 6703 15466
rect 5533 15408 5538 15464
rect 5594 15408 6642 15464
rect 6698 15408 6703 15464
rect 5533 15406 6703 15408
rect 5533 15403 5599 15406
rect 6637 15403 6703 15406
rect 6862 15404 6868 15468
rect 6932 15466 6938 15468
rect 8886 15466 8892 15468
rect 6932 15406 8892 15466
rect 6932 15404 6938 15406
rect 8886 15404 8892 15406
rect 8956 15404 8962 15468
rect 9254 15404 9260 15468
rect 9324 15466 9330 15468
rect 9489 15466 9555 15469
rect 9806 15466 9812 15468
rect 9324 15464 9812 15466
rect 9324 15408 9494 15464
rect 9550 15408 9812 15464
rect 9324 15406 9812 15408
rect 9324 15404 9330 15406
rect 6870 15330 6930 15404
rect 4616 15270 6930 15330
rect 8894 15330 8954 15404
rect 9489 15403 9555 15406
rect 9806 15404 9812 15406
rect 9876 15404 9882 15468
rect 9990 15404 9996 15468
rect 10060 15466 10066 15468
rect 10133 15466 10199 15469
rect 10060 15464 10199 15466
rect 10060 15408 10138 15464
rect 10194 15408 10199 15464
rect 10060 15406 10199 15408
rect 10060 15404 10066 15406
rect 10133 15403 10199 15406
rect 10358 15404 10364 15468
rect 10428 15466 10434 15468
rect 10869 15466 10935 15469
rect 10428 15464 10935 15466
rect 10428 15408 10874 15464
rect 10930 15408 10935 15464
rect 10428 15406 10935 15408
rect 10428 15404 10434 15406
rect 10869 15403 10935 15406
rect 10593 15330 10659 15333
rect 8894 15328 10659 15330
rect 8894 15272 10598 15328
rect 10654 15272 10659 15328
rect 8894 15270 10659 15272
rect 10593 15267 10659 15270
rect 11830 15268 11836 15332
rect 11900 15330 11906 15332
rect 11973 15330 12039 15333
rect 11900 15328 12039 15330
rect 11900 15272 11978 15328
rect 12034 15272 12039 15328
rect 11900 15270 12039 15272
rect 11900 15268 11906 15270
rect 11973 15267 12039 15270
rect 3409 15264 3729 15265
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 15199 3729 15200
rect 8340 15264 8660 15265
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 15199 8660 15200
rect 13270 15264 13590 15265
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13270 15199 13590 15200
rect 3182 15132 3188 15196
rect 3252 15132 3258 15196
rect 6913 15194 6979 15197
rect 3880 15192 6979 15194
rect 3880 15136 6918 15192
rect 6974 15136 6979 15192
rect 3880 15134 6979 15136
rect 2497 15058 2563 15061
rect 3880 15058 3940 15134
rect 6913 15131 6979 15134
rect 8937 15194 9003 15197
rect 9489 15194 9555 15197
rect 8937 15192 9555 15194
rect 8937 15136 8942 15192
rect 8998 15136 9494 15192
rect 9550 15136 9555 15192
rect 8937 15134 9555 15136
rect 8937 15131 9003 15134
rect 9489 15131 9555 15134
rect 9622 15132 9628 15196
rect 9692 15194 9698 15196
rect 10317 15194 10383 15197
rect 9692 15192 10383 15194
rect 9692 15136 10322 15192
rect 10378 15136 10383 15192
rect 9692 15134 10383 15136
rect 9692 15132 9698 15134
rect 10317 15131 10383 15134
rect 11053 15194 11119 15197
rect 11646 15194 11652 15196
rect 11053 15192 11652 15194
rect 11053 15136 11058 15192
rect 11114 15136 11652 15192
rect 11053 15134 11652 15136
rect 11053 15131 11119 15134
rect 11646 15132 11652 15134
rect 11716 15132 11722 15196
rect 2497 15056 3940 15058
rect 2497 15000 2502 15056
rect 2558 15000 3940 15056
rect 2497 14998 3940 15000
rect 4429 15058 4495 15061
rect 11789 15058 11855 15061
rect 4429 15056 11855 15058
rect 4429 15000 4434 15056
rect 4490 15000 11794 15056
rect 11850 15000 11855 15056
rect 4429 14998 11855 15000
rect 2497 14995 2563 14998
rect 4429 14995 4495 14998
rect 11789 14995 11855 14998
rect 12014 14996 12020 15060
rect 12084 15058 12090 15060
rect 13813 15058 13879 15061
rect 12084 15056 13879 15058
rect 12084 15000 13818 15056
rect 13874 15000 13879 15056
rect 12084 14998 13879 15000
rect 12084 14996 12090 14998
rect 13813 14995 13879 14998
rect 2589 14922 2655 14925
rect 13813 14922 13879 14925
rect 2589 14920 13879 14922
rect 2589 14864 2594 14920
rect 2650 14864 13818 14920
rect 13874 14864 13879 14920
rect 2589 14862 13879 14864
rect 2589 14859 2655 14862
rect 13813 14859 13879 14862
rect 0 14786 480 14816
rect 3049 14786 3115 14789
rect 0 14784 3115 14786
rect 0 14728 3054 14784
rect 3110 14728 3115 14784
rect 0 14726 3115 14728
rect 0 14696 480 14726
rect 3049 14723 3115 14726
rect 4613 14788 4679 14789
rect 4613 14784 4660 14788
rect 4724 14786 4730 14788
rect 6453 14786 6519 14789
rect 7005 14786 7071 14789
rect 7189 14788 7255 14789
rect 7189 14786 7236 14788
rect 4613 14728 4618 14784
rect 4613 14724 4660 14728
rect 4724 14726 4770 14786
rect 6453 14784 7071 14786
rect 6453 14728 6458 14784
rect 6514 14728 7010 14784
rect 7066 14728 7071 14784
rect 6453 14726 7071 14728
rect 7144 14784 7236 14786
rect 7144 14728 7194 14784
rect 7144 14726 7236 14728
rect 4724 14724 4730 14726
rect 4613 14723 4679 14724
rect 6453 14723 6519 14726
rect 7005 14723 7071 14726
rect 7189 14724 7236 14726
rect 7300 14724 7306 14788
rect 8477 14786 8543 14789
rect 9070 14786 9076 14788
rect 8477 14784 9076 14786
rect 8477 14728 8482 14784
rect 8538 14728 9076 14784
rect 8477 14726 9076 14728
rect 7189 14723 7255 14724
rect 8477 14723 8543 14726
rect 9070 14724 9076 14726
rect 9140 14724 9146 14788
rect 9305 14786 9371 14789
rect 10409 14786 10475 14789
rect 9305 14784 10475 14786
rect 9305 14728 9310 14784
rect 9366 14728 10414 14784
rect 10470 14728 10475 14784
rect 9305 14726 10475 14728
rect 9305 14723 9371 14726
rect 10409 14723 10475 14726
rect 11973 14786 12039 14789
rect 14641 14786 14707 14789
rect 11973 14784 14707 14786
rect 11973 14728 11978 14784
rect 12034 14728 14646 14784
rect 14702 14728 14707 14784
rect 11973 14726 14707 14728
rect 11973 14723 12039 14726
rect 14641 14723 14707 14726
rect 5874 14720 6194 14721
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6194 14720
rect 5874 14655 6194 14656
rect 10805 14720 11125 14721
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10805 14655 11125 14656
rect 4245 14650 4311 14653
rect 7189 14650 7255 14653
rect 9121 14650 9187 14653
rect 4245 14648 5642 14650
rect 4245 14592 4250 14648
rect 4306 14592 5642 14648
rect 4245 14590 5642 14592
rect 4245 14587 4311 14590
rect 4429 14514 4495 14517
rect 5257 14514 5323 14517
rect 4429 14512 5323 14514
rect 4429 14456 4434 14512
rect 4490 14456 5262 14512
rect 5318 14456 5323 14512
rect 4429 14454 5323 14456
rect 5582 14514 5642 14590
rect 7189 14648 9187 14650
rect 7189 14592 7194 14648
rect 7250 14592 9126 14648
rect 9182 14592 9187 14648
rect 7189 14590 9187 14592
rect 7189 14587 7255 14590
rect 9121 14587 9187 14590
rect 9673 14650 9739 14653
rect 9857 14650 9923 14653
rect 10501 14652 10567 14653
rect 10501 14650 10548 14652
rect 9673 14648 9923 14650
rect 9673 14592 9678 14648
rect 9734 14592 9862 14648
rect 9918 14592 9923 14648
rect 9673 14590 9923 14592
rect 10456 14648 10548 14650
rect 10456 14592 10506 14648
rect 10456 14590 10548 14592
rect 9673 14587 9739 14590
rect 9857 14587 9923 14590
rect 10501 14588 10548 14590
rect 10612 14588 10618 14652
rect 11421 14650 11487 14653
rect 12985 14650 13051 14653
rect 11421 14648 13051 14650
rect 11421 14592 11426 14648
rect 11482 14592 12990 14648
rect 13046 14592 13051 14648
rect 11421 14590 13051 14592
rect 10501 14587 10567 14588
rect 11421 14587 11487 14590
rect 12985 14587 13051 14590
rect 12985 14516 13051 14517
rect 12014 14514 12020 14516
rect 5582 14454 12020 14514
rect 4429 14451 4495 14454
rect 5257 14451 5323 14454
rect 12014 14452 12020 14454
rect 12084 14452 12090 14516
rect 12934 14514 12940 14516
rect 12894 14454 12940 14514
rect 13004 14512 13051 14516
rect 14089 14514 14155 14517
rect 13046 14456 13051 14512
rect 12934 14452 12940 14454
rect 13004 14452 13051 14456
rect 12985 14451 13051 14452
rect 13310 14512 14155 14514
rect 13310 14456 14094 14512
rect 14150 14456 14155 14512
rect 13310 14454 14155 14456
rect 2957 14380 3023 14381
rect 2957 14376 3004 14380
rect 3068 14378 3074 14380
rect 3785 14378 3851 14381
rect 8661 14378 8727 14381
rect 2957 14320 2962 14376
rect 2957 14316 3004 14320
rect 3068 14318 3114 14378
rect 3785 14376 8727 14378
rect 3785 14320 3790 14376
rect 3846 14320 8666 14376
rect 8722 14320 8727 14376
rect 3785 14318 8727 14320
rect 3068 14316 3074 14318
rect 2957 14315 3023 14316
rect 3785 14315 3851 14318
rect 8661 14315 8727 14318
rect 9121 14378 9187 14381
rect 13310 14378 13370 14454
rect 14089 14451 14155 14454
rect 13629 14380 13695 14381
rect 13629 14378 13676 14380
rect 9121 14376 13370 14378
rect 9121 14320 9126 14376
rect 9182 14320 13370 14376
rect 9121 14318 13370 14320
rect 13584 14376 13676 14378
rect 13584 14320 13634 14376
rect 13584 14318 13676 14320
rect 9121 14315 9187 14318
rect 13629 14316 13676 14318
rect 13740 14316 13746 14380
rect 13629 14315 13695 14316
rect 3877 14242 3943 14245
rect 5901 14242 5967 14245
rect 3877 14240 5967 14242
rect 3877 14184 3882 14240
rect 3938 14184 5906 14240
rect 5962 14184 5967 14240
rect 3877 14182 5967 14184
rect 3877 14179 3943 14182
rect 5901 14179 5967 14182
rect 8937 14242 9003 14245
rect 12985 14242 13051 14245
rect 8937 14240 13051 14242
rect 8937 14184 8942 14240
rect 8998 14184 12990 14240
rect 13046 14184 13051 14240
rect 8937 14182 13051 14184
rect 8937 14179 9003 14182
rect 12985 14179 13051 14182
rect 3409 14176 3729 14177
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 14111 3729 14112
rect 8340 14176 8660 14177
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 14111 8660 14112
rect 13270 14176 13590 14177
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 14111 13590 14112
rect 7189 14106 7255 14109
rect 3926 14104 7255 14106
rect 3926 14048 7194 14104
rect 7250 14048 7255 14104
rect 3926 14046 7255 14048
rect 3182 13908 3188 13972
rect 3252 13970 3258 13972
rect 3926 13970 3986 14046
rect 7189 14043 7255 14046
rect 9121 14106 9187 14109
rect 9254 14106 9260 14108
rect 9121 14104 9260 14106
rect 9121 14048 9126 14104
rect 9182 14048 9260 14104
rect 9121 14046 9260 14048
rect 9121 14043 9187 14046
rect 9254 14044 9260 14046
rect 9324 14044 9330 14108
rect 11421 14106 11487 14109
rect 9676 14104 11487 14106
rect 9676 14048 11426 14104
rect 11482 14048 11487 14104
rect 9676 14046 11487 14048
rect 3252 13910 3986 13970
rect 3252 13908 3258 13910
rect 4286 13908 4292 13972
rect 4356 13970 4362 13972
rect 4981 13970 5047 13973
rect 4356 13968 5047 13970
rect 4356 13912 4986 13968
rect 5042 13912 5047 13968
rect 4356 13910 5047 13912
rect 4356 13908 4362 13910
rect 4981 13907 5047 13910
rect 6545 13970 6611 13973
rect 9676 13970 9736 14046
rect 11421 14043 11487 14046
rect 6545 13968 9736 13970
rect 6545 13912 6550 13968
rect 6606 13912 9736 13968
rect 6545 13910 9736 13912
rect 6545 13907 6611 13910
rect 9806 13908 9812 13972
rect 9876 13970 9882 13972
rect 12433 13970 12499 13973
rect 9876 13968 12499 13970
rect 9876 13912 12438 13968
rect 12494 13912 12499 13968
rect 9876 13910 12499 13912
rect 9876 13908 9882 13910
rect 12433 13907 12499 13910
rect 13629 13970 13695 13973
rect 16520 13970 17000 14000
rect 13629 13968 17000 13970
rect 13629 13912 13634 13968
rect 13690 13912 17000 13968
rect 13629 13910 17000 13912
rect 13629 13907 13695 13910
rect 16520 13880 17000 13910
rect 0 13834 480 13864
rect 3877 13834 3943 13837
rect 4613 13834 4679 13837
rect 0 13832 3943 13834
rect 0 13776 3882 13832
rect 3938 13776 3943 13832
rect 0 13774 3943 13776
rect 0 13744 480 13774
rect 3877 13771 3943 13774
rect 4064 13832 4679 13834
rect 4064 13776 4618 13832
rect 4674 13776 4679 13832
rect 4064 13774 4679 13776
rect 4064 13701 4124 13774
rect 4613 13771 4679 13774
rect 7005 13834 7071 13837
rect 12249 13834 12315 13837
rect 13905 13834 13971 13837
rect 7005 13832 12128 13834
rect 7005 13776 7010 13832
rect 7066 13776 12128 13832
rect 7005 13774 12128 13776
rect 7005 13771 7071 13774
rect 3417 13698 3483 13701
rect 4061 13698 4127 13701
rect 3417 13696 4127 13698
rect 3417 13640 3422 13696
rect 3478 13640 4066 13696
rect 4122 13640 4127 13696
rect 3417 13638 4127 13640
rect 3417 13635 3483 13638
rect 4061 13635 4127 13638
rect 4245 13698 4311 13701
rect 5533 13698 5599 13701
rect 4245 13696 5599 13698
rect 4245 13640 4250 13696
rect 4306 13640 5538 13696
rect 5594 13640 5599 13696
rect 4245 13638 5599 13640
rect 4245 13635 4311 13638
rect 5533 13635 5599 13638
rect 6637 13698 6703 13701
rect 11329 13698 11395 13701
rect 11462 13698 11468 13700
rect 6637 13696 10656 13698
rect 6637 13640 6642 13696
rect 6698 13640 10656 13696
rect 6637 13638 10656 13640
rect 6637 13635 6703 13638
rect 5874 13632 6194 13633
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6194 13632
rect 5874 13567 6194 13568
rect 10596 13565 10656 13638
rect 11329 13696 11468 13698
rect 11329 13640 11334 13696
rect 11390 13640 11468 13696
rect 11329 13638 11468 13640
rect 11329 13635 11395 13638
rect 11462 13636 11468 13638
rect 11532 13636 11538 13700
rect 12068 13698 12128 13774
rect 12249 13832 13971 13834
rect 12249 13776 12254 13832
rect 12310 13776 13910 13832
rect 13966 13776 13971 13832
rect 12249 13774 13971 13776
rect 12249 13771 12315 13774
rect 13905 13771 13971 13774
rect 13813 13698 13879 13701
rect 12068 13696 13879 13698
rect 12068 13640 13818 13696
rect 13874 13640 13879 13696
rect 12068 13638 13879 13640
rect 13813 13635 13879 13638
rect 10805 13632 11125 13633
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10805 13567 11125 13568
rect 4153 13562 4219 13565
rect 5441 13562 5507 13565
rect 4153 13560 5507 13562
rect 4153 13504 4158 13560
rect 4214 13504 5446 13560
rect 5502 13504 5507 13560
rect 4153 13502 5507 13504
rect 4153 13499 4219 13502
rect 5441 13499 5507 13502
rect 6729 13562 6795 13565
rect 8385 13562 8451 13565
rect 6729 13560 8451 13562
rect 6729 13504 6734 13560
rect 6790 13504 8390 13560
rect 8446 13504 8451 13560
rect 6729 13502 8451 13504
rect 6729 13499 6795 13502
rect 8385 13499 8451 13502
rect 8753 13562 8819 13565
rect 10409 13562 10475 13565
rect 8753 13560 10475 13562
rect 8753 13504 8758 13560
rect 8814 13504 10414 13560
rect 10470 13504 10475 13560
rect 8753 13502 10475 13504
rect 8753 13499 8819 13502
rect 10409 13499 10475 13502
rect 10593 13560 10659 13565
rect 10593 13504 10598 13560
rect 10654 13504 10659 13560
rect 10593 13499 10659 13504
rect 11329 13562 11395 13565
rect 12566 13562 12572 13564
rect 11329 13560 12572 13562
rect 11329 13504 11334 13560
rect 11390 13504 12572 13560
rect 11329 13502 12572 13504
rect 11329 13499 11395 13502
rect 12566 13500 12572 13502
rect 12636 13562 12642 13564
rect 13261 13562 13327 13565
rect 12636 13560 13327 13562
rect 12636 13504 13266 13560
rect 13322 13504 13327 13560
rect 12636 13502 13327 13504
rect 12636 13500 12642 13502
rect 13261 13499 13327 13502
rect 4705 13426 4771 13429
rect 5022 13426 5028 13428
rect 4705 13424 5028 13426
rect 4705 13368 4710 13424
rect 4766 13368 5028 13424
rect 4705 13366 5028 13368
rect 4705 13363 4771 13366
rect 5022 13364 5028 13366
rect 5092 13364 5098 13428
rect 7189 13426 7255 13429
rect 11421 13426 11487 13429
rect 11973 13428 12039 13429
rect 12157 13428 12223 13429
rect 11973 13426 12020 13428
rect 7189 13424 11487 13426
rect 7189 13368 7194 13424
rect 7250 13368 11426 13424
rect 11482 13368 11487 13424
rect 7189 13366 11487 13368
rect 11928 13424 12020 13426
rect 11928 13368 11978 13424
rect 11928 13366 12020 13368
rect 7189 13363 7255 13366
rect 11421 13363 11487 13366
rect 11973 13364 12020 13366
rect 12084 13364 12090 13428
rect 12157 13424 12204 13428
rect 12268 13426 12274 13428
rect 12157 13368 12162 13424
rect 12157 13364 12204 13368
rect 12268 13366 12314 13426
rect 12268 13364 12274 13366
rect 12566 13364 12572 13428
rect 12636 13426 12642 13428
rect 13445 13426 13511 13429
rect 12636 13424 13511 13426
rect 12636 13368 13450 13424
rect 13506 13368 13511 13424
rect 12636 13366 13511 13368
rect 12636 13364 12642 13366
rect 11973 13363 12039 13364
rect 12157 13363 12223 13364
rect 13445 13363 13511 13366
rect 13997 13428 14063 13429
rect 13997 13424 14044 13428
rect 14108 13426 14114 13428
rect 13997 13368 14002 13424
rect 13997 13364 14044 13368
rect 14108 13366 14154 13426
rect 14108 13364 14114 13366
rect 13997 13363 14063 13364
rect 1577 13290 1643 13293
rect 13997 13290 14063 13293
rect 1577 13288 14063 13290
rect 1577 13232 1582 13288
rect 1638 13232 14002 13288
rect 14058 13232 14063 13288
rect 1577 13230 14063 13232
rect 1577 13227 1643 13230
rect 13997 13227 14063 13230
rect 7925 13154 7991 13157
rect 8150 13154 8156 13156
rect 7925 13152 8156 13154
rect 7925 13096 7930 13152
rect 7986 13096 8156 13152
rect 7925 13094 8156 13096
rect 7925 13091 7991 13094
rect 8150 13092 8156 13094
rect 8220 13092 8226 13156
rect 8753 13154 8819 13157
rect 11421 13154 11487 13157
rect 8753 13152 11487 13154
rect 8753 13096 8758 13152
rect 8814 13096 11426 13152
rect 11482 13096 11487 13152
rect 8753 13094 11487 13096
rect 8753 13091 8819 13094
rect 11421 13091 11487 13094
rect 11646 13092 11652 13156
rect 11716 13154 11722 13156
rect 12341 13154 12407 13157
rect 11716 13152 12407 13154
rect 11716 13096 12346 13152
rect 12402 13096 12407 13152
rect 11716 13094 12407 13096
rect 11716 13092 11722 13094
rect 12341 13091 12407 13094
rect 3409 13088 3729 13089
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3409 13023 3729 13024
rect 8340 13088 8660 13089
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 13023 8660 13024
rect 13270 13088 13590 13089
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 13023 13590 13024
rect 4102 12956 4108 13020
rect 4172 13018 4178 13020
rect 5809 13018 5875 13021
rect 4172 13016 5875 13018
rect 4172 12960 5814 13016
rect 5870 12960 5875 13016
rect 4172 12958 5875 12960
rect 4172 12956 4178 12958
rect 5809 12955 5875 12958
rect 8886 12956 8892 13020
rect 8956 13018 8962 13020
rect 9673 13018 9739 13021
rect 8956 13016 9739 13018
rect 8956 12960 9678 13016
rect 9734 12960 9739 13016
rect 8956 12958 9739 12960
rect 8956 12956 8962 12958
rect 9673 12955 9739 12958
rect 9949 13018 10015 13021
rect 10174 13018 10180 13020
rect 9949 13016 10180 13018
rect 9949 12960 9954 13016
rect 10010 12960 10180 13016
rect 9949 12958 10180 12960
rect 9949 12955 10015 12958
rect 10174 12956 10180 12958
rect 10244 12956 10250 13020
rect 10409 13018 10475 13021
rect 11145 13018 11211 13021
rect 10409 13016 11211 13018
rect 10409 12960 10414 13016
rect 10470 12960 11150 13016
rect 11206 12960 11211 13016
rect 10409 12958 11211 12960
rect 10409 12955 10475 12958
rect 11145 12955 11211 12958
rect 11278 12956 11284 13020
rect 11348 13018 11354 13020
rect 11605 13018 11671 13021
rect 11348 13016 11671 13018
rect 11348 12960 11610 13016
rect 11666 12960 11671 13016
rect 11348 12958 11671 12960
rect 11348 12956 11354 12958
rect 11605 12955 11671 12958
rect 13721 13018 13787 13021
rect 13854 13018 13860 13020
rect 13721 13016 13860 13018
rect 13721 12960 13726 13016
rect 13782 12960 13860 13016
rect 13721 12958 13860 12960
rect 13721 12955 13787 12958
rect 13854 12956 13860 12958
rect 13924 12956 13930 13020
rect 0 12882 480 12912
rect 2865 12882 2931 12885
rect 7189 12882 7255 12885
rect 0 12880 2931 12882
rect 0 12824 2870 12880
rect 2926 12824 2931 12880
rect 0 12822 2931 12824
rect 0 12792 480 12822
rect 2865 12819 2931 12822
rect 5582 12880 7255 12882
rect 5582 12824 7194 12880
rect 7250 12824 7255 12880
rect 5582 12822 7255 12824
rect 2497 12746 2563 12749
rect 5582 12746 5642 12822
rect 7189 12819 7255 12822
rect 7833 12882 7899 12885
rect 13077 12882 13143 12885
rect 7833 12880 13143 12882
rect 7833 12824 7838 12880
rect 7894 12824 13082 12880
rect 13138 12824 13143 12880
rect 7833 12822 13143 12824
rect 7833 12819 7899 12822
rect 13077 12819 13143 12822
rect 2497 12744 5642 12746
rect 2497 12688 2502 12744
rect 2558 12688 5642 12744
rect 2497 12686 5642 12688
rect 5809 12746 5875 12749
rect 6453 12746 6519 12749
rect 11789 12746 11855 12749
rect 5809 12744 11855 12746
rect 5809 12688 5814 12744
rect 5870 12688 6458 12744
rect 6514 12688 11794 12744
rect 11850 12688 11855 12744
rect 5809 12686 11855 12688
rect 2497 12683 2563 12686
rect 5809 12683 5875 12686
rect 6453 12683 6519 12686
rect 11789 12683 11855 12686
rect 5390 12548 5396 12612
rect 5460 12610 5466 12612
rect 5625 12610 5691 12613
rect 5460 12608 5691 12610
rect 5460 12552 5630 12608
rect 5686 12552 5691 12608
rect 5460 12550 5691 12552
rect 5460 12548 5466 12550
rect 5625 12547 5691 12550
rect 9213 12610 9279 12613
rect 11237 12610 11303 12613
rect 12801 12610 12867 12613
rect 9213 12608 10380 12610
rect 9213 12552 9218 12608
rect 9274 12552 10380 12608
rect 9213 12550 10380 12552
rect 9213 12547 9279 12550
rect 5874 12544 6194 12545
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6194 12544
rect 5874 12479 6194 12480
rect 2313 12474 2379 12477
rect 5349 12474 5415 12477
rect 2313 12472 5415 12474
rect 2313 12416 2318 12472
rect 2374 12416 5354 12472
rect 5410 12416 5415 12472
rect 2313 12414 5415 12416
rect 2313 12411 2379 12414
rect 5349 12411 5415 12414
rect 6453 12474 6519 12477
rect 6862 12474 6868 12476
rect 6453 12472 6868 12474
rect 6453 12416 6458 12472
rect 6514 12416 6868 12472
rect 6453 12414 6868 12416
rect 6453 12411 6519 12414
rect 6862 12412 6868 12414
rect 6932 12412 6938 12476
rect 7833 12474 7899 12477
rect 9673 12474 9739 12477
rect 7833 12472 9739 12474
rect 7833 12416 7838 12472
rect 7894 12416 9678 12472
rect 9734 12416 9739 12472
rect 7833 12414 9739 12416
rect 7833 12411 7899 12414
rect 9673 12411 9739 12414
rect 9806 12412 9812 12476
rect 9876 12474 9882 12476
rect 10133 12474 10199 12477
rect 9876 12472 10199 12474
rect 9876 12416 10138 12472
rect 10194 12416 10199 12472
rect 9876 12414 10199 12416
rect 9876 12412 9882 12414
rect 10133 12411 10199 12414
rect 3141 12340 3207 12341
rect 3141 12338 3188 12340
rect 3096 12336 3188 12338
rect 3096 12280 3146 12336
rect 3096 12278 3188 12280
rect 3141 12276 3188 12278
rect 3252 12276 3258 12340
rect 6913 12338 6979 12341
rect 9581 12338 9647 12341
rect 6913 12336 9647 12338
rect 6913 12280 6918 12336
rect 6974 12280 9586 12336
rect 9642 12280 9647 12336
rect 6913 12278 9647 12280
rect 10320 12338 10380 12550
rect 11237 12608 12867 12610
rect 11237 12552 11242 12608
rect 11298 12552 12806 12608
rect 12862 12552 12867 12608
rect 11237 12550 12867 12552
rect 11237 12547 11303 12550
rect 12801 12547 12867 12550
rect 10805 12544 11125 12545
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10805 12479 11125 12480
rect 14181 12474 14247 12477
rect 11240 12472 14247 12474
rect 11240 12416 14186 12472
rect 14242 12416 14247 12472
rect 11240 12414 14247 12416
rect 11240 12338 11300 12414
rect 14181 12411 14247 12414
rect 10320 12278 11300 12338
rect 3141 12275 3207 12276
rect 6913 12275 6979 12278
rect 9581 12275 9647 12278
rect 12382 12276 12388 12340
rect 12452 12338 12458 12340
rect 13721 12338 13787 12341
rect 12452 12336 13787 12338
rect 12452 12280 13726 12336
rect 13782 12280 13787 12336
rect 12452 12278 13787 12280
rect 12452 12276 12458 12278
rect 13721 12275 13787 12278
rect 2773 12202 2839 12205
rect 4889 12202 4955 12205
rect 7281 12202 7347 12205
rect 2773 12200 4768 12202
rect 2773 12144 2778 12200
rect 2834 12144 4768 12200
rect 2773 12142 4768 12144
rect 2773 12139 2839 12142
rect 4708 12066 4768 12142
rect 4889 12200 7347 12202
rect 4889 12144 4894 12200
rect 4950 12144 7286 12200
rect 7342 12144 7347 12200
rect 4889 12142 7347 12144
rect 4889 12139 4955 12142
rect 7281 12139 7347 12142
rect 7465 12202 7531 12205
rect 14273 12202 14339 12205
rect 7465 12200 14339 12202
rect 7465 12144 7470 12200
rect 7526 12144 14278 12200
rect 14334 12144 14339 12200
rect 7465 12142 14339 12144
rect 7465 12139 7531 12142
rect 14273 12139 14339 12142
rect 7833 12068 7899 12069
rect 6494 12066 6500 12068
rect 4708 12006 6500 12066
rect 6494 12004 6500 12006
rect 6564 12004 6570 12068
rect 7782 12004 7788 12068
rect 7852 12066 7899 12068
rect 8845 12066 8911 12069
rect 9213 12066 9279 12069
rect 7852 12064 7944 12066
rect 7894 12008 7944 12064
rect 7852 12006 7944 12008
rect 8845 12064 9279 12066
rect 8845 12008 8850 12064
rect 8906 12008 9218 12064
rect 9274 12008 9279 12064
rect 8845 12006 9279 12008
rect 7852 12004 7899 12006
rect 7833 12003 7899 12004
rect 8845 12003 8911 12006
rect 9213 12003 9279 12006
rect 10542 12004 10548 12068
rect 10612 12066 10618 12068
rect 10869 12066 10935 12069
rect 12709 12066 12775 12069
rect 12893 12066 12959 12069
rect 10612 12064 12959 12066
rect 10612 12008 10874 12064
rect 10930 12008 12714 12064
rect 12770 12008 12898 12064
rect 12954 12008 12959 12064
rect 10612 12006 12959 12008
rect 10612 12004 10618 12006
rect 10869 12003 10935 12006
rect 12709 12003 12775 12006
rect 12893 12003 12959 12006
rect 3409 12000 3729 12001
rect 0 11930 480 11960
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 11935 3729 11936
rect 8340 12000 8660 12001
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 11935 8660 11936
rect 13270 12000 13590 12001
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 11935 13590 11936
rect 1853 11930 1919 11933
rect 0 11928 1919 11930
rect 0 11872 1858 11928
rect 1914 11872 1919 11928
rect 0 11870 1919 11872
rect 0 11840 480 11870
rect 1853 11867 1919 11870
rect 4061 11930 4127 11933
rect 5717 11930 5783 11933
rect 8109 11930 8175 11933
rect 4061 11928 8175 11930
rect 4061 11872 4066 11928
rect 4122 11872 5722 11928
rect 5778 11872 8114 11928
rect 8170 11872 8175 11928
rect 4061 11870 8175 11872
rect 4061 11867 4127 11870
rect 5717 11867 5783 11870
rect 8109 11867 8175 11870
rect 8886 11868 8892 11932
rect 8956 11930 8962 11932
rect 8956 11870 13186 11930
rect 8956 11868 8962 11870
rect 5441 11794 5507 11797
rect 10961 11794 11027 11797
rect 5441 11792 11027 11794
rect 5441 11736 5446 11792
rect 5502 11736 10966 11792
rect 11022 11736 11027 11792
rect 5441 11734 11027 11736
rect 5441 11731 5507 11734
rect 10961 11731 11027 11734
rect 11329 11794 11395 11797
rect 11646 11794 11652 11796
rect 11329 11792 11652 11794
rect 11329 11736 11334 11792
rect 11390 11736 11652 11792
rect 11329 11734 11652 11736
rect 11329 11731 11395 11734
rect 11646 11732 11652 11734
rect 11716 11732 11722 11796
rect 13126 11794 13186 11870
rect 13905 11794 13971 11797
rect 13126 11792 13971 11794
rect 13126 11736 13910 11792
rect 13966 11736 13971 11792
rect 13126 11734 13971 11736
rect 13905 11731 13971 11734
rect 2313 11658 2379 11661
rect 8886 11658 8892 11660
rect 2313 11656 8892 11658
rect 2313 11600 2318 11656
rect 2374 11600 8892 11656
rect 2313 11598 8892 11600
rect 2313 11595 2379 11598
rect 8886 11596 8892 11598
rect 8956 11596 8962 11660
rect 9622 11596 9628 11660
rect 9692 11658 9698 11660
rect 9990 11658 9996 11660
rect 9692 11598 9996 11658
rect 9692 11596 9698 11598
rect 9990 11596 9996 11598
rect 10060 11596 10066 11660
rect 13629 11658 13695 11661
rect 10596 11656 13695 11658
rect 10596 11600 13634 11656
rect 13690 11600 13695 11656
rect 10596 11598 13695 11600
rect 6269 11522 6335 11525
rect 10596 11522 10656 11598
rect 13629 11595 13695 11598
rect 11329 11524 11395 11525
rect 6269 11520 10656 11522
rect 6269 11464 6274 11520
rect 6330 11464 10656 11520
rect 6269 11462 10656 11464
rect 6269 11459 6335 11462
rect 11278 11460 11284 11524
rect 11348 11522 11395 11524
rect 12709 11522 12775 11525
rect 14181 11524 14247 11525
rect 13854 11522 13860 11524
rect 11348 11520 11440 11522
rect 11390 11464 11440 11520
rect 11348 11462 11440 11464
rect 12709 11520 13860 11522
rect 12709 11464 12714 11520
rect 12770 11464 13860 11520
rect 12709 11462 13860 11464
rect 11348 11460 11395 11462
rect 11329 11459 11395 11460
rect 12709 11459 12775 11462
rect 13854 11460 13860 11462
rect 13924 11460 13930 11524
rect 14181 11522 14228 11524
rect 14136 11520 14228 11522
rect 14136 11464 14186 11520
rect 14136 11462 14228 11464
rect 14181 11460 14228 11462
rect 14292 11460 14298 11524
rect 14181 11459 14247 11460
rect 5874 11456 6194 11457
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6194 11456
rect 5874 11391 6194 11392
rect 10805 11456 11125 11457
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 11391 11125 11392
rect 5441 11388 5507 11389
rect 5390 11324 5396 11388
rect 5460 11386 5507 11388
rect 6729 11386 6795 11389
rect 8201 11386 8267 11389
rect 5460 11384 5552 11386
rect 5502 11328 5552 11384
rect 5460 11326 5552 11328
rect 6729 11384 8267 11386
rect 6729 11328 6734 11384
rect 6790 11328 8206 11384
rect 8262 11328 8267 11384
rect 6729 11326 8267 11328
rect 5460 11324 5507 11326
rect 5441 11323 5507 11324
rect 6729 11323 6795 11326
rect 8201 11323 8267 11326
rect 9029 11386 9095 11389
rect 10225 11386 10291 11389
rect 9029 11384 10291 11386
rect 9029 11328 9034 11384
rect 9090 11328 10230 11384
rect 10286 11328 10291 11384
rect 9029 11326 10291 11328
rect 9029 11323 9095 11326
rect 10225 11323 10291 11326
rect 10501 11388 10567 11389
rect 10501 11384 10548 11388
rect 10612 11386 10618 11388
rect 10501 11328 10506 11384
rect 10501 11324 10548 11328
rect 10612 11326 10658 11386
rect 10612 11324 10618 11326
rect 11278 11324 11284 11388
rect 11348 11386 11354 11388
rect 12750 11386 12756 11388
rect 11348 11326 12756 11386
rect 11348 11324 11354 11326
rect 12750 11324 12756 11326
rect 12820 11324 12826 11388
rect 10501 11323 10567 11324
rect 1945 11250 2011 11253
rect 14273 11250 14339 11253
rect 1945 11248 14339 11250
rect 1945 11192 1950 11248
rect 2006 11192 14278 11248
rect 14334 11192 14339 11248
rect 1945 11190 14339 11192
rect 1945 11187 2011 11190
rect 14273 11187 14339 11190
rect 3182 11052 3188 11116
rect 3252 11114 3258 11116
rect 3693 11114 3759 11117
rect 5349 11114 5415 11117
rect 9673 11114 9739 11117
rect 3252 11112 5274 11114
rect 3252 11056 3698 11112
rect 3754 11056 5274 11112
rect 3252 11054 5274 11056
rect 3252 11052 3258 11054
rect 3693 11051 3759 11054
rect 0 10978 480 11008
rect 2998 10978 3004 10980
rect 0 10918 3004 10978
rect 0 10888 480 10918
rect 2998 10916 3004 10918
rect 3068 10916 3074 10980
rect 5214 10978 5274 11054
rect 5349 11112 9739 11114
rect 5349 11056 5354 11112
rect 5410 11056 9678 11112
rect 9734 11056 9739 11112
rect 5349 11054 9739 11056
rect 5349 11051 5415 11054
rect 9673 11051 9739 11054
rect 10041 11114 10107 11117
rect 10174 11114 10180 11116
rect 10041 11112 10180 11114
rect 10041 11056 10046 11112
rect 10102 11056 10180 11112
rect 10041 11054 10180 11056
rect 10041 11051 10107 11054
rect 10174 11052 10180 11054
rect 10244 11052 10250 11116
rect 14549 11114 14615 11117
rect 12022 11112 14615 11114
rect 12022 11056 14554 11112
rect 14610 11056 14615 11112
rect 12022 11054 14615 11056
rect 6913 10978 6979 10981
rect 9029 10978 9095 10981
rect 12022 10978 12082 11054
rect 14549 11051 14615 11054
rect 5214 10976 8172 10978
rect 5214 10920 6918 10976
rect 6974 10920 8172 10976
rect 5214 10918 8172 10920
rect 6913 10915 6979 10918
rect 3409 10912 3729 10913
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 10847 3729 10848
rect 5390 10780 5396 10844
rect 5460 10842 5466 10844
rect 7230 10842 7236 10844
rect 5460 10782 7236 10842
rect 5460 10780 5466 10782
rect 7230 10780 7236 10782
rect 7300 10842 7306 10844
rect 7465 10842 7531 10845
rect 7300 10840 7531 10842
rect 7300 10784 7470 10840
rect 7526 10784 7531 10840
rect 7300 10782 7531 10784
rect 7300 10780 7306 10782
rect 7465 10779 7531 10782
rect 3601 10706 3667 10709
rect 8112 10706 8172 10918
rect 9029 10976 12082 10978
rect 9029 10920 9034 10976
rect 9090 10920 12082 10976
rect 9029 10918 12082 10920
rect 9029 10915 9095 10918
rect 12382 10916 12388 10980
rect 12452 10978 12458 10980
rect 12893 10978 12959 10981
rect 12452 10976 12959 10978
rect 12452 10920 12898 10976
rect 12954 10920 12959 10976
rect 12452 10918 12959 10920
rect 12452 10916 12458 10918
rect 12893 10915 12959 10918
rect 8340 10912 8660 10913
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 10847 8660 10848
rect 13270 10912 13590 10913
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 10847 13590 10848
rect 9765 10842 9831 10845
rect 11053 10842 11119 10845
rect 9765 10840 11119 10842
rect 9765 10784 9770 10840
rect 9826 10784 11058 10840
rect 11114 10784 11119 10840
rect 9765 10782 11119 10784
rect 9765 10779 9831 10782
rect 11053 10779 11119 10782
rect 9305 10706 9371 10709
rect 3601 10704 8034 10706
rect 3601 10648 3606 10704
rect 3662 10648 8034 10704
rect 3601 10646 8034 10648
rect 8112 10704 9371 10706
rect 8112 10648 9310 10704
rect 9366 10648 9371 10704
rect 8112 10646 9371 10648
rect 3601 10643 3667 10646
rect 1853 10570 1919 10573
rect 7833 10570 7899 10573
rect 1853 10568 7899 10570
rect 1853 10512 1858 10568
rect 1914 10512 7838 10568
rect 7894 10512 7899 10568
rect 1853 10510 7899 10512
rect 7974 10570 8034 10646
rect 9305 10643 9371 10646
rect 10501 10706 10567 10709
rect 12934 10706 12940 10708
rect 10501 10704 12940 10706
rect 10501 10648 10506 10704
rect 10562 10648 12940 10704
rect 10501 10646 12940 10648
rect 10501 10643 10567 10646
rect 12934 10644 12940 10646
rect 13004 10644 13010 10708
rect 9806 10570 9812 10572
rect 7974 10510 9812 10570
rect 1853 10507 1919 10510
rect 7833 10507 7899 10510
rect 9806 10508 9812 10510
rect 9876 10570 9882 10572
rect 12566 10570 12572 10572
rect 9876 10510 12572 10570
rect 9876 10508 9882 10510
rect 12566 10508 12572 10510
rect 12636 10508 12642 10572
rect 12934 10508 12940 10572
rect 13004 10570 13010 10572
rect 13077 10570 13143 10573
rect 13004 10568 13143 10570
rect 13004 10512 13082 10568
rect 13138 10512 13143 10568
rect 13004 10510 13143 10512
rect 13004 10508 13010 10510
rect 13077 10507 13143 10510
rect 13261 10570 13327 10573
rect 14038 10570 14044 10572
rect 13261 10568 14044 10570
rect 13261 10512 13266 10568
rect 13322 10512 14044 10568
rect 13261 10510 14044 10512
rect 13261 10507 13327 10510
rect 14038 10508 14044 10510
rect 14108 10570 14114 10572
rect 15193 10570 15259 10573
rect 14108 10568 15259 10570
rect 14108 10512 15198 10568
rect 15254 10512 15259 10568
rect 14108 10510 15259 10512
rect 14108 10508 14114 10510
rect 15193 10507 15259 10510
rect 2998 10372 3004 10436
rect 3068 10434 3074 10436
rect 4061 10434 4127 10437
rect 3068 10432 4127 10434
rect 3068 10376 4066 10432
rect 4122 10376 4127 10432
rect 3068 10374 4127 10376
rect 3068 10372 3074 10374
rect 4061 10371 4127 10374
rect 8150 10372 8156 10436
rect 8220 10434 8226 10436
rect 8937 10434 9003 10437
rect 8220 10432 9003 10434
rect 8220 10376 8942 10432
rect 8998 10376 9003 10432
rect 8220 10374 9003 10376
rect 8220 10372 8226 10374
rect 8937 10371 9003 10374
rect 9622 10372 9628 10436
rect 9692 10434 9698 10436
rect 10409 10434 10475 10437
rect 9692 10432 10475 10434
rect 9692 10376 10414 10432
rect 10470 10376 10475 10432
rect 9692 10374 10475 10376
rect 9692 10372 9698 10374
rect 10409 10371 10475 10374
rect 12893 10434 12959 10437
rect 14222 10434 14228 10436
rect 12893 10432 14228 10434
rect 12893 10376 12898 10432
rect 12954 10376 14228 10432
rect 12893 10374 14228 10376
rect 12893 10371 12959 10374
rect 14222 10372 14228 10374
rect 14292 10372 14298 10436
rect 5874 10368 6194 10369
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6194 10368
rect 5874 10303 6194 10304
rect 10805 10368 11125 10369
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10805 10303 11125 10304
rect 2497 10298 2563 10301
rect 4889 10298 4955 10301
rect 2497 10296 4955 10298
rect 2497 10240 2502 10296
rect 2558 10240 4894 10296
rect 4950 10240 4955 10296
rect 2497 10238 4955 10240
rect 2497 10235 2563 10238
rect 4889 10235 4955 10238
rect 6494 10236 6500 10300
rect 6564 10298 6570 10300
rect 9029 10298 9095 10301
rect 6564 10296 9095 10298
rect 6564 10240 9034 10296
rect 9090 10240 9095 10296
rect 6564 10238 9095 10240
rect 6564 10236 6570 10238
rect 9029 10235 9095 10238
rect 9622 10236 9628 10300
rect 9692 10298 9698 10300
rect 9949 10298 10015 10301
rect 9692 10296 10015 10298
rect 9692 10240 9954 10296
rect 10010 10240 10015 10296
rect 9692 10238 10015 10240
rect 9692 10236 9698 10238
rect 9949 10235 10015 10238
rect 1393 10162 1459 10165
rect 3601 10162 3667 10165
rect 9438 10162 9444 10164
rect 1393 10160 3667 10162
rect 1393 10104 1398 10160
rect 1454 10104 3606 10160
rect 3662 10104 3667 10160
rect 1393 10102 3667 10104
rect 1393 10099 1459 10102
rect 3601 10099 3667 10102
rect 3742 10102 9444 10162
rect 0 10026 480 10056
rect 565 10026 631 10029
rect 0 10024 631 10026
rect 0 9968 570 10024
rect 626 9968 631 10024
rect 0 9966 631 9968
rect 0 9936 480 9966
rect 565 9963 631 9966
rect 2681 10026 2747 10029
rect 3742 10026 3802 10102
rect 9438 10100 9444 10102
rect 9508 10162 9514 10164
rect 12893 10162 12959 10165
rect 9508 10160 12959 10162
rect 9508 10104 12898 10160
rect 12954 10104 12959 10160
rect 9508 10102 12959 10104
rect 9508 10100 9514 10102
rect 12893 10099 12959 10102
rect 4061 10028 4127 10029
rect 4061 10026 4108 10028
rect 2681 10024 3802 10026
rect 2681 9968 2686 10024
rect 2742 9968 3802 10024
rect 2681 9966 3802 9968
rect 4016 10024 4108 10026
rect 4016 9968 4066 10024
rect 4016 9966 4108 9968
rect 2681 9963 2747 9966
rect 4061 9964 4108 9966
rect 4172 9964 4178 10028
rect 4521 10026 4587 10029
rect 6678 10026 6684 10028
rect 4521 10024 6684 10026
rect 4521 9968 4526 10024
rect 4582 9968 6684 10024
rect 4521 9966 6684 9968
rect 4061 9963 4127 9964
rect 4521 9963 4587 9966
rect 6678 9964 6684 9966
rect 6748 9964 6754 10028
rect 14181 10026 14247 10029
rect 6824 10024 14247 10026
rect 6824 9968 14186 10024
rect 14242 9968 14247 10024
rect 6824 9966 14247 9968
rect 4613 9890 4679 9893
rect 5349 9890 5415 9893
rect 6824 9890 6884 9966
rect 14181 9963 14247 9966
rect 4613 9888 6884 9890
rect 4613 9832 4618 9888
rect 4674 9832 5354 9888
rect 5410 9832 6884 9888
rect 4613 9830 6884 9832
rect 4613 9827 4679 9830
rect 5349 9827 5415 9830
rect 9070 9828 9076 9892
rect 9140 9890 9146 9892
rect 9213 9890 9279 9893
rect 9140 9888 9279 9890
rect 9140 9832 9218 9888
rect 9274 9832 9279 9888
rect 9140 9830 9279 9832
rect 9140 9828 9146 9830
rect 9213 9827 9279 9830
rect 15469 9890 15535 9893
rect 16520 9890 17000 9920
rect 15469 9888 17000 9890
rect 15469 9832 15474 9888
rect 15530 9832 17000 9888
rect 15469 9830 17000 9832
rect 15469 9827 15535 9830
rect 3409 9824 3729 9825
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 9759 3729 9760
rect 8340 9824 8660 9825
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 9759 8660 9760
rect 13270 9824 13590 9825
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 16520 9800 17000 9830
rect 13270 9759 13590 9760
rect 4889 9754 4955 9757
rect 5993 9754 6059 9757
rect 4889 9752 6059 9754
rect 4889 9696 4894 9752
rect 4950 9696 5998 9752
rect 6054 9696 6059 9752
rect 4889 9694 6059 9696
rect 4889 9691 4955 9694
rect 5993 9691 6059 9694
rect 9121 9754 9187 9757
rect 9254 9754 9260 9756
rect 9121 9752 9260 9754
rect 9121 9696 9126 9752
rect 9182 9696 9260 9752
rect 9121 9694 9260 9696
rect 9121 9691 9187 9694
rect 9254 9692 9260 9694
rect 9324 9692 9330 9756
rect 3601 9618 3667 9621
rect 6269 9618 6335 9621
rect 3601 9616 6335 9618
rect 3601 9560 3606 9616
rect 3662 9560 6274 9616
rect 6330 9560 6335 9616
rect 3601 9558 6335 9560
rect 3601 9555 3667 9558
rect 6269 9555 6335 9558
rect 6637 9618 6703 9621
rect 13813 9618 13879 9621
rect 13997 9620 14063 9621
rect 13997 9618 14044 9620
rect 6637 9616 13879 9618
rect 6637 9560 6642 9616
rect 6698 9560 13818 9616
rect 13874 9560 13879 9616
rect 6637 9558 13879 9560
rect 13952 9616 14044 9618
rect 13952 9560 14002 9616
rect 13952 9558 14044 9560
rect 6637 9555 6703 9558
rect 13813 9555 13879 9558
rect 13997 9556 14044 9558
rect 14108 9556 14114 9620
rect 13997 9555 14063 9556
rect 1669 9482 1735 9485
rect 12934 9482 12940 9484
rect 1669 9480 12940 9482
rect 1669 9424 1674 9480
rect 1730 9424 12940 9480
rect 1669 9422 12940 9424
rect 1669 9419 1735 9422
rect 12934 9420 12940 9422
rect 13004 9482 13010 9484
rect 13445 9482 13511 9485
rect 13004 9480 13511 9482
rect 13004 9424 13450 9480
rect 13506 9424 13511 9480
rect 13004 9422 13511 9424
rect 13004 9420 13010 9422
rect 13445 9419 13511 9422
rect 8109 9346 8175 9349
rect 10501 9346 10567 9349
rect 8109 9344 10567 9346
rect 8109 9288 8114 9344
rect 8170 9288 10506 9344
rect 10562 9288 10567 9344
rect 8109 9286 10567 9288
rect 8109 9283 8175 9286
rect 10501 9283 10567 9286
rect 12433 9346 12499 9349
rect 13854 9346 13860 9348
rect 12433 9344 13860 9346
rect 12433 9288 12438 9344
rect 12494 9288 13860 9344
rect 12433 9286 13860 9288
rect 12433 9283 12499 9286
rect 13854 9284 13860 9286
rect 13924 9284 13930 9348
rect 5874 9280 6194 9281
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6194 9280
rect 5874 9215 6194 9216
rect 10805 9280 11125 9281
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 9215 11125 9216
rect 9581 9210 9647 9213
rect 7836 9208 9647 9210
rect 7836 9152 9586 9208
rect 9642 9152 9647 9208
rect 7836 9150 9647 9152
rect 0 9074 480 9104
rect 2773 9074 2839 9077
rect 7836 9074 7896 9150
rect 9581 9147 9647 9150
rect 11462 9148 11468 9212
rect 11532 9210 11538 9212
rect 13629 9210 13695 9213
rect 11532 9208 13695 9210
rect 11532 9152 13634 9208
rect 13690 9152 13695 9208
rect 11532 9150 13695 9152
rect 11532 9148 11538 9150
rect 13629 9147 13695 9150
rect 0 9072 2839 9074
rect 0 9016 2778 9072
rect 2834 9016 2839 9072
rect 0 9014 2839 9016
rect 0 8984 480 9014
rect 2773 9011 2839 9014
rect 4846 9014 7896 9074
rect 2037 8938 2103 8941
rect 4846 8938 4906 9014
rect 7966 9012 7972 9076
rect 8036 9074 8042 9076
rect 14457 9074 14523 9077
rect 8036 9072 14523 9074
rect 8036 9016 14462 9072
rect 14518 9016 14523 9072
rect 8036 9014 14523 9016
rect 8036 9012 8042 9014
rect 14457 9011 14523 9014
rect 2037 8936 4906 8938
rect 2037 8880 2042 8936
rect 2098 8880 4906 8936
rect 2037 8878 4906 8880
rect 5073 8938 5139 8941
rect 12566 8938 12572 8940
rect 5073 8936 12572 8938
rect 5073 8880 5078 8936
rect 5134 8880 12572 8936
rect 5073 8878 12572 8880
rect 2037 8875 2103 8878
rect 5073 8875 5139 8878
rect 12566 8876 12572 8878
rect 12636 8876 12642 8940
rect 5533 8802 5599 8805
rect 8201 8802 8267 8805
rect 5533 8800 8267 8802
rect 5533 8744 5538 8800
rect 5594 8744 8206 8800
rect 8262 8744 8267 8800
rect 5533 8742 8267 8744
rect 5533 8739 5599 8742
rect 8201 8739 8267 8742
rect 9070 8740 9076 8804
rect 9140 8802 9146 8804
rect 12014 8802 12020 8804
rect 9140 8742 12020 8802
rect 9140 8740 9146 8742
rect 12014 8740 12020 8742
rect 12084 8802 12090 8804
rect 12525 8802 12591 8805
rect 12084 8800 12591 8802
rect 12084 8744 12530 8800
rect 12586 8744 12591 8800
rect 12084 8742 12591 8744
rect 12084 8740 12090 8742
rect 12525 8739 12591 8742
rect 3409 8736 3729 8737
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 8671 3729 8672
rect 8340 8736 8660 8737
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8340 8671 8660 8672
rect 13270 8736 13590 8737
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 8671 13590 8672
rect 6862 8604 6868 8668
rect 6932 8666 6938 8668
rect 8845 8666 8911 8669
rect 11881 8666 11947 8669
rect 12014 8666 12020 8668
rect 6932 8606 7298 8666
rect 6932 8604 6938 8606
rect 2957 8530 3023 8533
rect 7097 8530 7163 8533
rect 2957 8528 7163 8530
rect 2957 8472 2962 8528
rect 3018 8472 7102 8528
rect 7158 8472 7163 8528
rect 2957 8470 7163 8472
rect 7238 8530 7298 8606
rect 8845 8664 12020 8666
rect 8845 8608 8850 8664
rect 8906 8608 11886 8664
rect 11942 8608 12020 8664
rect 8845 8606 12020 8608
rect 8845 8603 8911 8606
rect 11881 8603 11947 8606
rect 12014 8604 12020 8606
rect 12084 8604 12090 8668
rect 15009 8530 15075 8533
rect 7238 8528 15075 8530
rect 7238 8472 15014 8528
rect 15070 8472 15075 8528
rect 7238 8470 15075 8472
rect 2957 8467 3023 8470
rect 7097 8467 7163 8470
rect 15009 8467 15075 8470
rect 4153 8394 4219 8397
rect 4153 8392 7160 8394
rect 4153 8336 4158 8392
rect 4214 8336 7160 8392
rect 4153 8334 7160 8336
rect 4153 8331 4219 8334
rect 7100 8258 7160 8334
rect 7230 8332 7236 8396
rect 7300 8394 7306 8396
rect 15009 8394 15075 8397
rect 7300 8392 15075 8394
rect 7300 8336 15014 8392
rect 15070 8336 15075 8392
rect 7300 8334 15075 8336
rect 7300 8332 7306 8334
rect 15009 8331 15075 8334
rect 7414 8258 7420 8260
rect 7100 8198 7420 8258
rect 7414 8196 7420 8198
rect 7484 8258 7490 8260
rect 8845 8258 8911 8261
rect 7484 8256 8911 8258
rect 7484 8200 8850 8256
rect 8906 8200 8911 8256
rect 7484 8198 8911 8200
rect 7484 8196 7490 8198
rect 8845 8195 8911 8198
rect 9857 8258 9923 8261
rect 12341 8260 12407 8261
rect 9990 8258 9996 8260
rect 9857 8256 9996 8258
rect 9857 8200 9862 8256
rect 9918 8200 9996 8256
rect 9857 8198 9996 8200
rect 9857 8195 9923 8198
rect 9990 8196 9996 8198
rect 10060 8196 10066 8260
rect 12341 8256 12388 8260
rect 12452 8258 12458 8260
rect 12341 8200 12346 8256
rect 12341 8196 12388 8200
rect 12452 8198 12498 8258
rect 12452 8196 12458 8198
rect 12341 8195 12407 8196
rect 5874 8192 6194 8193
rect 0 8122 480 8152
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6194 8192
rect 5874 8127 6194 8128
rect 10805 8192 11125 8193
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 8127 11125 8128
rect 3049 8122 3115 8125
rect 0 8120 3115 8122
rect 0 8064 3054 8120
rect 3110 8064 3115 8120
rect 0 8062 3115 8064
rect 0 8032 480 8062
rect 3049 8059 3115 8062
rect 7281 8122 7347 8125
rect 8845 8122 8911 8125
rect 7281 8120 8911 8122
rect 7281 8064 7286 8120
rect 7342 8064 8850 8120
rect 8906 8064 8911 8120
rect 7281 8062 8911 8064
rect 7281 8059 7347 8062
rect 8845 8059 8911 8062
rect 3785 7986 3851 7989
rect 12249 7986 12315 7989
rect 3785 7984 12315 7986
rect 3785 7928 3790 7984
rect 3846 7928 12254 7984
rect 12310 7928 12315 7984
rect 3785 7926 12315 7928
rect 3785 7923 3851 7926
rect 12249 7923 12315 7926
rect 12525 7986 12591 7989
rect 12750 7986 12756 7988
rect 12525 7984 12756 7986
rect 12525 7928 12530 7984
rect 12586 7928 12756 7984
rect 12525 7926 12756 7928
rect 12525 7923 12591 7926
rect 12750 7924 12756 7926
rect 12820 7924 12826 7988
rect 1761 7850 1827 7853
rect 12750 7850 12756 7852
rect 1761 7848 12756 7850
rect 1761 7792 1766 7848
rect 1822 7792 12756 7848
rect 1761 7790 12756 7792
rect 1761 7787 1827 7790
rect 12750 7788 12756 7790
rect 12820 7788 12826 7852
rect 6545 7714 6611 7717
rect 7281 7714 7347 7717
rect 6545 7712 7347 7714
rect 6545 7656 6550 7712
rect 6606 7656 7286 7712
rect 7342 7656 7347 7712
rect 6545 7654 7347 7656
rect 6545 7651 6611 7654
rect 7281 7651 7347 7654
rect 7557 7714 7623 7717
rect 8109 7714 8175 7717
rect 7557 7712 8175 7714
rect 7557 7656 7562 7712
rect 7618 7656 8114 7712
rect 8170 7656 8175 7712
rect 7557 7654 8175 7656
rect 7557 7651 7623 7654
rect 8109 7651 8175 7654
rect 10174 7652 10180 7716
rect 10244 7714 10250 7716
rect 13077 7714 13143 7717
rect 10244 7712 13143 7714
rect 10244 7656 13082 7712
rect 13138 7656 13143 7712
rect 10244 7654 13143 7656
rect 10244 7652 10250 7654
rect 13077 7651 13143 7654
rect 3409 7648 3729 7649
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 7583 3729 7584
rect 8340 7648 8660 7649
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 7583 8660 7584
rect 13270 7648 13590 7649
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13270 7583 13590 7584
rect 5165 7578 5231 7581
rect 8201 7578 8267 7581
rect 5165 7576 8267 7578
rect 5165 7520 5170 7576
rect 5226 7520 8206 7576
rect 8262 7520 8267 7576
rect 5165 7518 8267 7520
rect 5165 7515 5231 7518
rect 8201 7515 8267 7518
rect 9254 7516 9260 7580
rect 9324 7578 9330 7580
rect 10685 7578 10751 7581
rect 9324 7576 10751 7578
rect 9324 7520 10690 7576
rect 10746 7520 10751 7576
rect 9324 7518 10751 7520
rect 9324 7516 9330 7518
rect 10685 7515 10751 7518
rect 5993 7442 6059 7445
rect 7741 7442 7807 7445
rect 11881 7442 11947 7445
rect 5993 7440 6700 7442
rect 5993 7384 5998 7440
rect 6054 7384 6700 7440
rect 5993 7382 6700 7384
rect 5993 7379 6059 7382
rect 1945 7306 2011 7309
rect 6640 7306 6700 7382
rect 7741 7440 11947 7442
rect 7741 7384 7746 7440
rect 7802 7384 11886 7440
rect 11942 7384 11947 7440
rect 7741 7382 11947 7384
rect 7741 7379 7807 7382
rect 11881 7379 11947 7382
rect 12249 7442 12315 7445
rect 13721 7442 13787 7445
rect 12249 7440 13787 7442
rect 12249 7384 12254 7440
rect 12310 7384 13726 7440
rect 13782 7384 13787 7440
rect 12249 7382 13787 7384
rect 12249 7379 12315 7382
rect 13721 7379 13787 7382
rect 10961 7306 11027 7309
rect 1945 7304 6562 7306
rect 1945 7248 1950 7304
rect 2006 7248 6562 7304
rect 1945 7246 6562 7248
rect 6640 7304 11027 7306
rect 6640 7248 10966 7304
rect 11022 7248 11027 7304
rect 6640 7246 11027 7248
rect 1945 7243 2011 7246
rect 0 7170 480 7200
rect 5073 7170 5139 7173
rect 0 7168 5139 7170
rect 0 7112 5078 7168
rect 5134 7112 5139 7168
rect 0 7110 5139 7112
rect 6502 7170 6562 7246
rect 10961 7243 11027 7246
rect 12617 7306 12683 7309
rect 13905 7306 13971 7309
rect 12617 7304 13971 7306
rect 12617 7248 12622 7304
rect 12678 7248 13910 7304
rect 13966 7248 13971 7304
rect 12617 7246 13971 7248
rect 12617 7243 12683 7246
rect 13905 7243 13971 7246
rect 14181 7308 14247 7309
rect 14181 7304 14228 7308
rect 14292 7306 14298 7308
rect 14181 7248 14186 7304
rect 14181 7244 14228 7248
rect 14292 7246 14338 7306
rect 14292 7244 14298 7246
rect 14181 7243 14247 7244
rect 9254 7170 9260 7172
rect 6502 7110 9260 7170
rect 0 7080 480 7110
rect 5073 7107 5139 7110
rect 9254 7108 9260 7110
rect 9324 7108 9330 7172
rect 11329 7170 11395 7173
rect 12525 7170 12591 7173
rect 11329 7168 12591 7170
rect 11329 7112 11334 7168
rect 11390 7112 12530 7168
rect 12586 7112 12591 7168
rect 11329 7110 12591 7112
rect 11329 7107 11395 7110
rect 12525 7107 12591 7110
rect 5874 7104 6194 7105
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6194 7104
rect 5874 7039 6194 7040
rect 10805 7104 11125 7105
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 7039 11125 7040
rect 10133 7034 10199 7037
rect 10501 7034 10567 7037
rect 10133 7032 10567 7034
rect 10133 6976 10138 7032
rect 10194 6976 10506 7032
rect 10562 6976 10567 7032
rect 10133 6974 10567 6976
rect 10133 6971 10199 6974
rect 10501 6971 10567 6974
rect 11881 7034 11947 7037
rect 12617 7034 12683 7037
rect 11881 7032 12683 7034
rect 11881 6976 11886 7032
rect 11942 6976 12622 7032
rect 12678 6976 12683 7032
rect 11881 6974 12683 6976
rect 11881 6971 11947 6974
rect 12617 6971 12683 6974
rect 2589 6898 2655 6901
rect 5625 6898 5691 6901
rect 2589 6896 5691 6898
rect 2589 6840 2594 6896
rect 2650 6840 5630 6896
rect 5686 6840 5691 6896
rect 2589 6838 5691 6840
rect 2589 6835 2655 6838
rect 5625 6835 5691 6838
rect 9581 6898 9647 6901
rect 11881 6898 11947 6901
rect 9581 6896 11947 6898
rect 9581 6840 9586 6896
rect 9642 6840 11886 6896
rect 11942 6840 11947 6896
rect 9581 6838 11947 6840
rect 9581 6835 9647 6838
rect 11881 6835 11947 6838
rect 12249 6898 12315 6901
rect 12249 6896 12772 6898
rect 12249 6840 12254 6896
rect 12310 6840 12772 6896
rect 12249 6838 12772 6840
rect 12249 6835 12315 6838
rect 2497 6762 2563 6765
rect 6729 6762 6795 6765
rect 2497 6760 6795 6762
rect 2497 6704 2502 6760
rect 2558 6704 6734 6760
rect 6790 6704 6795 6760
rect 2497 6702 6795 6704
rect 2497 6699 2563 6702
rect 6729 6699 6795 6702
rect 7465 6762 7531 6765
rect 7465 6760 11162 6762
rect 7465 6704 7470 6760
rect 7526 6704 11162 6760
rect 7465 6702 11162 6704
rect 7465 6699 7531 6702
rect 9029 6626 9095 6629
rect 9397 6626 9463 6629
rect 9029 6624 9463 6626
rect 9029 6568 9034 6624
rect 9090 6568 9402 6624
rect 9458 6568 9463 6624
rect 9029 6566 9463 6568
rect 9029 6563 9095 6566
rect 9397 6563 9463 6566
rect 9949 6626 10015 6629
rect 10777 6626 10843 6629
rect 9949 6624 10843 6626
rect 9949 6568 9954 6624
rect 10010 6568 10782 6624
rect 10838 6568 10843 6624
rect 9949 6566 10843 6568
rect 11102 6626 11162 6702
rect 11278 6700 11284 6764
rect 11348 6762 11354 6764
rect 12525 6762 12591 6765
rect 11348 6760 12591 6762
rect 11348 6704 12530 6760
rect 12586 6704 12591 6760
rect 11348 6702 12591 6704
rect 12712 6762 12772 6838
rect 13118 6836 13124 6900
rect 13188 6898 13194 6900
rect 13721 6898 13787 6901
rect 13188 6896 13787 6898
rect 13188 6840 13726 6896
rect 13782 6840 13787 6896
rect 13188 6838 13787 6840
rect 13188 6836 13194 6838
rect 13721 6835 13787 6838
rect 13997 6762 14063 6765
rect 12712 6760 14063 6762
rect 12712 6704 14002 6760
rect 14058 6704 14063 6760
rect 12712 6702 14063 6704
rect 11348 6700 11354 6702
rect 12525 6699 12591 6702
rect 13997 6699 14063 6702
rect 11973 6626 12039 6629
rect 11102 6624 12039 6626
rect 11102 6568 11978 6624
rect 12034 6568 12039 6624
rect 11102 6566 12039 6568
rect 9949 6563 10015 6566
rect 10777 6563 10843 6566
rect 11973 6563 12039 6566
rect 3409 6560 3729 6561
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 6495 3729 6496
rect 8340 6560 8660 6561
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 6495 8660 6496
rect 13270 6560 13590 6561
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 6495 13590 6496
rect 5809 6490 5875 6493
rect 7649 6490 7715 6493
rect 5809 6488 7715 6490
rect 5809 6432 5814 6488
rect 5870 6432 7654 6488
rect 7710 6432 7715 6488
rect 5809 6430 7715 6432
rect 5809 6427 5875 6430
rect 7649 6427 7715 6430
rect 9213 6490 9279 6493
rect 12382 6490 12388 6492
rect 9213 6488 12388 6490
rect 9213 6432 9218 6488
rect 9274 6432 12388 6488
rect 9213 6430 12388 6432
rect 9213 6427 9279 6430
rect 12382 6428 12388 6430
rect 12452 6428 12458 6492
rect 3785 6354 3851 6357
rect 7005 6354 7071 6357
rect 3785 6352 7071 6354
rect 3785 6296 3790 6352
rect 3846 6296 7010 6352
rect 7066 6296 7071 6352
rect 3785 6294 7071 6296
rect 3785 6291 3851 6294
rect 7005 6291 7071 6294
rect 9029 6354 9095 6357
rect 15009 6354 15075 6357
rect 9029 6352 15075 6354
rect 9029 6296 9034 6352
rect 9090 6296 15014 6352
rect 15070 6296 15075 6352
rect 9029 6294 15075 6296
rect 9029 6291 9095 6294
rect 15009 6291 15075 6294
rect 0 6218 480 6248
rect 1209 6218 1275 6221
rect 0 6216 1275 6218
rect 0 6160 1214 6216
rect 1270 6160 1275 6216
rect 0 6158 1275 6160
rect 0 6128 480 6158
rect 1209 6155 1275 6158
rect 1853 6218 1919 6221
rect 12893 6218 12959 6221
rect 1853 6216 12959 6218
rect 1853 6160 1858 6216
rect 1914 6160 12898 6216
rect 12954 6160 12959 6216
rect 1853 6158 12959 6160
rect 1853 6155 1919 6158
rect 12893 6155 12959 6158
rect 3325 6082 3391 6085
rect 4102 6082 4108 6084
rect 3325 6080 4108 6082
rect 3325 6024 3330 6080
rect 3386 6024 4108 6080
rect 3325 6022 4108 6024
rect 3325 6019 3391 6022
rect 4102 6020 4108 6022
rect 4172 6020 4178 6084
rect 8201 6082 8267 6085
rect 8201 6080 9552 6082
rect 8201 6024 8206 6080
rect 8262 6024 9552 6080
rect 8201 6022 9552 6024
rect 8201 6019 8267 6022
rect 5874 6016 6194 6017
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6194 6016
rect 5874 5951 6194 5952
rect 6310 5884 6316 5948
rect 6380 5946 6386 5948
rect 9029 5946 9095 5949
rect 6380 5944 9095 5946
rect 6380 5888 9034 5944
rect 9090 5888 9095 5944
rect 6380 5886 9095 5888
rect 9492 5946 9552 6022
rect 9622 6020 9628 6084
rect 9692 6082 9698 6084
rect 10409 6082 10475 6085
rect 9692 6080 10475 6082
rect 9692 6024 10414 6080
rect 10470 6024 10475 6080
rect 9692 6022 10475 6024
rect 9692 6020 9698 6022
rect 10409 6019 10475 6022
rect 12341 6082 12407 6085
rect 13445 6082 13511 6085
rect 12341 6080 13511 6082
rect 12341 6024 12346 6080
rect 12402 6024 13450 6080
rect 13506 6024 13511 6080
rect 12341 6022 13511 6024
rect 12341 6019 12407 6022
rect 13445 6019 13511 6022
rect 10805 6016 11125 6017
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 5951 11125 5952
rect 10501 5946 10567 5949
rect 12985 5946 13051 5949
rect 9492 5944 10567 5946
rect 9492 5888 10506 5944
rect 10562 5888 10567 5944
rect 9492 5886 10567 5888
rect 6380 5884 6386 5886
rect 9029 5883 9095 5886
rect 10501 5883 10567 5886
rect 11286 5944 13051 5946
rect 11286 5888 12990 5944
rect 13046 5888 13051 5944
rect 11286 5886 13051 5888
rect 1853 5810 1919 5813
rect 4153 5810 4219 5813
rect 1853 5808 4219 5810
rect 1853 5752 1858 5808
rect 1914 5752 4158 5808
rect 4214 5752 4219 5808
rect 1853 5750 4219 5752
rect 1853 5747 1919 5750
rect 4153 5747 4219 5750
rect 4429 5810 4495 5813
rect 8150 5810 8156 5812
rect 4429 5808 8156 5810
rect 4429 5752 4434 5808
rect 4490 5752 8156 5808
rect 4429 5750 8156 5752
rect 4429 5747 4495 5750
rect 8150 5748 8156 5750
rect 8220 5748 8226 5812
rect 10869 5810 10935 5813
rect 11286 5810 11346 5886
rect 12985 5883 13051 5886
rect 13537 5946 13603 5949
rect 14038 5946 14044 5948
rect 13537 5944 14044 5946
rect 13537 5888 13542 5944
rect 13598 5888 14044 5944
rect 13537 5886 14044 5888
rect 13537 5883 13603 5886
rect 14038 5884 14044 5886
rect 14108 5884 14114 5948
rect 14733 5946 14799 5949
rect 16520 5946 17000 5976
rect 14733 5944 17000 5946
rect 14733 5888 14738 5944
rect 14794 5888 17000 5944
rect 14733 5886 17000 5888
rect 14733 5883 14799 5886
rect 16520 5856 17000 5886
rect 13169 5810 13235 5813
rect 8342 5750 10794 5810
rect 2773 5674 2839 5677
rect 5165 5674 5231 5677
rect 8342 5674 8402 5750
rect 2773 5672 3940 5674
rect 2773 5616 2778 5672
rect 2834 5616 3940 5672
rect 2773 5614 3940 5616
rect 2773 5611 2839 5614
rect 3880 5538 3940 5614
rect 5165 5672 8402 5674
rect 5165 5616 5170 5672
rect 5226 5616 8402 5672
rect 5165 5614 8402 5616
rect 9029 5674 9095 5677
rect 10358 5674 10364 5676
rect 9029 5672 10364 5674
rect 9029 5616 9034 5672
rect 9090 5616 10364 5672
rect 9029 5614 10364 5616
rect 5165 5611 5231 5614
rect 9029 5611 9095 5614
rect 10358 5612 10364 5614
rect 10428 5612 10434 5676
rect 10734 5674 10794 5750
rect 10869 5808 11346 5810
rect 10869 5752 10874 5808
rect 10930 5752 11346 5808
rect 10869 5750 11346 5752
rect 11424 5808 13235 5810
rect 11424 5752 13174 5808
rect 13230 5752 13235 5808
rect 11424 5750 13235 5752
rect 10869 5747 10935 5750
rect 11424 5674 11484 5750
rect 13169 5747 13235 5750
rect 10734 5614 11484 5674
rect 12065 5674 12131 5677
rect 12341 5674 12407 5677
rect 12065 5672 12407 5674
rect 12065 5616 12070 5672
rect 12126 5616 12346 5672
rect 12402 5616 12407 5672
rect 12065 5614 12407 5616
rect 12065 5611 12131 5614
rect 12341 5611 12407 5614
rect 12709 5674 12775 5677
rect 13629 5674 13695 5677
rect 12709 5672 13695 5674
rect 12709 5616 12714 5672
rect 12770 5616 13634 5672
rect 13690 5616 13695 5672
rect 12709 5614 13695 5616
rect 12709 5611 12775 5614
rect 13629 5611 13695 5614
rect 7925 5538 7991 5541
rect 8109 5538 8175 5541
rect 3880 5536 8175 5538
rect 3880 5480 7930 5536
rect 7986 5480 8114 5536
rect 8170 5480 8175 5536
rect 3880 5478 8175 5480
rect 7925 5475 7991 5478
rect 8109 5475 8175 5478
rect 9765 5538 9831 5541
rect 10225 5538 10291 5541
rect 10358 5538 10364 5540
rect 9765 5536 10364 5538
rect 9765 5480 9770 5536
rect 9826 5480 10230 5536
rect 10286 5480 10364 5536
rect 9765 5478 10364 5480
rect 9765 5475 9831 5478
rect 10225 5475 10291 5478
rect 10358 5476 10364 5478
rect 10428 5476 10434 5540
rect 10593 5538 10659 5541
rect 10777 5538 10843 5541
rect 13077 5538 13143 5541
rect 10593 5536 13143 5538
rect 10593 5480 10598 5536
rect 10654 5480 10782 5536
rect 10838 5480 13082 5536
rect 13138 5480 13143 5536
rect 10593 5478 13143 5480
rect 10593 5475 10659 5478
rect 10777 5475 10843 5478
rect 13077 5475 13143 5478
rect 3409 5472 3729 5473
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 5407 3729 5408
rect 8340 5472 8660 5473
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 5407 8660 5408
rect 13270 5472 13590 5473
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 5407 13590 5408
rect 7557 5402 7623 5405
rect 12617 5402 12683 5405
rect 7008 5400 7623 5402
rect 7008 5344 7562 5400
rect 7618 5344 7623 5400
rect 7008 5342 7623 5344
rect 0 5266 480 5296
rect 7008 5269 7068 5342
rect 7557 5339 7623 5342
rect 8894 5400 12683 5402
rect 8894 5344 12622 5400
rect 12678 5344 12683 5400
rect 8894 5342 12683 5344
rect 0 5206 1962 5266
rect 0 5176 480 5206
rect 1902 5130 1962 5206
rect 7005 5264 7071 5269
rect 7005 5208 7010 5264
rect 7066 5208 7071 5264
rect 7005 5203 7071 5208
rect 7782 5204 7788 5268
rect 7852 5266 7858 5268
rect 8477 5266 8543 5269
rect 7852 5264 8543 5266
rect 7852 5208 8482 5264
rect 8538 5208 8543 5264
rect 7852 5206 8543 5208
rect 7852 5204 7858 5206
rect 8477 5203 8543 5206
rect 2037 5130 2103 5133
rect 1902 5128 2103 5130
rect 1902 5072 2042 5128
rect 2098 5072 2103 5128
rect 1902 5070 2103 5072
rect 2037 5067 2103 5070
rect 4061 5130 4127 5133
rect 6637 5130 6703 5133
rect 4061 5128 6703 5130
rect 4061 5072 4066 5128
rect 4122 5072 6642 5128
rect 6698 5072 6703 5128
rect 4061 5070 6703 5072
rect 4061 5067 4127 5070
rect 6637 5067 6703 5070
rect 7649 5130 7715 5133
rect 8894 5130 8954 5342
rect 12617 5339 12683 5342
rect 9438 5204 9444 5268
rect 9508 5266 9514 5268
rect 11145 5266 11211 5269
rect 14641 5266 14707 5269
rect 9508 5264 11211 5266
rect 9508 5208 11150 5264
rect 11206 5208 11211 5264
rect 9508 5206 11211 5208
rect 9508 5204 9514 5206
rect 11145 5203 11211 5206
rect 11424 5264 14707 5266
rect 11424 5208 14646 5264
rect 14702 5208 14707 5264
rect 11424 5206 14707 5208
rect 9949 5130 10015 5133
rect 11424 5130 11484 5206
rect 14641 5203 14707 5206
rect 13721 5130 13787 5133
rect 7649 5128 8954 5130
rect 7649 5072 7654 5128
rect 7710 5072 8954 5128
rect 7649 5070 8954 5072
rect 9078 5128 10015 5130
rect 9078 5072 9954 5128
rect 10010 5072 10015 5128
rect 9078 5070 10015 5072
rect 7649 5067 7715 5070
rect 4286 4932 4292 4996
rect 4356 4994 4362 4996
rect 5349 4994 5415 4997
rect 4356 4992 5415 4994
rect 4356 4936 5354 4992
rect 5410 4936 5415 4992
rect 4356 4934 5415 4936
rect 4356 4932 4362 4934
rect 5349 4931 5415 4934
rect 6637 4994 6703 4997
rect 9078 4994 9138 5070
rect 9949 5067 10015 5070
rect 10596 5070 11484 5130
rect 11608 5128 13787 5130
rect 11608 5072 13726 5128
rect 13782 5072 13787 5128
rect 11608 5070 13787 5072
rect 10596 4994 10656 5070
rect 6637 4992 9138 4994
rect 6637 4936 6642 4992
rect 6698 4936 9138 4992
rect 6637 4934 9138 4936
rect 9216 4934 10656 4994
rect 6637 4931 6703 4934
rect 5874 4928 6194 4929
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6194 4928
rect 5874 4863 6194 4864
rect 3509 4858 3575 4861
rect 5717 4858 5783 4861
rect 3509 4856 5783 4858
rect 3509 4800 3514 4856
rect 3570 4800 5722 4856
rect 5778 4800 5783 4856
rect 3509 4798 5783 4800
rect 3509 4795 3575 4798
rect 5717 4795 5783 4798
rect 7046 4796 7052 4860
rect 7116 4858 7122 4860
rect 9216 4858 9276 4934
rect 11278 4932 11284 4996
rect 11348 4994 11354 4996
rect 11608 4994 11668 5070
rect 13721 5067 13787 5070
rect 11348 4934 11668 4994
rect 11348 4932 11354 4934
rect 12750 4932 12756 4996
rect 12820 4994 12826 4996
rect 13261 4994 13327 4997
rect 12820 4992 13327 4994
rect 12820 4936 13266 4992
rect 13322 4936 13327 4992
rect 12820 4934 13327 4936
rect 12820 4932 12826 4934
rect 13261 4931 13327 4934
rect 10805 4928 11125 4929
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 4863 11125 4864
rect 7116 4798 9276 4858
rect 7116 4796 7122 4798
rect 9438 4796 9444 4860
rect 9508 4858 9514 4860
rect 9765 4858 9831 4861
rect 9508 4856 9831 4858
rect 9508 4800 9770 4856
rect 9826 4800 9831 4856
rect 10174 4827 10180 4860
rect 10133 4824 10180 4827
rect 9508 4798 9831 4800
rect 9508 4796 9514 4798
rect 9765 4795 9831 4798
rect 10122 4822 10180 4824
rect 10122 4766 10138 4822
rect 10244 4796 10250 4860
rect 13445 4858 13511 4861
rect 14038 4858 14044 4860
rect 13445 4856 14044 4858
rect 13445 4800 13450 4856
rect 13506 4800 14044 4856
rect 13445 4798 14044 4800
rect 10194 4766 10242 4796
rect 13445 4795 13511 4798
rect 14038 4796 14044 4798
rect 14108 4796 14114 4860
rect 10122 4764 10242 4766
rect 10133 4761 10199 4764
rect 4613 4722 4679 4725
rect 4981 4722 5047 4725
rect 9990 4722 9996 4724
rect 4613 4720 9996 4722
rect 4613 4664 4618 4720
rect 4674 4664 4986 4720
rect 5042 4664 9996 4720
rect 4613 4662 9996 4664
rect 4613 4659 4679 4662
rect 4981 4659 5047 4662
rect 9990 4660 9996 4662
rect 10060 4660 10066 4724
rect 10317 4722 10383 4725
rect 15101 4722 15167 4725
rect 10317 4720 15167 4722
rect 10317 4664 10322 4720
rect 10378 4664 15106 4720
rect 15162 4664 15167 4720
rect 10317 4662 15167 4664
rect 10317 4659 10383 4662
rect 15101 4659 15167 4662
rect 2957 4586 3023 4589
rect 11053 4586 11119 4589
rect 2957 4584 11119 4586
rect 2957 4528 2962 4584
rect 3018 4528 11058 4584
rect 11114 4528 11119 4584
rect 2957 4526 11119 4528
rect 2957 4523 3023 4526
rect 11053 4523 11119 4526
rect 11237 4586 11303 4589
rect 11513 4586 11579 4589
rect 11237 4584 11579 4586
rect 11237 4528 11242 4584
rect 11298 4528 11518 4584
rect 11574 4528 11579 4584
rect 11237 4526 11579 4528
rect 11237 4523 11303 4526
rect 11513 4523 11579 4526
rect 11646 4524 11652 4588
rect 11716 4586 11722 4588
rect 12525 4586 12591 4589
rect 12709 4588 12775 4589
rect 12709 4586 12756 4588
rect 11716 4584 12591 4586
rect 11716 4528 12530 4584
rect 12586 4528 12591 4584
rect 11716 4526 12591 4528
rect 12664 4584 12756 4586
rect 12664 4528 12714 4584
rect 12664 4526 12756 4528
rect 11716 4524 11722 4526
rect 12525 4523 12591 4526
rect 12709 4524 12756 4526
rect 12820 4524 12826 4588
rect 15009 4586 15075 4589
rect 13126 4584 15075 4586
rect 13126 4528 15014 4584
rect 15070 4528 15075 4584
rect 13126 4526 15075 4528
rect 12709 4523 12775 4524
rect 5349 4450 5415 4453
rect 7005 4450 7071 4453
rect 5349 4448 7071 4450
rect 5349 4392 5354 4448
rect 5410 4392 7010 4448
rect 7066 4392 7071 4448
rect 5349 4390 7071 4392
rect 5349 4387 5415 4390
rect 7005 4387 7071 4390
rect 9254 4388 9260 4452
rect 9324 4450 9330 4452
rect 11278 4450 11284 4452
rect 9324 4390 11284 4450
rect 9324 4388 9330 4390
rect 11278 4388 11284 4390
rect 11348 4388 11354 4452
rect 11646 4388 11652 4452
rect 11716 4450 11722 4452
rect 11789 4450 11855 4453
rect 11716 4448 11855 4450
rect 11716 4392 11794 4448
rect 11850 4392 11855 4448
rect 11716 4390 11855 4392
rect 11716 4388 11722 4390
rect 11789 4387 11855 4390
rect 12014 4388 12020 4452
rect 12084 4450 12090 4452
rect 12709 4450 12775 4453
rect 12084 4448 12775 4450
rect 12084 4392 12714 4448
rect 12770 4392 12775 4448
rect 12084 4390 12775 4392
rect 12084 4388 12090 4390
rect 12709 4387 12775 4390
rect 3409 4384 3729 4385
rect 0 4314 480 4344
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 4319 3729 4320
rect 8340 4384 8660 4385
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 4319 8660 4320
rect 1117 4314 1183 4317
rect 0 4312 1183 4314
rect 0 4256 1122 4312
rect 1178 4256 1183 4312
rect 0 4254 1183 4256
rect 0 4224 480 4254
rect 1117 4251 1183 4254
rect 3969 4314 4035 4317
rect 4705 4314 4771 4317
rect 3969 4312 4771 4314
rect 3969 4256 3974 4312
rect 4030 4256 4710 4312
rect 4766 4256 4771 4312
rect 3969 4254 4771 4256
rect 3969 4251 4035 4254
rect 4705 4251 4771 4254
rect 5073 4314 5139 4317
rect 5809 4314 5875 4317
rect 5073 4312 5875 4314
rect 5073 4256 5078 4312
rect 5134 4256 5814 4312
rect 5870 4256 5875 4312
rect 5073 4254 5875 4256
rect 5073 4251 5139 4254
rect 5809 4251 5875 4254
rect 5993 4314 6059 4317
rect 7925 4314 7991 4317
rect 5993 4312 7991 4314
rect 5993 4256 5998 4312
rect 6054 4256 7930 4312
rect 7986 4256 7991 4312
rect 5993 4254 7991 4256
rect 5993 4251 6059 4254
rect 7925 4251 7991 4254
rect 8886 4252 8892 4316
rect 8956 4314 8962 4316
rect 13126 4314 13186 4526
rect 15009 4523 15075 4526
rect 13270 4384 13590 4385
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13270 4319 13590 4320
rect 8956 4254 13186 4314
rect 8956 4252 8962 4254
rect 4102 4116 4108 4180
rect 4172 4178 4178 4180
rect 7465 4178 7531 4181
rect 4172 4176 7531 4178
rect 4172 4120 7470 4176
rect 7526 4120 7531 4176
rect 4172 4118 7531 4120
rect 4172 4116 4178 4118
rect 7465 4115 7531 4118
rect 7598 4116 7604 4180
rect 7668 4178 7674 4180
rect 8293 4178 8359 4181
rect 7668 4176 8359 4178
rect 7668 4120 8298 4176
rect 8354 4120 8359 4176
rect 7668 4118 8359 4120
rect 7668 4116 7674 4118
rect 8293 4115 8359 4118
rect 9029 4178 9095 4181
rect 9581 4178 9647 4181
rect 9029 4176 9647 4178
rect 9029 4120 9034 4176
rect 9090 4120 9586 4176
rect 9642 4120 9647 4176
rect 9029 4118 9647 4120
rect 9029 4115 9095 4118
rect 9581 4115 9647 4118
rect 10358 4116 10364 4180
rect 10428 4178 10434 4180
rect 10428 4118 12128 4178
rect 10428 4116 10434 4118
rect 2681 4042 2747 4045
rect 11881 4044 11947 4045
rect 2681 4040 11346 4042
rect 2681 3984 2686 4040
rect 2742 3984 11346 4040
rect 2681 3982 11346 3984
rect 2681 3979 2747 3982
rect 6361 3906 6427 3909
rect 6637 3906 6703 3909
rect 6821 3908 6887 3909
rect 6821 3906 6868 3908
rect 6361 3904 6703 3906
rect 6361 3848 6366 3904
rect 6422 3848 6642 3904
rect 6698 3848 6703 3904
rect 6361 3846 6703 3848
rect 6776 3904 6868 3906
rect 6776 3848 6826 3904
rect 6776 3846 6868 3848
rect 6361 3843 6427 3846
rect 6637 3843 6703 3846
rect 6821 3844 6868 3846
rect 6932 3844 6938 3908
rect 7005 3906 7071 3909
rect 10041 3906 10107 3909
rect 7005 3904 10107 3906
rect 7005 3848 7010 3904
rect 7066 3848 10046 3904
rect 10102 3848 10107 3904
rect 7005 3846 10107 3848
rect 6821 3843 6887 3844
rect 7005 3843 7071 3846
rect 10041 3843 10107 3846
rect 10358 3844 10364 3908
rect 10428 3906 10434 3908
rect 10593 3906 10659 3909
rect 10428 3904 10659 3906
rect 10428 3848 10598 3904
rect 10654 3848 10659 3904
rect 10428 3846 10659 3848
rect 11286 3906 11346 3982
rect 11830 3980 11836 4044
rect 11900 4042 11947 4044
rect 12068 4042 12128 4118
rect 12566 4116 12572 4180
rect 12636 4178 12642 4180
rect 12709 4178 12775 4181
rect 12636 4176 12775 4178
rect 12636 4120 12714 4176
rect 12770 4120 12775 4176
rect 12636 4118 12775 4120
rect 12636 4116 12642 4118
rect 12709 4115 12775 4118
rect 13118 4116 13124 4180
rect 13188 4178 13194 4180
rect 13629 4178 13695 4181
rect 13188 4176 13695 4178
rect 13188 4120 13634 4176
rect 13690 4120 13695 4176
rect 13188 4118 13695 4120
rect 13188 4116 13194 4118
rect 13629 4115 13695 4118
rect 14457 4042 14523 4045
rect 11900 4040 11992 4042
rect 11942 3984 11992 4040
rect 11900 3982 11992 3984
rect 12068 4040 14523 4042
rect 12068 3984 14462 4040
rect 14518 3984 14523 4040
rect 12068 3982 14523 3984
rect 11900 3980 11947 3982
rect 11881 3979 11947 3980
rect 14457 3979 14523 3982
rect 14641 3906 14707 3909
rect 11286 3904 14707 3906
rect 11286 3848 14646 3904
rect 14702 3848 14707 3904
rect 11286 3846 14707 3848
rect 10428 3844 10434 3846
rect 10593 3843 10659 3846
rect 14641 3843 14707 3846
rect 5874 3840 6194 3841
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6194 3840
rect 5874 3775 6194 3776
rect 10805 3840 11125 3841
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10805 3775 11125 3776
rect 3601 3770 3667 3773
rect 5390 3770 5396 3772
rect 3601 3768 5396 3770
rect 3601 3712 3606 3768
rect 3662 3712 5396 3768
rect 3601 3710 5396 3712
rect 3601 3707 3667 3710
rect 5390 3708 5396 3710
rect 5460 3708 5466 3772
rect 6637 3770 6703 3773
rect 10225 3770 10291 3773
rect 10593 3770 10659 3773
rect 6637 3768 10104 3770
rect 6637 3712 6642 3768
rect 6698 3712 10104 3768
rect 6637 3710 10104 3712
rect 6637 3707 6703 3710
rect 3233 3634 3299 3637
rect 4470 3634 4476 3636
rect 3233 3632 4476 3634
rect 3233 3576 3238 3632
rect 3294 3576 4476 3632
rect 3233 3574 4476 3576
rect 3233 3571 3299 3574
rect 4470 3572 4476 3574
rect 4540 3572 4546 3636
rect 4797 3634 4863 3637
rect 9765 3634 9831 3637
rect 4797 3632 9831 3634
rect 4797 3576 4802 3632
rect 4858 3576 9770 3632
rect 9826 3576 9831 3632
rect 4797 3574 9831 3576
rect 10044 3634 10104 3710
rect 10225 3768 10659 3770
rect 10225 3712 10230 3768
rect 10286 3712 10598 3768
rect 10654 3712 10659 3768
rect 10225 3710 10659 3712
rect 10225 3707 10291 3710
rect 10593 3707 10659 3710
rect 11421 3770 11487 3773
rect 12157 3770 12223 3773
rect 11421 3768 12223 3770
rect 11421 3712 11426 3768
rect 11482 3712 12162 3768
rect 12218 3712 12223 3768
rect 11421 3710 12223 3712
rect 11421 3707 11487 3710
rect 12157 3707 12223 3710
rect 11830 3634 11836 3636
rect 10044 3574 11836 3634
rect 4797 3571 4863 3574
rect 9765 3571 9831 3574
rect 11830 3572 11836 3574
rect 11900 3572 11906 3636
rect 12014 3572 12020 3636
rect 12084 3634 12090 3636
rect 12617 3634 12683 3637
rect 12084 3632 12683 3634
rect 12084 3576 12622 3632
rect 12678 3576 12683 3632
rect 12084 3574 12683 3576
rect 12084 3572 12090 3574
rect 12617 3571 12683 3574
rect 12750 3572 12756 3636
rect 12820 3634 12826 3636
rect 13261 3634 13327 3637
rect 13854 3634 13860 3636
rect 12820 3632 13860 3634
rect 12820 3576 13266 3632
rect 13322 3576 13860 3632
rect 12820 3574 13860 3576
rect 12820 3572 12826 3574
rect 13261 3571 13327 3574
rect 13854 3572 13860 3574
rect 13924 3572 13930 3636
rect 1025 3498 1091 3501
rect 8477 3498 8543 3501
rect 9121 3500 9187 3501
rect 1025 3496 8543 3498
rect 1025 3440 1030 3496
rect 1086 3440 8482 3496
rect 8538 3440 8543 3496
rect 1025 3438 8543 3440
rect 1025 3435 1091 3438
rect 8477 3435 8543 3438
rect 9070 3436 9076 3500
rect 9140 3498 9187 3500
rect 9397 3498 9463 3501
rect 13813 3498 13879 3501
rect 9140 3496 9232 3498
rect 9182 3440 9232 3496
rect 9140 3438 9232 3440
rect 9397 3496 9736 3498
rect 9397 3440 9402 3496
rect 9458 3464 9736 3496
rect 9814 3496 13879 3498
rect 9814 3464 13818 3496
rect 9458 3440 13818 3464
rect 13874 3440 13879 3496
rect 9397 3438 13879 3440
rect 9140 3436 9187 3438
rect 9121 3435 9187 3436
rect 9397 3435 9463 3438
rect 9676 3404 9874 3438
rect 13813 3435 13879 3438
rect 0 3362 480 3392
rect 3049 3362 3115 3365
rect 0 3360 3115 3362
rect 0 3304 3054 3360
rect 3110 3304 3115 3360
rect 0 3302 3115 3304
rect 0 3272 480 3302
rect 3049 3299 3115 3302
rect 3969 3362 4035 3365
rect 6085 3362 6151 3365
rect 6913 3362 6979 3365
rect 3969 3360 6979 3362
rect 3969 3304 3974 3360
rect 4030 3304 6090 3360
rect 6146 3304 6918 3360
rect 6974 3304 6979 3360
rect 3969 3302 6979 3304
rect 3969 3299 4035 3302
rect 6085 3299 6151 3302
rect 6913 3299 6979 3302
rect 10593 3362 10659 3365
rect 11513 3362 11579 3365
rect 11881 3364 11947 3365
rect 11830 3362 11836 3364
rect 10593 3360 11579 3362
rect 10593 3304 10598 3360
rect 10654 3304 11518 3360
rect 11574 3304 11579 3360
rect 10593 3302 11579 3304
rect 11790 3302 11836 3362
rect 11900 3360 11947 3364
rect 11942 3304 11947 3360
rect 10593 3299 10659 3302
rect 11513 3299 11579 3302
rect 11830 3300 11836 3302
rect 11900 3300 11947 3304
rect 11881 3299 11947 3300
rect 3409 3296 3729 3297
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 3231 3729 3232
rect 8340 3296 8660 3297
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 3231 8660 3232
rect 13270 3296 13590 3297
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 13270 3231 13590 3232
rect 5441 3226 5507 3229
rect 7189 3226 7255 3229
rect 5441 3224 7255 3226
rect 5441 3168 5446 3224
rect 5502 3168 7194 3224
rect 7250 3168 7255 3224
rect 5441 3166 7255 3168
rect 5441 3163 5507 3166
rect 7189 3163 7255 3166
rect 7373 3226 7439 3229
rect 7925 3226 7991 3229
rect 7373 3224 7991 3226
rect 7373 3168 7378 3224
rect 7434 3168 7930 3224
rect 7986 3168 7991 3224
rect 7373 3166 7991 3168
rect 7373 3163 7439 3166
rect 7925 3163 7991 3166
rect 8894 3166 12772 3226
rect 3049 3090 3115 3093
rect 8894 3090 8954 3166
rect 3049 3088 8954 3090
rect 3049 3032 3054 3088
rect 3110 3032 8954 3088
rect 3049 3030 8954 3032
rect 3049 3027 3115 3030
rect 9622 3028 9628 3092
rect 9692 3090 9698 3092
rect 10225 3090 10291 3093
rect 9692 3088 10291 3090
rect 9692 3032 10230 3088
rect 10286 3032 10291 3088
rect 9692 3030 10291 3032
rect 9692 3028 9698 3030
rect 10225 3027 10291 3030
rect 10869 3090 10935 3093
rect 11697 3090 11763 3093
rect 10869 3088 11763 3090
rect 10869 3032 10874 3088
rect 10930 3032 11702 3088
rect 11758 3032 11763 3088
rect 10869 3030 11763 3032
rect 10869 3027 10935 3030
rect 11697 3027 11763 3030
rect 12382 3028 12388 3092
rect 12452 3090 12458 3092
rect 12525 3090 12591 3093
rect 12452 3088 12591 3090
rect 12452 3032 12530 3088
rect 12586 3032 12591 3088
rect 12452 3030 12591 3032
rect 12712 3090 12772 3166
rect 15009 3090 15075 3093
rect 12712 3088 15075 3090
rect 12712 3032 15014 3088
rect 15070 3032 15075 3088
rect 12712 3030 15075 3032
rect 12452 3028 12458 3030
rect 12525 3027 12591 3030
rect 15009 3027 15075 3030
rect 3182 2892 3188 2956
rect 3252 2954 3258 2956
rect 3417 2954 3483 2957
rect 4245 2956 4311 2957
rect 4245 2954 4292 2956
rect 3252 2952 3483 2954
rect 3252 2896 3422 2952
rect 3478 2896 3483 2952
rect 3252 2894 3483 2896
rect 4200 2952 4292 2954
rect 4200 2896 4250 2952
rect 4200 2894 4292 2896
rect 3252 2892 3258 2894
rect 3417 2891 3483 2894
rect 4245 2892 4292 2894
rect 4356 2892 4362 2956
rect 5349 2954 5415 2957
rect 7833 2956 7899 2957
rect 7598 2954 7604 2956
rect 5349 2952 7604 2954
rect 5349 2896 5354 2952
rect 5410 2896 7604 2952
rect 5349 2894 7604 2896
rect 4245 2891 4311 2892
rect 5349 2891 5415 2894
rect 7598 2892 7604 2894
rect 7668 2892 7674 2956
rect 7782 2892 7788 2956
rect 7852 2954 7899 2956
rect 8017 2954 8083 2957
rect 8569 2954 8635 2957
rect 14733 2954 14799 2957
rect 7852 2952 7944 2954
rect 7894 2896 7944 2952
rect 7852 2894 7944 2896
rect 8017 2952 8635 2954
rect 8017 2896 8022 2952
rect 8078 2896 8574 2952
rect 8630 2896 8635 2952
rect 8017 2894 8635 2896
rect 7852 2892 7899 2894
rect 7833 2891 7899 2892
rect 8017 2891 8083 2894
rect 8569 2891 8635 2894
rect 9676 2952 14799 2954
rect 9676 2896 14738 2952
rect 14794 2896 14799 2952
rect 9676 2894 14799 2896
rect 4337 2818 4403 2821
rect 5717 2818 5783 2821
rect 4337 2816 5783 2818
rect 4337 2760 4342 2816
rect 4398 2760 5722 2816
rect 5778 2760 5783 2816
rect 4337 2758 5783 2760
rect 4337 2755 4403 2758
rect 5717 2755 5783 2758
rect 6678 2756 6684 2820
rect 6748 2818 6754 2820
rect 7189 2818 7255 2821
rect 6748 2816 7255 2818
rect 6748 2760 7194 2816
rect 7250 2760 7255 2816
rect 6748 2758 7255 2760
rect 6748 2756 6754 2758
rect 7189 2755 7255 2758
rect 7557 2818 7623 2821
rect 9676 2818 9736 2894
rect 14733 2891 14799 2894
rect 7557 2816 9736 2818
rect 7557 2760 7562 2816
rect 7618 2760 9736 2816
rect 7557 2758 9736 2760
rect 7557 2755 7623 2758
rect 9806 2756 9812 2820
rect 9876 2818 9882 2820
rect 10593 2818 10659 2821
rect 9876 2816 10659 2818
rect 9876 2760 10598 2816
rect 10654 2760 10659 2816
rect 9876 2758 10659 2760
rect 9876 2756 9882 2758
rect 10593 2755 10659 2758
rect 11513 2818 11579 2821
rect 12198 2818 12204 2820
rect 11513 2816 12204 2818
rect 11513 2760 11518 2816
rect 11574 2760 12204 2816
rect 11513 2758 12204 2760
rect 11513 2755 11579 2758
rect 12198 2756 12204 2758
rect 12268 2818 12274 2820
rect 14825 2818 14891 2821
rect 12268 2816 14891 2818
rect 12268 2760 14830 2816
rect 14886 2760 14891 2816
rect 12268 2758 14891 2760
rect 12268 2756 12274 2758
rect 14825 2755 14891 2758
rect 5874 2752 6194 2753
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6194 2752
rect 5874 2687 6194 2688
rect 10805 2752 11125 2753
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10805 2687 11125 2688
rect 2865 2682 2931 2685
rect 4654 2682 4660 2684
rect 2865 2680 4660 2682
rect 2865 2624 2870 2680
rect 2926 2624 4660 2680
rect 2865 2622 4660 2624
rect 2865 2619 2931 2622
rect 4654 2620 4660 2622
rect 4724 2620 4730 2684
rect 7925 2682 7991 2685
rect 10041 2684 10107 2685
rect 9806 2682 9812 2684
rect 7925 2680 9812 2682
rect 7925 2624 7930 2680
rect 7986 2624 9812 2680
rect 7925 2622 9812 2624
rect 7925 2619 7991 2622
rect 9806 2620 9812 2622
rect 9876 2620 9882 2684
rect 9990 2682 9996 2684
rect 9950 2622 9996 2682
rect 10060 2680 10107 2684
rect 10102 2624 10107 2680
rect 9990 2620 9996 2622
rect 10060 2620 10107 2624
rect 10174 2620 10180 2684
rect 10244 2682 10250 2684
rect 10317 2682 10383 2685
rect 10244 2680 10383 2682
rect 10244 2624 10322 2680
rect 10378 2624 10383 2680
rect 10244 2622 10383 2624
rect 10244 2620 10250 2622
rect 10041 2619 10107 2620
rect 10317 2619 10383 2622
rect 11237 2682 11303 2685
rect 15561 2682 15627 2685
rect 11237 2680 15627 2682
rect 11237 2624 11242 2680
rect 11298 2624 15566 2680
rect 15622 2624 15627 2680
rect 11237 2622 15627 2624
rect 11237 2619 11303 2622
rect 15561 2619 15627 2622
rect 1669 2546 1735 2549
rect 5441 2546 5507 2549
rect 1669 2544 5507 2546
rect 1669 2488 1674 2544
rect 1730 2488 5446 2544
rect 5502 2488 5507 2544
rect 1669 2486 5507 2488
rect 1669 2483 1735 2486
rect 5441 2483 5507 2486
rect 5625 2546 5691 2549
rect 6310 2546 6316 2548
rect 5625 2544 6316 2546
rect 5625 2488 5630 2544
rect 5686 2488 6316 2544
rect 5625 2486 6316 2488
rect 5625 2483 5691 2486
rect 6310 2484 6316 2486
rect 6380 2484 6386 2548
rect 6453 2546 6519 2549
rect 7465 2548 7531 2549
rect 8017 2548 8083 2549
rect 7230 2546 7236 2548
rect 6453 2544 7236 2546
rect 6453 2488 6458 2544
rect 6514 2488 7236 2544
rect 6453 2486 7236 2488
rect 6453 2483 6519 2486
rect 7230 2484 7236 2486
rect 7300 2484 7306 2548
rect 7414 2484 7420 2548
rect 7484 2546 7531 2548
rect 7484 2544 7576 2546
rect 7526 2488 7576 2544
rect 7484 2486 7576 2488
rect 7484 2484 7531 2486
rect 7966 2484 7972 2548
rect 8036 2546 8083 2548
rect 8477 2546 8543 2549
rect 10133 2546 10199 2549
rect 11462 2546 11468 2548
rect 8036 2544 8128 2546
rect 8078 2488 8128 2544
rect 8036 2486 8128 2488
rect 8477 2544 11468 2546
rect 8477 2488 8482 2544
rect 8538 2488 10138 2544
rect 10194 2488 11468 2544
rect 8477 2486 11468 2488
rect 8036 2484 8083 2486
rect 7465 2483 7531 2484
rect 8017 2483 8083 2484
rect 8477 2483 8543 2486
rect 10133 2483 10199 2486
rect 11462 2484 11468 2486
rect 11532 2484 11538 2548
rect 11697 2546 11763 2549
rect 13721 2546 13787 2549
rect 11697 2544 13787 2546
rect 11697 2488 11702 2544
rect 11758 2488 13726 2544
rect 13782 2488 13787 2544
rect 11697 2486 13787 2488
rect 11697 2483 11763 2486
rect 13721 2483 13787 2486
rect 0 2410 480 2440
rect 4797 2410 4863 2413
rect 7097 2410 7163 2413
rect 0 2350 3986 2410
rect 0 2320 480 2350
rect 3926 2274 3986 2350
rect 4797 2408 7163 2410
rect 4797 2352 4802 2408
rect 4858 2352 7102 2408
rect 7158 2352 7163 2408
rect 4797 2350 7163 2352
rect 4797 2347 4863 2350
rect 7097 2347 7163 2350
rect 9949 2410 10015 2413
rect 12433 2410 12499 2413
rect 9949 2408 12499 2410
rect 9949 2352 9954 2408
rect 10010 2352 12438 2408
rect 12494 2352 12499 2408
rect 9949 2350 12499 2352
rect 9949 2347 10015 2350
rect 12433 2347 12499 2350
rect 12985 2410 13051 2413
rect 13118 2410 13124 2412
rect 12985 2408 13124 2410
rect 12985 2352 12990 2408
rect 13046 2352 13124 2408
rect 12985 2350 13124 2352
rect 12985 2347 13051 2350
rect 13118 2348 13124 2350
rect 13188 2348 13194 2412
rect 6494 2274 6500 2276
rect 3926 2214 6500 2274
rect 6494 2212 6500 2214
rect 6564 2274 6570 2276
rect 6729 2274 6795 2277
rect 6564 2272 6795 2274
rect 6564 2216 6734 2272
rect 6790 2216 6795 2272
rect 6564 2214 6795 2216
rect 6564 2212 6570 2214
rect 6729 2211 6795 2214
rect 10409 2274 10475 2277
rect 12566 2274 12572 2276
rect 10409 2272 12572 2274
rect 10409 2216 10414 2272
rect 10470 2216 12572 2272
rect 10409 2214 12572 2216
rect 10409 2211 10475 2214
rect 12566 2212 12572 2214
rect 12636 2212 12642 2276
rect 3409 2208 3729 2209
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2143 3729 2144
rect 8340 2208 8660 2209
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2143 8660 2144
rect 13270 2208 13590 2209
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2143 13590 2144
rect 4981 2138 5047 2141
rect 7833 2138 7899 2141
rect 4981 2136 7899 2138
rect 4981 2080 4986 2136
rect 5042 2080 7838 2136
rect 7894 2080 7899 2136
rect 4981 2078 7899 2080
rect 4981 2075 5047 2078
rect 7833 2075 7899 2078
rect 9489 2138 9555 2141
rect 11646 2138 11652 2140
rect 9489 2136 11652 2138
rect 9489 2080 9494 2136
rect 9550 2080 11652 2136
rect 9489 2078 11652 2080
rect 9489 2075 9555 2078
rect 11646 2076 11652 2078
rect 11716 2076 11722 2140
rect 1209 2002 1275 2005
rect 7925 2002 7991 2005
rect 1209 2000 7991 2002
rect 1209 1944 1214 2000
rect 1270 1944 7930 2000
rect 7986 1944 7991 2000
rect 1209 1942 7991 1944
rect 1209 1939 1275 1942
rect 7925 1939 7991 1942
rect 8150 1940 8156 2004
rect 8220 2002 8226 2004
rect 11881 2002 11947 2005
rect 8220 2000 11947 2002
rect 8220 1944 11886 2000
rect 11942 1944 11947 2000
rect 8220 1942 11947 1944
rect 8220 1940 8226 1942
rect 11881 1939 11947 1942
rect 12893 2002 12959 2005
rect 16520 2002 17000 2032
rect 12893 2000 17000 2002
rect 12893 1944 12898 2000
rect 12954 1944 17000 2000
rect 12893 1942 17000 1944
rect 12893 1939 12959 1942
rect 16520 1912 17000 1942
rect 4061 1866 4127 1869
rect 13670 1866 13676 1868
rect 4061 1864 13676 1866
rect 4061 1808 4066 1864
rect 4122 1808 13676 1864
rect 4061 1806 13676 1808
rect 4061 1803 4127 1806
rect 13670 1804 13676 1806
rect 13740 1804 13746 1868
rect 3877 1730 3943 1733
rect 8886 1730 8892 1732
rect 3877 1728 8892 1730
rect 3877 1672 3882 1728
rect 3938 1672 8892 1728
rect 3877 1670 8892 1672
rect 3877 1667 3943 1670
rect 8886 1668 8892 1670
rect 8956 1668 8962 1732
rect 3509 1594 3575 1597
rect 7046 1594 7052 1596
rect 3509 1592 7052 1594
rect 3509 1536 3514 1592
rect 3570 1536 7052 1592
rect 3509 1534 7052 1536
rect 3509 1531 3575 1534
rect 7046 1532 7052 1534
rect 7116 1532 7122 1596
rect 7598 1532 7604 1596
rect 7668 1594 7674 1596
rect 14549 1594 14615 1597
rect 7668 1592 14615 1594
rect 7668 1536 14554 1592
rect 14610 1536 14615 1592
rect 7668 1534 14615 1536
rect 7668 1532 7674 1534
rect 14549 1531 14615 1534
rect 0 1458 480 1488
rect 2773 1458 2839 1461
rect 0 1456 2839 1458
rect 0 1400 2778 1456
rect 2834 1400 2839 1456
rect 0 1398 2839 1400
rect 0 1368 480 1398
rect 2773 1395 2839 1398
rect 3233 1458 3299 1461
rect 10542 1458 10548 1460
rect 3233 1456 10548 1458
rect 3233 1400 3238 1456
rect 3294 1400 10548 1456
rect 3233 1398 10548 1400
rect 3233 1395 3299 1398
rect 10542 1396 10548 1398
rect 10612 1396 10618 1460
rect 12617 1458 12683 1461
rect 14038 1458 14044 1460
rect 12617 1456 14044 1458
rect 12617 1400 12622 1456
rect 12678 1400 14044 1456
rect 12617 1398 14044 1400
rect 12617 1395 12683 1398
rect 14038 1396 14044 1398
rect 14108 1396 14114 1460
rect 8477 1322 8543 1325
rect 12750 1322 12756 1324
rect 8477 1320 12756 1322
rect 8477 1264 8482 1320
rect 8538 1264 12756 1320
rect 8477 1262 12756 1264
rect 8477 1259 8543 1262
rect 12750 1260 12756 1262
rect 12820 1260 12826 1324
rect 12934 1260 12940 1324
rect 13004 1322 13010 1324
rect 13445 1322 13511 1325
rect 13004 1320 13511 1322
rect 13004 1264 13450 1320
rect 13506 1264 13511 1320
rect 13004 1262 13511 1264
rect 13004 1260 13010 1262
rect 13445 1259 13511 1262
rect 4337 1186 4403 1189
rect 9438 1186 9444 1188
rect 4337 1184 9444 1186
rect 4337 1128 4342 1184
rect 4398 1128 9444 1184
rect 4337 1126 9444 1128
rect 4337 1123 4403 1126
rect 9438 1124 9444 1126
rect 9508 1124 9514 1188
rect 0 506 480 536
rect 3141 506 3207 509
rect 0 504 3207 506
rect 0 448 3146 504
rect 3202 448 3207 504
rect 0 446 3207 448
rect 0 416 480 446
rect 3141 443 3207 446
<< via3 >>
rect 3417 17436 3481 17440
rect 3417 17380 3421 17436
rect 3421 17380 3477 17436
rect 3477 17380 3481 17436
rect 3417 17376 3481 17380
rect 3497 17436 3561 17440
rect 3497 17380 3501 17436
rect 3501 17380 3557 17436
rect 3557 17380 3561 17436
rect 3497 17376 3561 17380
rect 3577 17436 3641 17440
rect 3577 17380 3581 17436
rect 3581 17380 3637 17436
rect 3637 17380 3641 17436
rect 3577 17376 3641 17380
rect 3657 17436 3721 17440
rect 3657 17380 3661 17436
rect 3661 17380 3717 17436
rect 3717 17380 3721 17436
rect 3657 17376 3721 17380
rect 8348 17436 8412 17440
rect 8348 17380 8352 17436
rect 8352 17380 8408 17436
rect 8408 17380 8412 17436
rect 8348 17376 8412 17380
rect 8428 17436 8492 17440
rect 8428 17380 8432 17436
rect 8432 17380 8488 17436
rect 8488 17380 8492 17436
rect 8428 17376 8492 17380
rect 8508 17436 8572 17440
rect 8508 17380 8512 17436
rect 8512 17380 8568 17436
rect 8568 17380 8572 17436
rect 8508 17376 8572 17380
rect 8588 17436 8652 17440
rect 8588 17380 8592 17436
rect 8592 17380 8648 17436
rect 8648 17380 8652 17436
rect 8588 17376 8652 17380
rect 13278 17436 13342 17440
rect 13278 17380 13282 17436
rect 13282 17380 13338 17436
rect 13338 17380 13342 17436
rect 13278 17376 13342 17380
rect 13358 17436 13422 17440
rect 13358 17380 13362 17436
rect 13362 17380 13418 17436
rect 13418 17380 13422 17436
rect 13358 17376 13422 17380
rect 13438 17436 13502 17440
rect 13438 17380 13442 17436
rect 13442 17380 13498 17436
rect 13498 17380 13502 17436
rect 13438 17376 13502 17380
rect 13518 17436 13582 17440
rect 13518 17380 13522 17436
rect 13522 17380 13578 17436
rect 13578 17380 13582 17436
rect 13518 17376 13582 17380
rect 12756 17036 12820 17100
rect 12204 16900 12268 16964
rect 5882 16892 5946 16896
rect 5882 16836 5886 16892
rect 5886 16836 5942 16892
rect 5942 16836 5946 16892
rect 5882 16832 5946 16836
rect 5962 16892 6026 16896
rect 5962 16836 5966 16892
rect 5966 16836 6022 16892
rect 6022 16836 6026 16892
rect 5962 16832 6026 16836
rect 6042 16892 6106 16896
rect 6042 16836 6046 16892
rect 6046 16836 6102 16892
rect 6102 16836 6106 16892
rect 6042 16832 6106 16836
rect 6122 16892 6186 16896
rect 6122 16836 6126 16892
rect 6126 16836 6182 16892
rect 6182 16836 6186 16892
rect 6122 16832 6186 16836
rect 10813 16892 10877 16896
rect 10813 16836 10817 16892
rect 10817 16836 10873 16892
rect 10873 16836 10877 16892
rect 10813 16832 10877 16836
rect 10893 16892 10957 16896
rect 10893 16836 10897 16892
rect 10897 16836 10953 16892
rect 10953 16836 10957 16892
rect 10893 16832 10957 16836
rect 10973 16892 11037 16896
rect 10973 16836 10977 16892
rect 10977 16836 11033 16892
rect 11033 16836 11037 16892
rect 10973 16832 11037 16836
rect 11053 16892 11117 16896
rect 11053 16836 11057 16892
rect 11057 16836 11113 16892
rect 11113 16836 11117 16892
rect 11053 16832 11117 16836
rect 5028 16764 5092 16828
rect 9260 16628 9324 16692
rect 13124 16628 13188 16692
rect 12756 16492 12820 16556
rect 4292 16416 4356 16420
rect 4292 16360 4342 16416
rect 4342 16360 4356 16416
rect 4292 16356 4356 16360
rect 7788 16356 7852 16420
rect 11468 16356 11532 16420
rect 3417 16348 3481 16352
rect 3417 16292 3421 16348
rect 3421 16292 3477 16348
rect 3477 16292 3481 16348
rect 3417 16288 3481 16292
rect 3497 16348 3561 16352
rect 3497 16292 3501 16348
rect 3501 16292 3557 16348
rect 3557 16292 3561 16348
rect 3497 16288 3561 16292
rect 3577 16348 3641 16352
rect 3577 16292 3581 16348
rect 3581 16292 3637 16348
rect 3637 16292 3641 16348
rect 3577 16288 3641 16292
rect 3657 16348 3721 16352
rect 3657 16292 3661 16348
rect 3661 16292 3717 16348
rect 3717 16292 3721 16348
rect 3657 16288 3721 16292
rect 8348 16348 8412 16352
rect 8348 16292 8352 16348
rect 8352 16292 8408 16348
rect 8408 16292 8412 16348
rect 8348 16288 8412 16292
rect 8428 16348 8492 16352
rect 8428 16292 8432 16348
rect 8432 16292 8488 16348
rect 8488 16292 8492 16348
rect 8428 16288 8492 16292
rect 8508 16348 8572 16352
rect 8508 16292 8512 16348
rect 8512 16292 8568 16348
rect 8568 16292 8572 16348
rect 8508 16288 8572 16292
rect 8588 16348 8652 16352
rect 8588 16292 8592 16348
rect 8592 16292 8648 16348
rect 8648 16292 8652 16348
rect 8588 16288 8652 16292
rect 13278 16348 13342 16352
rect 13278 16292 13282 16348
rect 13282 16292 13338 16348
rect 13338 16292 13342 16348
rect 13278 16288 13342 16292
rect 13358 16348 13422 16352
rect 13358 16292 13362 16348
rect 13362 16292 13418 16348
rect 13418 16292 13422 16348
rect 13358 16288 13422 16292
rect 13438 16348 13502 16352
rect 13438 16292 13442 16348
rect 13442 16292 13498 16348
rect 13498 16292 13502 16348
rect 13438 16288 13502 16292
rect 13518 16348 13582 16352
rect 13518 16292 13522 16348
rect 13522 16292 13578 16348
rect 13578 16292 13582 16348
rect 13518 16288 13582 16292
rect 7604 16220 7668 16284
rect 3004 15812 3068 15876
rect 9444 15872 9508 15876
rect 9444 15816 9458 15872
rect 9458 15816 9508 15872
rect 9444 15812 9508 15816
rect 10180 15812 10244 15876
rect 5882 15804 5946 15808
rect 5882 15748 5886 15804
rect 5886 15748 5942 15804
rect 5942 15748 5946 15804
rect 5882 15744 5946 15748
rect 5962 15804 6026 15808
rect 5962 15748 5966 15804
rect 5966 15748 6022 15804
rect 6022 15748 6026 15804
rect 5962 15744 6026 15748
rect 6042 15804 6106 15808
rect 6042 15748 6046 15804
rect 6046 15748 6102 15804
rect 6102 15748 6106 15804
rect 6042 15744 6106 15748
rect 6122 15804 6186 15808
rect 6122 15748 6126 15804
rect 6126 15748 6182 15804
rect 6182 15748 6186 15804
rect 6122 15744 6186 15748
rect 10813 15804 10877 15808
rect 10813 15748 10817 15804
rect 10817 15748 10873 15804
rect 10873 15748 10877 15804
rect 10813 15744 10877 15748
rect 10893 15804 10957 15808
rect 10893 15748 10897 15804
rect 10897 15748 10953 15804
rect 10953 15748 10957 15804
rect 10893 15744 10957 15748
rect 10973 15804 11037 15808
rect 10973 15748 10977 15804
rect 10977 15748 11033 15804
rect 11033 15748 11037 15804
rect 10973 15744 11037 15748
rect 11053 15804 11117 15808
rect 11053 15748 11057 15804
rect 11057 15748 11113 15804
rect 11113 15748 11117 15804
rect 11053 15744 11117 15748
rect 5396 15676 5460 15740
rect 12572 15676 12636 15740
rect 12388 15540 12452 15604
rect 4476 15268 4540 15332
rect 6868 15404 6932 15468
rect 8892 15404 8956 15468
rect 9260 15404 9324 15468
rect 9812 15404 9876 15468
rect 9996 15404 10060 15468
rect 10364 15404 10428 15468
rect 11836 15268 11900 15332
rect 3417 15260 3481 15264
rect 3417 15204 3421 15260
rect 3421 15204 3477 15260
rect 3477 15204 3481 15260
rect 3417 15200 3481 15204
rect 3497 15260 3561 15264
rect 3497 15204 3501 15260
rect 3501 15204 3557 15260
rect 3557 15204 3561 15260
rect 3497 15200 3561 15204
rect 3577 15260 3641 15264
rect 3577 15204 3581 15260
rect 3581 15204 3637 15260
rect 3637 15204 3641 15260
rect 3577 15200 3641 15204
rect 3657 15260 3721 15264
rect 3657 15204 3661 15260
rect 3661 15204 3717 15260
rect 3717 15204 3721 15260
rect 3657 15200 3721 15204
rect 8348 15260 8412 15264
rect 8348 15204 8352 15260
rect 8352 15204 8408 15260
rect 8408 15204 8412 15260
rect 8348 15200 8412 15204
rect 8428 15260 8492 15264
rect 8428 15204 8432 15260
rect 8432 15204 8488 15260
rect 8488 15204 8492 15260
rect 8428 15200 8492 15204
rect 8508 15260 8572 15264
rect 8508 15204 8512 15260
rect 8512 15204 8568 15260
rect 8568 15204 8572 15260
rect 8508 15200 8572 15204
rect 8588 15260 8652 15264
rect 8588 15204 8592 15260
rect 8592 15204 8648 15260
rect 8648 15204 8652 15260
rect 8588 15200 8652 15204
rect 13278 15260 13342 15264
rect 13278 15204 13282 15260
rect 13282 15204 13338 15260
rect 13338 15204 13342 15260
rect 13278 15200 13342 15204
rect 13358 15260 13422 15264
rect 13358 15204 13362 15260
rect 13362 15204 13418 15260
rect 13418 15204 13422 15260
rect 13358 15200 13422 15204
rect 13438 15260 13502 15264
rect 13438 15204 13442 15260
rect 13442 15204 13498 15260
rect 13498 15204 13502 15260
rect 13438 15200 13502 15204
rect 13518 15260 13582 15264
rect 13518 15204 13522 15260
rect 13522 15204 13578 15260
rect 13578 15204 13582 15260
rect 13518 15200 13582 15204
rect 3188 15132 3252 15196
rect 9628 15132 9692 15196
rect 11652 15132 11716 15196
rect 12020 14996 12084 15060
rect 4660 14784 4724 14788
rect 4660 14728 4674 14784
rect 4674 14728 4724 14784
rect 4660 14724 4724 14728
rect 7236 14784 7300 14788
rect 7236 14728 7250 14784
rect 7250 14728 7300 14784
rect 7236 14724 7300 14728
rect 9076 14724 9140 14788
rect 5882 14716 5946 14720
rect 5882 14660 5886 14716
rect 5886 14660 5942 14716
rect 5942 14660 5946 14716
rect 5882 14656 5946 14660
rect 5962 14716 6026 14720
rect 5962 14660 5966 14716
rect 5966 14660 6022 14716
rect 6022 14660 6026 14716
rect 5962 14656 6026 14660
rect 6042 14716 6106 14720
rect 6042 14660 6046 14716
rect 6046 14660 6102 14716
rect 6102 14660 6106 14716
rect 6042 14656 6106 14660
rect 6122 14716 6186 14720
rect 6122 14660 6126 14716
rect 6126 14660 6182 14716
rect 6182 14660 6186 14716
rect 6122 14656 6186 14660
rect 10813 14716 10877 14720
rect 10813 14660 10817 14716
rect 10817 14660 10873 14716
rect 10873 14660 10877 14716
rect 10813 14656 10877 14660
rect 10893 14716 10957 14720
rect 10893 14660 10897 14716
rect 10897 14660 10953 14716
rect 10953 14660 10957 14716
rect 10893 14656 10957 14660
rect 10973 14716 11037 14720
rect 10973 14660 10977 14716
rect 10977 14660 11033 14716
rect 11033 14660 11037 14716
rect 10973 14656 11037 14660
rect 11053 14716 11117 14720
rect 11053 14660 11057 14716
rect 11057 14660 11113 14716
rect 11113 14660 11117 14716
rect 11053 14656 11117 14660
rect 10548 14648 10612 14652
rect 10548 14592 10562 14648
rect 10562 14592 10612 14648
rect 10548 14588 10612 14592
rect 12020 14452 12084 14516
rect 12940 14512 13004 14516
rect 12940 14456 12990 14512
rect 12990 14456 13004 14512
rect 12940 14452 13004 14456
rect 3004 14376 3068 14380
rect 3004 14320 3018 14376
rect 3018 14320 3068 14376
rect 3004 14316 3068 14320
rect 13676 14376 13740 14380
rect 13676 14320 13690 14376
rect 13690 14320 13740 14376
rect 13676 14316 13740 14320
rect 3417 14172 3481 14176
rect 3417 14116 3421 14172
rect 3421 14116 3477 14172
rect 3477 14116 3481 14172
rect 3417 14112 3481 14116
rect 3497 14172 3561 14176
rect 3497 14116 3501 14172
rect 3501 14116 3557 14172
rect 3557 14116 3561 14172
rect 3497 14112 3561 14116
rect 3577 14172 3641 14176
rect 3577 14116 3581 14172
rect 3581 14116 3637 14172
rect 3637 14116 3641 14172
rect 3577 14112 3641 14116
rect 3657 14172 3721 14176
rect 3657 14116 3661 14172
rect 3661 14116 3717 14172
rect 3717 14116 3721 14172
rect 3657 14112 3721 14116
rect 8348 14172 8412 14176
rect 8348 14116 8352 14172
rect 8352 14116 8408 14172
rect 8408 14116 8412 14172
rect 8348 14112 8412 14116
rect 8428 14172 8492 14176
rect 8428 14116 8432 14172
rect 8432 14116 8488 14172
rect 8488 14116 8492 14172
rect 8428 14112 8492 14116
rect 8508 14172 8572 14176
rect 8508 14116 8512 14172
rect 8512 14116 8568 14172
rect 8568 14116 8572 14172
rect 8508 14112 8572 14116
rect 8588 14172 8652 14176
rect 8588 14116 8592 14172
rect 8592 14116 8648 14172
rect 8648 14116 8652 14172
rect 8588 14112 8652 14116
rect 13278 14172 13342 14176
rect 13278 14116 13282 14172
rect 13282 14116 13338 14172
rect 13338 14116 13342 14172
rect 13278 14112 13342 14116
rect 13358 14172 13422 14176
rect 13358 14116 13362 14172
rect 13362 14116 13418 14172
rect 13418 14116 13422 14172
rect 13358 14112 13422 14116
rect 13438 14172 13502 14176
rect 13438 14116 13442 14172
rect 13442 14116 13498 14172
rect 13498 14116 13502 14172
rect 13438 14112 13502 14116
rect 13518 14172 13582 14176
rect 13518 14116 13522 14172
rect 13522 14116 13578 14172
rect 13578 14116 13582 14172
rect 13518 14112 13582 14116
rect 3188 13908 3252 13972
rect 9260 14044 9324 14108
rect 4292 13908 4356 13972
rect 9812 13908 9876 13972
rect 5882 13628 5946 13632
rect 5882 13572 5886 13628
rect 5886 13572 5942 13628
rect 5942 13572 5946 13628
rect 5882 13568 5946 13572
rect 5962 13628 6026 13632
rect 5962 13572 5966 13628
rect 5966 13572 6022 13628
rect 6022 13572 6026 13628
rect 5962 13568 6026 13572
rect 6042 13628 6106 13632
rect 6042 13572 6046 13628
rect 6046 13572 6102 13628
rect 6102 13572 6106 13628
rect 6042 13568 6106 13572
rect 6122 13628 6186 13632
rect 6122 13572 6126 13628
rect 6126 13572 6182 13628
rect 6182 13572 6186 13628
rect 6122 13568 6186 13572
rect 11468 13636 11532 13700
rect 10813 13628 10877 13632
rect 10813 13572 10817 13628
rect 10817 13572 10873 13628
rect 10873 13572 10877 13628
rect 10813 13568 10877 13572
rect 10893 13628 10957 13632
rect 10893 13572 10897 13628
rect 10897 13572 10953 13628
rect 10953 13572 10957 13628
rect 10893 13568 10957 13572
rect 10973 13628 11037 13632
rect 10973 13572 10977 13628
rect 10977 13572 11033 13628
rect 11033 13572 11037 13628
rect 10973 13568 11037 13572
rect 11053 13628 11117 13632
rect 11053 13572 11057 13628
rect 11057 13572 11113 13628
rect 11113 13572 11117 13628
rect 11053 13568 11117 13572
rect 12572 13500 12636 13564
rect 5028 13364 5092 13428
rect 12020 13424 12084 13428
rect 12020 13368 12034 13424
rect 12034 13368 12084 13424
rect 12020 13364 12084 13368
rect 12204 13424 12268 13428
rect 12204 13368 12218 13424
rect 12218 13368 12268 13424
rect 12204 13364 12268 13368
rect 12572 13364 12636 13428
rect 14044 13424 14108 13428
rect 14044 13368 14058 13424
rect 14058 13368 14108 13424
rect 14044 13364 14108 13368
rect 8156 13092 8220 13156
rect 11652 13092 11716 13156
rect 3417 13084 3481 13088
rect 3417 13028 3421 13084
rect 3421 13028 3477 13084
rect 3477 13028 3481 13084
rect 3417 13024 3481 13028
rect 3497 13084 3561 13088
rect 3497 13028 3501 13084
rect 3501 13028 3557 13084
rect 3557 13028 3561 13084
rect 3497 13024 3561 13028
rect 3577 13084 3641 13088
rect 3577 13028 3581 13084
rect 3581 13028 3637 13084
rect 3637 13028 3641 13084
rect 3577 13024 3641 13028
rect 3657 13084 3721 13088
rect 3657 13028 3661 13084
rect 3661 13028 3717 13084
rect 3717 13028 3721 13084
rect 3657 13024 3721 13028
rect 8348 13084 8412 13088
rect 8348 13028 8352 13084
rect 8352 13028 8408 13084
rect 8408 13028 8412 13084
rect 8348 13024 8412 13028
rect 8428 13084 8492 13088
rect 8428 13028 8432 13084
rect 8432 13028 8488 13084
rect 8488 13028 8492 13084
rect 8428 13024 8492 13028
rect 8508 13084 8572 13088
rect 8508 13028 8512 13084
rect 8512 13028 8568 13084
rect 8568 13028 8572 13084
rect 8508 13024 8572 13028
rect 8588 13084 8652 13088
rect 8588 13028 8592 13084
rect 8592 13028 8648 13084
rect 8648 13028 8652 13084
rect 8588 13024 8652 13028
rect 13278 13084 13342 13088
rect 13278 13028 13282 13084
rect 13282 13028 13338 13084
rect 13338 13028 13342 13084
rect 13278 13024 13342 13028
rect 13358 13084 13422 13088
rect 13358 13028 13362 13084
rect 13362 13028 13418 13084
rect 13418 13028 13422 13084
rect 13358 13024 13422 13028
rect 13438 13084 13502 13088
rect 13438 13028 13442 13084
rect 13442 13028 13498 13084
rect 13498 13028 13502 13084
rect 13438 13024 13502 13028
rect 13518 13084 13582 13088
rect 13518 13028 13522 13084
rect 13522 13028 13578 13084
rect 13578 13028 13582 13084
rect 13518 13024 13582 13028
rect 4108 12956 4172 13020
rect 8892 12956 8956 13020
rect 10180 12956 10244 13020
rect 11284 12956 11348 13020
rect 13860 12956 13924 13020
rect 5396 12548 5460 12612
rect 5882 12540 5946 12544
rect 5882 12484 5886 12540
rect 5886 12484 5942 12540
rect 5942 12484 5946 12540
rect 5882 12480 5946 12484
rect 5962 12540 6026 12544
rect 5962 12484 5966 12540
rect 5966 12484 6022 12540
rect 6022 12484 6026 12540
rect 5962 12480 6026 12484
rect 6042 12540 6106 12544
rect 6042 12484 6046 12540
rect 6046 12484 6102 12540
rect 6102 12484 6106 12540
rect 6042 12480 6106 12484
rect 6122 12540 6186 12544
rect 6122 12484 6126 12540
rect 6126 12484 6182 12540
rect 6182 12484 6186 12540
rect 6122 12480 6186 12484
rect 6868 12412 6932 12476
rect 9812 12412 9876 12476
rect 3188 12336 3252 12340
rect 3188 12280 3202 12336
rect 3202 12280 3252 12336
rect 3188 12276 3252 12280
rect 10813 12540 10877 12544
rect 10813 12484 10817 12540
rect 10817 12484 10873 12540
rect 10873 12484 10877 12540
rect 10813 12480 10877 12484
rect 10893 12540 10957 12544
rect 10893 12484 10897 12540
rect 10897 12484 10953 12540
rect 10953 12484 10957 12540
rect 10893 12480 10957 12484
rect 10973 12540 11037 12544
rect 10973 12484 10977 12540
rect 10977 12484 11033 12540
rect 11033 12484 11037 12540
rect 10973 12480 11037 12484
rect 11053 12540 11117 12544
rect 11053 12484 11057 12540
rect 11057 12484 11113 12540
rect 11113 12484 11117 12540
rect 11053 12480 11117 12484
rect 12388 12276 12452 12340
rect 6500 12004 6564 12068
rect 7788 12064 7852 12068
rect 7788 12008 7838 12064
rect 7838 12008 7852 12064
rect 7788 12004 7852 12008
rect 10548 12004 10612 12068
rect 3417 11996 3481 12000
rect 3417 11940 3421 11996
rect 3421 11940 3477 11996
rect 3477 11940 3481 11996
rect 3417 11936 3481 11940
rect 3497 11996 3561 12000
rect 3497 11940 3501 11996
rect 3501 11940 3557 11996
rect 3557 11940 3561 11996
rect 3497 11936 3561 11940
rect 3577 11996 3641 12000
rect 3577 11940 3581 11996
rect 3581 11940 3637 11996
rect 3637 11940 3641 11996
rect 3577 11936 3641 11940
rect 3657 11996 3721 12000
rect 3657 11940 3661 11996
rect 3661 11940 3717 11996
rect 3717 11940 3721 11996
rect 3657 11936 3721 11940
rect 8348 11996 8412 12000
rect 8348 11940 8352 11996
rect 8352 11940 8408 11996
rect 8408 11940 8412 11996
rect 8348 11936 8412 11940
rect 8428 11996 8492 12000
rect 8428 11940 8432 11996
rect 8432 11940 8488 11996
rect 8488 11940 8492 11996
rect 8428 11936 8492 11940
rect 8508 11996 8572 12000
rect 8508 11940 8512 11996
rect 8512 11940 8568 11996
rect 8568 11940 8572 11996
rect 8508 11936 8572 11940
rect 8588 11996 8652 12000
rect 8588 11940 8592 11996
rect 8592 11940 8648 11996
rect 8648 11940 8652 11996
rect 8588 11936 8652 11940
rect 13278 11996 13342 12000
rect 13278 11940 13282 11996
rect 13282 11940 13338 11996
rect 13338 11940 13342 11996
rect 13278 11936 13342 11940
rect 13358 11996 13422 12000
rect 13358 11940 13362 11996
rect 13362 11940 13418 11996
rect 13418 11940 13422 11996
rect 13358 11936 13422 11940
rect 13438 11996 13502 12000
rect 13438 11940 13442 11996
rect 13442 11940 13498 11996
rect 13498 11940 13502 11996
rect 13438 11936 13502 11940
rect 13518 11996 13582 12000
rect 13518 11940 13522 11996
rect 13522 11940 13578 11996
rect 13578 11940 13582 11996
rect 13518 11936 13582 11940
rect 8892 11868 8956 11932
rect 11652 11732 11716 11796
rect 8892 11596 8956 11660
rect 9628 11596 9692 11660
rect 9996 11596 10060 11660
rect 11284 11520 11348 11524
rect 11284 11464 11334 11520
rect 11334 11464 11348 11520
rect 11284 11460 11348 11464
rect 13860 11460 13924 11524
rect 14228 11520 14292 11524
rect 14228 11464 14242 11520
rect 14242 11464 14292 11520
rect 14228 11460 14292 11464
rect 5882 11452 5946 11456
rect 5882 11396 5886 11452
rect 5886 11396 5942 11452
rect 5942 11396 5946 11452
rect 5882 11392 5946 11396
rect 5962 11452 6026 11456
rect 5962 11396 5966 11452
rect 5966 11396 6022 11452
rect 6022 11396 6026 11452
rect 5962 11392 6026 11396
rect 6042 11452 6106 11456
rect 6042 11396 6046 11452
rect 6046 11396 6102 11452
rect 6102 11396 6106 11452
rect 6042 11392 6106 11396
rect 6122 11452 6186 11456
rect 6122 11396 6126 11452
rect 6126 11396 6182 11452
rect 6182 11396 6186 11452
rect 6122 11392 6186 11396
rect 10813 11452 10877 11456
rect 10813 11396 10817 11452
rect 10817 11396 10873 11452
rect 10873 11396 10877 11452
rect 10813 11392 10877 11396
rect 10893 11452 10957 11456
rect 10893 11396 10897 11452
rect 10897 11396 10953 11452
rect 10953 11396 10957 11452
rect 10893 11392 10957 11396
rect 10973 11452 11037 11456
rect 10973 11396 10977 11452
rect 10977 11396 11033 11452
rect 11033 11396 11037 11452
rect 10973 11392 11037 11396
rect 11053 11452 11117 11456
rect 11053 11396 11057 11452
rect 11057 11396 11113 11452
rect 11113 11396 11117 11452
rect 11053 11392 11117 11396
rect 5396 11384 5460 11388
rect 5396 11328 5446 11384
rect 5446 11328 5460 11384
rect 5396 11324 5460 11328
rect 10548 11384 10612 11388
rect 10548 11328 10562 11384
rect 10562 11328 10612 11384
rect 10548 11324 10612 11328
rect 11284 11324 11348 11388
rect 12756 11324 12820 11388
rect 3188 11052 3252 11116
rect 3004 10916 3068 10980
rect 10180 11052 10244 11116
rect 3417 10908 3481 10912
rect 3417 10852 3421 10908
rect 3421 10852 3477 10908
rect 3477 10852 3481 10908
rect 3417 10848 3481 10852
rect 3497 10908 3561 10912
rect 3497 10852 3501 10908
rect 3501 10852 3557 10908
rect 3557 10852 3561 10908
rect 3497 10848 3561 10852
rect 3577 10908 3641 10912
rect 3577 10852 3581 10908
rect 3581 10852 3637 10908
rect 3637 10852 3641 10908
rect 3577 10848 3641 10852
rect 3657 10908 3721 10912
rect 3657 10852 3661 10908
rect 3661 10852 3717 10908
rect 3717 10852 3721 10908
rect 3657 10848 3721 10852
rect 5396 10780 5460 10844
rect 7236 10780 7300 10844
rect 12388 10916 12452 10980
rect 8348 10908 8412 10912
rect 8348 10852 8352 10908
rect 8352 10852 8408 10908
rect 8408 10852 8412 10908
rect 8348 10848 8412 10852
rect 8428 10908 8492 10912
rect 8428 10852 8432 10908
rect 8432 10852 8488 10908
rect 8488 10852 8492 10908
rect 8428 10848 8492 10852
rect 8508 10908 8572 10912
rect 8508 10852 8512 10908
rect 8512 10852 8568 10908
rect 8568 10852 8572 10908
rect 8508 10848 8572 10852
rect 8588 10908 8652 10912
rect 8588 10852 8592 10908
rect 8592 10852 8648 10908
rect 8648 10852 8652 10908
rect 8588 10848 8652 10852
rect 13278 10908 13342 10912
rect 13278 10852 13282 10908
rect 13282 10852 13338 10908
rect 13338 10852 13342 10908
rect 13278 10848 13342 10852
rect 13358 10908 13422 10912
rect 13358 10852 13362 10908
rect 13362 10852 13418 10908
rect 13418 10852 13422 10908
rect 13358 10848 13422 10852
rect 13438 10908 13502 10912
rect 13438 10852 13442 10908
rect 13442 10852 13498 10908
rect 13498 10852 13502 10908
rect 13438 10848 13502 10852
rect 13518 10908 13582 10912
rect 13518 10852 13522 10908
rect 13522 10852 13578 10908
rect 13578 10852 13582 10908
rect 13518 10848 13582 10852
rect 12940 10644 13004 10708
rect 9812 10508 9876 10572
rect 12572 10508 12636 10572
rect 12940 10508 13004 10572
rect 14044 10508 14108 10572
rect 3004 10372 3068 10436
rect 8156 10372 8220 10436
rect 9628 10372 9692 10436
rect 14228 10372 14292 10436
rect 5882 10364 5946 10368
rect 5882 10308 5886 10364
rect 5886 10308 5942 10364
rect 5942 10308 5946 10364
rect 5882 10304 5946 10308
rect 5962 10364 6026 10368
rect 5962 10308 5966 10364
rect 5966 10308 6022 10364
rect 6022 10308 6026 10364
rect 5962 10304 6026 10308
rect 6042 10364 6106 10368
rect 6042 10308 6046 10364
rect 6046 10308 6102 10364
rect 6102 10308 6106 10364
rect 6042 10304 6106 10308
rect 6122 10364 6186 10368
rect 6122 10308 6126 10364
rect 6126 10308 6182 10364
rect 6182 10308 6186 10364
rect 6122 10304 6186 10308
rect 10813 10364 10877 10368
rect 10813 10308 10817 10364
rect 10817 10308 10873 10364
rect 10873 10308 10877 10364
rect 10813 10304 10877 10308
rect 10893 10364 10957 10368
rect 10893 10308 10897 10364
rect 10897 10308 10953 10364
rect 10953 10308 10957 10364
rect 10893 10304 10957 10308
rect 10973 10364 11037 10368
rect 10973 10308 10977 10364
rect 10977 10308 11033 10364
rect 11033 10308 11037 10364
rect 10973 10304 11037 10308
rect 11053 10364 11117 10368
rect 11053 10308 11057 10364
rect 11057 10308 11113 10364
rect 11113 10308 11117 10364
rect 11053 10304 11117 10308
rect 6500 10236 6564 10300
rect 9628 10236 9692 10300
rect 9444 10100 9508 10164
rect 4108 10024 4172 10028
rect 4108 9968 4122 10024
rect 4122 9968 4172 10024
rect 4108 9964 4172 9968
rect 6684 9964 6748 10028
rect 9076 9828 9140 9892
rect 3417 9820 3481 9824
rect 3417 9764 3421 9820
rect 3421 9764 3477 9820
rect 3477 9764 3481 9820
rect 3417 9760 3481 9764
rect 3497 9820 3561 9824
rect 3497 9764 3501 9820
rect 3501 9764 3557 9820
rect 3557 9764 3561 9820
rect 3497 9760 3561 9764
rect 3577 9820 3641 9824
rect 3577 9764 3581 9820
rect 3581 9764 3637 9820
rect 3637 9764 3641 9820
rect 3577 9760 3641 9764
rect 3657 9820 3721 9824
rect 3657 9764 3661 9820
rect 3661 9764 3717 9820
rect 3717 9764 3721 9820
rect 3657 9760 3721 9764
rect 8348 9820 8412 9824
rect 8348 9764 8352 9820
rect 8352 9764 8408 9820
rect 8408 9764 8412 9820
rect 8348 9760 8412 9764
rect 8428 9820 8492 9824
rect 8428 9764 8432 9820
rect 8432 9764 8488 9820
rect 8488 9764 8492 9820
rect 8428 9760 8492 9764
rect 8508 9820 8572 9824
rect 8508 9764 8512 9820
rect 8512 9764 8568 9820
rect 8568 9764 8572 9820
rect 8508 9760 8572 9764
rect 8588 9820 8652 9824
rect 8588 9764 8592 9820
rect 8592 9764 8648 9820
rect 8648 9764 8652 9820
rect 8588 9760 8652 9764
rect 13278 9820 13342 9824
rect 13278 9764 13282 9820
rect 13282 9764 13338 9820
rect 13338 9764 13342 9820
rect 13278 9760 13342 9764
rect 13358 9820 13422 9824
rect 13358 9764 13362 9820
rect 13362 9764 13418 9820
rect 13418 9764 13422 9820
rect 13358 9760 13422 9764
rect 13438 9820 13502 9824
rect 13438 9764 13442 9820
rect 13442 9764 13498 9820
rect 13498 9764 13502 9820
rect 13438 9760 13502 9764
rect 13518 9820 13582 9824
rect 13518 9764 13522 9820
rect 13522 9764 13578 9820
rect 13578 9764 13582 9820
rect 13518 9760 13582 9764
rect 9260 9692 9324 9756
rect 14044 9616 14108 9620
rect 14044 9560 14058 9616
rect 14058 9560 14108 9616
rect 14044 9556 14108 9560
rect 12940 9420 13004 9484
rect 13860 9284 13924 9348
rect 5882 9276 5946 9280
rect 5882 9220 5886 9276
rect 5886 9220 5942 9276
rect 5942 9220 5946 9276
rect 5882 9216 5946 9220
rect 5962 9276 6026 9280
rect 5962 9220 5966 9276
rect 5966 9220 6022 9276
rect 6022 9220 6026 9276
rect 5962 9216 6026 9220
rect 6042 9276 6106 9280
rect 6042 9220 6046 9276
rect 6046 9220 6102 9276
rect 6102 9220 6106 9276
rect 6042 9216 6106 9220
rect 6122 9276 6186 9280
rect 6122 9220 6126 9276
rect 6126 9220 6182 9276
rect 6182 9220 6186 9276
rect 6122 9216 6186 9220
rect 10813 9276 10877 9280
rect 10813 9220 10817 9276
rect 10817 9220 10873 9276
rect 10873 9220 10877 9276
rect 10813 9216 10877 9220
rect 10893 9276 10957 9280
rect 10893 9220 10897 9276
rect 10897 9220 10953 9276
rect 10953 9220 10957 9276
rect 10893 9216 10957 9220
rect 10973 9276 11037 9280
rect 10973 9220 10977 9276
rect 10977 9220 11033 9276
rect 11033 9220 11037 9276
rect 10973 9216 11037 9220
rect 11053 9276 11117 9280
rect 11053 9220 11057 9276
rect 11057 9220 11113 9276
rect 11113 9220 11117 9276
rect 11053 9216 11117 9220
rect 11468 9148 11532 9212
rect 7972 9012 8036 9076
rect 12572 8876 12636 8940
rect 9076 8740 9140 8804
rect 12020 8740 12084 8804
rect 3417 8732 3481 8736
rect 3417 8676 3421 8732
rect 3421 8676 3477 8732
rect 3477 8676 3481 8732
rect 3417 8672 3481 8676
rect 3497 8732 3561 8736
rect 3497 8676 3501 8732
rect 3501 8676 3557 8732
rect 3557 8676 3561 8732
rect 3497 8672 3561 8676
rect 3577 8732 3641 8736
rect 3577 8676 3581 8732
rect 3581 8676 3637 8732
rect 3637 8676 3641 8732
rect 3577 8672 3641 8676
rect 3657 8732 3721 8736
rect 3657 8676 3661 8732
rect 3661 8676 3717 8732
rect 3717 8676 3721 8732
rect 3657 8672 3721 8676
rect 8348 8732 8412 8736
rect 8348 8676 8352 8732
rect 8352 8676 8408 8732
rect 8408 8676 8412 8732
rect 8348 8672 8412 8676
rect 8428 8732 8492 8736
rect 8428 8676 8432 8732
rect 8432 8676 8488 8732
rect 8488 8676 8492 8732
rect 8428 8672 8492 8676
rect 8508 8732 8572 8736
rect 8508 8676 8512 8732
rect 8512 8676 8568 8732
rect 8568 8676 8572 8732
rect 8508 8672 8572 8676
rect 8588 8732 8652 8736
rect 8588 8676 8592 8732
rect 8592 8676 8648 8732
rect 8648 8676 8652 8732
rect 8588 8672 8652 8676
rect 13278 8732 13342 8736
rect 13278 8676 13282 8732
rect 13282 8676 13338 8732
rect 13338 8676 13342 8732
rect 13278 8672 13342 8676
rect 13358 8732 13422 8736
rect 13358 8676 13362 8732
rect 13362 8676 13418 8732
rect 13418 8676 13422 8732
rect 13358 8672 13422 8676
rect 13438 8732 13502 8736
rect 13438 8676 13442 8732
rect 13442 8676 13498 8732
rect 13498 8676 13502 8732
rect 13438 8672 13502 8676
rect 13518 8732 13582 8736
rect 13518 8676 13522 8732
rect 13522 8676 13578 8732
rect 13578 8676 13582 8732
rect 13518 8672 13582 8676
rect 6868 8604 6932 8668
rect 12020 8604 12084 8668
rect 7236 8332 7300 8396
rect 7420 8196 7484 8260
rect 9996 8196 10060 8260
rect 12388 8256 12452 8260
rect 12388 8200 12402 8256
rect 12402 8200 12452 8256
rect 12388 8196 12452 8200
rect 5882 8188 5946 8192
rect 5882 8132 5886 8188
rect 5886 8132 5942 8188
rect 5942 8132 5946 8188
rect 5882 8128 5946 8132
rect 5962 8188 6026 8192
rect 5962 8132 5966 8188
rect 5966 8132 6022 8188
rect 6022 8132 6026 8188
rect 5962 8128 6026 8132
rect 6042 8188 6106 8192
rect 6042 8132 6046 8188
rect 6046 8132 6102 8188
rect 6102 8132 6106 8188
rect 6042 8128 6106 8132
rect 6122 8188 6186 8192
rect 6122 8132 6126 8188
rect 6126 8132 6182 8188
rect 6182 8132 6186 8188
rect 6122 8128 6186 8132
rect 10813 8188 10877 8192
rect 10813 8132 10817 8188
rect 10817 8132 10873 8188
rect 10873 8132 10877 8188
rect 10813 8128 10877 8132
rect 10893 8188 10957 8192
rect 10893 8132 10897 8188
rect 10897 8132 10953 8188
rect 10953 8132 10957 8188
rect 10893 8128 10957 8132
rect 10973 8188 11037 8192
rect 10973 8132 10977 8188
rect 10977 8132 11033 8188
rect 11033 8132 11037 8188
rect 10973 8128 11037 8132
rect 11053 8188 11117 8192
rect 11053 8132 11057 8188
rect 11057 8132 11113 8188
rect 11113 8132 11117 8188
rect 11053 8128 11117 8132
rect 12756 7924 12820 7988
rect 12756 7788 12820 7852
rect 10180 7652 10244 7716
rect 3417 7644 3481 7648
rect 3417 7588 3421 7644
rect 3421 7588 3477 7644
rect 3477 7588 3481 7644
rect 3417 7584 3481 7588
rect 3497 7644 3561 7648
rect 3497 7588 3501 7644
rect 3501 7588 3557 7644
rect 3557 7588 3561 7644
rect 3497 7584 3561 7588
rect 3577 7644 3641 7648
rect 3577 7588 3581 7644
rect 3581 7588 3637 7644
rect 3637 7588 3641 7644
rect 3577 7584 3641 7588
rect 3657 7644 3721 7648
rect 3657 7588 3661 7644
rect 3661 7588 3717 7644
rect 3717 7588 3721 7644
rect 3657 7584 3721 7588
rect 8348 7644 8412 7648
rect 8348 7588 8352 7644
rect 8352 7588 8408 7644
rect 8408 7588 8412 7644
rect 8348 7584 8412 7588
rect 8428 7644 8492 7648
rect 8428 7588 8432 7644
rect 8432 7588 8488 7644
rect 8488 7588 8492 7644
rect 8428 7584 8492 7588
rect 8508 7644 8572 7648
rect 8508 7588 8512 7644
rect 8512 7588 8568 7644
rect 8568 7588 8572 7644
rect 8508 7584 8572 7588
rect 8588 7644 8652 7648
rect 8588 7588 8592 7644
rect 8592 7588 8648 7644
rect 8648 7588 8652 7644
rect 8588 7584 8652 7588
rect 13278 7644 13342 7648
rect 13278 7588 13282 7644
rect 13282 7588 13338 7644
rect 13338 7588 13342 7644
rect 13278 7584 13342 7588
rect 13358 7644 13422 7648
rect 13358 7588 13362 7644
rect 13362 7588 13418 7644
rect 13418 7588 13422 7644
rect 13358 7584 13422 7588
rect 13438 7644 13502 7648
rect 13438 7588 13442 7644
rect 13442 7588 13498 7644
rect 13498 7588 13502 7644
rect 13438 7584 13502 7588
rect 13518 7644 13582 7648
rect 13518 7588 13522 7644
rect 13522 7588 13578 7644
rect 13578 7588 13582 7644
rect 13518 7584 13582 7588
rect 9260 7516 9324 7580
rect 14228 7304 14292 7308
rect 14228 7248 14242 7304
rect 14242 7248 14292 7304
rect 14228 7244 14292 7248
rect 9260 7108 9324 7172
rect 5882 7100 5946 7104
rect 5882 7044 5886 7100
rect 5886 7044 5942 7100
rect 5942 7044 5946 7100
rect 5882 7040 5946 7044
rect 5962 7100 6026 7104
rect 5962 7044 5966 7100
rect 5966 7044 6022 7100
rect 6022 7044 6026 7100
rect 5962 7040 6026 7044
rect 6042 7100 6106 7104
rect 6042 7044 6046 7100
rect 6046 7044 6102 7100
rect 6102 7044 6106 7100
rect 6042 7040 6106 7044
rect 6122 7100 6186 7104
rect 6122 7044 6126 7100
rect 6126 7044 6182 7100
rect 6182 7044 6186 7100
rect 6122 7040 6186 7044
rect 10813 7100 10877 7104
rect 10813 7044 10817 7100
rect 10817 7044 10873 7100
rect 10873 7044 10877 7100
rect 10813 7040 10877 7044
rect 10893 7100 10957 7104
rect 10893 7044 10897 7100
rect 10897 7044 10953 7100
rect 10953 7044 10957 7100
rect 10893 7040 10957 7044
rect 10973 7100 11037 7104
rect 10973 7044 10977 7100
rect 10977 7044 11033 7100
rect 11033 7044 11037 7100
rect 10973 7040 11037 7044
rect 11053 7100 11117 7104
rect 11053 7044 11057 7100
rect 11057 7044 11113 7100
rect 11113 7044 11117 7100
rect 11053 7040 11117 7044
rect 11284 6700 11348 6764
rect 13124 6836 13188 6900
rect 3417 6556 3481 6560
rect 3417 6500 3421 6556
rect 3421 6500 3477 6556
rect 3477 6500 3481 6556
rect 3417 6496 3481 6500
rect 3497 6556 3561 6560
rect 3497 6500 3501 6556
rect 3501 6500 3557 6556
rect 3557 6500 3561 6556
rect 3497 6496 3561 6500
rect 3577 6556 3641 6560
rect 3577 6500 3581 6556
rect 3581 6500 3637 6556
rect 3637 6500 3641 6556
rect 3577 6496 3641 6500
rect 3657 6556 3721 6560
rect 3657 6500 3661 6556
rect 3661 6500 3717 6556
rect 3717 6500 3721 6556
rect 3657 6496 3721 6500
rect 8348 6556 8412 6560
rect 8348 6500 8352 6556
rect 8352 6500 8408 6556
rect 8408 6500 8412 6556
rect 8348 6496 8412 6500
rect 8428 6556 8492 6560
rect 8428 6500 8432 6556
rect 8432 6500 8488 6556
rect 8488 6500 8492 6556
rect 8428 6496 8492 6500
rect 8508 6556 8572 6560
rect 8508 6500 8512 6556
rect 8512 6500 8568 6556
rect 8568 6500 8572 6556
rect 8508 6496 8572 6500
rect 8588 6556 8652 6560
rect 8588 6500 8592 6556
rect 8592 6500 8648 6556
rect 8648 6500 8652 6556
rect 8588 6496 8652 6500
rect 13278 6556 13342 6560
rect 13278 6500 13282 6556
rect 13282 6500 13338 6556
rect 13338 6500 13342 6556
rect 13278 6496 13342 6500
rect 13358 6556 13422 6560
rect 13358 6500 13362 6556
rect 13362 6500 13418 6556
rect 13418 6500 13422 6556
rect 13358 6496 13422 6500
rect 13438 6556 13502 6560
rect 13438 6500 13442 6556
rect 13442 6500 13498 6556
rect 13498 6500 13502 6556
rect 13438 6496 13502 6500
rect 13518 6556 13582 6560
rect 13518 6500 13522 6556
rect 13522 6500 13578 6556
rect 13578 6500 13582 6556
rect 13518 6496 13582 6500
rect 12388 6428 12452 6492
rect 4108 6020 4172 6084
rect 5882 6012 5946 6016
rect 5882 5956 5886 6012
rect 5886 5956 5942 6012
rect 5942 5956 5946 6012
rect 5882 5952 5946 5956
rect 5962 6012 6026 6016
rect 5962 5956 5966 6012
rect 5966 5956 6022 6012
rect 6022 5956 6026 6012
rect 5962 5952 6026 5956
rect 6042 6012 6106 6016
rect 6042 5956 6046 6012
rect 6046 5956 6102 6012
rect 6102 5956 6106 6012
rect 6042 5952 6106 5956
rect 6122 6012 6186 6016
rect 6122 5956 6126 6012
rect 6126 5956 6182 6012
rect 6182 5956 6186 6012
rect 6122 5952 6186 5956
rect 6316 5884 6380 5948
rect 9628 6020 9692 6084
rect 10813 6012 10877 6016
rect 10813 5956 10817 6012
rect 10817 5956 10873 6012
rect 10873 5956 10877 6012
rect 10813 5952 10877 5956
rect 10893 6012 10957 6016
rect 10893 5956 10897 6012
rect 10897 5956 10953 6012
rect 10953 5956 10957 6012
rect 10893 5952 10957 5956
rect 10973 6012 11037 6016
rect 10973 5956 10977 6012
rect 10977 5956 11033 6012
rect 11033 5956 11037 6012
rect 10973 5952 11037 5956
rect 11053 6012 11117 6016
rect 11053 5956 11057 6012
rect 11057 5956 11113 6012
rect 11113 5956 11117 6012
rect 11053 5952 11117 5956
rect 8156 5748 8220 5812
rect 14044 5884 14108 5948
rect 10364 5612 10428 5676
rect 10364 5476 10428 5540
rect 3417 5468 3481 5472
rect 3417 5412 3421 5468
rect 3421 5412 3477 5468
rect 3477 5412 3481 5468
rect 3417 5408 3481 5412
rect 3497 5468 3561 5472
rect 3497 5412 3501 5468
rect 3501 5412 3557 5468
rect 3557 5412 3561 5468
rect 3497 5408 3561 5412
rect 3577 5468 3641 5472
rect 3577 5412 3581 5468
rect 3581 5412 3637 5468
rect 3637 5412 3641 5468
rect 3577 5408 3641 5412
rect 3657 5468 3721 5472
rect 3657 5412 3661 5468
rect 3661 5412 3717 5468
rect 3717 5412 3721 5468
rect 3657 5408 3721 5412
rect 8348 5468 8412 5472
rect 8348 5412 8352 5468
rect 8352 5412 8408 5468
rect 8408 5412 8412 5468
rect 8348 5408 8412 5412
rect 8428 5468 8492 5472
rect 8428 5412 8432 5468
rect 8432 5412 8488 5468
rect 8488 5412 8492 5468
rect 8428 5408 8492 5412
rect 8508 5468 8572 5472
rect 8508 5412 8512 5468
rect 8512 5412 8568 5468
rect 8568 5412 8572 5468
rect 8508 5408 8572 5412
rect 8588 5468 8652 5472
rect 8588 5412 8592 5468
rect 8592 5412 8648 5468
rect 8648 5412 8652 5468
rect 8588 5408 8652 5412
rect 13278 5468 13342 5472
rect 13278 5412 13282 5468
rect 13282 5412 13338 5468
rect 13338 5412 13342 5468
rect 13278 5408 13342 5412
rect 13358 5468 13422 5472
rect 13358 5412 13362 5468
rect 13362 5412 13418 5468
rect 13418 5412 13422 5468
rect 13358 5408 13422 5412
rect 13438 5468 13502 5472
rect 13438 5412 13442 5468
rect 13442 5412 13498 5468
rect 13498 5412 13502 5468
rect 13438 5408 13502 5412
rect 13518 5468 13582 5472
rect 13518 5412 13522 5468
rect 13522 5412 13578 5468
rect 13578 5412 13582 5468
rect 13518 5408 13582 5412
rect 7788 5204 7852 5268
rect 9444 5204 9508 5268
rect 4292 4932 4356 4996
rect 5882 4924 5946 4928
rect 5882 4868 5886 4924
rect 5886 4868 5942 4924
rect 5942 4868 5946 4924
rect 5882 4864 5946 4868
rect 5962 4924 6026 4928
rect 5962 4868 5966 4924
rect 5966 4868 6022 4924
rect 6022 4868 6026 4924
rect 5962 4864 6026 4868
rect 6042 4924 6106 4928
rect 6042 4868 6046 4924
rect 6046 4868 6102 4924
rect 6102 4868 6106 4924
rect 6042 4864 6106 4868
rect 6122 4924 6186 4928
rect 6122 4868 6126 4924
rect 6126 4868 6182 4924
rect 6182 4868 6186 4924
rect 6122 4864 6186 4868
rect 7052 4796 7116 4860
rect 11284 4932 11348 4996
rect 12756 4932 12820 4996
rect 10813 4924 10877 4928
rect 10813 4868 10817 4924
rect 10817 4868 10873 4924
rect 10873 4868 10877 4924
rect 10813 4864 10877 4868
rect 10893 4924 10957 4928
rect 10893 4868 10897 4924
rect 10897 4868 10953 4924
rect 10953 4868 10957 4924
rect 10893 4864 10957 4868
rect 10973 4924 11037 4928
rect 10973 4868 10977 4924
rect 10977 4868 11033 4924
rect 11033 4868 11037 4924
rect 10973 4864 11037 4868
rect 11053 4924 11117 4928
rect 11053 4868 11057 4924
rect 11057 4868 11113 4924
rect 11113 4868 11117 4924
rect 11053 4864 11117 4868
rect 9444 4796 9508 4860
rect 10180 4822 10244 4860
rect 10180 4796 10194 4822
rect 10194 4796 10244 4822
rect 14044 4796 14108 4860
rect 9996 4660 10060 4724
rect 11652 4524 11716 4588
rect 12756 4584 12820 4588
rect 12756 4528 12770 4584
rect 12770 4528 12820 4584
rect 12756 4524 12820 4528
rect 9260 4388 9324 4452
rect 11284 4388 11348 4452
rect 11652 4388 11716 4452
rect 12020 4388 12084 4452
rect 3417 4380 3481 4384
rect 3417 4324 3421 4380
rect 3421 4324 3477 4380
rect 3477 4324 3481 4380
rect 3417 4320 3481 4324
rect 3497 4380 3561 4384
rect 3497 4324 3501 4380
rect 3501 4324 3557 4380
rect 3557 4324 3561 4380
rect 3497 4320 3561 4324
rect 3577 4380 3641 4384
rect 3577 4324 3581 4380
rect 3581 4324 3637 4380
rect 3637 4324 3641 4380
rect 3577 4320 3641 4324
rect 3657 4380 3721 4384
rect 3657 4324 3661 4380
rect 3661 4324 3717 4380
rect 3717 4324 3721 4380
rect 3657 4320 3721 4324
rect 8348 4380 8412 4384
rect 8348 4324 8352 4380
rect 8352 4324 8408 4380
rect 8408 4324 8412 4380
rect 8348 4320 8412 4324
rect 8428 4380 8492 4384
rect 8428 4324 8432 4380
rect 8432 4324 8488 4380
rect 8488 4324 8492 4380
rect 8428 4320 8492 4324
rect 8508 4380 8572 4384
rect 8508 4324 8512 4380
rect 8512 4324 8568 4380
rect 8568 4324 8572 4380
rect 8508 4320 8572 4324
rect 8588 4380 8652 4384
rect 8588 4324 8592 4380
rect 8592 4324 8648 4380
rect 8648 4324 8652 4380
rect 8588 4320 8652 4324
rect 8892 4252 8956 4316
rect 13278 4380 13342 4384
rect 13278 4324 13282 4380
rect 13282 4324 13338 4380
rect 13338 4324 13342 4380
rect 13278 4320 13342 4324
rect 13358 4380 13422 4384
rect 13358 4324 13362 4380
rect 13362 4324 13418 4380
rect 13418 4324 13422 4380
rect 13358 4320 13422 4324
rect 13438 4380 13502 4384
rect 13438 4324 13442 4380
rect 13442 4324 13498 4380
rect 13498 4324 13502 4380
rect 13438 4320 13502 4324
rect 13518 4380 13582 4384
rect 13518 4324 13522 4380
rect 13522 4324 13578 4380
rect 13578 4324 13582 4380
rect 13518 4320 13582 4324
rect 4108 4116 4172 4180
rect 7604 4116 7668 4180
rect 10364 4116 10428 4180
rect 6868 3904 6932 3908
rect 6868 3848 6882 3904
rect 6882 3848 6932 3904
rect 6868 3844 6932 3848
rect 10364 3844 10428 3908
rect 11836 4040 11900 4044
rect 12572 4116 12636 4180
rect 13124 4116 13188 4180
rect 11836 3984 11886 4040
rect 11886 3984 11900 4040
rect 11836 3980 11900 3984
rect 5882 3836 5946 3840
rect 5882 3780 5886 3836
rect 5886 3780 5942 3836
rect 5942 3780 5946 3836
rect 5882 3776 5946 3780
rect 5962 3836 6026 3840
rect 5962 3780 5966 3836
rect 5966 3780 6022 3836
rect 6022 3780 6026 3836
rect 5962 3776 6026 3780
rect 6042 3836 6106 3840
rect 6042 3780 6046 3836
rect 6046 3780 6102 3836
rect 6102 3780 6106 3836
rect 6042 3776 6106 3780
rect 6122 3836 6186 3840
rect 6122 3780 6126 3836
rect 6126 3780 6182 3836
rect 6182 3780 6186 3836
rect 6122 3776 6186 3780
rect 10813 3836 10877 3840
rect 10813 3780 10817 3836
rect 10817 3780 10873 3836
rect 10873 3780 10877 3836
rect 10813 3776 10877 3780
rect 10893 3836 10957 3840
rect 10893 3780 10897 3836
rect 10897 3780 10953 3836
rect 10953 3780 10957 3836
rect 10893 3776 10957 3780
rect 10973 3836 11037 3840
rect 10973 3780 10977 3836
rect 10977 3780 11033 3836
rect 11033 3780 11037 3836
rect 10973 3776 11037 3780
rect 11053 3836 11117 3840
rect 11053 3780 11057 3836
rect 11057 3780 11113 3836
rect 11113 3780 11117 3836
rect 11053 3776 11117 3780
rect 5396 3708 5460 3772
rect 4476 3572 4540 3636
rect 11836 3572 11900 3636
rect 12020 3572 12084 3636
rect 12756 3572 12820 3636
rect 13860 3572 13924 3636
rect 9076 3496 9140 3500
rect 9076 3440 9126 3496
rect 9126 3440 9140 3496
rect 9076 3436 9140 3440
rect 11836 3360 11900 3364
rect 11836 3304 11886 3360
rect 11886 3304 11900 3360
rect 11836 3300 11900 3304
rect 3417 3292 3481 3296
rect 3417 3236 3421 3292
rect 3421 3236 3477 3292
rect 3477 3236 3481 3292
rect 3417 3232 3481 3236
rect 3497 3292 3561 3296
rect 3497 3236 3501 3292
rect 3501 3236 3557 3292
rect 3557 3236 3561 3292
rect 3497 3232 3561 3236
rect 3577 3292 3641 3296
rect 3577 3236 3581 3292
rect 3581 3236 3637 3292
rect 3637 3236 3641 3292
rect 3577 3232 3641 3236
rect 3657 3292 3721 3296
rect 3657 3236 3661 3292
rect 3661 3236 3717 3292
rect 3717 3236 3721 3292
rect 3657 3232 3721 3236
rect 8348 3292 8412 3296
rect 8348 3236 8352 3292
rect 8352 3236 8408 3292
rect 8408 3236 8412 3292
rect 8348 3232 8412 3236
rect 8428 3292 8492 3296
rect 8428 3236 8432 3292
rect 8432 3236 8488 3292
rect 8488 3236 8492 3292
rect 8428 3232 8492 3236
rect 8508 3292 8572 3296
rect 8508 3236 8512 3292
rect 8512 3236 8568 3292
rect 8568 3236 8572 3292
rect 8508 3232 8572 3236
rect 8588 3292 8652 3296
rect 8588 3236 8592 3292
rect 8592 3236 8648 3292
rect 8648 3236 8652 3292
rect 8588 3232 8652 3236
rect 13278 3292 13342 3296
rect 13278 3236 13282 3292
rect 13282 3236 13338 3292
rect 13338 3236 13342 3292
rect 13278 3232 13342 3236
rect 13358 3292 13422 3296
rect 13358 3236 13362 3292
rect 13362 3236 13418 3292
rect 13418 3236 13422 3292
rect 13358 3232 13422 3236
rect 13438 3292 13502 3296
rect 13438 3236 13442 3292
rect 13442 3236 13498 3292
rect 13498 3236 13502 3292
rect 13438 3232 13502 3236
rect 13518 3292 13582 3296
rect 13518 3236 13522 3292
rect 13522 3236 13578 3292
rect 13578 3236 13582 3292
rect 13518 3232 13582 3236
rect 9628 3028 9692 3092
rect 12388 3028 12452 3092
rect 3188 2892 3252 2956
rect 4292 2952 4356 2956
rect 4292 2896 4306 2952
rect 4306 2896 4356 2952
rect 4292 2892 4356 2896
rect 7604 2892 7668 2956
rect 7788 2952 7852 2956
rect 7788 2896 7838 2952
rect 7838 2896 7852 2952
rect 7788 2892 7852 2896
rect 6684 2756 6748 2820
rect 9812 2756 9876 2820
rect 12204 2756 12268 2820
rect 5882 2748 5946 2752
rect 5882 2692 5886 2748
rect 5886 2692 5942 2748
rect 5942 2692 5946 2748
rect 5882 2688 5946 2692
rect 5962 2748 6026 2752
rect 5962 2692 5966 2748
rect 5966 2692 6022 2748
rect 6022 2692 6026 2748
rect 5962 2688 6026 2692
rect 6042 2748 6106 2752
rect 6042 2692 6046 2748
rect 6046 2692 6102 2748
rect 6102 2692 6106 2748
rect 6042 2688 6106 2692
rect 6122 2748 6186 2752
rect 6122 2692 6126 2748
rect 6126 2692 6182 2748
rect 6182 2692 6186 2748
rect 6122 2688 6186 2692
rect 10813 2748 10877 2752
rect 10813 2692 10817 2748
rect 10817 2692 10873 2748
rect 10873 2692 10877 2748
rect 10813 2688 10877 2692
rect 10893 2748 10957 2752
rect 10893 2692 10897 2748
rect 10897 2692 10953 2748
rect 10953 2692 10957 2748
rect 10893 2688 10957 2692
rect 10973 2748 11037 2752
rect 10973 2692 10977 2748
rect 10977 2692 11033 2748
rect 11033 2692 11037 2748
rect 10973 2688 11037 2692
rect 11053 2748 11117 2752
rect 11053 2692 11057 2748
rect 11057 2692 11113 2748
rect 11113 2692 11117 2748
rect 11053 2688 11117 2692
rect 4660 2620 4724 2684
rect 9812 2620 9876 2684
rect 9996 2680 10060 2684
rect 9996 2624 10046 2680
rect 10046 2624 10060 2680
rect 9996 2620 10060 2624
rect 10180 2620 10244 2684
rect 6316 2484 6380 2548
rect 7236 2484 7300 2548
rect 7420 2544 7484 2548
rect 7420 2488 7470 2544
rect 7470 2488 7484 2544
rect 7420 2484 7484 2488
rect 7972 2544 8036 2548
rect 7972 2488 8022 2544
rect 8022 2488 8036 2544
rect 7972 2484 8036 2488
rect 11468 2484 11532 2548
rect 13124 2348 13188 2412
rect 6500 2212 6564 2276
rect 12572 2212 12636 2276
rect 3417 2204 3481 2208
rect 3417 2148 3421 2204
rect 3421 2148 3477 2204
rect 3477 2148 3481 2204
rect 3417 2144 3481 2148
rect 3497 2204 3561 2208
rect 3497 2148 3501 2204
rect 3501 2148 3557 2204
rect 3557 2148 3561 2204
rect 3497 2144 3561 2148
rect 3577 2204 3641 2208
rect 3577 2148 3581 2204
rect 3581 2148 3637 2204
rect 3637 2148 3641 2204
rect 3577 2144 3641 2148
rect 3657 2204 3721 2208
rect 3657 2148 3661 2204
rect 3661 2148 3717 2204
rect 3717 2148 3721 2204
rect 3657 2144 3721 2148
rect 8348 2204 8412 2208
rect 8348 2148 8352 2204
rect 8352 2148 8408 2204
rect 8408 2148 8412 2204
rect 8348 2144 8412 2148
rect 8428 2204 8492 2208
rect 8428 2148 8432 2204
rect 8432 2148 8488 2204
rect 8488 2148 8492 2204
rect 8428 2144 8492 2148
rect 8508 2204 8572 2208
rect 8508 2148 8512 2204
rect 8512 2148 8568 2204
rect 8568 2148 8572 2204
rect 8508 2144 8572 2148
rect 8588 2204 8652 2208
rect 8588 2148 8592 2204
rect 8592 2148 8648 2204
rect 8648 2148 8652 2204
rect 8588 2144 8652 2148
rect 13278 2204 13342 2208
rect 13278 2148 13282 2204
rect 13282 2148 13338 2204
rect 13338 2148 13342 2204
rect 13278 2144 13342 2148
rect 13358 2204 13422 2208
rect 13358 2148 13362 2204
rect 13362 2148 13418 2204
rect 13418 2148 13422 2204
rect 13358 2144 13422 2148
rect 13438 2204 13502 2208
rect 13438 2148 13442 2204
rect 13442 2148 13498 2204
rect 13498 2148 13502 2204
rect 13438 2144 13502 2148
rect 13518 2204 13582 2208
rect 13518 2148 13522 2204
rect 13522 2148 13578 2204
rect 13578 2148 13582 2204
rect 13518 2144 13582 2148
rect 11652 2076 11716 2140
rect 8156 1940 8220 2004
rect 13676 1804 13740 1868
rect 8892 1668 8956 1732
rect 7052 1532 7116 1596
rect 7604 1532 7668 1596
rect 10548 1396 10612 1460
rect 14044 1396 14108 1460
rect 12756 1260 12820 1324
rect 12940 1260 13004 1324
rect 9444 1124 9508 1188
<< metal4 >>
rect 3409 17440 3729 17456
rect 3409 17376 3417 17440
rect 3481 17376 3497 17440
rect 3561 17376 3577 17440
rect 3641 17376 3657 17440
rect 3721 17376 3729 17440
rect 3409 16352 3729 17376
rect 5874 16896 6195 17456
rect 5874 16832 5882 16896
rect 5946 16832 5962 16896
rect 6026 16832 6042 16896
rect 6106 16832 6122 16896
rect 6186 16832 6195 16896
rect 5027 16828 5093 16829
rect 5027 16764 5028 16828
rect 5092 16764 5093 16828
rect 5027 16763 5093 16764
rect 4291 16420 4357 16421
rect 4291 16356 4292 16420
rect 4356 16356 4357 16420
rect 4291 16355 4357 16356
rect 3409 16288 3417 16352
rect 3481 16288 3497 16352
rect 3561 16288 3577 16352
rect 3641 16288 3657 16352
rect 3721 16288 3729 16352
rect 3003 15876 3069 15877
rect 3003 15812 3004 15876
rect 3068 15812 3069 15876
rect 3003 15811 3069 15812
rect 3006 14381 3066 15811
rect 3409 15264 3729 16288
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3187 15196 3253 15197
rect 3187 15132 3188 15196
rect 3252 15132 3253 15196
rect 3187 15131 3253 15132
rect 3003 14380 3069 14381
rect 3003 14316 3004 14380
rect 3068 14316 3069 14380
rect 3003 14315 3069 14316
rect 3190 13973 3250 15131
rect 3409 14176 3729 15200
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3187 13972 3253 13973
rect 3187 13908 3188 13972
rect 3252 13908 3253 13972
rect 3187 13907 3253 13908
rect 3190 12341 3250 13907
rect 3409 13088 3729 14112
rect 4294 13973 4354 16355
rect 4475 15332 4541 15333
rect 4475 15268 4476 15332
rect 4540 15268 4541 15332
rect 4475 15267 4541 15268
rect 4291 13972 4357 13973
rect 4291 13908 4292 13972
rect 4356 13908 4357 13972
rect 4291 13907 4357 13908
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3187 12340 3253 12341
rect 3187 12276 3188 12340
rect 3252 12276 3253 12340
rect 3187 12275 3253 12276
rect 3409 12000 3729 13024
rect 4107 13020 4173 13021
rect 4107 12956 4108 13020
rect 4172 12956 4173 13020
rect 4107 12955 4173 12956
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3187 11116 3253 11117
rect 3187 11052 3188 11116
rect 3252 11052 3253 11116
rect 3187 11051 3253 11052
rect 3003 10980 3069 10981
rect 3003 10916 3004 10980
rect 3068 10916 3069 10980
rect 3003 10915 3069 10916
rect 3006 10437 3066 10915
rect 3003 10436 3069 10437
rect 3003 10372 3004 10436
rect 3068 10372 3069 10436
rect 3003 10371 3069 10372
rect 3190 2957 3250 11051
rect 3409 10912 3729 11936
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 9824 3729 10848
rect 4110 10029 4170 12955
rect 4107 10028 4173 10029
rect 4107 9964 4108 10028
rect 4172 9964 4173 10028
rect 4107 9963 4173 9964
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 8736 3729 9760
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 7648 3729 8672
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 6560 3729 7584
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 5472 3729 6496
rect 4107 6084 4173 6085
rect 4107 6020 4108 6084
rect 4172 6020 4173 6084
rect 4107 6019 4173 6020
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 4384 3729 5408
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 3296 3729 4320
rect 4110 4181 4170 6019
rect 4291 4996 4357 4997
rect 4291 4932 4292 4996
rect 4356 4932 4357 4996
rect 4291 4931 4357 4932
rect 4107 4180 4173 4181
rect 4107 4116 4108 4180
rect 4172 4116 4173 4180
rect 4107 4115 4173 4116
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3187 2956 3253 2957
rect 3187 2892 3188 2956
rect 3252 2892 3253 2956
rect 3187 2891 3253 2892
rect 3409 2208 3729 3232
rect 4294 2957 4354 4931
rect 4478 3637 4538 15267
rect 4659 14788 4725 14789
rect 4659 14724 4660 14788
rect 4724 14724 4725 14788
rect 4659 14723 4725 14724
rect 4475 3636 4541 3637
rect 4475 3572 4476 3636
rect 4540 3572 4541 3636
rect 4475 3571 4541 3572
rect 4291 2956 4357 2957
rect 4291 2892 4292 2956
rect 4356 2892 4357 2956
rect 4291 2891 4357 2892
rect 4662 2685 4722 14723
rect 5030 13429 5090 16763
rect 5874 15808 6195 16832
rect 8340 17440 8660 17456
rect 8340 17376 8348 17440
rect 8412 17376 8428 17440
rect 8492 17376 8508 17440
rect 8572 17376 8588 17440
rect 8652 17376 8660 17440
rect 7787 16420 7853 16421
rect 7787 16356 7788 16420
rect 7852 16356 7853 16420
rect 7787 16355 7853 16356
rect 7603 16284 7669 16285
rect 7603 16220 7604 16284
rect 7668 16220 7669 16284
rect 7603 16219 7669 16220
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6195 15808
rect 5395 15740 5461 15741
rect 5395 15676 5396 15740
rect 5460 15676 5461 15740
rect 5395 15675 5461 15676
rect 5027 13428 5093 13429
rect 5027 13364 5028 13428
rect 5092 13364 5093 13428
rect 5027 13363 5093 13364
rect 5398 12613 5458 15675
rect 5874 14720 6195 15744
rect 6867 15468 6933 15469
rect 6867 15404 6868 15468
rect 6932 15404 6933 15468
rect 6867 15403 6933 15404
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6195 14720
rect 5874 13632 6195 14656
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6195 13632
rect 5395 12612 5461 12613
rect 5395 12548 5396 12612
rect 5460 12548 5461 12612
rect 5395 12547 5461 12548
rect 5398 11389 5458 12547
rect 5874 12544 6195 13568
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6195 12544
rect 5874 11456 6195 12480
rect 6870 12477 6930 15403
rect 7235 14788 7301 14789
rect 7235 14724 7236 14788
rect 7300 14724 7301 14788
rect 7235 14723 7301 14724
rect 6867 12476 6933 12477
rect 6867 12412 6868 12476
rect 6932 12412 6933 12476
rect 6867 12411 6933 12412
rect 6499 12068 6565 12069
rect 6499 12004 6500 12068
rect 6564 12004 6565 12068
rect 6499 12003 6565 12004
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6195 11456
rect 5395 11388 5461 11389
rect 5395 11324 5396 11388
rect 5460 11324 5461 11388
rect 5395 11323 5461 11324
rect 5395 10844 5461 10845
rect 5395 10780 5396 10844
rect 5460 10780 5461 10844
rect 5395 10779 5461 10780
rect 5398 3773 5458 10779
rect 5874 10368 6195 11392
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6195 10368
rect 5874 9280 6195 10304
rect 6502 10301 6562 12003
rect 7238 10845 7298 14723
rect 7235 10844 7301 10845
rect 7235 10780 7236 10844
rect 7300 10780 7301 10844
rect 7235 10779 7301 10780
rect 6499 10300 6565 10301
rect 6499 10236 6500 10300
rect 6564 10236 6565 10300
rect 6499 10235 6565 10236
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6195 9280
rect 5874 8192 6195 9216
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6195 8192
rect 5874 7104 6195 8128
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6195 7104
rect 5874 6016 6195 7040
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6195 6016
rect 5874 4928 6195 5952
rect 6315 5948 6381 5949
rect 6315 5884 6316 5948
rect 6380 5884 6381 5948
rect 6315 5883 6381 5884
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6195 4928
rect 5874 3840 6195 4864
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6195 3840
rect 5395 3772 5461 3773
rect 5395 3708 5396 3772
rect 5460 3708 5461 3772
rect 5395 3707 5461 3708
rect 5874 2752 6195 3776
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6195 2752
rect 4659 2684 4725 2685
rect 4659 2620 4660 2684
rect 4724 2620 4725 2684
rect 4659 2619 4725 2620
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2128 3729 2144
rect 5874 2128 6195 2688
rect 6318 2549 6378 5883
rect 6315 2548 6381 2549
rect 6315 2484 6316 2548
rect 6380 2484 6381 2548
rect 6315 2483 6381 2484
rect 6502 2277 6562 10235
rect 6683 10028 6749 10029
rect 6683 9964 6684 10028
rect 6748 9964 6749 10028
rect 6683 9963 6749 9964
rect 6686 2821 6746 9963
rect 6867 8668 6933 8669
rect 6867 8604 6868 8668
rect 6932 8604 6933 8668
rect 6867 8603 6933 8604
rect 6870 3909 6930 8603
rect 7235 8396 7301 8397
rect 7235 8332 7236 8396
rect 7300 8332 7301 8396
rect 7235 8331 7301 8332
rect 7051 4860 7117 4861
rect 7051 4796 7052 4860
rect 7116 4796 7117 4860
rect 7051 4795 7117 4796
rect 6867 3908 6933 3909
rect 6867 3844 6868 3908
rect 6932 3844 6933 3908
rect 6867 3843 6933 3844
rect 6683 2820 6749 2821
rect 6683 2756 6684 2820
rect 6748 2756 6749 2820
rect 6683 2755 6749 2756
rect 6499 2276 6565 2277
rect 6499 2212 6500 2276
rect 6564 2212 6565 2276
rect 6499 2211 6565 2212
rect 7054 1597 7114 4795
rect 7238 2549 7298 8331
rect 7419 8260 7485 8261
rect 7419 8196 7420 8260
rect 7484 8196 7485 8260
rect 7419 8195 7485 8196
rect 7422 2549 7482 8195
rect 7606 4181 7666 16219
rect 7790 12069 7850 16355
rect 8340 16352 8660 17376
rect 10805 16896 11125 17456
rect 13270 17440 13590 17456
rect 13270 17376 13278 17440
rect 13342 17376 13358 17440
rect 13422 17376 13438 17440
rect 13502 17376 13518 17440
rect 13582 17376 13590 17440
rect 12755 17100 12821 17101
rect 12755 17036 12756 17100
rect 12820 17036 12821 17100
rect 12755 17035 12821 17036
rect 12203 16964 12269 16965
rect 12203 16900 12204 16964
rect 12268 16900 12269 16964
rect 12203 16899 12269 16900
rect 10805 16832 10813 16896
rect 10877 16832 10893 16896
rect 10957 16832 10973 16896
rect 11037 16832 11053 16896
rect 11117 16832 11125 16896
rect 9259 16692 9325 16693
rect 9259 16628 9260 16692
rect 9324 16628 9325 16692
rect 9259 16627 9325 16628
rect 8340 16288 8348 16352
rect 8412 16288 8428 16352
rect 8492 16288 8508 16352
rect 8572 16288 8588 16352
rect 8652 16288 8660 16352
rect 8340 15264 8660 16288
rect 9262 15469 9322 16627
rect 9443 15876 9509 15877
rect 9443 15812 9444 15876
rect 9508 15812 9509 15876
rect 9443 15811 9509 15812
rect 10179 15876 10245 15877
rect 10179 15812 10180 15876
rect 10244 15812 10245 15876
rect 10179 15811 10245 15812
rect 8891 15468 8957 15469
rect 8891 15404 8892 15468
rect 8956 15404 8957 15468
rect 8891 15403 8957 15404
rect 9259 15468 9325 15469
rect 9259 15404 9260 15468
rect 9324 15404 9325 15468
rect 9259 15403 9325 15404
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 14176 8660 15200
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8155 13156 8221 13157
rect 8155 13092 8156 13156
rect 8220 13092 8221 13156
rect 8155 13091 8221 13092
rect 7787 12068 7853 12069
rect 7787 12004 7788 12068
rect 7852 12004 7853 12068
rect 7787 12003 7853 12004
rect 8158 10437 8218 13091
rect 8340 13088 8660 14112
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 12000 8660 13024
rect 8894 13021 8954 15403
rect 9075 14788 9141 14789
rect 9075 14724 9076 14788
rect 9140 14724 9141 14788
rect 9075 14723 9141 14724
rect 8891 13020 8957 13021
rect 8891 12956 8892 13020
rect 8956 12956 8957 13020
rect 8891 12955 8957 12956
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 10912 8660 11936
rect 8891 11932 8957 11933
rect 8891 11868 8892 11932
rect 8956 11868 8957 11932
rect 8891 11867 8957 11868
rect 8894 11661 8954 11867
rect 8891 11660 8957 11661
rect 8891 11596 8892 11660
rect 8956 11596 8957 11660
rect 8891 11595 8957 11596
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8155 10436 8221 10437
rect 8155 10372 8156 10436
rect 8220 10372 8221 10436
rect 8155 10371 8221 10372
rect 8340 9824 8660 10848
rect 9078 9893 9138 14723
rect 9259 14108 9325 14109
rect 9259 14044 9260 14108
rect 9324 14044 9325 14108
rect 9259 14043 9325 14044
rect 9075 9892 9141 9893
rect 9075 9828 9076 9892
rect 9140 9828 9141 9892
rect 9075 9827 9141 9828
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 7971 9076 8037 9077
rect 7971 9012 7972 9076
rect 8036 9012 8037 9076
rect 7971 9011 8037 9012
rect 7787 5268 7853 5269
rect 7787 5204 7788 5268
rect 7852 5204 7853 5268
rect 7787 5203 7853 5204
rect 7603 4180 7669 4181
rect 7603 4116 7604 4180
rect 7668 4116 7669 4180
rect 7603 4115 7669 4116
rect 7790 2957 7850 5203
rect 7603 2956 7669 2957
rect 7603 2892 7604 2956
rect 7668 2892 7669 2956
rect 7603 2891 7669 2892
rect 7787 2956 7853 2957
rect 7787 2892 7788 2956
rect 7852 2892 7853 2956
rect 7787 2891 7853 2892
rect 7235 2548 7301 2549
rect 7235 2484 7236 2548
rect 7300 2484 7301 2548
rect 7235 2483 7301 2484
rect 7419 2548 7485 2549
rect 7419 2484 7420 2548
rect 7484 2484 7485 2548
rect 7419 2483 7485 2484
rect 7606 1597 7666 2891
rect 7974 2549 8034 9011
rect 8340 8736 8660 9760
rect 9262 9757 9322 14043
rect 9446 10165 9506 15811
rect 9811 15468 9877 15469
rect 9811 15404 9812 15468
rect 9876 15404 9877 15468
rect 9811 15403 9877 15404
rect 9995 15468 10061 15469
rect 9995 15404 9996 15468
rect 10060 15404 10061 15468
rect 9995 15403 10061 15404
rect 9627 15196 9693 15197
rect 9627 15132 9628 15196
rect 9692 15132 9693 15196
rect 9627 15131 9693 15132
rect 9630 11661 9690 15131
rect 9814 13973 9874 15403
rect 9811 13972 9877 13973
rect 9811 13908 9812 13972
rect 9876 13908 9877 13972
rect 9811 13907 9877 13908
rect 9811 12476 9877 12477
rect 9811 12412 9812 12476
rect 9876 12412 9877 12476
rect 9811 12411 9877 12412
rect 9627 11660 9693 11661
rect 9627 11596 9628 11660
rect 9692 11596 9693 11660
rect 9627 11595 9693 11596
rect 9814 11114 9874 12411
rect 9998 11794 10058 15403
rect 10182 13698 10242 15811
rect 10805 15808 11125 16832
rect 11467 16420 11533 16421
rect 11467 16356 11468 16420
rect 11532 16356 11533 16420
rect 11467 16355 11533 16356
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10363 15468 10429 15469
rect 10363 15404 10364 15468
rect 10428 15404 10429 15468
rect 10363 15403 10429 15404
rect 10182 13638 10288 13698
rect 10228 13290 10288 13638
rect 10182 13230 10288 13290
rect 10182 13021 10242 13230
rect 10179 13020 10245 13021
rect 10179 12956 10180 13020
rect 10244 12956 10245 13020
rect 10179 12955 10245 12956
rect 9998 11734 10242 11794
rect 9995 11660 10061 11661
rect 9995 11596 9996 11660
rect 10060 11596 10061 11660
rect 9995 11595 10061 11596
rect 9630 11054 9874 11114
rect 9630 10437 9690 11054
rect 9998 10842 10058 11595
rect 10182 11117 10242 11734
rect 10179 11116 10245 11117
rect 10179 11052 10180 11116
rect 10244 11052 10245 11116
rect 10179 11051 10245 11052
rect 9998 10782 10242 10842
rect 9811 10572 9877 10573
rect 9811 10508 9812 10572
rect 9876 10508 9877 10572
rect 9811 10507 9877 10508
rect 9627 10436 9693 10437
rect 9627 10372 9628 10436
rect 9692 10372 9693 10436
rect 9627 10371 9693 10372
rect 9627 10300 9693 10301
rect 9627 10236 9628 10300
rect 9692 10236 9693 10300
rect 9627 10235 9693 10236
rect 9443 10164 9509 10165
rect 9443 10100 9444 10164
rect 9508 10100 9509 10164
rect 9443 10099 9509 10100
rect 9259 9756 9325 9757
rect 9259 9692 9260 9756
rect 9324 9692 9325 9756
rect 9259 9691 9325 9692
rect 9075 8804 9141 8805
rect 9075 8740 9076 8804
rect 9140 8740 9141 8804
rect 9075 8739 9141 8740
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8340 7648 8660 8672
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 6560 8660 7584
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8155 5812 8221 5813
rect 8155 5748 8156 5812
rect 8220 5748 8221 5812
rect 8155 5747 8221 5748
rect 7971 2548 8037 2549
rect 7971 2484 7972 2548
rect 8036 2484 8037 2548
rect 7971 2483 8037 2484
rect 8158 2005 8218 5747
rect 8340 5472 8660 6496
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 4384 8660 5408
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 3296 8660 4320
rect 8891 4316 8957 4317
rect 8891 4252 8892 4316
rect 8956 4252 8957 4316
rect 8891 4251 8957 4252
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 2208 8660 3232
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2128 8660 2144
rect 8155 2004 8221 2005
rect 8155 1940 8156 2004
rect 8220 1940 8221 2004
rect 8155 1939 8221 1940
rect 8894 1733 8954 4251
rect 9078 3501 9138 8739
rect 9259 7580 9325 7581
rect 9259 7516 9260 7580
rect 9324 7516 9325 7580
rect 9259 7515 9325 7516
rect 9262 7173 9322 7515
rect 9259 7172 9325 7173
rect 9259 7108 9260 7172
rect 9324 7108 9325 7172
rect 9259 7107 9325 7108
rect 9262 5946 9322 7107
rect 9630 6085 9690 10235
rect 9627 6084 9693 6085
rect 9627 6020 9628 6084
rect 9692 6020 9693 6084
rect 9627 6019 9693 6020
rect 9262 5886 9690 5946
rect 9443 5268 9509 5269
rect 9443 5204 9444 5268
rect 9508 5204 9509 5268
rect 9443 5203 9509 5204
rect 9446 4861 9506 5203
rect 9443 4860 9509 4861
rect 9443 4796 9444 4860
rect 9508 4796 9509 4860
rect 9443 4795 9509 4796
rect 9259 4452 9325 4453
rect 9259 4388 9260 4452
rect 9324 4388 9325 4452
rect 9259 4387 9325 4388
rect 9262 3634 9322 4387
rect 9262 3574 9368 3634
rect 9075 3500 9141 3501
rect 9075 3436 9076 3500
rect 9140 3436 9141 3500
rect 9308 3498 9368 3574
rect 9308 3438 9506 3498
rect 9075 3435 9141 3436
rect 8891 1732 8957 1733
rect 8891 1668 8892 1732
rect 8956 1668 8957 1732
rect 8891 1667 8957 1668
rect 7051 1596 7117 1597
rect 7051 1532 7052 1596
rect 7116 1532 7117 1596
rect 7051 1531 7117 1532
rect 7603 1596 7669 1597
rect 7603 1532 7604 1596
rect 7668 1532 7669 1596
rect 7603 1531 7669 1532
rect 9446 1189 9506 3438
rect 9630 3093 9690 5886
rect 9627 3092 9693 3093
rect 9627 3028 9628 3092
rect 9692 3028 9693 3092
rect 9627 3027 9693 3028
rect 9814 2821 9874 10507
rect 9995 8260 10061 8261
rect 9995 8196 9996 8260
rect 10060 8196 10061 8260
rect 9995 8195 10061 8196
rect 9998 4725 10058 8195
rect 10182 7717 10242 10782
rect 10179 7716 10245 7717
rect 10179 7652 10180 7716
rect 10244 7652 10245 7716
rect 10179 7651 10245 7652
rect 10182 4861 10242 7651
rect 10366 5677 10426 15403
rect 10805 14720 11125 15744
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10547 14652 10613 14653
rect 10547 14588 10548 14652
rect 10612 14588 10613 14652
rect 10547 14587 10613 14588
rect 10550 12069 10610 14587
rect 10805 13632 11125 14656
rect 11470 13701 11530 16355
rect 11835 15332 11901 15333
rect 11835 15268 11836 15332
rect 11900 15268 11901 15332
rect 11835 15267 11901 15268
rect 11651 15196 11717 15197
rect 11651 15132 11652 15196
rect 11716 15132 11717 15196
rect 11651 15131 11717 15132
rect 11467 13700 11533 13701
rect 11467 13636 11468 13700
rect 11532 13636 11533 13700
rect 11467 13635 11533 13636
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10805 12544 11125 13568
rect 11283 13020 11349 13021
rect 11283 12956 11284 13020
rect 11348 12956 11349 13020
rect 11283 12955 11349 12956
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10547 12068 10613 12069
rect 10547 12004 10548 12068
rect 10612 12004 10613 12068
rect 10547 12003 10613 12004
rect 10805 11456 11125 12480
rect 11286 11525 11346 12955
rect 11283 11524 11349 11525
rect 11283 11460 11284 11524
rect 11348 11460 11349 11524
rect 11283 11459 11349 11460
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10547 11388 10613 11389
rect 10547 11324 10548 11388
rect 10612 11324 10613 11388
rect 10547 11323 10613 11324
rect 10363 5676 10429 5677
rect 10363 5612 10364 5676
rect 10428 5612 10429 5676
rect 10363 5611 10429 5612
rect 10363 5540 10429 5541
rect 10363 5476 10364 5540
rect 10428 5476 10429 5540
rect 10363 5475 10429 5476
rect 10179 4860 10245 4861
rect 10179 4796 10180 4860
rect 10244 4796 10245 4860
rect 10179 4795 10245 4796
rect 9995 4724 10061 4725
rect 9995 4660 9996 4724
rect 10060 4660 10061 4724
rect 9995 4659 10061 4660
rect 9811 2820 9877 2821
rect 9811 2756 9812 2820
rect 9876 2756 9877 2820
rect 9811 2755 9877 2756
rect 9998 2685 10058 4659
rect 10182 2685 10242 4795
rect 10366 4181 10426 5475
rect 10363 4180 10429 4181
rect 10363 4116 10364 4180
rect 10428 4116 10429 4180
rect 10363 4115 10429 4116
rect 10363 3908 10429 3909
rect 10363 3844 10364 3908
rect 10428 3844 10429 3908
rect 10363 3843 10429 3844
rect 9811 2684 9877 2685
rect 9811 2620 9812 2684
rect 9876 2620 9877 2684
rect 9811 2619 9877 2620
rect 9995 2684 10061 2685
rect 9995 2620 9996 2684
rect 10060 2620 10061 2684
rect 9995 2619 10061 2620
rect 10179 2684 10245 2685
rect 10179 2620 10180 2684
rect 10244 2620 10245 2684
rect 10179 2619 10245 2620
rect 9814 2546 9874 2619
rect 10366 2546 10426 3843
rect 9814 2486 10426 2546
rect 10550 1461 10610 11323
rect 10805 10368 11125 11392
rect 11283 11388 11349 11389
rect 11283 11324 11284 11388
rect 11348 11324 11349 11388
rect 11283 11323 11349 11324
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10805 9280 11125 10304
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 8192 11125 9216
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 7104 11125 8128
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 6016 11125 7040
rect 11286 6765 11346 11323
rect 11470 9213 11530 13635
rect 11654 13157 11714 15131
rect 11651 13156 11717 13157
rect 11651 13092 11652 13156
rect 11716 13092 11717 13156
rect 11651 13091 11717 13092
rect 11651 11796 11717 11797
rect 11651 11732 11652 11796
rect 11716 11732 11717 11796
rect 11651 11731 11717 11732
rect 11467 9212 11533 9213
rect 11467 9148 11468 9212
rect 11532 9148 11533 9212
rect 11467 9147 11533 9148
rect 11283 6764 11349 6765
rect 11283 6700 11284 6764
rect 11348 6700 11349 6764
rect 11283 6699 11349 6700
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 4928 11125 5952
rect 11286 5130 11346 6699
rect 11286 5070 11530 5130
rect 11283 4996 11349 4997
rect 11283 4932 11284 4996
rect 11348 4932 11349 4996
rect 11283 4931 11349 4932
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 3840 11125 4864
rect 11286 4453 11346 4931
rect 11283 4452 11349 4453
rect 11283 4388 11284 4452
rect 11348 4388 11349 4452
rect 11283 4387 11349 4388
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10805 2752 11125 3776
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10805 2128 11125 2688
rect 11470 2549 11530 5070
rect 11654 4589 11714 11731
rect 11651 4588 11717 4589
rect 11651 4524 11652 4588
rect 11716 4524 11717 4588
rect 11651 4523 11717 4524
rect 11651 4452 11717 4453
rect 11651 4388 11652 4452
rect 11716 4388 11717 4452
rect 11651 4387 11717 4388
rect 11467 2548 11533 2549
rect 11467 2484 11468 2548
rect 11532 2484 11533 2548
rect 11467 2483 11533 2484
rect 11654 2141 11714 4387
rect 11838 4045 11898 15267
rect 12019 15060 12085 15061
rect 12019 14996 12020 15060
rect 12084 14996 12085 15060
rect 12019 14995 12085 14996
rect 12022 14517 12082 14995
rect 12019 14516 12085 14517
rect 12019 14452 12020 14516
rect 12084 14452 12085 14516
rect 12019 14451 12085 14452
rect 12206 14378 12266 16899
rect 12758 16557 12818 17035
rect 13123 16692 13189 16693
rect 13123 16628 13124 16692
rect 13188 16628 13189 16692
rect 13123 16627 13189 16628
rect 12755 16556 12821 16557
rect 12755 16492 12756 16556
rect 12820 16492 12821 16556
rect 12755 16491 12821 16492
rect 12571 15740 12637 15741
rect 12571 15676 12572 15740
rect 12636 15676 12637 15740
rect 12571 15675 12637 15676
rect 12387 15604 12453 15605
rect 12387 15540 12388 15604
rect 12452 15540 12453 15604
rect 12387 15539 12453 15540
rect 12022 14318 12266 14378
rect 12022 13429 12082 14318
rect 12019 13428 12085 13429
rect 12019 13364 12020 13428
rect 12084 13364 12085 13428
rect 12019 13363 12085 13364
rect 12203 13428 12269 13429
rect 12203 13364 12204 13428
rect 12268 13364 12269 13428
rect 12203 13363 12269 13364
rect 12022 8805 12082 13363
rect 12019 8804 12085 8805
rect 12019 8740 12020 8804
rect 12084 8740 12085 8804
rect 12019 8739 12085 8740
rect 12019 8668 12085 8669
rect 12019 8604 12020 8668
rect 12084 8604 12085 8668
rect 12019 8603 12085 8604
rect 12022 4453 12082 8603
rect 12019 4452 12085 4453
rect 12019 4388 12020 4452
rect 12084 4388 12085 4452
rect 12019 4387 12085 4388
rect 11835 4044 11901 4045
rect 11835 3980 11836 4044
rect 11900 3980 11901 4044
rect 11835 3979 11901 3980
rect 12022 3637 12082 4387
rect 11835 3636 11901 3637
rect 11835 3572 11836 3636
rect 11900 3572 11901 3636
rect 11835 3571 11901 3572
rect 12019 3636 12085 3637
rect 12019 3572 12020 3636
rect 12084 3572 12085 3636
rect 12019 3571 12085 3572
rect 11838 3365 11898 3571
rect 11835 3364 11901 3365
rect 11835 3300 11836 3364
rect 11900 3300 11901 3364
rect 11835 3299 11901 3300
rect 12206 2821 12266 13363
rect 12390 12341 12450 15539
rect 12574 13565 12634 15675
rect 12571 13564 12637 13565
rect 12571 13500 12572 13564
rect 12636 13500 12637 13564
rect 12571 13499 12637 13500
rect 12571 13428 12637 13429
rect 12571 13364 12572 13428
rect 12636 13364 12637 13428
rect 12571 13363 12637 13364
rect 12387 12340 12453 12341
rect 12387 12276 12388 12340
rect 12452 12276 12453 12340
rect 12387 12275 12453 12276
rect 12387 10980 12453 10981
rect 12387 10916 12388 10980
rect 12452 10916 12453 10980
rect 12387 10915 12453 10916
rect 12390 8261 12450 10915
rect 12574 10573 12634 13363
rect 12758 11389 12818 16491
rect 12939 14516 13005 14517
rect 12939 14452 12940 14516
rect 13004 14452 13005 14516
rect 12939 14451 13005 14452
rect 12755 11388 12821 11389
rect 12755 11324 12756 11388
rect 12820 11324 12821 11388
rect 12755 11323 12821 11324
rect 12942 10709 13002 14451
rect 12939 10708 13005 10709
rect 12939 10644 12940 10708
rect 13004 10644 13005 10708
rect 12939 10643 13005 10644
rect 12571 10572 12637 10573
rect 12571 10508 12572 10572
rect 12636 10508 12637 10572
rect 12571 10507 12637 10508
rect 12939 10572 13005 10573
rect 12939 10508 12940 10572
rect 13004 10508 13005 10572
rect 12939 10507 13005 10508
rect 12942 9754 13002 10507
rect 12758 9694 13002 9754
rect 12571 8940 12637 8941
rect 12571 8876 12572 8940
rect 12636 8876 12637 8940
rect 12571 8875 12637 8876
rect 12387 8260 12453 8261
rect 12387 8196 12388 8260
rect 12452 8196 12453 8260
rect 12387 8195 12453 8196
rect 12387 6492 12453 6493
rect 12387 6428 12388 6492
rect 12452 6428 12453 6492
rect 12387 6427 12453 6428
rect 12390 3093 12450 6427
rect 12574 4181 12634 8875
rect 12758 7989 12818 9694
rect 12939 9484 13005 9485
rect 12939 9420 12940 9484
rect 13004 9420 13005 9484
rect 12939 9419 13005 9420
rect 12755 7988 12821 7989
rect 12755 7924 12756 7988
rect 12820 7924 12821 7988
rect 12755 7923 12821 7924
rect 12755 7852 12821 7853
rect 12755 7788 12756 7852
rect 12820 7788 12821 7852
rect 12755 7787 12821 7788
rect 12758 4997 12818 7787
rect 12755 4996 12821 4997
rect 12755 4932 12756 4996
rect 12820 4932 12821 4996
rect 12755 4931 12821 4932
rect 12755 4588 12821 4589
rect 12755 4524 12756 4588
rect 12820 4524 12821 4588
rect 12755 4523 12821 4524
rect 12571 4180 12637 4181
rect 12571 4116 12572 4180
rect 12636 4116 12637 4180
rect 12571 4115 12637 4116
rect 12758 4042 12818 4523
rect 12574 3982 12818 4042
rect 12387 3092 12453 3093
rect 12387 3028 12388 3092
rect 12452 3028 12453 3092
rect 12387 3027 12453 3028
rect 12203 2820 12269 2821
rect 12203 2756 12204 2820
rect 12268 2756 12269 2820
rect 12203 2755 12269 2756
rect 12574 2277 12634 3982
rect 12755 3636 12821 3637
rect 12755 3572 12756 3636
rect 12820 3572 12821 3636
rect 12755 3571 12821 3572
rect 12571 2276 12637 2277
rect 12571 2212 12572 2276
rect 12636 2212 12637 2276
rect 12571 2211 12637 2212
rect 11651 2140 11717 2141
rect 11651 2076 11652 2140
rect 11716 2076 11717 2140
rect 11651 2075 11717 2076
rect 10547 1460 10613 1461
rect 10547 1396 10548 1460
rect 10612 1396 10613 1460
rect 10547 1395 10613 1396
rect 12758 1325 12818 3571
rect 12942 1325 13002 9419
rect 13126 6901 13186 16627
rect 13270 16352 13590 17376
rect 13270 16288 13278 16352
rect 13342 16288 13358 16352
rect 13422 16288 13438 16352
rect 13502 16288 13518 16352
rect 13582 16288 13590 16352
rect 13270 15264 13590 16288
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13270 14176 13590 15200
rect 13675 14380 13741 14381
rect 13675 14316 13676 14380
rect 13740 14316 13741 14380
rect 13675 14315 13741 14316
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 13088 13590 14112
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 12000 13590 13024
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 10912 13590 11936
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 9824 13590 10848
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 13270 8736 13590 9760
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 7648 13590 8672
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13123 6900 13189 6901
rect 13123 6836 13124 6900
rect 13188 6836 13189 6900
rect 13123 6835 13189 6836
rect 13270 6560 13590 7584
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 5472 13590 6496
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 4384 13590 5408
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13123 4180 13189 4181
rect 13123 4116 13124 4180
rect 13188 4116 13189 4180
rect 13123 4115 13189 4116
rect 13126 2413 13186 4115
rect 13270 3296 13590 4320
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 13123 2412 13189 2413
rect 13123 2348 13124 2412
rect 13188 2348 13189 2412
rect 13123 2347 13189 2348
rect 13270 2208 13590 3232
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2128 13590 2144
rect 13678 1869 13738 14315
rect 14043 13428 14109 13429
rect 14043 13364 14044 13428
rect 14108 13364 14109 13428
rect 14043 13363 14109 13364
rect 13859 13020 13925 13021
rect 13859 12956 13860 13020
rect 13924 12956 13925 13020
rect 13859 12955 13925 12956
rect 13862 11525 13922 12955
rect 13859 11524 13925 11525
rect 13859 11460 13860 11524
rect 13924 11460 13925 11524
rect 13859 11459 13925 11460
rect 14046 10573 14106 13363
rect 14227 11524 14293 11525
rect 14227 11460 14228 11524
rect 14292 11460 14293 11524
rect 14227 11459 14293 11460
rect 14043 10572 14109 10573
rect 14043 10508 14044 10572
rect 14108 10508 14109 10572
rect 14043 10507 14109 10508
rect 14230 10437 14290 11459
rect 14227 10436 14293 10437
rect 14227 10372 14228 10436
rect 14292 10372 14293 10436
rect 14227 10371 14293 10372
rect 14043 9620 14109 9621
rect 14043 9556 14044 9620
rect 14108 9556 14109 9620
rect 14043 9555 14109 9556
rect 13859 9348 13925 9349
rect 13859 9284 13860 9348
rect 13924 9284 13925 9348
rect 13859 9283 13925 9284
rect 13862 3637 13922 9283
rect 14046 5949 14106 9555
rect 14230 7309 14290 10371
rect 14227 7308 14293 7309
rect 14227 7244 14228 7308
rect 14292 7244 14293 7308
rect 14227 7243 14293 7244
rect 14043 5948 14109 5949
rect 14043 5884 14044 5948
rect 14108 5884 14109 5948
rect 14043 5883 14109 5884
rect 14043 4860 14109 4861
rect 14043 4796 14044 4860
rect 14108 4796 14109 4860
rect 14043 4795 14109 4796
rect 13859 3636 13925 3637
rect 13859 3572 13860 3636
rect 13924 3572 13925 3636
rect 13859 3571 13925 3572
rect 13675 1868 13741 1869
rect 13675 1804 13676 1868
rect 13740 1804 13741 1868
rect 13675 1803 13741 1804
rect 14046 1461 14106 4795
rect 14043 1460 14109 1461
rect 14043 1396 14044 1460
rect 14108 1396 14109 1460
rect 14043 1395 14109 1396
rect 12755 1324 12821 1325
rect 12755 1260 12756 1324
rect 12820 1260 12821 1324
rect 12755 1259 12821 1260
rect 12939 1324 13005 1325
rect 12939 1260 12940 1324
rect 13004 1260 13005 1324
rect 12939 1259 13005 1260
rect 9443 1188 9509 1189
rect 9443 1124 9444 1188
rect 9508 1124 9509 1188
rect 9443 1123 9509 1124
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 2852 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2852 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1606821651
transform 1 0 1564 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606821651
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14
timestamp 1606821651
transform 1 0 2392 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _21_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3680 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 4048 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_1_
timestamp 1606821651
transform 1 0 4324 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1606821651
transform 1 0 3496 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1606821651
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1606821651
transform 1 0 5520 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 5980 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1606821651
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1606821651
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6348 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1606821651
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_1_
timestamp 1606821651
transform 1 0 8188 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 8556 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1606821651
transform 1 0 7636 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72
timestamp 1606821651
transform 1 0 7728 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76
timestamp 1606821651
transform 1 0 8096 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_80
timestamp 1606821651
transform 1 0 8464 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_1_
timestamp 1606821651
transform 1 0 9200 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1606821651
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1606821651
transform 1 0 10396 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1606821651
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 9384 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_86
timestamp 1606821651
transform 1 0 9016 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103
timestamp 1606821651
transform 1 0 10580 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_87
timestamp 1606821651
transform 1 0 9108 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_97
timestamp 1606821651
transform 1 0 10028 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 11776 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1606821651
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1606821651
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1606821651
transform 1 0 11224 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1606821651
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1606821651
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1606821651
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_119
timestamp 1606821651
transform 1 0 12052 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 13616 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 13524 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1606821651
transform 1 0 14444 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_131
timestamp 1606821651
transform 1 0 13156 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1606821651
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_132
timestamp 1606821651
transform 1 0 13248 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_142
timestamp 1606821651
transform 1 0 14168 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1606821651
transform 1 0 14536 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606821651
transform -1 0 15824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606821651
transform -1 0 15824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1606821651
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 15272 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151
timestamp 1606821651
transform 1 0 14996 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156
timestamp 1606821651
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_150
timestamp 1606821651
transform 1 0 14904 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 1380 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1606821651
transform 1 0 2852 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606821651
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1606821651
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_28
timestamp 1606821651
transform 1 0 3680 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_41
timestamp 1606821651
transform 1 0 4876 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_2_
timestamp 1606821651
transform 1 0 4968 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5796 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6624 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1606821651
transform 1 0 7452 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1606821651
transform 1 0 8280 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1606821651
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_87
timestamp 1606821651
transform 1 0 9108 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1606821651
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_102
timestamp 1606821651
transform 1 0 10488 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1606821651
transform 1 0 11684 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1606821651
transform 1 0 10856 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1606821651
transform 1 0 12052 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1606821651
transform 1 0 14444 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13248 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_128
timestamp 1606821651
transform 1 0 12880 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1606821651
transform 1 0 14076 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606821651
transform -1 0 15824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1606821651
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1606821651
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_154
timestamp 1606821651
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2576 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1606821651
transform 1 0 1564 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606821651
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1606821651
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_14
timestamp 1606821651
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 4876 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1606821651
transform 1 0 4048 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1606821651
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5520 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1606821651
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_47
timestamp 1606821651
transform 1 0 5428 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1606821651
transform 1 0 6348 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1606821651
transform 1 0 8004 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_71
timestamp 1606821651
transform 1 0 7636 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_2_
timestamp 1606821651
transform 1 0 10396 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1606821651
transform 1 0 8832 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 10028 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_93
timestamp 1606821651
transform 1 0 9660 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_100
timestamp 1606821651
transform 1 0 10304 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1606821651
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1606821651
transform 1 0 11224 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606821651
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp 1606821651
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1606821651
transform 1 0 13616 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_132
timestamp 1606821651
transform 1 0 13248 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_145
timestamp 1606821651
transform 1 0 14444 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1606821651
transform 1 0 14812 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606821651
transform -1 0 15824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_153
timestamp 1606821651
transform 1 0 15180 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 1380 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1606821651
transform 1 0 2852 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606821651
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606821651
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_28
timestamp 1606821651
transform 1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_41
timestamp 1606821651
transform 1 0 4876 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6440 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1606821651
transform 1 0 5244 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_54
timestamp 1606821651
transform 1 0 6072 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1606821651
transform 1 0 8280 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_74
timestamp 1606821651
transform 1 0 7912 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1606821651
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606821651
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_87
timestamp 1606821651
transform 1 0 9108 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1606821651
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_102
timestamp 1606821651
transform 1 0 10488 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10856 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12052 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_115
timestamp 1606821651
transform 1 0 11684 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1606821651
transform 1 0 14444 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1606821651
transform 1 0 13248 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_128
timestamp 1606821651
transform 1 0 12880 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1606821651
transform 1 0 14076 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606821651
transform -1 0 15824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606821651
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1606821651
transform 1 0 14812 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1606821651
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1606821651
transform 1 0 1380 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1606821651
transform 1 0 2484 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606821651
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_12
timestamp 1606821651
transform 1 0 2208 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 4876 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1606821651
transform 1 0 3680 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_24
timestamp 1606821651
transform 1 0 3312 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_37
timestamp 1606821651
transform 1 0 4508 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606821651
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1606821651
transform 1 0 6348 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_62 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6808 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7360 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1606821651
transform 1 0 9200 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1606821651
transform 1 0 10396 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_84
timestamp 1606821651
transform 1 0 8832 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_97
timestamp 1606821651
transform 1 0 10028 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1606821651
transform 1 0 11592 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l4_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606821651
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_110
timestamp 1606821651
transform 1 0 11224 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1606821651
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1606821651
transform 1 0 13616 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_132
timestamp 1606821651
transform 1 0 13248 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_145
timestamp 1606821651
transform 1 0 14444 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1606821651
transform 1 0 14812 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606821651
transform -1 0 15824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_153
timestamp 1606821651
transform 1 0 15180 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1606821651
transform 1 0 1748 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1606821651
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606821651
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606821651
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1606821651
transform 1 0 1564 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1606821651
transform 1 0 1840 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1606821651
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_17
timestamp 1606821651
transform 1 0 2668 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_14
timestamp 1606821651
transform 1 0 2392 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1606821651
transform 1 0 2760 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 4876 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 3036 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1606821651
transform 1 0 4508 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606821651
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606821651
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1606821651
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_36
timestamp 1606821651
transform 1 0 4416 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_37
timestamp 1606821651
transform 1 0 4508 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 5704 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606821651
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_46
timestamp 1606821651
transform 1 0 5336 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1606821651
transform 1 0 6348 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 8648 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7636 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_66
timestamp 1606821651
transform 1 0 7176 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_70
timestamp 1606821651
transform 1 0 7544 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_78
timestamp 1606821651
transform 1 0 8280 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1606821651
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1606821651
transform 1 0 10488 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606821651
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_87
timestamp 1606821651
transform 1 0 9108 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1606821651
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_102
timestamp 1606821651
transform 1 0 10488 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_98
timestamp 1606821651
transform 1 0 10120 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1606821651
transform 1 0 11684 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1606821651
transform 1 0 10856 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12052 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1606821651
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606821651
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_115
timestamp 1606821651
transform 1 0 11684 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_111
timestamp 1606821651
transform 1 0 11316 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1606821651
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1606821651
transform 1 0 14444 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_3_
timestamp 1606821651
transform 1 0 13248 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_0_
timestamp 1606821651
transform 1 0 13616 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1606821651
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_128
timestamp 1606821651
transform 1 0 12880 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp 1606821651
transform 1 0 14076 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_134
timestamp 1606821651
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_145
timestamp 1606821651
transform 1 0 14444 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1606821651
transform 1 0 14812 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606821651
transform -1 0 15824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606821651
transform -1 0 15824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606821651
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1606821651
transform 1 0 14812 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1606821651
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_153
timestamp 1606821651
transform 1 0 15180 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2116 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1564 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606821651
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1606821651
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1606821651
transform 1 0 4508 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606821651
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606821651
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_32
timestamp 1606821651
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_36
timestamp 1606821651
transform 1 0 4416 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5704 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_46
timestamp 1606821651
transform 1 0 5336 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7544 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_66
timestamp 1606821651
transform 1 0 7176 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1606821651
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606821651
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_86
timestamp 1606821651
transform 1 0 9016 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_102
timestamp 1606821651
transform 1 0 10488 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10856 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1606821651
transform 1 0 12052 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_115
timestamp 1606821651
transform 1 0 11684 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1606821651
transform 1 0 14444 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1606821651
transform 1 0 13248 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_128
timestamp 1606821651
transform 1 0 12880 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1606821651
transform 1 0 14076 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606821651
transform -1 0 15824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606821651
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1606821651
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_154
timestamp 1606821651
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1606821651
transform 1 0 1840 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606821651
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1606821651
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1606821651
transform 1 0 1748 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_17
timestamp 1606821651
transform 1 0 2668 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4876 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 3036 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_37
timestamp 1606821651
transform 1 0 4508 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 6808 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606821651
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1606821651
transform 1 0 6348 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 8648 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_78
timestamp 1606821651
transform 1 0 8280 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1606821651
transform 1 0 10488 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_98
timestamp 1606821651
transform 1 0 10120 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1606821651
transform 1 0 11684 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606821651
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_111
timestamp 1606821651
transform 1 0 11316 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1606821651
transform 1 0 11960 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13616 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_132
timestamp 1606821651
transform 1 0 13248 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_145
timestamp 1606821651
transform 1 0 14444 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1606821651
transform 1 0 14812 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606821651
transform -1 0 15824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_153
timestamp 1606821651
transform 1 0 15180 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1606821651
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 2116 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606821651
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_7
timestamp 1606821651
transform 1 0 1748 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1606821651
transform 1 0 4508 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606821651
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1606821651
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_32
timestamp 1606821651
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_36
timestamp 1606821651
transform 1 0 4416 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5428 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_46
timestamp 1606821651
transform 1 0 5336 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7268 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_63
timestamp 1606821651
transform 1 0 6900 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_83
timestamp 1606821651
transform 1 0 8740 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9660 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606821651
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 9108 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1606821651
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1606821651
transform 1 0 11500 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_109
timestamp 1606821651
transform 1 0 11132 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_122
timestamp 1606821651
transform 1 0 12328 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12696 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1606821651
transform 1 0 13892 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1606821651
transform 1 0 13524 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606821651
transform -1 0 15824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606821651
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_148
timestamp 1606821651
transform 1 0 14720 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1606821651
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_154
timestamp 1606821651
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1606821651
transform 1 0 2208 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1606821651
transform 1 0 1380 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606821651
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 4876 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 3036 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_37
timestamp 1606821651
transform 1 0 4508 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6808 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606821651
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1606821651
transform 1 0 6348 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 8648 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_78
timestamp 1606821651
transform 1 0 8280 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10488 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_98
timestamp 1606821651
transform 1 0 10120 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1606821651
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606821651
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_118
timestamp 1606821651
transform 1 0 11960 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1606821651
transform 1 0 13616 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_132
timestamp 1606821651
transform 1 0 13248 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_145
timestamp 1606821651
transform 1 0 14444 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1606821651
transform 1 0 14812 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606821651
transform -1 0 15824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_153
timestamp 1606821651
transform 1 0 15180 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1606821651
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 2116 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606821651
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_7
timestamp 1606821651
transform 1 0 1748 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 4232 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606821651
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1606821651
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1606821651
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5704 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7544 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_66
timestamp 1606821651
transform 1 0 7176 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 9660 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606821651
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_86
timestamp 1606821651
transform 1 0 9016 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 11500 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_109
timestamp 1606821651
transform 1 0 11132 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1606821651
transform 1 0 13340 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_129
timestamp 1606821651
transform 1 0 12972 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_142
timestamp 1606821651
transform 1 0 14168 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1606821651
transform 1 0 14536 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606821651
transform -1 0 15824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606821651
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1606821651
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_154
timestamp 1606821651
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1606821651
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 2116 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1606821651
transform 1 0 1840 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606821651
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606821651
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1606821651
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1606821651
transform 1 0 1748 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_17
timestamp 1606821651
transform 1 0 2668 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_7
timestamp 1606821651
transform 1 0 1748 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 3036 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 4048 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606821651
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 4876 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_37
timestamp 1606821651
transform 1 0 4508 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1606821651
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5888 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 5244 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606821651
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_44
timestamp 1606821651
transform 1 0 5152 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_62
timestamp 1606821651
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_48
timestamp 1606821651
transform 1 0 5520 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7728 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 7176 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_14_68
timestamp 1606821651
transform 1 0 7360 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10488 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 9016 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606821651
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_88
timestamp 1606821651
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11500 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1606821651
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606821651
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_118
timestamp 1606821651
transform 1 0 11960 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_109
timestamp 1606821651
transform 1 0 11132 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_122
timestamp 1606821651
transform 1 0 12328 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1606821651
transform 1 0 13892 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1606821651
transform 1 0 13616 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1606821651
transform 1 0 12696 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_132
timestamp 1606821651
transform 1 0 13248 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_145
timestamp 1606821651
transform 1 0 14444 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_135
timestamp 1606821651
transform 1 0 13524 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1606821651
transform 1 0 14812 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606821651
transform -1 0 15824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606821651
transform -1 0 15824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606821651
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_153
timestamp 1606821651
transform 1 0 15180 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_148
timestamp 1606821651
transform 1 0 14720 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1606821651
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_154
timestamp 1606821651
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1606821651
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1606821651
transform 1 0 1840 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606821651
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1606821651
transform 1 0 1748 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_17
timestamp 1606821651
transform 1 0 2668 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 4876 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 3036 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_37
timestamp 1606821651
transform 1 0 4508 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606821651
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1606821651
transform 1 0 6348 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8648 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_78
timestamp 1606821651
transform 1 0 8280 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10488 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_98
timestamp 1606821651
transform 1 0 10120 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1606821651
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606821651
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1606821651
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13616 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_132
timestamp 1606821651
transform 1 0 13248 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_145
timestamp 1606821651
transform 1 0 14444 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1606821651
transform 1 0 14812 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606821651
transform -1 0 15824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1606821651
transform 1 0 15180 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 2116 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1564 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606821651
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1606821651
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 4048 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606821651
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1606821651
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 6348 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 6072 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_48
timestamp 1606821651
transform 1 0 5520 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1606821651
transform 1 0 8188 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_73
timestamp 1606821651
transform 1 0 7820 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1606821651
transform 1 0 8464 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1606821651
transform 1 0 8832 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9660 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606821651
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_87
timestamp 1606821651
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1606821651
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1606821651
transform 1 0 11500 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_109
timestamp 1606821651
transform 1 0 11132 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_122
timestamp 1606821651
transform 1 0 12328 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12696 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1606821651
transform 1 0 13892 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_135
timestamp 1606821651
transform 1 0 13524 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606821651
transform -1 0 15824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606821651
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_148
timestamp 1606821651
transform 1 0 14720 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1606821651
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1606821651
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1606821651
transform 1 0 1840 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606821651
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1606821651
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1606821651
transform 1 0 1748 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_17
timestamp 1606821651
transform 1 0 2668 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 3036 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4876 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_37
timestamp 1606821651
transform 1 0 4508 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6808 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606821651
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1606821651
transform 1 0 6348 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 8648 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_78
timestamp 1606821651
transform 1 0 8280 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10488 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_98
timestamp 1606821651
transform 1 0 10120 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1606821651
transform 1 0 11684 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606821651
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_111
timestamp 1606821651
transform 1 0 11316 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1606821651
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1606821651
transform 1 0 13616 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_132
timestamp 1606821651
transform 1 0 13248 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_145
timestamp 1606821651
transform 1 0 14444 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1606821651
transform 1 0 14812 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606821651
transform -1 0 15824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_153
timestamp 1606821651
transform 1 0 15180 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1606821651
transform 1 0 1656 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606821651
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1606821651
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1606821651
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4692 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606821651
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1606821651
transform 1 0 4324 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1606821651
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_37
timestamp 1606821651
transform 1 0 4508 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1606821651
transform 1 0 5888 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_48
timestamp 1606821651
transform 1 0 5520 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_61
timestamp 1606821651
transform 1 0 6716 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1606821651
transform 1 0 8280 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1606821651
transform 1 0 7084 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_74
timestamp 1606821651
transform 1 0 7912 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_81
timestamp 1606821651
transform 1 0 8556 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1606821651
transform 1 0 8924 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1606821651
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606821651
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_88
timestamp 1606821651
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_102
timestamp 1606821651
transform 1 0 10488 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1606821651
transform 1 0 10856 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12052 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_115
timestamp 1606821651
transform 1 0 11684 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1606821651
transform 1 0 14444 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1606821651
transform 1 0 13248 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_128
timestamp 1606821651
transform 1 0 12880 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1606821651
transform 1 0 14076 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606821651
transform -1 0 15824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606821651
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_149
timestamp 1606821651
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_154
timestamp 1606821651
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1606821651
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1606821651
transform 1 0 1748 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1606821651
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606821651
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606821651
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1606821651
transform 1 0 1564 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1606821651
transform 1 0 1840 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_14
timestamp 1606821651
transform 1 0 2392 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_17
timestamp 1606821651
transform 1 0 2668 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1606821651
transform 1 0 2760 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 3036 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4876 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 4048 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606821651
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_37
timestamp 1606821651
transform 1 0 4508 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1606821651
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_38
timestamp 1606821651
transform 1 0 4600 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1606821651
transform 1 0 5152 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5796 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606821651
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1606821651
transform 1 0 6348 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_62
timestamp 1606821651
transform 1 0 6808 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_47
timestamp 1606821651
transform 1 0 5428 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6900 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1606821651
transform 1 0 8740 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1606821651
transform 1 0 7636 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_19_79
timestamp 1606821651
transform 1 0 8372 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_67
timestamp 1606821651
transform 1 0 7268 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1606821651
transform 1 0 8464 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1606821651
transform 1 0 8832 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1606821651
transform 1 0 9936 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9660 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1606821651
transform 1 0 10580 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606821651
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_92
timestamp 1606821651
transform 1 0 9568 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_99
timestamp 1606821651
transform 1 0 10212 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_87
timestamp 1606821651
transform 1 0 9108 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1606821651
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1606821651
transform 1 0 11500 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606821651
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 11776 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_112
timestamp 1606821651
transform 1 0 11408 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_119
timestamp 1606821651
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_109
timestamp 1606821651
transform 1 0 11132 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_122
timestamp 1606821651
transform 1 0 12328 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1606821651
transform 1 0 12696 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13616 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1606821651
transform 1 0 13892 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_19_132
timestamp 1606821651
transform 1 0 13248 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_145
timestamp 1606821651
transform 1 0 14444 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1606821651
transform 1 0 13524 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1606821651
transform 1 0 14812 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606821651
transform -1 0 15824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606821651
transform -1 0 15824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606821651
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp 1606821651
transform 1 0 15180 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_148
timestamp 1606821651
transform 1 0 14720 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1606821651
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1606821651
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1606821651
transform 1 0 2484 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1564 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606821651
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1606821651
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_11
timestamp 1606821651
transform 1 0 2116 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4876 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1606821651
transform 1 0 3680 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_24
timestamp 1606821651
transform 1 0 3312 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_37
timestamp 1606821651
transform 1 0 4508 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606821651
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1606821651
transform 1 0 6348 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_62
timestamp 1606821651
transform 1 0 6808 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1606821651
transform 1 0 8464 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1606821651
transform 1 0 7268 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_66
timestamp 1606821651
transform 1 0 7176 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_76
timestamp 1606821651
transform 1 0 8096 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_83
timestamp 1606821651
transform 1 0 8740 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9108 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_21_103
timestamp 1606821651
transform 1 0 10580 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1606821651
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1606821651
transform 1 0 11040 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606821651
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_107
timestamp 1606821651
transform 1 0 10948 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_117
timestamp 1606821651
transform 1 0 11868 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1606821651
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 13708 0 1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_21_132
timestamp 1606821651
transform 1 0 13248 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_136
timestamp 1606821651
transform 1 0 13616 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606821651
transform -1 0 15824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_150
timestamp 1606821651
transform 1 0 14904 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_156
timestamp 1606821651
transform 1 0 15456 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1606821651
transform 1 0 2760 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1606821651
transform 1 0 1564 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606821651
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1606821651
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_14
timestamp 1606821651
transform 1 0 2392 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1606821651
transform 1 0 4140 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606821651
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1606821651
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_32
timestamp 1606821651
transform 1 0 4048 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 6808 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 5336 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 6256 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_42
timestamp 1606821651
transform 1 0 4968 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_52
timestamp 1606821651
transform 1 0 5888 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_59
timestamp 1606821651
transform 1 0 6532 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1606821651
transform 1 0 8648 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_78
timestamp 1606821651
transform 1 0 8280 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 10212 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606821651
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_85
timestamp 1606821651
transform 1 0 8924 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_93
timestamp 1606821651
transform 1 0 9660 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_102
timestamp 1606821651
transform 1 0 10488 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1606821651
transform 1 0 12052 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1606821651
transform 1 0 10856 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_115
timestamp 1606821651
transform 1 0 11684 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1606821651
transform 1 0 14444 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1606821651
transform 1 0 13248 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1606821651
transform 1 0 13064 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_128
timestamp 1606821651
transform 1 0 12880 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1606821651
transform 1 0 14076 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606821651
transform -1 0 15824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606821651
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_149
timestamp 1606821651
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_154
timestamp 1606821651
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1606821651
transform 1 0 1932 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606821651
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1606821651
transform 1 0 1380 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_18
timestamp 1606821651
transform 1 0 2760 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4324 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1606821651
transform 1 0 3128 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_31
timestamp 1606821651
transform 1 0 3956 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 6808 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606821651
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 5520 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 6164 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_44
timestamp 1606821651
transform 1 0 5152 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1606821651
transform 1 0 5796 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_58
timestamp 1606821651
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8648 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_78
timestamp 1606821651
transform 1 0 8280 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 9844 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_91
timestamp 1606821651
transform 1 0 9476 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_98 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 10120 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1606821651
transform 1 0 11040 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1606821651
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606821651
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_106
timestamp 1606821651
transform 1 0 10856 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_117
timestamp 1606821651
transform 1 0 11868 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1606821651
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1606821651
transform 1 0 14352 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1606821651
transform 1 0 13616 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_132
timestamp 1606821651
transform 1 0 13248 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_140
timestamp 1606821651
transform 1 0 13984 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606821651
transform -1 0 15824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_148
timestamp 1606821651
transform 1 0 14720 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_156
timestamp 1606821651
transform 1 0 15456 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1840 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1606821651
transform 1 0 2760 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606821651
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1606821651
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1606821651
transform 1 0 1748 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_14
timestamp 1606821651
transform 1 0 2392 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4140 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606821651
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1606821651
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_32
timestamp 1606821651
transform 1 0 4048 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1606821651
transform 1 0 5336 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1606821651
transform 1 0 6532 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_42
timestamp 1606821651
transform 1 0 4968 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_55
timestamp 1606821651
transform 1 0 6164 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1606821651
transform 1 0 7728 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_68
timestamp 1606821651
transform 1 0 7360 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_81
timestamp 1606821651
transform 1 0 8556 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1606821651
transform 1 0 8924 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1606821651
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606821651
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_88
timestamp 1606821651
transform 1 0 9200 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_102
timestamp 1606821651
transform 1 0 10488 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10856 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12052 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_115
timestamp 1606821651
transform 1 0 11684 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1606821651
transform 1 0 13984 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1606821651
transform 1 0 13248 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_128
timestamp 1606821651
transform 1 0 12880 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1606821651
transform 1 0 13616 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_144
timestamp 1606821651
transform 1 0 14352 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606821651
transform -1 0 15824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606821651
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1606821651
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_154
timestamp 1606821651
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1606821651
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2208 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606821651
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_7
timestamp 1606821651
transform 1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_11
timestamp 1606821651
transform 1 0 2116 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_18
timestamp 1606821651
transform 1 0 2760 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1606821651
transform 1 0 4324 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1606821651
transform 1 0 3128 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_31
timestamp 1606821651
transform 1 0 3956 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1606821651
transform 1 0 5520 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606821651
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_44
timestamp 1606821651
transform 1 0 5152 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1606821651
transform 1 0 6348 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_62
timestamp 1606821651
transform 1 0 6808 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1606821651
transform 1 0 8096 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6900 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_72
timestamp 1606821651
transform 1 0 7728 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_80
timestamp 1606821651
transform 1 0 8464 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1606821651
transform 1 0 9200 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1606821651
transform 1 0 10396 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 8832 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_87
timestamp 1606821651
transform 1 0 9108 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_97
timestamp 1606821651
transform 1 0 10028 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1606821651
transform 1 0 11592 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606821651
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_110
timestamp 1606821651
transform 1 0 11224 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_118
timestamp 1606821651
transform 1 0 11960 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1606821651
transform 1 0 13616 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1606821651
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_134
timestamp 1606821651
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_140
timestamp 1606821651
transform 1 0 13984 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01
timestamp 1606821651
transform 1 0 14628 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606821651
transform -1 0 15824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_146
timestamp 1606821651
transform 1 0 14536 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_153
timestamp 1606821651
transform 1 0 15180 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1606821651
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1606821651
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606821651
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606821651
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1564 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1606821651
transform 1 0 1748 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_11
timestamp 1606821651
transform 1 0 2116 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1840 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_14
timestamp 1606821651
transform 1 0 2392 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2760 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2484 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_30
timestamp 1606821651
transform 1 0 3864 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_24
timestamp 1606821651
transform 1 0 3312 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_26_28
timestamp 1606821651
transform 1 0 3680 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_21
timestamp 1606821651
transform 1 0 3036 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 3404 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606821651
transform 1 0 3956 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606821651
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_32
timestamp 1606821651
transform 1 0 4048 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_32
timestamp 1606821651
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1606821651
transform 1 0 4416 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 4324 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1606821651
transform 1 0 6164 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1606821651
transform 1 0 5612 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606821651
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_51
timestamp 1606821651
transform 1 0 5796 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_59
timestamp 1606821651
transform 1 0 6532 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_45
timestamp 1606821651
transform 1 0 5244 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_58
timestamp 1606821651
transform 1 0 6440 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1606821651
transform 1 0 8096 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6900 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1606821651
transform 1 0 7176 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1606821651
transform 1 0 8372 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_72
timestamp 1606821651
transform 1 0 7728 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_63
timestamp 1606821651
transform 1 0 6900 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_75
timestamp 1606821651
transform 1 0 8004 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_92
timestamp 1606821651
transform 1 0 9568 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_88
timestamp 1606821651
transform 1 0 9200 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1606821651
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_85
timestamp 1606821651
transform 1 0 8924 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606821651
transform 1 0 9660 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606821651
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1606821651
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_103
timestamp 1606821651
transform 1 0 10580 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_102
timestamp 1606821651
transform 1 0 10488 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1606821651
transform 1 0 9752 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1606821651
transform 1 0 10948 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1606821651
transform 1 0 10856 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_111
timestamp 1606821651
transform 1 0 11316 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_110
timestamp 1606821651
transform 1 0 11224 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_118
timestamp 1606821651
transform 1 0 11960 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1606821651
transform 1 0 11592 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1606821651
transform 1 0 11684 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp 1606821651
transform 1 0 12420 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_119
timestamp 1606821651
transform 1 0 12052 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1606821651
transform 1 0 12328 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606821651
transform 1 0 12512 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1606821651
transform 1 0 12604 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1606821651
transform 1 0 13800 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1606821651
transform 1 0 13064 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606821651
transform 1 0 13432 0 1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_26_126
timestamp 1606821651
transform 1 0 12696 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_134
timestamp 1606821651
transform 1 0 13432 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_142
timestamp 1606821651
transform 1 0 14168 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_129
timestamp 1606821651
transform 1 0 12972 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_133
timestamp 1606821651
transform 1 0 13340 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1606821651
transform 1 0 14536 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606821651
transform -1 0 15824 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606821651
transform -1 0 15824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606821651
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606821651
transform 1 0 15364 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_149
timestamp 1606821651
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_154
timestamp 1606821651
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_147
timestamp 1606821651
transform 1 0 14628 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_156
timestamp 1606821651
transform 1 0 15456 0 1 16864
box -38 -48 130 592
<< labels >>
rlabel metal2 s 202 19520 258 20000 6 IO_ISOL_N
port 0 nsew default input
rlabel metal3 s 0 1368 480 1488 6 ccff_head
port 1 nsew default input
rlabel metal3 s 16520 1912 17000 2032 6 ccff_tail
port 2 nsew default tristate
rlabel metal2 s 8482 0 8538 480 6 chany_bottom_in[0]
port 3 nsew default input
rlabel metal2 s 12622 0 12678 480 6 chany_bottom_in[10]
port 4 nsew default input
rlabel metal2 s 12990 0 13046 480 6 chany_bottom_in[11]
port 5 nsew default input
rlabel metal2 s 13450 0 13506 480 6 chany_bottom_in[12]
port 6 nsew default input
rlabel metal2 s 13818 0 13874 480 6 chany_bottom_in[13]
port 7 nsew default input
rlabel metal2 s 14278 0 14334 480 6 chany_bottom_in[14]
port 8 nsew default input
rlabel metal2 s 14646 0 14702 480 6 chany_bottom_in[15]
port 9 nsew default input
rlabel metal2 s 15106 0 15162 480 6 chany_bottom_in[16]
port 10 nsew default input
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_in[17]
port 11 nsew default input
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_in[18]
port 12 nsew default input
rlabel metal2 s 16302 0 16358 480 6 chany_bottom_in[19]
port 13 nsew default input
rlabel metal2 s 8850 0 8906 480 6 chany_bottom_in[1]
port 14 nsew default input
rlabel metal2 s 9310 0 9366 480 6 chany_bottom_in[2]
port 15 nsew default input
rlabel metal2 s 9678 0 9734 480 6 chany_bottom_in[3]
port 16 nsew default input
rlabel metal2 s 10138 0 10194 480 6 chany_bottom_in[4]
port 17 nsew default input
rlabel metal2 s 10506 0 10562 480 6 chany_bottom_in[5]
port 18 nsew default input
rlabel metal2 s 10966 0 11022 480 6 chany_bottom_in[6]
port 19 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[7]
port 20 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_in[8]
port 21 nsew default input
rlabel metal2 s 12162 0 12218 480 6 chany_bottom_in[9]
port 22 nsew default input
rlabel metal2 s 202 0 258 480 6 chany_bottom_out[0]
port 23 nsew default tristate
rlabel metal2 s 4342 0 4398 480 6 chany_bottom_out[10]
port 24 nsew default tristate
rlabel metal2 s 4710 0 4766 480 6 chany_bottom_out[11]
port 25 nsew default tristate
rlabel metal2 s 5170 0 5226 480 6 chany_bottom_out[12]
port 26 nsew default tristate
rlabel metal2 s 5538 0 5594 480 6 chany_bottom_out[13]
port 27 nsew default tristate
rlabel metal2 s 5998 0 6054 480 6 chany_bottom_out[14]
port 28 nsew default tristate
rlabel metal2 s 6366 0 6422 480 6 chany_bottom_out[15]
port 29 nsew default tristate
rlabel metal2 s 6826 0 6882 480 6 chany_bottom_out[16]
port 30 nsew default tristate
rlabel metal2 s 7194 0 7250 480 6 chany_bottom_out[17]
port 31 nsew default tristate
rlabel metal2 s 7654 0 7710 480 6 chany_bottom_out[18]
port 32 nsew default tristate
rlabel metal2 s 8022 0 8078 480 6 chany_bottom_out[19]
port 33 nsew default tristate
rlabel metal2 s 570 0 626 480 6 chany_bottom_out[1]
port 34 nsew default tristate
rlabel metal2 s 1030 0 1086 480 6 chany_bottom_out[2]
port 35 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_out[3]
port 36 nsew default tristate
rlabel metal2 s 1858 0 1914 480 6 chany_bottom_out[4]
port 37 nsew default tristate
rlabel metal2 s 2226 0 2282 480 6 chany_bottom_out[5]
port 38 nsew default tristate
rlabel metal2 s 2686 0 2742 480 6 chany_bottom_out[6]
port 39 nsew default tristate
rlabel metal2 s 3054 0 3110 480 6 chany_bottom_out[7]
port 40 nsew default tristate
rlabel metal2 s 3514 0 3570 480 6 chany_bottom_out[8]
port 41 nsew default tristate
rlabel metal2 s 3882 0 3938 480 6 chany_bottom_out[9]
port 42 nsew default tristate
rlabel metal2 s 8666 19520 8722 20000 6 chany_top_in[0]
port 43 nsew default input
rlabel metal2 s 12714 19520 12770 20000 6 chany_top_in[10]
port 44 nsew default input
rlabel metal2 s 13082 19520 13138 20000 6 chany_top_in[11]
port 45 nsew default input
rlabel metal2 s 13542 19520 13598 20000 6 chany_top_in[12]
port 46 nsew default input
rlabel metal2 s 13910 19520 13966 20000 6 chany_top_in[13]
port 47 nsew default input
rlabel metal2 s 14370 19520 14426 20000 6 chany_top_in[14]
port 48 nsew default input
rlabel metal2 s 14738 19520 14794 20000 6 chany_top_in[15]
port 49 nsew default input
rlabel metal2 s 15106 19520 15162 20000 6 chany_top_in[16]
port 50 nsew default input
rlabel metal2 s 15566 19520 15622 20000 6 chany_top_in[17]
port 51 nsew default input
rlabel metal2 s 15934 19520 15990 20000 6 chany_top_in[18]
port 52 nsew default input
rlabel metal2 s 16394 19520 16450 20000 6 chany_top_in[19]
port 53 nsew default input
rlabel metal2 s 9034 19520 9090 20000 6 chany_top_in[1]
port 54 nsew default input
rlabel metal2 s 9494 19520 9550 20000 6 chany_top_in[2]
port 55 nsew default input
rlabel metal2 s 9862 19520 9918 20000 6 chany_top_in[3]
port 56 nsew default input
rlabel metal2 s 10322 19520 10378 20000 6 chany_top_in[4]
port 57 nsew default input
rlabel metal2 s 10690 19520 10746 20000 6 chany_top_in[5]
port 58 nsew default input
rlabel metal2 s 11058 19520 11114 20000 6 chany_top_in[6]
port 59 nsew default input
rlabel metal2 s 11518 19520 11574 20000 6 chany_top_in[7]
port 60 nsew default input
rlabel metal2 s 11886 19520 11942 20000 6 chany_top_in[8]
port 61 nsew default input
rlabel metal2 s 12346 19520 12402 20000 6 chany_top_in[9]
port 62 nsew default input
rlabel metal2 s 570 19520 626 20000 6 chany_top_out[0]
port 63 nsew default tristate
rlabel metal2 s 4618 19520 4674 20000 6 chany_top_out[10]
port 64 nsew default tristate
rlabel metal2 s 4986 19520 5042 20000 6 chany_top_out[11]
port 65 nsew default tristate
rlabel metal2 s 5446 19520 5502 20000 6 chany_top_out[12]
port 66 nsew default tristate
rlabel metal2 s 5814 19520 5870 20000 6 chany_top_out[13]
port 67 nsew default tristate
rlabel metal2 s 6274 19520 6330 20000 6 chany_top_out[14]
port 68 nsew default tristate
rlabel metal2 s 6642 19520 6698 20000 6 chany_top_out[15]
port 69 nsew default tristate
rlabel metal2 s 7010 19520 7066 20000 6 chany_top_out[16]
port 70 nsew default tristate
rlabel metal2 s 7470 19520 7526 20000 6 chany_top_out[17]
port 71 nsew default tristate
rlabel metal2 s 7838 19520 7894 20000 6 chany_top_out[18]
port 72 nsew default tristate
rlabel metal2 s 8298 19520 8354 20000 6 chany_top_out[19]
port 73 nsew default tristate
rlabel metal2 s 938 19520 994 20000 6 chany_top_out[1]
port 74 nsew default tristate
rlabel metal2 s 1398 19520 1454 20000 6 chany_top_out[2]
port 75 nsew default tristate
rlabel metal2 s 1766 19520 1822 20000 6 chany_top_out[3]
port 76 nsew default tristate
rlabel metal2 s 2226 19520 2282 20000 6 chany_top_out[4]
port 77 nsew default tristate
rlabel metal2 s 2594 19520 2650 20000 6 chany_top_out[5]
port 78 nsew default tristate
rlabel metal2 s 2962 19520 3018 20000 6 chany_top_out[6]
port 79 nsew default tristate
rlabel metal2 s 3422 19520 3478 20000 6 chany_top_out[7]
port 80 nsew default tristate
rlabel metal2 s 3790 19520 3846 20000 6 chany_top_out[8]
port 81 nsew default tristate
rlabel metal2 s 4250 19520 4306 20000 6 chany_top_out[9]
port 82 nsew default tristate
rlabel metal3 s 16520 9800 17000 9920 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 83 nsew default tristate
rlabel metal3 s 16520 13880 17000 14000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 84 nsew default input
rlabel metal3 s 16520 17824 17000 17944 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 85 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 left_grid_pin_16_
port 86 nsew default tristate
rlabel metal3 s 0 4224 480 4344 6 left_grid_pin_17_
port 87 nsew default tristate
rlabel metal3 s 0 5176 480 5296 6 left_grid_pin_18_
port 88 nsew default tristate
rlabel metal3 s 0 6128 480 6248 6 left_grid_pin_19_
port 89 nsew default tristate
rlabel metal3 s 0 7080 480 7200 6 left_grid_pin_20_
port 90 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 left_grid_pin_21_
port 91 nsew default tristate
rlabel metal3 s 0 8984 480 9104 6 left_grid_pin_22_
port 92 nsew default tristate
rlabel metal3 s 0 9936 480 10056 6 left_grid_pin_23_
port 93 nsew default tristate
rlabel metal3 s 0 10888 480 11008 6 left_grid_pin_24_
port 94 nsew default tristate
rlabel metal3 s 0 11840 480 11960 6 left_grid_pin_25_
port 95 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 left_grid_pin_26_
port 96 nsew default tristate
rlabel metal3 s 0 13744 480 13864 6 left_grid_pin_27_
port 97 nsew default tristate
rlabel metal3 s 0 14696 480 14816 6 left_grid_pin_28_
port 98 nsew default tristate
rlabel metal3 s 0 15648 480 15768 6 left_grid_pin_29_
port 99 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 left_grid_pin_30_
port 100 nsew default tristate
rlabel metal3 s 0 17552 480 17672 6 left_grid_pin_31_
port 101 nsew default tristate
rlabel metal3 s 0 18504 480 18624 6 left_width_0_height_0__pin_0_
port 102 nsew default input
rlabel metal3 s 0 416 480 536 6 left_width_0_height_0__pin_1_lower
port 103 nsew default tristate
rlabel metal3 s 0 19456 480 19576 6 left_width_0_height_0__pin_1_upper
port 104 nsew default tristate
rlabel metal2 s 16762 19520 16818 20000 6 prog_clk_0_N_out
port 105 nsew default tristate
rlabel metal2 s 16762 0 16818 480 6 prog_clk_0_S_out
port 106 nsew default tristate
rlabel metal3 s 0 2320 480 2440 6 prog_clk_0_W_in
port 107 nsew default input
rlabel metal3 s 16520 5856 17000 5976 6 right_grid_pin_0_
port 108 nsew default tristate
rlabel metal4 s 3409 2128 3729 17456 6 VPWR
port 109 nsew default input
rlabel metal4 s 5875 2128 6195 17456 6 VGND
port 110 nsew default input
<< properties >>
string FIXED_BBOX 0 0 17000 20000
<< end >>
