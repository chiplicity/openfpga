magic
tech sky130A
magscale 1 2
timestamp 1605122599
<< locali >>
rect 12081 26163 12115 26537
rect 12541 26163 12575 26469
rect 12265 26095 12299 26129
rect 11839 26061 12299 26095
rect 13369 26095 13403 26333
rect 13921 25755 13955 26265
rect 16589 26163 16623 26333
rect 17325 25823 17359 26469
rect 17417 25755 17451 26537
rect 16405 25143 16439 25449
rect 17049 25143 17083 25449
rect 17509 25279 17543 25449
rect 25053 24599 25087 24769
rect 25605 23511 25639 23613
rect 14289 21879 14323 21981
rect 22569 21947 22603 22049
rect 17693 21471 17727 21573
rect 22477 20247 22511 20485
rect 857 12359 891 15521
rect 949 9707 983 19125
rect 9873 18071 9907 18241
rect 15853 18071 15887 18377
rect 19257 18241 19349 18275
rect 19257 18071 19291 18241
rect 2513 17051 2547 17221
rect 2697 16507 2731 16677
rect 24409 16439 24443 16677
rect 24777 16575 24811 16745
rect 16129 15351 16163 15589
rect 9689 14807 9723 15113
rect 15577 14875 15611 15045
rect 17601 14807 17635 15045
rect 22109 14807 22143 15113
rect 2237 14331 2271 14501
rect 13645 13719 13679 14025
rect 21833 13719 21867 13957
rect 8401 12699 8435 12869
rect 12633 12155 12667 12325
rect 19441 12087 19475 12257
rect 24501 11747 24535 11849
rect 5549 9911 5583 10013
rect 17141 9911 17175 10081
rect 22845 9911 22879 10217
rect 21281 9367 21315 9537
rect 14841 6647 14875 6817
rect 14933 6647 14967 6885
rect 2513 5015 2547 5321
<< viali >>
rect 12081 26537 12115 26571
rect 17417 26537 17451 26571
rect 12541 26469 12575 26503
rect 17325 26469 17359 26503
rect 12081 26129 12115 26163
rect 12265 26129 12299 26163
rect 12541 26129 12575 26163
rect 13369 26333 13403 26367
rect 11805 26061 11839 26095
rect 16589 26333 16623 26367
rect 13369 26061 13403 26095
rect 13921 26265 13955 26299
rect 16589 26129 16623 26163
rect 17325 25789 17359 25823
rect 13921 25721 13955 25755
rect 17417 25721 17451 25755
rect 10517 25449 10551 25483
rect 11621 25449 11655 25483
rect 13921 25449 13955 25483
rect 15209 25449 15243 25483
rect 15485 25449 15519 25483
rect 15945 25449 15979 25483
rect 16405 25449 16439 25483
rect 16865 25449 16899 25483
rect 17049 25449 17083 25483
rect 17325 25449 17359 25483
rect 17509 25449 17543 25483
rect 21925 25449 21959 25483
rect 10333 25313 10367 25347
rect 11437 25313 11471 25347
rect 12817 25313 12851 25347
rect 13553 25313 13587 25347
rect 14105 25313 14139 25347
rect 15853 25313 15887 25347
rect 13001 25245 13035 25279
rect 14381 25245 14415 25279
rect 16037 25245 16071 25279
rect 10241 25177 10275 25211
rect 11253 25177 11287 25211
rect 11989 25177 12023 25211
rect 17141 25313 17175 25347
rect 18889 25313 18923 25347
rect 19993 25313 20027 25347
rect 21741 25313 21775 25347
rect 22845 25313 22879 25347
rect 24501 25313 24535 25347
rect 24593 25313 24627 25347
rect 17509 25245 17543 25279
rect 24685 25245 24719 25279
rect 19073 25177 19107 25211
rect 20177 25177 20211 25211
rect 23029 25177 23063 25211
rect 9413 25109 9447 25143
rect 10885 25109 10919 25143
rect 12449 25109 12483 25143
rect 14841 25109 14875 25143
rect 16405 25109 16439 25143
rect 16589 25109 16623 25143
rect 17049 25109 17083 25143
rect 17693 25109 17727 25143
rect 23857 25109 23891 25143
rect 24133 25109 24167 25143
rect 1593 24905 1627 24939
rect 9229 24905 9263 24939
rect 14657 24905 14691 24939
rect 20361 24905 20395 24939
rect 25605 24905 25639 24939
rect 9689 24837 9723 24871
rect 10333 24837 10367 24871
rect 22661 24837 22695 24871
rect 12265 24769 12299 24803
rect 13645 24769 13679 24803
rect 15393 24769 15427 24803
rect 16865 24769 16899 24803
rect 18521 24769 18555 24803
rect 24501 24769 24535 24803
rect 25053 24769 25087 24803
rect 1409 24701 1443 24735
rect 9045 24701 9079 24735
rect 10149 24701 10183 24735
rect 11253 24701 11287 24735
rect 18337 24701 18371 24735
rect 20177 24701 20211 24735
rect 20729 24701 20763 24735
rect 21281 24701 21315 24735
rect 22477 24701 22511 24735
rect 24225 24701 24259 24735
rect 12909 24633 12943 24667
rect 13461 24633 13495 24667
rect 14289 24633 14323 24667
rect 15209 24633 15243 24667
rect 15853 24633 15887 24667
rect 16681 24633 16715 24667
rect 24317 24633 24351 24667
rect 25421 24701 25455 24735
rect 25973 24701 26007 24735
rect 2053 24565 2087 24599
rect 8677 24565 8711 24599
rect 10057 24565 10091 24599
rect 10793 24565 10827 24599
rect 11161 24565 11195 24599
rect 11437 24565 11471 24599
rect 11897 24565 11931 24599
rect 13001 24565 13035 24599
rect 13369 24565 13403 24599
rect 14749 24565 14783 24599
rect 15117 24565 15151 24599
rect 16129 24565 16163 24599
rect 16313 24565 16347 24599
rect 16773 24565 16807 24599
rect 17325 24565 17359 24599
rect 17785 24565 17819 24599
rect 19073 24565 19107 24599
rect 19993 24565 20027 24599
rect 21097 24565 21131 24599
rect 21465 24565 21499 24599
rect 21925 24565 21959 24599
rect 23029 24565 23063 24599
rect 23489 24565 23523 24599
rect 23857 24565 23891 24599
rect 24869 24565 24903 24599
rect 25053 24565 25087 24599
rect 25329 24565 25363 24599
rect 1593 24361 1627 24395
rect 7573 24361 7607 24395
rect 8677 24361 8711 24395
rect 11345 24361 11379 24395
rect 13461 24361 13495 24395
rect 13829 24361 13863 24395
rect 14841 24361 14875 24395
rect 15761 24361 15795 24395
rect 16865 24361 16899 24395
rect 18061 24361 18095 24395
rect 21373 24361 21407 24395
rect 17325 24293 17359 24327
rect 21465 24293 21499 24327
rect 1409 24225 1443 24259
rect 7389 24225 7423 24259
rect 8493 24225 8527 24259
rect 10241 24225 10275 24259
rect 11713 24225 11747 24259
rect 11805 24225 11839 24259
rect 15669 24225 15703 24259
rect 17233 24225 17267 24259
rect 18889 24225 18923 24259
rect 22201 24225 22235 24259
rect 23489 24225 23523 24259
rect 25053 24225 25087 24259
rect 11897 24157 11931 24191
rect 13921 24157 13955 24191
rect 14105 24157 14139 24191
rect 15853 24157 15887 24191
rect 17417 24157 17451 24191
rect 18429 24157 18463 24191
rect 19073 24157 19107 24191
rect 21557 24157 21591 24191
rect 22569 24157 22603 24191
rect 23581 24157 23615 24191
rect 23673 24157 23707 24191
rect 25145 24157 25179 24191
rect 25237 24157 25271 24191
rect 10425 24089 10459 24123
rect 11253 24089 11287 24123
rect 24501 24089 24535 24123
rect 8401 24021 8435 24055
rect 9045 24021 9079 24055
rect 9413 24021 9447 24055
rect 9873 24021 9907 24055
rect 10793 24021 10827 24055
rect 12725 24021 12759 24055
rect 13093 24021 13127 24055
rect 15301 24021 15335 24055
rect 16313 24021 16347 24055
rect 16773 24021 16807 24055
rect 19625 24021 19659 24055
rect 21005 24021 21039 24055
rect 22845 24021 22879 24055
rect 23121 24021 23155 24055
rect 24133 24021 24167 24055
rect 24685 24021 24719 24055
rect 1593 23817 1627 23851
rect 2697 23817 2731 23851
rect 8033 23817 8067 23851
rect 9137 23817 9171 23851
rect 9505 23817 9539 23851
rect 10241 23817 10275 23851
rect 10793 23817 10827 23851
rect 13277 23817 13311 23851
rect 15209 23817 15243 23851
rect 16221 23817 16255 23851
rect 18061 23817 18095 23851
rect 20361 23817 20395 23851
rect 20729 23817 20763 23851
rect 21925 23817 21959 23851
rect 22661 23817 22695 23851
rect 25421 23817 25455 23851
rect 8493 23749 8527 23783
rect 17049 23749 17083 23783
rect 17417 23749 17451 23783
rect 19073 23749 19107 23783
rect 24685 23749 24719 23783
rect 11437 23681 11471 23715
rect 12817 23681 12851 23715
rect 13829 23681 13863 23715
rect 15853 23681 15887 23715
rect 18613 23681 18647 23715
rect 19901 23681 19935 23715
rect 21373 23681 21407 23715
rect 21557 23681 21591 23715
rect 23489 23681 23523 23715
rect 24317 23681 24351 23715
rect 25145 23681 25179 23715
rect 1409 23613 1443 23647
rect 2513 23613 2547 23647
rect 3065 23613 3099 23647
rect 7849 23613 7883 23647
rect 8953 23613 8987 23647
rect 11161 23613 11195 23647
rect 13645 23613 13679 23647
rect 14381 23613 14415 23647
rect 15669 23613 15703 23647
rect 16865 23613 16899 23647
rect 17785 23613 17819 23647
rect 18429 23613 18463 23647
rect 18521 23613 18555 23647
rect 19625 23613 19659 23647
rect 21281 23613 21315 23647
rect 22477 23613 22511 23647
rect 25237 23613 25271 23647
rect 25605 23613 25639 23647
rect 8769 23545 8803 23579
rect 10701 23545 10735 23579
rect 11253 23545 11287 23579
rect 13185 23545 13219 23579
rect 14749 23545 14783 23579
rect 15577 23545 15611 23579
rect 24133 23545 24167 23579
rect 26249 23545 26283 23579
rect 2053 23477 2087 23511
rect 7481 23477 7515 23511
rect 9873 23477 9907 23511
rect 11805 23477 11839 23511
rect 12265 23477 12299 23511
rect 13737 23477 13771 23511
rect 15025 23477 15059 23511
rect 16773 23477 16807 23511
rect 19533 23477 19567 23511
rect 20913 23477 20947 23511
rect 22385 23477 22419 23511
rect 23029 23477 23063 23511
rect 23673 23477 23707 23511
rect 24041 23477 24075 23511
rect 25605 23477 25639 23511
rect 25881 23477 25915 23511
rect 7205 23273 7239 23307
rect 11621 23273 11655 23307
rect 15117 23273 15151 23307
rect 16681 23273 16715 23307
rect 17325 23273 17359 23307
rect 18153 23273 18187 23307
rect 18429 23273 18463 23307
rect 21189 23273 21223 23307
rect 23489 23273 23523 23307
rect 25237 23273 25271 23307
rect 7849 23205 7883 23239
rect 14749 23205 14783 23239
rect 15669 23205 15703 23239
rect 25605 23205 25639 23239
rect 2145 23137 2179 23171
rect 7573 23137 7607 23171
rect 9505 23137 9539 23171
rect 10425 23137 10459 23171
rect 10517 23137 10551 23171
rect 11989 23137 12023 23171
rect 13553 23137 13587 23171
rect 14197 23137 14231 23171
rect 15761 23137 15795 23171
rect 17233 23137 17267 23171
rect 18797 23137 18831 23171
rect 19625 23137 19659 23171
rect 22293 23137 22327 23171
rect 23857 23137 23891 23171
rect 25053 23137 25087 23171
rect 1685 23069 1719 23103
rect 2329 23069 2363 23103
rect 10609 23069 10643 23103
rect 12081 23069 12115 23103
rect 12173 23069 12207 23103
rect 12725 23069 12759 23103
rect 13645 23069 13679 23103
rect 13737 23069 13771 23103
rect 15945 23069 15979 23103
rect 16405 23069 16439 23103
rect 17417 23069 17451 23103
rect 18889 23069 18923 23103
rect 18981 23069 19015 23103
rect 22385 23069 22419 23103
rect 22477 23069 22511 23103
rect 23949 23069 23983 23103
rect 24133 23069 24167 23103
rect 9137 23001 9171 23035
rect 10057 23001 10091 23035
rect 11437 23001 11471 23035
rect 24685 23001 24719 23035
rect 6929 22933 6963 22967
rect 8677 22933 8711 22967
rect 9965 22933 9999 22967
rect 13001 22933 13035 22967
rect 13185 22933 13219 22967
rect 15301 22933 15335 22967
rect 16865 22933 16899 22967
rect 20361 22933 20395 22967
rect 20729 22933 20763 22967
rect 21465 22933 21499 22967
rect 21925 22933 21959 22967
rect 23213 22933 23247 22967
rect 1593 22729 1627 22763
rect 4629 22729 4663 22763
rect 9045 22729 9079 22763
rect 10149 22729 10183 22763
rect 11713 22729 11747 22763
rect 13277 22729 13311 22763
rect 15485 22729 15519 22763
rect 17417 22729 17451 22763
rect 19625 22729 19659 22763
rect 21833 22729 21867 22763
rect 25053 22729 25087 22763
rect 25605 22729 25639 22763
rect 8953 22661 8987 22695
rect 20729 22661 20763 22695
rect 23857 22661 23891 22695
rect 7757 22593 7791 22627
rect 9505 22593 9539 22627
rect 9597 22593 9631 22627
rect 11161 22593 11195 22627
rect 13737 22593 13771 22627
rect 13921 22593 13955 22627
rect 14473 22593 14507 22627
rect 16589 22593 16623 22627
rect 18521 22593 18555 22627
rect 18613 22593 18647 22627
rect 20177 22593 20211 22627
rect 22477 22593 22511 22627
rect 24501 22593 24535 22627
rect 1409 22525 1443 22559
rect 4445 22525 4479 22559
rect 4997 22525 5031 22559
rect 7113 22525 7147 22559
rect 7665 22525 7699 22559
rect 9413 22525 9447 22559
rect 11069 22525 11103 22559
rect 13185 22525 13219 22559
rect 13645 22525 13679 22559
rect 14933 22525 14967 22559
rect 16497 22525 16531 22559
rect 19073 22525 19107 22559
rect 25421 22525 25455 22559
rect 25973 22525 26007 22559
rect 5549 22457 5583 22491
rect 5917 22457 5951 22491
rect 6285 22457 6319 22491
rect 7573 22457 7607 22491
rect 12817 22457 12851 22491
rect 18429 22457 18463 22491
rect 19993 22457 20027 22491
rect 22201 22457 22235 22491
rect 23121 22457 23155 22491
rect 24225 22457 24259 22491
rect 2053 22389 2087 22423
rect 2421 22389 2455 22423
rect 6653 22389 6687 22423
rect 7205 22389 7239 22423
rect 8217 22389 8251 22423
rect 10425 22389 10459 22423
rect 10609 22389 10643 22423
rect 10977 22389 11011 22423
rect 11989 22389 12023 22423
rect 14749 22389 14783 22423
rect 15117 22389 15151 22423
rect 15853 22389 15887 22423
rect 16037 22389 16071 22423
rect 16405 22389 16439 22423
rect 17141 22389 17175 22423
rect 17785 22389 17819 22423
rect 18061 22389 18095 22423
rect 19441 22389 19475 22423
rect 20085 22389 20119 22423
rect 21281 22389 21315 22423
rect 21649 22389 21683 22423
rect 22293 22389 22327 22423
rect 23489 22389 23523 22423
rect 24317 22389 24351 22423
rect 4445 22185 4479 22219
rect 4813 22185 4847 22219
rect 13461 22185 13495 22219
rect 14473 22185 14507 22219
rect 15117 22185 15151 22219
rect 21649 22185 21683 22219
rect 23857 22185 23891 22219
rect 5365 22117 5399 22151
rect 12265 22117 12299 22151
rect 13829 22117 13863 22151
rect 17785 22117 17819 22151
rect 18613 22117 18647 22151
rect 23673 22117 23707 22151
rect 1409 22049 1443 22083
rect 5089 22049 5123 22083
rect 7380 22049 7414 22083
rect 9505 22049 9539 22083
rect 9956 22049 9990 22083
rect 11713 22049 11747 22083
rect 13001 22049 13035 22083
rect 16304 22049 16338 22083
rect 20729 22049 20763 22083
rect 22017 22049 22051 22083
rect 22569 22049 22603 22083
rect 23397 22049 23431 22083
rect 24225 22049 24259 22083
rect 25605 22049 25639 22083
rect 7113 21981 7147 22015
rect 9689 21981 9723 22015
rect 12357 21981 12391 22015
rect 12541 21981 12575 22015
rect 13921 21981 13955 22015
rect 14105 21981 14139 22015
rect 14289 21981 14323 22015
rect 15577 21981 15611 22015
rect 16037 21981 16071 22015
rect 18705 21981 18739 22015
rect 18797 21981 18831 22015
rect 19717 21981 19751 22015
rect 21189 21981 21223 22015
rect 22109 21981 22143 22015
rect 22293 21981 22327 22015
rect 1593 21913 1627 21947
rect 8493 21913 8527 21947
rect 11897 21913 11931 21947
rect 24317 21981 24351 22015
rect 24409 21981 24443 22015
rect 25237 21981 25271 22015
rect 18245 21913 18279 21947
rect 21557 21913 21591 21947
rect 22569 21913 22603 21947
rect 5917 21845 5951 21879
rect 6561 21845 6595 21879
rect 6929 21845 6963 21879
rect 9045 21845 9079 21879
rect 11069 21845 11103 21879
rect 13277 21845 13311 21879
rect 14289 21845 14323 21879
rect 15945 21845 15979 21879
rect 17417 21845 17451 21879
rect 18153 21845 18187 21879
rect 19257 21845 19291 21879
rect 20361 21845 20395 21879
rect 22661 21845 22695 21879
rect 24869 21845 24903 21879
rect 1593 21641 1627 21675
rect 3985 21641 4019 21675
rect 4997 21641 5031 21675
rect 6653 21641 6687 21675
rect 7113 21641 7147 21675
rect 10793 21641 10827 21675
rect 12725 21641 12759 21675
rect 14749 21641 14783 21675
rect 15393 21641 15427 21675
rect 19073 21641 19107 21675
rect 20269 21641 20303 21675
rect 20453 21641 20487 21675
rect 21833 21641 21867 21675
rect 22017 21641 22051 21675
rect 23029 21641 23063 21675
rect 25605 21641 25639 21675
rect 4629 21573 4663 21607
rect 16957 21573 16991 21607
rect 17693 21573 17727 21607
rect 17785 21573 17819 21607
rect 19809 21573 19843 21607
rect 2053 21505 2087 21539
rect 4353 21505 4387 21539
rect 5825 21505 5859 21539
rect 11989 21505 12023 21539
rect 18613 21505 18647 21539
rect 19441 21505 19475 21539
rect 20913 21505 20947 21539
rect 21097 21505 21131 21539
rect 21557 21505 21591 21539
rect 22569 21505 22603 21539
rect 24501 21505 24535 21539
rect 1409 21437 1443 21471
rect 2513 21437 2547 21471
rect 3065 21437 3099 21471
rect 6193 21437 6227 21471
rect 7205 21437 7239 21471
rect 7461 21437 7495 21471
rect 9413 21437 9447 21471
rect 13369 21437 13403 21471
rect 15577 21437 15611 21471
rect 15833 21437 15867 21471
rect 17693 21437 17727 21471
rect 18521 21437 18555 21471
rect 20821 21437 20855 21471
rect 22477 21437 22511 21471
rect 24225 21437 24259 21471
rect 25421 21437 25455 21471
rect 25973 21437 26007 21471
rect 5641 21369 5675 21403
rect 9658 21369 9692 21403
rect 13636 21369 13670 21403
rect 15025 21369 15059 21403
rect 24317 21369 24351 21403
rect 2329 21301 2363 21335
rect 2697 21301 2731 21335
rect 5181 21301 5215 21335
rect 5549 21301 5583 21335
rect 8585 21301 8619 21335
rect 8861 21301 8895 21335
rect 9321 21301 9355 21335
rect 11069 21301 11103 21335
rect 11529 21301 11563 21335
rect 13277 21301 13311 21335
rect 17417 21301 17451 21335
rect 18061 21301 18095 21335
rect 18429 21301 18463 21335
rect 22385 21301 22419 21335
rect 23489 21301 23523 21335
rect 23857 21301 23891 21335
rect 24961 21301 24995 21335
rect 25329 21301 25363 21335
rect 1593 21097 1627 21131
rect 2697 21097 2731 21131
rect 3157 21097 3191 21131
rect 3525 21097 3559 21131
rect 4905 21097 4939 21131
rect 6285 21097 6319 21131
rect 6929 21097 6963 21131
rect 8033 21097 8067 21131
rect 9873 21097 9907 21131
rect 13645 21097 13679 21131
rect 16405 21097 16439 21131
rect 16589 21097 16623 21131
rect 18153 21097 18187 21131
rect 19533 21097 19567 21131
rect 21005 21097 21039 21131
rect 23397 21097 23431 21131
rect 25145 21097 25179 21131
rect 2237 21029 2271 21063
rect 4445 21029 4479 21063
rect 6837 21029 6871 21063
rect 11060 21029 11094 21063
rect 12449 21029 12483 21063
rect 13093 21029 13127 21063
rect 14105 21029 14139 21063
rect 15577 21029 15611 21063
rect 1409 20961 1443 20995
rect 2513 20961 2547 20995
rect 5273 20961 5307 20995
rect 5365 20961 5399 20995
rect 7573 20961 7607 20995
rect 8401 20961 8435 20995
rect 8493 20961 8527 20995
rect 9689 20961 9723 20995
rect 10793 20961 10827 20995
rect 14013 20961 14047 20995
rect 15301 20961 15335 20995
rect 16957 20961 16991 20995
rect 18521 20961 18555 20995
rect 19717 20961 19751 20995
rect 21373 20961 21407 20995
rect 23765 20961 23799 20995
rect 23857 20961 23891 20995
rect 24777 20961 24811 20995
rect 24961 20961 24995 20995
rect 5457 20893 5491 20927
rect 7021 20893 7055 20927
rect 7941 20893 7975 20927
rect 8585 20893 8619 20927
rect 9413 20893 9447 20927
rect 14289 20893 14323 20927
rect 17049 20893 17083 20927
rect 17233 20893 17267 20927
rect 18613 20893 18647 20927
rect 18797 20893 18831 20927
rect 21465 20893 21499 20927
rect 21649 20893 21683 20927
rect 22937 20893 22971 20927
rect 23949 20893 23983 20927
rect 4813 20825 4847 20859
rect 6469 20825 6503 20859
rect 10609 20825 10643 20859
rect 13461 20825 13495 20859
rect 14749 20825 14783 20859
rect 16129 20825 16163 20859
rect 18061 20825 18095 20859
rect 19901 20825 19935 20859
rect 22109 20825 22143 20859
rect 23305 20825 23339 20859
rect 3893 20757 3927 20791
rect 6009 20757 6043 20791
rect 9137 20757 9171 20791
rect 10333 20757 10367 20791
rect 12173 20757 12207 20791
rect 15117 20757 15151 20791
rect 17601 20757 17635 20791
rect 19165 20757 19199 20791
rect 20545 20757 20579 20791
rect 22385 20757 22419 20791
rect 24409 20757 24443 20791
rect 2697 20553 2731 20587
rect 5181 20553 5215 20587
rect 6837 20553 6871 20587
rect 8125 20553 8159 20587
rect 8585 20553 8619 20587
rect 10149 20553 10183 20587
rect 13737 20553 13771 20587
rect 14197 20553 14231 20587
rect 14381 20553 14415 20587
rect 16405 20553 16439 20587
rect 21005 20553 21039 20587
rect 24961 20553 24995 20587
rect 25421 20553 25455 20587
rect 2053 20485 2087 20519
rect 9597 20485 9631 20519
rect 15485 20485 15519 20519
rect 18061 20485 18095 20519
rect 19165 20485 19199 20519
rect 22477 20485 22511 20519
rect 5733 20417 5767 20451
rect 7297 20417 7331 20451
rect 7389 20417 7423 20451
rect 8493 20417 8527 20451
rect 9229 20417 9263 20451
rect 10701 20417 10735 20451
rect 13001 20417 13035 20451
rect 14841 20417 14875 20451
rect 14933 20417 14967 20451
rect 16221 20417 16255 20451
rect 16957 20417 16991 20451
rect 18613 20417 18647 20451
rect 20177 20417 20211 20451
rect 20729 20417 20763 20451
rect 21741 20417 21775 20451
rect 22201 20417 22235 20451
rect 1409 20349 1443 20383
rect 2513 20349 2547 20383
rect 3433 20349 3467 20383
rect 3617 20349 3651 20383
rect 4169 20349 4203 20383
rect 5641 20349 5675 20383
rect 6653 20349 6687 20383
rect 10609 20349 10643 20383
rect 18429 20349 18463 20383
rect 18521 20349 18555 20383
rect 19993 20349 20027 20383
rect 21557 20349 21591 20383
rect 3157 20281 3191 20315
rect 4629 20281 4663 20315
rect 5549 20281 5583 20315
rect 8953 20281 8987 20315
rect 12265 20281 12299 20315
rect 12909 20281 12943 20315
rect 16865 20281 16899 20315
rect 22661 20417 22695 20451
rect 24133 20417 24167 20451
rect 24317 20417 24351 20451
rect 25237 20349 25271 20383
rect 25789 20349 25823 20383
rect 24041 20281 24075 20315
rect 1593 20213 1627 20247
rect 2421 20213 2455 20247
rect 3801 20213 3835 20247
rect 4997 20213 5031 20247
rect 6193 20213 6227 20247
rect 7205 20213 7239 20247
rect 9045 20213 9079 20247
rect 9965 20213 9999 20247
rect 10517 20213 10551 20247
rect 11253 20213 11287 20247
rect 11529 20213 11563 20247
rect 12449 20213 12483 20247
rect 12817 20213 12851 20247
rect 14749 20213 14783 20247
rect 15945 20213 15979 20247
rect 16773 20213 16807 20247
rect 17417 20213 17451 20247
rect 17877 20213 17911 20247
rect 19441 20213 19475 20247
rect 19625 20213 19659 20247
rect 20085 20213 20119 20247
rect 21189 20213 21223 20247
rect 21649 20213 21683 20247
rect 22477 20213 22511 20247
rect 23029 20213 23063 20247
rect 23489 20213 23523 20247
rect 23673 20213 23707 20247
rect 4261 20009 4295 20043
rect 4721 20009 4755 20043
rect 5733 20009 5767 20043
rect 7573 20009 7607 20043
rect 8033 20009 8067 20043
rect 9873 20009 9907 20043
rect 11069 20009 11103 20043
rect 11529 20009 11563 20043
rect 12541 20009 12575 20043
rect 14381 20009 14415 20043
rect 15117 20009 15151 20043
rect 15301 20009 15335 20043
rect 18521 20009 18555 20043
rect 18981 20009 19015 20043
rect 20085 20009 20119 20043
rect 22477 20009 22511 20043
rect 24041 20009 24075 20043
rect 25053 20009 25087 20043
rect 1961 19941 1995 19975
rect 9413 19941 9447 19975
rect 11437 19941 11471 19975
rect 14657 19941 14691 19975
rect 16221 19941 16255 19975
rect 21373 19941 21407 19975
rect 24409 19941 24443 19975
rect 1685 19873 1719 19907
rect 4629 19873 4663 19907
rect 5365 19873 5399 19907
rect 5825 19873 5859 19907
rect 6092 19873 6126 19907
rect 8401 19873 8435 19907
rect 10057 19873 10091 19907
rect 12909 19873 12943 19907
rect 13268 19873 13302 19907
rect 16313 19873 16347 19907
rect 16569 19873 16603 19907
rect 18889 19873 18923 19907
rect 21281 19873 21315 19907
rect 22845 19873 22879 19907
rect 25421 19873 25455 19907
rect 3709 19805 3743 19839
rect 4905 19805 4939 19839
rect 8493 19805 8527 19839
rect 8677 19805 8711 19839
rect 11621 19805 11655 19839
rect 13001 19805 13035 19839
rect 19073 19805 19107 19839
rect 21557 19805 21591 19839
rect 22937 19805 22971 19839
rect 23121 19805 23155 19839
rect 24501 19805 24535 19839
rect 24685 19805 24719 19839
rect 7941 19737 7975 19771
rect 12081 19737 12115 19771
rect 22385 19737 22419 19771
rect 2421 19669 2455 19703
rect 2881 19669 2915 19703
rect 3249 19669 3283 19703
rect 7205 19669 7239 19703
rect 9137 19669 9171 19703
rect 10885 19669 10919 19703
rect 15853 19669 15887 19703
rect 17693 19669 17727 19703
rect 18245 19669 18279 19703
rect 19717 19669 19751 19703
rect 20361 19669 20395 19703
rect 20913 19669 20947 19703
rect 21925 19669 21959 19703
rect 23765 19669 23799 19703
rect 25789 19669 25823 19703
rect 4721 19465 4755 19499
rect 8401 19465 8435 19499
rect 10793 19465 10827 19499
rect 11805 19465 11839 19499
rect 12449 19465 12483 19499
rect 15669 19465 15703 19499
rect 18061 19465 18095 19499
rect 22477 19465 22511 19499
rect 23673 19465 23707 19499
rect 2605 19329 2639 19363
rect 4261 19329 4295 19363
rect 5825 19329 5859 19363
rect 7481 19329 7515 19363
rect 11437 19329 11471 19363
rect 12173 19329 12207 19363
rect 13001 19329 13035 19363
rect 14565 19329 14599 19363
rect 15761 19329 15795 19363
rect 18613 19329 18647 19363
rect 20177 19329 20211 19363
rect 21741 19329 21775 19363
rect 24317 19329 24351 19363
rect 3525 19261 3559 19295
rect 4077 19261 4111 19295
rect 5641 19261 5675 19295
rect 6653 19261 6687 19295
rect 7297 19261 7331 19295
rect 8585 19261 8619 19295
rect 10241 19261 10275 19295
rect 12909 19261 12943 19295
rect 13921 19261 13955 19295
rect 14473 19261 14507 19295
rect 15301 19261 15335 19295
rect 16017 19261 16051 19295
rect 17417 19261 17451 19295
rect 18429 19261 18463 19295
rect 19073 19261 19107 19295
rect 19533 19261 19567 19295
rect 19993 19261 20027 19295
rect 21005 19261 21039 19295
rect 21557 19261 21591 19295
rect 22937 19261 22971 19295
rect 24133 19261 24167 19295
rect 25053 19261 25087 19295
rect 25237 19261 25271 19295
rect 25789 19261 25823 19295
rect 26249 19261 26283 19295
rect 5549 19193 5583 19227
rect 7205 19193 7239 19227
rect 8830 19193 8864 19227
rect 10701 19193 10735 19227
rect 11161 19193 11195 19227
rect 11253 19193 11287 19227
rect 14381 19193 14415 19227
rect 21649 19193 21683 19227
rect 24041 19193 24075 19227
rect 949 19125 983 19159
rect 1869 19125 1903 19159
rect 2053 19125 2087 19159
rect 2421 19125 2455 19159
rect 2513 19125 2547 19159
rect 3065 19125 3099 19159
rect 3617 19125 3651 19159
rect 3985 19125 4019 19159
rect 4997 19125 5031 19159
rect 5181 19125 5215 19159
rect 6193 19125 6227 19159
rect 6837 19125 6871 19159
rect 8033 19125 8067 19159
rect 9965 19125 9999 19159
rect 12817 19125 12851 19159
rect 13461 19125 13495 19159
rect 14013 19125 14047 19159
rect 17141 19125 17175 19159
rect 17785 19125 17819 19159
rect 18521 19125 18555 19159
rect 19625 19125 19659 19159
rect 20085 19125 20119 19159
rect 20729 19125 20763 19159
rect 21189 19125 21223 19159
rect 23397 19125 23431 19159
rect 24777 19125 24811 19159
rect 25421 19125 25455 19159
rect 857 15521 891 15555
rect 857 12325 891 12359
rect 2329 18921 2363 18955
rect 2789 18921 2823 18955
rect 2881 18921 2915 18955
rect 3709 18921 3743 18955
rect 4261 18921 4295 18955
rect 4721 18921 4755 18955
rect 5365 18921 5399 18955
rect 5733 18921 5767 18955
rect 8309 18921 8343 18955
rect 8953 18921 8987 18955
rect 11161 18921 11195 18955
rect 14197 18921 14231 18955
rect 15853 18921 15887 18955
rect 16589 18921 16623 18955
rect 21925 18921 21959 18955
rect 22937 18921 22971 18955
rect 23673 18921 23707 18955
rect 24041 18921 24075 18955
rect 24501 18921 24535 18955
rect 25053 18921 25087 18955
rect 6377 18853 6411 18887
rect 8585 18853 8619 18887
rect 11529 18853 11563 18887
rect 13062 18853 13096 18887
rect 14473 18853 14507 18887
rect 19349 18853 19383 18887
rect 22385 18853 22419 18887
rect 24409 18853 24443 18887
rect 25421 18853 25455 18887
rect 4077 18785 4111 18819
rect 5181 18785 5215 18819
rect 6929 18785 6963 18819
rect 7196 18785 7230 18819
rect 12817 18785 12851 18819
rect 15669 18785 15703 18819
rect 16773 18785 16807 18819
rect 17029 18785 17063 18819
rect 19441 18785 19475 18819
rect 21281 18785 21315 18819
rect 22845 18785 22879 18819
rect 3065 18717 3099 18751
rect 5825 18717 5859 18751
rect 6009 18717 6043 18751
rect 11621 18717 11655 18751
rect 11713 18717 11747 18751
rect 19533 18717 19567 18751
rect 21373 18717 21407 18751
rect 21557 18717 21591 18751
rect 23121 18717 23155 18751
rect 24593 18717 24627 18751
rect 15485 18649 15519 18683
rect 20913 18649 20947 18683
rect 22477 18649 22511 18683
rect 1961 18581 1995 18615
rect 2421 18581 2455 18615
rect 6837 18581 6871 18615
rect 9321 18581 9355 18615
rect 9873 18581 9907 18615
rect 10333 18581 10367 18615
rect 10885 18581 10919 18615
rect 12541 18581 12575 18615
rect 14841 18581 14875 18615
rect 16313 18581 16347 18615
rect 18153 18581 18187 18615
rect 18521 18581 18555 18615
rect 18981 18581 19015 18615
rect 20085 18581 20119 18615
rect 20729 18581 20763 18615
rect 25881 18581 25915 18615
rect 3065 18377 3099 18411
rect 4629 18377 4663 18411
rect 5089 18377 5123 18411
rect 6285 18377 6319 18411
rect 13461 18377 13495 18411
rect 14013 18377 14047 18411
rect 15669 18377 15703 18411
rect 15853 18377 15887 18411
rect 16221 18377 16255 18411
rect 18061 18377 18095 18411
rect 19625 18377 19659 18411
rect 23673 18377 23707 18411
rect 3433 18309 3467 18343
rect 7021 18309 7055 18343
rect 2605 18241 2639 18275
rect 4261 18241 4295 18275
rect 5733 18241 5767 18275
rect 7481 18241 7515 18275
rect 7573 18241 7607 18275
rect 8493 18241 8527 18275
rect 9045 18241 9079 18275
rect 9137 18241 9171 18275
rect 9873 18241 9907 18275
rect 10057 18241 10091 18275
rect 13001 18241 13035 18275
rect 14565 18241 14599 18275
rect 3985 18173 4019 18207
rect 4077 18173 4111 18207
rect 6653 18173 6687 18207
rect 8953 18173 8987 18207
rect 2421 18105 2455 18139
rect 5549 18105 5583 18139
rect 7389 18105 7423 18139
rect 10149 18173 10183 18207
rect 10416 18173 10450 18207
rect 11805 18173 11839 18207
rect 14473 18173 14507 18207
rect 12909 18105 12943 18139
rect 24685 18309 24719 18343
rect 16773 18241 16807 18275
rect 18705 18241 18739 18275
rect 19349 18241 19383 18275
rect 19533 18241 19567 18275
rect 20269 18241 20303 18275
rect 21833 18241 21867 18275
rect 24133 18241 24167 18275
rect 24225 18241 24259 18275
rect 25513 18241 25547 18275
rect 26341 18241 26375 18275
rect 16037 18105 16071 18139
rect 16681 18105 16715 18139
rect 17785 18105 17819 18139
rect 18429 18105 18463 18139
rect 21649 18173 21683 18207
rect 24041 18173 24075 18207
rect 25237 18173 25271 18207
rect 25973 18173 26007 18207
rect 19993 18105 20027 18139
rect 20085 18105 20119 18139
rect 20729 18105 20763 18139
rect 21557 18105 21591 18139
rect 22937 18105 22971 18139
rect 1869 18037 1903 18071
rect 2053 18037 2087 18071
rect 2513 18037 2547 18071
rect 3617 18037 3651 18071
rect 5181 18037 5215 18071
rect 5641 18037 5675 18071
rect 8033 18037 8067 18071
rect 8585 18037 8619 18071
rect 9689 18037 9723 18071
rect 9873 18037 9907 18071
rect 11529 18037 11563 18071
rect 12173 18037 12207 18071
rect 12449 18037 12483 18071
rect 12817 18037 12851 18071
rect 13921 18037 13955 18071
rect 14381 18037 14415 18071
rect 15117 18037 15151 18071
rect 15853 18037 15887 18071
rect 16589 18037 16623 18071
rect 17417 18037 17451 18071
rect 18521 18037 18555 18071
rect 19073 18037 19107 18071
rect 19257 18037 19291 18071
rect 21005 18037 21039 18071
rect 21189 18037 21223 18071
rect 22569 18037 22603 18071
rect 23397 18037 23431 18071
rect 25145 18037 25179 18071
rect 2421 17833 2455 17867
rect 4353 17833 4387 17867
rect 4537 17833 4571 17867
rect 7757 17833 7791 17867
rect 8493 17833 8527 17867
rect 8861 17833 8895 17867
rect 10701 17833 10735 17867
rect 13645 17833 13679 17867
rect 14197 17833 14231 17867
rect 15117 17833 15151 17867
rect 15301 17833 15335 17867
rect 15761 17833 15795 17867
rect 16405 17833 16439 17867
rect 16865 17833 16899 17867
rect 19073 17833 19107 17867
rect 20177 17833 20211 17867
rect 20729 17833 20763 17867
rect 22477 17833 22511 17867
rect 23305 17833 23339 17867
rect 24225 17833 24259 17867
rect 25421 17833 25455 17867
rect 2789 17765 2823 17799
rect 4905 17765 4939 17799
rect 9689 17765 9723 17799
rect 10609 17765 10643 17799
rect 11161 17765 11195 17799
rect 11805 17765 11839 17799
rect 12541 17765 12575 17799
rect 19625 17765 19659 17799
rect 21189 17765 21223 17799
rect 24869 17765 24903 17799
rect 6357 17697 6391 17731
rect 8309 17697 8343 17731
rect 9229 17697 9263 17731
rect 11069 17697 11103 17731
rect 13001 17697 13035 17731
rect 15669 17697 15703 17731
rect 17141 17697 17175 17731
rect 17408 17697 17442 17731
rect 19349 17697 19383 17731
rect 21649 17697 21683 17731
rect 23213 17697 23247 17731
rect 24777 17697 24811 17731
rect 2881 17629 2915 17663
rect 3065 17629 3099 17663
rect 4997 17629 5031 17663
rect 5089 17629 5123 17663
rect 5917 17629 5951 17663
rect 6101 17629 6135 17663
rect 11345 17629 11379 17663
rect 13093 17629 13127 17663
rect 13185 17629 13219 17663
rect 15853 17629 15887 17663
rect 21741 17629 21775 17663
rect 21833 17629 21867 17663
rect 23397 17629 23431 17663
rect 24961 17629 24995 17663
rect 12173 17561 12207 17595
rect 22845 17561 22879 17595
rect 24409 17561 24443 17595
rect 25789 17561 25823 17595
rect 1685 17493 1719 17527
rect 2145 17493 2179 17527
rect 3617 17493 3651 17527
rect 5641 17493 5675 17527
rect 7481 17493 7515 17527
rect 8125 17493 8159 17527
rect 10149 17493 10183 17527
rect 12633 17493 12667 17527
rect 14013 17493 14047 17527
rect 14749 17493 14783 17527
rect 18521 17493 18555 17527
rect 21281 17493 21315 17527
rect 23949 17493 23983 17527
rect 26249 17493 26283 17527
rect 1593 17289 1627 17323
rect 2605 17289 2639 17323
rect 5825 17289 5859 17323
rect 7021 17289 7055 17323
rect 8125 17289 8159 17323
rect 9505 17289 9539 17323
rect 11069 17289 11103 17323
rect 14841 17289 14875 17323
rect 18061 17289 18095 17323
rect 19165 17289 19199 17323
rect 19625 17289 19659 17323
rect 25053 17289 25087 17323
rect 26341 17289 26375 17323
rect 2513 17221 2547 17255
rect 4261 17221 4295 17255
rect 6193 17221 6227 17255
rect 11345 17221 11379 17255
rect 17141 17221 17175 17255
rect 24777 17221 24811 17255
rect 2237 17153 2271 17187
rect 3709 17153 3743 17187
rect 4629 17153 4663 17187
rect 5181 17153 5215 17187
rect 5273 17153 5307 17187
rect 8033 17153 8067 17187
rect 8769 17153 8803 17187
rect 11713 17153 11747 17187
rect 13553 17153 13587 17187
rect 17877 17153 17911 17187
rect 18705 17153 18739 17187
rect 19533 17153 19567 17187
rect 20177 17153 20211 17187
rect 22385 17153 22419 17187
rect 24317 17153 24351 17187
rect 25421 17153 25455 17187
rect 3065 17085 3099 17119
rect 5089 17085 5123 17119
rect 6837 17085 6871 17119
rect 7389 17085 7423 17119
rect 8493 17085 8527 17119
rect 9689 17085 9723 17119
rect 9945 17085 9979 17119
rect 13369 17085 13403 17119
rect 14473 17085 14507 17119
rect 14657 17085 14691 17119
rect 15761 17085 15795 17119
rect 18521 17085 18555 17119
rect 23029 17085 23063 17119
rect 24133 17085 24167 17119
rect 25237 17085 25271 17119
rect 25973 17085 26007 17119
rect 1961 17017 1995 17051
rect 2513 17017 2547 17051
rect 9137 17017 9171 17051
rect 12265 17017 12299 17051
rect 12817 17017 12851 17051
rect 16028 17017 16062 17051
rect 17417 17017 17451 17051
rect 18429 17017 18463 17051
rect 19993 17017 20027 17051
rect 2053 16949 2087 16983
rect 3157 16949 3191 16983
rect 3525 16949 3559 16983
rect 3617 16949 3651 16983
rect 4721 16949 4755 16983
rect 6561 16949 6595 16983
rect 8585 16949 8619 16983
rect 12909 16949 12943 16983
rect 13277 16949 13311 16983
rect 14013 16949 14047 16983
rect 15301 16949 15335 16983
rect 20085 16949 20119 16983
rect 20913 16949 20947 16983
rect 21281 16949 21315 16983
rect 21649 16949 21683 16983
rect 21833 16949 21867 16983
rect 22201 16949 22235 16983
rect 22293 16949 22327 16983
rect 23397 16949 23431 16983
rect 23673 16949 23707 16983
rect 24041 16949 24075 16983
rect 2973 16745 3007 16779
rect 3893 16745 3927 16779
rect 5641 16745 5675 16779
rect 6009 16745 6043 16779
rect 7205 16745 7239 16779
rect 7665 16745 7699 16779
rect 8401 16745 8435 16779
rect 8677 16745 8711 16779
rect 9045 16745 9079 16779
rect 9413 16745 9447 16779
rect 11069 16745 11103 16779
rect 11345 16745 11379 16779
rect 13737 16745 13771 16779
rect 14381 16745 14415 16779
rect 14657 16745 14691 16779
rect 16681 16745 16715 16779
rect 17233 16745 17267 16779
rect 17509 16745 17543 16779
rect 19901 16745 19935 16779
rect 20361 16745 20395 16779
rect 21281 16745 21315 16779
rect 23121 16745 23155 16779
rect 24777 16745 24811 16779
rect 24961 16745 24995 16779
rect 1777 16677 1811 16711
rect 2421 16677 2455 16711
rect 2697 16677 2731 16711
rect 2881 16677 2915 16711
rect 12326 16677 12360 16711
rect 15025 16677 15059 16711
rect 18788 16677 18822 16711
rect 21618 16677 21652 16711
rect 24041 16677 24075 16711
rect 24409 16677 24443 16711
rect 24593 16677 24627 16711
rect 1869 16541 1903 16575
rect 2053 16541 2087 16575
rect 4445 16609 4479 16643
rect 4537 16609 4571 16643
rect 5457 16609 5491 16643
rect 6653 16609 6687 16643
rect 7021 16609 7055 16643
rect 7573 16609 7607 16643
rect 9956 16609 9990 16643
rect 11805 16609 11839 16643
rect 15301 16609 15335 16643
rect 15568 16609 15602 16643
rect 18521 16609 18555 16643
rect 23949 16609 23983 16643
rect 4629 16541 4663 16575
rect 6101 16541 6135 16575
rect 6193 16541 6227 16575
rect 7757 16541 7791 16575
rect 9689 16541 9723 16575
rect 12081 16541 12115 16575
rect 21373 16541 21407 16575
rect 23489 16541 23523 16575
rect 24133 16541 24167 16575
rect 2697 16473 2731 16507
rect 13461 16473 13495 16507
rect 23581 16473 23615 16507
rect 25145 16609 25179 16643
rect 25421 16609 25455 16643
rect 24777 16541 24811 16575
rect 25881 16541 25915 16575
rect 26249 16541 26283 16575
rect 1409 16405 1443 16439
rect 3433 16405 3467 16439
rect 4077 16405 4111 16439
rect 5181 16405 5215 16439
rect 18153 16405 18187 16439
rect 20729 16405 20763 16439
rect 22753 16405 22787 16439
rect 24409 16405 24443 16439
rect 3893 16201 3927 16235
rect 6101 16201 6135 16235
rect 7941 16201 7975 16235
rect 10333 16201 10367 16235
rect 10517 16201 10551 16235
rect 11621 16201 11655 16235
rect 12081 16201 12115 16235
rect 13001 16201 13035 16235
rect 15761 16201 15795 16235
rect 17049 16201 17083 16235
rect 19073 16201 19107 16235
rect 21833 16201 21867 16235
rect 23397 16201 23431 16235
rect 23673 16201 23707 16235
rect 25421 16201 25455 16235
rect 26249 16201 26283 16235
rect 4445 16133 4479 16167
rect 15117 16133 15151 16167
rect 17509 16133 17543 16167
rect 21373 16133 21407 16167
rect 2053 16065 2087 16099
rect 4353 16065 4387 16099
rect 4997 16065 5031 16099
rect 7113 16065 7147 16099
rect 8309 16065 8343 16099
rect 10977 16065 11011 16099
rect 11069 16065 11103 16099
rect 13737 16065 13771 16099
rect 16405 16065 16439 16099
rect 16497 16065 16531 16099
rect 18705 16065 18739 16099
rect 19625 16065 19659 16099
rect 22477 16065 22511 16099
rect 24133 16065 24167 16099
rect 24317 16065 24351 16099
rect 24777 16065 24811 16099
rect 1777 15997 1811 16031
rect 2973 15997 3007 16031
rect 4813 15997 4847 16031
rect 6837 15997 6871 16031
rect 8565 15997 8599 16031
rect 15393 15997 15427 16031
rect 16313 15997 16347 16031
rect 17693 15997 17727 16031
rect 18429 15997 18463 16031
rect 25237 15997 25271 16031
rect 25789 15997 25823 16031
rect 3249 15929 3283 15963
rect 5733 15929 5767 15963
rect 10057 15929 10091 15963
rect 12449 15929 12483 15963
rect 14004 15929 14038 15963
rect 18521 15929 18555 15963
rect 19533 15929 19567 15963
rect 19870 15929 19904 15963
rect 21649 15929 21683 15963
rect 22293 15929 22327 15963
rect 24041 15929 24075 15963
rect 1409 15861 1443 15895
rect 1869 15861 1903 15895
rect 2513 15861 2547 15895
rect 2881 15861 2915 15895
rect 4905 15861 4939 15895
rect 6561 15861 6595 15895
rect 7665 15861 7699 15895
rect 9689 15861 9723 15895
rect 10885 15861 10919 15895
rect 13645 15861 13679 15895
rect 15945 15861 15979 15895
rect 17325 15861 17359 15895
rect 18061 15861 18095 15895
rect 21005 15861 21039 15895
rect 22201 15861 22235 15895
rect 23121 15861 23155 15895
rect 25053 15861 25087 15895
rect 6009 15657 6043 15691
rect 6561 15657 6595 15691
rect 9413 15657 9447 15691
rect 9873 15657 9907 15691
rect 10885 15657 10919 15691
rect 12449 15657 12483 15691
rect 14289 15657 14323 15691
rect 16313 15657 16347 15691
rect 21281 15657 21315 15691
rect 23029 15657 23063 15691
rect 23581 15657 23615 15691
rect 24041 15657 24075 15691
rect 25053 15657 25087 15691
rect 25329 15657 25363 15691
rect 6377 15589 6411 15623
rect 8401 15589 8435 15623
rect 13176 15589 13210 15623
rect 15669 15589 15703 15623
rect 16129 15589 16163 15623
rect 18061 15589 18095 15623
rect 23489 15589 23523 15623
rect 25697 15589 25731 15623
rect 26065 15589 26099 15623
rect 1777 15521 1811 15555
rect 4620 15521 4654 15555
rect 6929 15521 6963 15555
rect 7941 15521 7975 15555
rect 8125 15521 8159 15555
rect 9689 15521 9723 15555
rect 11253 15521 11287 15555
rect 12909 15521 12943 15555
rect 15761 15521 15795 15555
rect 1869 15453 1903 15487
rect 2053 15453 2087 15487
rect 4353 15453 4387 15487
rect 7021 15453 7055 15487
rect 7113 15453 7147 15487
rect 11345 15453 11379 15487
rect 11437 15453 11471 15487
rect 15945 15453 15979 15487
rect 3709 15385 3743 15419
rect 5733 15385 5767 15419
rect 14657 15385 14691 15419
rect 15301 15385 15335 15419
rect 17417 15521 17451 15555
rect 17509 15521 17543 15555
rect 18521 15521 18555 15555
rect 18880 15521 18914 15555
rect 20729 15521 20763 15555
rect 21640 15521 21674 15555
rect 23949 15521 23983 15555
rect 25145 15521 25179 15555
rect 17693 15453 17727 15487
rect 18613 15453 18647 15487
rect 20269 15453 20303 15487
rect 21373 15453 21407 15487
rect 24133 15453 24167 15487
rect 16865 15385 16899 15419
rect 22753 15385 22787 15419
rect 1409 15317 1443 15351
rect 2421 15317 2455 15351
rect 2973 15317 3007 15351
rect 3433 15317 3467 15351
rect 7665 15317 7699 15351
rect 8861 15317 8895 15351
rect 10333 15317 10367 15351
rect 10701 15317 10735 15351
rect 11897 15317 11931 15351
rect 15025 15317 15059 15351
rect 16129 15317 16163 15351
rect 17049 15317 17083 15351
rect 19993 15317 20027 15351
rect 24593 15317 24627 15351
rect 3709 15113 3743 15147
rect 6837 15113 6871 15147
rect 8401 15113 8435 15147
rect 9413 15113 9447 15147
rect 9689 15113 9723 15147
rect 9965 15113 9999 15147
rect 11437 15113 11471 15147
rect 11989 15113 12023 15147
rect 12817 15113 12851 15147
rect 13461 15113 13495 15147
rect 15025 15113 15059 15147
rect 16313 15113 16347 15147
rect 19165 15113 19199 15147
rect 19625 15113 19659 15147
rect 20729 15113 20763 15147
rect 22109 15113 22143 15147
rect 22753 15113 22787 15147
rect 23673 15113 23707 15147
rect 24685 15113 24719 15147
rect 25973 15113 26007 15147
rect 2421 15045 2455 15079
rect 6285 15045 6319 15079
rect 2973 14977 3007 15011
rect 4537 14977 4571 15011
rect 7297 14977 7331 15011
rect 7389 14977 7423 15011
rect 7941 14977 7975 15011
rect 9045 14977 9079 15011
rect 1685 14909 1719 14943
rect 2789 14909 2823 14943
rect 4804 14909 4838 14943
rect 7205 14909 7239 14943
rect 8309 14909 8343 14943
rect 8769 14909 8803 14943
rect 3985 14841 4019 14875
rect 6561 14841 6595 14875
rect 8861 14841 8895 14875
rect 11529 15045 11563 15079
rect 15577 15045 15611 15079
rect 16405 15045 16439 15079
rect 17601 15045 17635 15079
rect 21189 15045 21223 15079
rect 10517 14977 10551 15011
rect 14381 14977 14415 15011
rect 14473 14977 14507 15011
rect 15393 14977 15427 15011
rect 11069 14909 11103 14943
rect 11713 14909 11747 14943
rect 13737 14909 13771 14943
rect 14289 14909 14323 14943
rect 16865 14977 16899 15011
rect 17049 14977 17083 15011
rect 9873 14841 9907 14875
rect 10333 14841 10367 14875
rect 15577 14841 15611 14875
rect 15761 14841 15795 14875
rect 16773 14841 16807 14875
rect 18705 14977 18739 15011
rect 19533 14977 19567 15011
rect 20177 14977 20211 15011
rect 21649 14977 21683 15011
rect 21741 14977 21775 15011
rect 17877 14909 17911 14943
rect 18429 14909 18463 14943
rect 21097 14909 21131 14943
rect 18521 14841 18555 14875
rect 20085 14841 20119 14875
rect 23489 15045 23523 15079
rect 24317 14977 24351 15011
rect 25421 14977 25455 15011
rect 24041 14909 24075 14943
rect 25237 14909 25271 14943
rect 25053 14841 25087 14875
rect 1961 14773 1995 14807
rect 2881 14773 2915 14807
rect 4445 14773 4479 14807
rect 5917 14773 5951 14807
rect 9689 14773 9723 14807
rect 10425 14773 10459 14807
rect 12909 14773 12943 14807
rect 13921 14773 13955 14807
rect 17417 14773 17451 14807
rect 17601 14773 17635 14807
rect 18061 14773 18095 14807
rect 19993 14773 20027 14807
rect 21557 14773 21591 14807
rect 22109 14773 22143 14807
rect 22293 14773 22327 14807
rect 23121 14773 23155 14807
rect 24133 14773 24167 14807
rect 26341 14773 26375 14807
rect 2789 14569 2823 14603
rect 5733 14569 5767 14603
rect 6469 14569 6503 14603
rect 8493 14569 8527 14603
rect 10149 14569 10183 14603
rect 12541 14569 12575 14603
rect 14473 14569 14507 14603
rect 15117 14569 15151 14603
rect 15669 14569 15703 14603
rect 16865 14569 16899 14603
rect 18889 14569 18923 14603
rect 20269 14569 20303 14603
rect 20637 14569 20671 14603
rect 23857 14569 23891 14603
rect 25421 14569 25455 14603
rect 1869 14501 1903 14535
rect 2237 14501 2271 14535
rect 3801 14501 3835 14535
rect 6101 14501 6135 14535
rect 6990 14501 7024 14535
rect 10057 14501 10091 14535
rect 13185 14501 13219 14535
rect 15761 14501 15795 14535
rect 16497 14501 16531 14535
rect 17408 14501 17442 14535
rect 23765 14501 23799 14535
rect 24961 14501 24995 14535
rect 1777 14433 1811 14467
rect 1961 14365 1995 14399
rect 3433 14433 3467 14467
rect 4077 14433 4111 14467
rect 4344 14433 4378 14467
rect 6653 14433 6687 14467
rect 9137 14433 9171 14467
rect 11621 14433 11655 14467
rect 13277 14433 13311 14467
rect 17049 14433 17083 14467
rect 19617 14433 19651 14467
rect 19742 14433 19776 14467
rect 21905 14433 21939 14467
rect 24225 14433 24259 14467
rect 24317 14433 24351 14467
rect 2973 14365 3007 14399
rect 6745 14365 6779 14399
rect 10241 14365 10275 14399
rect 11713 14365 11747 14399
rect 11897 14365 11931 14399
rect 13369 14365 13403 14399
rect 15853 14365 15887 14399
rect 17141 14365 17175 14399
rect 19349 14365 19383 14399
rect 21649 14365 21683 14399
rect 23397 14365 23431 14399
rect 24501 14365 24535 14399
rect 2237 14297 2271 14331
rect 8769 14297 8803 14331
rect 9505 14297 9539 14331
rect 15301 14297 15335 14331
rect 19901 14297 19935 14331
rect 23029 14297 23063 14331
rect 1409 14229 1443 14263
rect 2421 14229 2455 14263
rect 5457 14229 5491 14263
rect 8125 14229 8159 14263
rect 8953 14229 8987 14263
rect 9689 14229 9723 14263
rect 10885 14229 10919 14263
rect 11253 14229 11287 14263
rect 12817 14229 12851 14263
rect 14013 14229 14047 14263
rect 18521 14229 18555 14263
rect 19441 14229 19475 14263
rect 21189 14229 21223 14263
rect 21557 14229 21591 14263
rect 25237 14229 25271 14263
rect 25973 14229 26007 14263
rect 26249 14229 26283 14263
rect 4813 14025 4847 14059
rect 4997 14025 5031 14059
rect 6193 14025 6227 14059
rect 6837 14025 6871 14059
rect 9965 14025 9999 14059
rect 10241 14025 10275 14059
rect 11897 14025 11931 14059
rect 12173 14025 12207 14059
rect 12449 14025 12483 14059
rect 13645 14025 13679 14059
rect 14013 14025 14047 14059
rect 15669 14025 15703 14059
rect 16405 14025 16439 14059
rect 17417 14025 17451 14059
rect 19441 14025 19475 14059
rect 19717 14025 19751 14059
rect 20913 14025 20947 14059
rect 22661 14025 22695 14059
rect 23029 14025 23063 14059
rect 23673 14025 23707 14059
rect 24685 14025 24719 14059
rect 4169 13957 4203 13991
rect 10793 13957 10827 13991
rect 13461 13957 13495 13991
rect 1685 13889 1719 13923
rect 5549 13889 5583 13923
rect 7389 13889 7423 13923
rect 7849 13889 7883 13923
rect 8493 13889 8527 13923
rect 11437 13889 11471 13923
rect 12909 13889 12943 13923
rect 13001 13889 13035 13923
rect 1501 13821 1535 13855
rect 2789 13821 2823 13855
rect 4537 13821 4571 13855
rect 6653 13821 6687 13855
rect 7297 13821 7331 13855
rect 8585 13821 8619 13855
rect 8852 13821 8886 13855
rect 10701 13821 10735 13855
rect 11253 13821 11287 13855
rect 2605 13753 2639 13787
rect 3034 13753 3068 13787
rect 7205 13753 7239 13787
rect 11161 13753 11195 13787
rect 15301 13957 15335 13991
rect 21833 13957 21867 13991
rect 21925 13957 21959 13991
rect 22385 13957 22419 13991
rect 14657 13889 14691 13923
rect 16313 13889 16347 13923
rect 17049 13889 17083 13923
rect 17785 13889 17819 13923
rect 21465 13889 21499 13923
rect 13921 13821 13955 13855
rect 14473 13821 14507 13855
rect 16865 13821 16899 13855
rect 18061 13821 18095 13855
rect 18328 13821 18362 13855
rect 20729 13821 20763 13855
rect 21373 13821 21407 13855
rect 16773 13753 16807 13787
rect 20453 13753 20487 13787
rect 21281 13753 21315 13787
rect 24225 13889 24259 13923
rect 25421 13889 25455 13923
rect 22477 13821 22511 13855
rect 25237 13821 25271 13855
rect 25973 13821 26007 13855
rect 24133 13753 24167 13787
rect 2237 13685 2271 13719
rect 5365 13685 5399 13719
rect 5457 13685 5491 13719
rect 12817 13685 12851 13719
rect 13645 13685 13679 13719
rect 14381 13685 14415 13719
rect 21833 13685 21867 13719
rect 23397 13685 23431 13719
rect 24041 13685 24075 13719
rect 25053 13685 25087 13719
rect 26341 13685 26375 13719
rect 2421 13481 2455 13515
rect 4445 13481 4479 13515
rect 5549 13481 5583 13515
rect 6377 13481 6411 13515
rect 6469 13481 6503 13515
rect 6929 13481 6963 13515
rect 8033 13481 8067 13515
rect 8401 13481 8435 13515
rect 9689 13481 9723 13515
rect 10149 13481 10183 13515
rect 10885 13481 10919 13515
rect 14657 13481 14691 13515
rect 16957 13481 16991 13515
rect 17325 13481 17359 13515
rect 18153 13481 18187 13515
rect 20269 13481 20303 13515
rect 22109 13481 22143 13515
rect 22753 13481 22787 13515
rect 25421 13481 25455 13515
rect 2789 13413 2823 13447
rect 8493 13413 8527 13447
rect 11682 13413 11716 13447
rect 13093 13413 13127 13447
rect 13461 13413 13495 13447
rect 14013 13413 14047 13447
rect 18880 13413 18914 13447
rect 21189 13413 21223 13447
rect 23029 13413 23063 13447
rect 25237 13413 25271 13447
rect 25881 13413 25915 13447
rect 26249 13413 26283 13447
rect 2881 13345 2915 13379
rect 5089 13345 5123 13379
rect 6837 13345 6871 13379
rect 9413 13345 9447 13379
rect 10057 13345 10091 13379
rect 11437 13345 11471 13379
rect 15568 13345 15602 13379
rect 17509 13345 17543 13379
rect 18613 13345 18647 13379
rect 22017 13345 22051 13379
rect 23213 13345 23247 13379
rect 23480 13345 23514 13379
rect 3065 13277 3099 13311
rect 3525 13277 3559 13311
rect 4537 13277 4571 13311
rect 4629 13277 4663 13311
rect 7113 13277 7147 13311
rect 8677 13277 8711 13311
rect 10241 13277 10275 13311
rect 14105 13277 14139 13311
rect 14289 13277 14323 13311
rect 15025 13277 15059 13311
rect 15301 13277 15335 13311
rect 22293 13277 22327 13311
rect 24869 13277 24903 13311
rect 4077 13209 4111 13243
rect 12817 13209 12851 13243
rect 13645 13209 13679 13243
rect 16681 13209 16715 13243
rect 21649 13209 21683 13243
rect 1685 13141 1719 13175
rect 2329 13141 2363 13175
rect 3801 13141 3835 13175
rect 5825 13141 5859 13175
rect 7481 13141 7515 13175
rect 7941 13141 7975 13175
rect 9137 13141 9171 13175
rect 11253 13141 11287 13175
rect 17693 13141 17727 13175
rect 18521 13141 18555 13175
rect 19993 13141 20027 13175
rect 20729 13141 20763 13175
rect 24593 13141 24627 13175
rect 1593 12937 1627 12971
rect 4721 12937 4755 12971
rect 5825 12937 5859 12971
rect 6193 12937 6227 12971
rect 9045 12937 9079 12971
rect 14197 12937 14231 12971
rect 16037 12937 16071 12971
rect 16773 12937 16807 12971
rect 17509 12937 17543 12971
rect 18429 12937 18463 12971
rect 19441 12937 19475 12971
rect 20269 12937 20303 12971
rect 21189 12937 21223 12971
rect 22201 12937 22235 12971
rect 22661 12937 22695 12971
rect 23305 12937 23339 12971
rect 25053 12937 25087 12971
rect 25329 12937 25363 12971
rect 25697 12937 25731 12971
rect 26065 12937 26099 12971
rect 26433 12937 26467 12971
rect 2697 12869 2731 12903
rect 3157 12869 3191 12903
rect 6469 12869 6503 12903
rect 8401 12869 8435 12903
rect 8585 12869 8619 12903
rect 10609 12869 10643 12903
rect 18245 12869 18279 12903
rect 19993 12869 20027 12903
rect 2145 12801 2179 12835
rect 3617 12801 3651 12835
rect 3801 12801 3835 12835
rect 4629 12801 4663 12835
rect 5181 12801 5215 12835
rect 5273 12801 5307 12835
rect 6837 12801 6871 12835
rect 3525 12733 3559 12767
rect 5089 12733 5123 12767
rect 9505 12801 9539 12835
rect 9597 12801 9631 12835
rect 10149 12801 10183 12835
rect 11069 12801 11103 12835
rect 11253 12801 11287 12835
rect 12449 12801 12483 12835
rect 16957 12801 16991 12835
rect 18889 12801 18923 12835
rect 19073 12801 19107 12835
rect 20729 12801 20763 12835
rect 21741 12801 21775 12835
rect 23673 12801 23707 12835
rect 8861 12733 8895 12767
rect 9413 12733 9447 12767
rect 14657 12733 14691 12767
rect 18797 12733 18831 12767
rect 20085 12733 20119 12767
rect 21649 12733 21683 12767
rect 2053 12665 2087 12699
rect 4261 12665 4295 12699
rect 7082 12665 7116 12699
rect 8401 12665 8435 12699
rect 12265 12665 12299 12699
rect 12716 12665 12750 12699
rect 14565 12665 14599 12699
rect 14924 12665 14958 12699
rect 16313 12665 16347 12699
rect 21005 12665 21039 12699
rect 21557 12665 21591 12699
rect 23918 12665 23952 12699
rect 1961 12597 1995 12631
rect 3065 12597 3099 12631
rect 8217 12597 8251 12631
rect 10517 12597 10551 12631
rect 10977 12597 11011 12631
rect 11713 12597 11747 12631
rect 13829 12597 13863 12631
rect 1685 12393 1719 12427
rect 3157 12393 3191 12427
rect 3525 12393 3559 12427
rect 3893 12393 3927 12427
rect 4261 12393 4295 12427
rect 4997 12393 5031 12427
rect 6377 12393 6411 12427
rect 8309 12393 8343 12427
rect 8677 12393 8711 12427
rect 9689 12393 9723 12427
rect 10149 12393 10183 12427
rect 16681 12393 16715 12427
rect 16957 12393 16991 12427
rect 17325 12393 17359 12427
rect 18521 12393 18555 12427
rect 23397 12393 23431 12427
rect 23765 12393 23799 12427
rect 24133 12393 24167 12427
rect 25329 12393 25363 12427
rect 26065 12393 26099 12427
rect 4721 12325 4755 12359
rect 6806 12325 6840 12359
rect 9505 12325 9539 12359
rect 12633 12325 12667 12359
rect 12725 12325 12759 12359
rect 15568 12325 15602 12359
rect 24685 12325 24719 12359
rect 1777 12257 1811 12291
rect 2033 12257 2067 12291
rect 5365 12257 5399 12291
rect 10057 12257 10091 12291
rect 11529 12257 11563 12291
rect 5457 12189 5491 12223
rect 5549 12189 5583 12223
rect 6561 12189 6595 12223
rect 10241 12189 10275 12223
rect 11621 12189 11655 12223
rect 11713 12189 11747 12223
rect 15301 12257 15335 12291
rect 17509 12257 17543 12291
rect 18981 12257 19015 12291
rect 19441 12257 19475 12291
rect 20729 12257 20763 12291
rect 20913 12257 20947 12291
rect 22284 12257 22318 12291
rect 24593 12257 24627 12291
rect 14473 12189 14507 12223
rect 19073 12189 19107 12223
rect 19257 12189 19291 12223
rect 12633 12121 12667 12155
rect 18613 12121 18647 12155
rect 22017 12189 22051 12223
rect 24777 12189 24811 12223
rect 20269 12121 20303 12155
rect 21097 12121 21131 12155
rect 6101 12053 6135 12087
rect 7941 12053 7975 12087
rect 9137 12053 9171 12087
rect 10701 12053 10735 12087
rect 11161 12053 11195 12087
rect 12541 12053 12575 12087
rect 14933 12053 14967 12087
rect 17693 12053 17727 12087
rect 18061 12053 18095 12087
rect 19441 12053 19475 12087
rect 19717 12053 19751 12087
rect 21649 12053 21683 12087
rect 24225 12053 24259 12087
rect 25605 12053 25639 12087
rect 3801 11849 3835 11883
rect 4353 11849 4387 11883
rect 6193 11849 6227 11883
rect 6561 11849 6595 11883
rect 7573 11849 7607 11883
rect 9781 11849 9815 11883
rect 10241 11849 10275 11883
rect 14657 11849 14691 11883
rect 16405 11849 16439 11883
rect 17509 11849 17543 11883
rect 20269 11849 20303 11883
rect 21833 11849 21867 11883
rect 23489 11849 23523 11883
rect 24501 11849 24535 11883
rect 24685 11849 24719 11883
rect 25421 11849 25455 11883
rect 5089 11781 5123 11815
rect 7849 11781 7883 11815
rect 14565 11781 14599 11815
rect 23673 11781 23707 11815
rect 2145 11713 2179 11747
rect 4721 11713 4755 11747
rect 5733 11713 5767 11747
rect 8033 11713 8067 11747
rect 10793 11713 10827 11747
rect 11621 11713 11655 11747
rect 12449 11713 12483 11747
rect 14197 11713 14231 11747
rect 15209 11713 15243 11747
rect 16957 11713 16991 11747
rect 20729 11713 20763 11747
rect 20821 11713 20855 11747
rect 22477 11713 22511 11747
rect 24133 11713 24167 11747
rect 24317 11713 24351 11747
rect 24501 11713 24535 11747
rect 25145 11713 25179 11747
rect 5641 11645 5675 11679
rect 8289 11645 8323 11679
rect 10149 11645 10183 11679
rect 10701 11645 10735 11679
rect 15117 11645 15151 11679
rect 18061 11645 18095 11679
rect 18317 11645 18351 11679
rect 20177 11645 20211 11679
rect 22937 11645 22971 11679
rect 24041 11645 24075 11679
rect 25237 11645 25271 11679
rect 2053 11577 2087 11611
rect 2412 11577 2446 11611
rect 5549 11577 5583 11611
rect 12716 11577 12750 11611
rect 16865 11577 16899 11611
rect 19717 11577 19751 11611
rect 21373 11577 21407 11611
rect 22293 11577 22327 11611
rect 25789 11577 25823 11611
rect 1685 11509 1719 11543
rect 3525 11509 3559 11543
rect 5181 11509 5215 11543
rect 6837 11509 6871 11543
rect 9413 11509 9447 11543
rect 10609 11509 10643 11543
rect 11253 11509 11287 11543
rect 12173 11509 12207 11543
rect 13829 11509 13863 11543
rect 15025 11509 15059 11543
rect 15945 11509 15979 11543
rect 16313 11509 16347 11543
rect 16773 11509 16807 11543
rect 19441 11509 19475 11543
rect 20637 11509 20671 11543
rect 21649 11509 21683 11543
rect 22201 11509 22235 11543
rect 26249 11509 26283 11543
rect 2973 11305 3007 11339
rect 4629 11305 4663 11339
rect 7297 11305 7331 11339
rect 8125 11305 8159 11339
rect 8493 11305 8527 11339
rect 8585 11305 8619 11339
rect 9413 11305 9447 11339
rect 9689 11305 9723 11339
rect 10701 11305 10735 11339
rect 12817 11305 12851 11339
rect 13645 11305 13679 11339
rect 14105 11305 14139 11339
rect 14657 11305 14691 11339
rect 15117 11305 15151 11339
rect 16681 11305 16715 11339
rect 20913 11305 20947 11339
rect 22017 11305 22051 11339
rect 23029 11305 23063 11339
rect 24961 11305 24995 11339
rect 25237 11305 25271 11339
rect 25973 11305 26007 11339
rect 4988 11237 5022 11271
rect 12081 11237 12115 11271
rect 13277 11237 13311 11271
rect 15568 11237 15602 11271
rect 23826 11237 23860 11271
rect 1593 11169 1627 11203
rect 1860 11169 1894 11203
rect 6377 11169 6411 11203
rect 6745 11169 6779 11203
rect 7389 11169 7423 11203
rect 10057 11169 10091 11203
rect 10149 11169 10183 11203
rect 12173 11169 12207 11203
rect 13185 11169 13219 11203
rect 14013 11169 14047 11203
rect 18236 11169 18270 11203
rect 19993 11169 20027 11203
rect 21281 11169 21315 11203
rect 22293 11169 22327 11203
rect 22477 11169 22511 11203
rect 3249 11101 3283 11135
rect 4721 11101 4755 11135
rect 7481 11101 7515 11135
rect 10241 11101 10275 11135
rect 11253 11101 11287 11135
rect 12265 11101 12299 11135
rect 13369 11101 13403 11135
rect 14197 11101 14231 11135
rect 15301 11101 15335 11135
rect 17969 11101 18003 11135
rect 21373 11101 21407 11135
rect 21465 11101 21499 11135
rect 23581 11101 23615 11135
rect 6929 11033 6963 11067
rect 9045 11033 9079 11067
rect 11713 11033 11747 11067
rect 16957 11033 16991 11067
rect 17417 11033 17451 11067
rect 17785 11033 17819 11067
rect 20269 11033 20303 11067
rect 20729 11033 20763 11067
rect 22661 11033 22695 11067
rect 3709 10965 3743 10999
rect 6101 10965 6135 10999
rect 11529 10965 11563 10999
rect 19349 10965 19383 10999
rect 23489 10965 23523 10999
rect 25605 10965 25639 10999
rect 2237 10761 2271 10795
rect 5917 10761 5951 10795
rect 8309 10761 8343 10795
rect 10333 10761 10367 10795
rect 13737 10761 13771 10795
rect 14105 10761 14139 10795
rect 16313 10761 16347 10795
rect 17509 10761 17543 10795
rect 18245 10761 18279 10795
rect 18981 10761 19015 10795
rect 20913 10761 20947 10795
rect 21189 10761 21223 10795
rect 23489 10761 23523 10795
rect 23673 10761 23707 10795
rect 24685 10761 24719 10795
rect 25973 10761 26007 10795
rect 5181 10693 5215 10727
rect 5549 10693 5583 10727
rect 11805 10693 11839 10727
rect 14841 10693 14875 10727
rect 21557 10693 21591 10727
rect 21741 10693 21775 10727
rect 22753 10693 22787 10727
rect 1777 10625 1811 10659
rect 2789 10625 2823 10659
rect 6653 10625 6687 10659
rect 7481 10625 7515 10659
rect 8953 10625 8987 10659
rect 10609 10625 10643 10659
rect 13001 10625 13035 10659
rect 15301 10625 15335 10659
rect 15485 10625 15519 10659
rect 16865 10625 16899 10659
rect 17049 10625 17083 10659
rect 22385 10625 22419 10659
rect 24225 10625 24259 10659
rect 25421 10625 25455 10659
rect 2605 10557 2639 10591
rect 3801 10557 3835 10591
rect 6285 10557 6319 10591
rect 7205 10557 7239 10591
rect 8585 10557 8619 10591
rect 9220 10557 9254 10591
rect 12265 10557 12299 10591
rect 12909 10557 12943 10591
rect 17785 10557 17819 10591
rect 18429 10557 18463 10591
rect 19533 10557 19567 10591
rect 22109 10557 22143 10591
rect 24041 10557 24075 10591
rect 25237 10557 25271 10591
rect 3709 10489 3743 10523
rect 4068 10489 4102 10523
rect 7297 10489 7331 10523
rect 7941 10489 7975 10523
rect 12817 10489 12851 10523
rect 16773 10489 16807 10523
rect 19778 10489 19812 10523
rect 25053 10489 25087 10523
rect 2145 10421 2179 10455
rect 2697 10421 2731 10455
rect 3249 10421 3283 10455
rect 6837 10421 6871 10455
rect 8401 10421 8435 10455
rect 11161 10421 11195 10455
rect 11345 10421 11379 10455
rect 12449 10421 12483 10455
rect 14381 10421 14415 10455
rect 15209 10421 15243 10455
rect 15853 10421 15887 10455
rect 16405 10421 16439 10455
rect 18613 10421 18647 10455
rect 19349 10421 19383 10455
rect 22201 10421 22235 10455
rect 24133 10421 24167 10455
rect 26341 10421 26375 10455
rect 1685 10217 1719 10251
rect 2329 10217 2363 10251
rect 2789 10217 2823 10251
rect 4629 10217 4663 10251
rect 4997 10217 5031 10251
rect 8309 10217 8343 10251
rect 8401 10217 8435 10251
rect 9505 10217 9539 10251
rect 10057 10217 10091 10251
rect 10149 10217 10183 10251
rect 10885 10217 10919 10251
rect 13645 10217 13679 10251
rect 13921 10217 13955 10251
rect 17233 10217 17267 10251
rect 17785 10217 17819 10251
rect 18245 10217 18279 10251
rect 19165 10217 19199 10251
rect 20913 10217 20947 10251
rect 22477 10217 22511 10251
rect 22845 10217 22879 10251
rect 24869 10217 24903 10251
rect 4537 10149 4571 10183
rect 6438 10149 6472 10183
rect 11713 10149 11747 10183
rect 15577 10149 15611 10183
rect 16589 10149 16623 10183
rect 18153 10149 18187 10183
rect 20729 10149 20763 10183
rect 21281 10149 21315 10183
rect 2881 10081 2915 10115
rect 3433 10081 3467 10115
rect 5089 10081 5123 10115
rect 5733 10081 5767 10115
rect 9045 10081 9079 10115
rect 12164 10081 12198 10115
rect 14105 10081 14139 10115
rect 16681 10081 16715 10115
rect 17141 10081 17175 10115
rect 17601 10081 17635 10115
rect 19533 10081 19567 10115
rect 19717 10081 19751 10115
rect 20361 10081 20395 10115
rect 2973 10013 3007 10047
rect 5273 10013 5307 10047
rect 5549 10013 5583 10047
rect 6193 10013 6227 10047
rect 10241 10013 10275 10047
rect 11897 10013 11931 10047
rect 14933 10013 14967 10047
rect 16129 10013 16163 10047
rect 16865 10013 16899 10047
rect 2421 9945 2455 9979
rect 13277 9945 13311 9979
rect 16221 9945 16255 9979
rect 18429 10013 18463 10047
rect 21373 10013 21407 10047
rect 21557 10013 21591 10047
rect 21925 10013 21959 10047
rect 18797 9945 18831 9979
rect 19901 9945 19935 9979
rect 22385 9945 22419 9979
rect 23756 10149 23790 10183
rect 23305 10013 23339 10047
rect 23489 10013 23523 10047
rect 25145 9945 25179 9979
rect 25513 9945 25547 9979
rect 3893 9877 3927 9911
rect 5549 9877 5583 9911
rect 6009 9877 6043 9911
rect 7573 9877 7607 9911
rect 7941 9877 7975 9911
rect 9689 9877 9723 9911
rect 11437 9877 11471 9911
rect 14289 9877 14323 9911
rect 17141 9877 17175 9911
rect 19349 9877 19383 9911
rect 22845 9877 22879 9911
rect 23029 9877 23063 9911
rect 25881 9877 25915 9911
rect 949 9673 983 9707
rect 4721 9673 4755 9707
rect 6193 9673 6227 9707
rect 14105 9673 14139 9707
rect 18337 9673 18371 9707
rect 21649 9673 21683 9707
rect 22753 9673 22787 9707
rect 23489 9673 23523 9707
rect 25053 9673 25087 9707
rect 1593 9605 1627 9639
rect 4997 9605 5031 9639
rect 8861 9605 8895 9639
rect 9321 9605 9355 9639
rect 9689 9605 9723 9639
rect 10701 9605 10735 9639
rect 14473 9605 14507 9639
rect 14657 9605 14691 9639
rect 16405 9605 16439 9639
rect 17509 9605 17543 9639
rect 17877 9605 17911 9639
rect 18521 9605 18555 9639
rect 20085 9605 20119 9639
rect 5641 9537 5675 9571
rect 5825 9537 5859 9571
rect 9781 9537 9815 9571
rect 11253 9537 11287 9571
rect 11437 9537 11471 9571
rect 12449 9537 12483 9571
rect 15209 9537 15243 9571
rect 16313 9537 16347 9571
rect 17049 9537 17083 9571
rect 18981 9537 19015 9571
rect 19073 9537 19107 9571
rect 20637 9537 20671 9571
rect 21281 9537 21315 9571
rect 22201 9537 22235 9571
rect 23121 9537 23155 9571
rect 1409 9469 1443 9503
rect 2697 9469 2731 9503
rect 6653 9469 6687 9503
rect 7481 9469 7515 9503
rect 10241 9469 10275 9503
rect 15117 9469 15151 9503
rect 19901 9469 19935 9503
rect 20453 9469 20487 9503
rect 2964 9401 2998 9435
rect 7389 9401 7423 9435
rect 7726 9401 7760 9435
rect 11161 9401 11195 9435
rect 12716 9401 12750 9435
rect 15025 9401 15059 9435
rect 16865 9401 16899 9435
rect 18889 9401 18923 9435
rect 23673 9469 23707 9503
rect 23940 9469 23974 9503
rect 21465 9401 21499 9435
rect 25329 9401 25363 9435
rect 25697 9401 25731 9435
rect 26065 9401 26099 9435
rect 2145 9333 2179 9367
rect 2421 9333 2455 9367
rect 4077 9333 4111 9367
rect 5181 9333 5215 9367
rect 5549 9333 5583 9367
rect 10793 9333 10827 9367
rect 11989 9333 12023 9367
rect 13829 9333 13863 9367
rect 15945 9333 15979 9367
rect 16773 9333 16807 9367
rect 19533 9333 19567 9367
rect 20545 9333 20579 9367
rect 21189 9333 21223 9367
rect 21281 9333 21315 9367
rect 22017 9333 22051 9367
rect 22109 9333 22143 9367
rect 1869 9129 1903 9163
rect 2421 9129 2455 9163
rect 4721 9129 4755 9163
rect 6561 9129 6595 9163
rect 9781 9129 9815 9163
rect 10333 9129 10367 9163
rect 12173 9129 12207 9163
rect 12817 9129 12851 9163
rect 14657 9129 14691 9163
rect 15117 9129 15151 9163
rect 15301 9129 15335 9163
rect 15669 9129 15703 9163
rect 16497 9129 16531 9163
rect 16865 9129 16899 9163
rect 17509 9129 17543 9163
rect 18613 9129 18647 9163
rect 18705 9129 18739 9163
rect 20177 9129 20211 9163
rect 24133 9129 24167 9163
rect 24869 9129 24903 9163
rect 25605 9129 25639 9163
rect 25881 9129 25915 9163
rect 26249 9129 26283 9163
rect 2881 9061 2915 9095
rect 5273 9061 5307 9095
rect 7389 9061 7423 9095
rect 9413 9061 9447 9095
rect 10701 9061 10735 9095
rect 11038 9061 11072 9095
rect 13369 9061 13403 9095
rect 22998 9061 23032 9095
rect 2789 8993 2823 9027
rect 5825 8993 5859 9027
rect 7481 8993 7515 9027
rect 13461 8993 13495 9027
rect 14013 8993 14047 9027
rect 19073 8993 19107 9027
rect 19717 8993 19751 9027
rect 20453 8993 20487 9027
rect 21281 8993 21315 9027
rect 24961 8993 24995 9027
rect 1409 8925 1443 8959
rect 2973 8925 3007 8959
rect 3433 8925 3467 8959
rect 5917 8925 5951 8959
rect 6009 8925 6043 8959
rect 7573 8925 7607 8959
rect 8585 8925 8619 8959
rect 10793 8925 10827 8959
rect 12541 8925 12575 8959
rect 13553 8925 13587 8959
rect 15761 8925 15795 8959
rect 15853 8925 15887 8959
rect 17601 8925 17635 8959
rect 17785 8925 17819 8959
rect 18245 8925 18279 8959
rect 19165 8925 19199 8959
rect 19349 8925 19383 8959
rect 21373 8925 21407 8959
rect 21465 8925 21499 8959
rect 22753 8925 22787 8959
rect 2237 8857 2271 8891
rect 3893 8857 3927 8891
rect 5457 8857 5491 8891
rect 7021 8857 7055 8891
rect 8125 8857 8159 8891
rect 4353 8789 4387 8823
rect 6837 8789 6871 8823
rect 8493 8789 8527 8823
rect 9137 8789 9171 8823
rect 13001 8789 13035 8823
rect 17141 8789 17175 8823
rect 20269 8789 20303 8823
rect 20913 8789 20947 8823
rect 22017 8789 22051 8823
rect 22293 8789 22327 8823
rect 24409 8789 24443 8823
rect 25145 8789 25179 8823
rect 5089 8585 5123 8619
rect 6285 8585 6319 8619
rect 6653 8585 6687 8619
rect 7941 8585 7975 8619
rect 8309 8585 8343 8619
rect 9965 8585 9999 8619
rect 13553 8585 13587 8619
rect 16313 8585 16347 8619
rect 17141 8585 17175 8619
rect 17785 8585 17819 8619
rect 19441 8585 19475 8619
rect 22201 8585 22235 8619
rect 22753 8585 22787 8619
rect 23673 8585 23707 8619
rect 24961 8585 24995 8619
rect 26157 8585 26191 8619
rect 6837 8517 6871 8551
rect 10793 8517 10827 8551
rect 14381 8517 14415 8551
rect 17233 8517 17267 8551
rect 20361 8517 20395 8551
rect 5549 8449 5583 8483
rect 5641 8449 5675 8483
rect 7389 8449 7423 8483
rect 9045 8449 9079 8483
rect 11253 8449 11287 8483
rect 11437 8449 11471 8483
rect 11805 8449 11839 8483
rect 13001 8449 13035 8483
rect 23121 8449 23155 8483
rect 24225 8449 24259 8483
rect 2881 8381 2915 8415
rect 4905 8381 4939 8415
rect 5457 8381 5491 8415
rect 7205 8381 7239 8415
rect 8769 8381 8803 8415
rect 9413 8381 9447 8415
rect 10149 8381 10183 8415
rect 10701 8381 10735 8415
rect 12265 8381 12299 8415
rect 12817 8381 12851 8415
rect 14933 8381 14967 8415
rect 15200 8381 15234 8415
rect 17417 8381 17451 8415
rect 18061 8381 18095 8415
rect 20545 8381 20579 8415
rect 20812 8381 20846 8415
rect 24041 8381 24075 8415
rect 25237 8381 25271 8415
rect 25789 8381 25823 8415
rect 1777 8313 1811 8347
rect 1869 8313 1903 8347
rect 3126 8313 3160 8347
rect 4629 8313 4663 8347
rect 7297 8313 7331 8347
rect 9781 8313 9815 8347
rect 12909 8313 12943 8347
rect 13829 8313 13863 8347
rect 14841 8313 14875 8347
rect 16773 8313 16807 8347
rect 18306 8313 18340 8347
rect 23489 8313 23523 8347
rect 2421 8245 2455 8279
rect 4261 8245 4295 8279
rect 8401 8245 8435 8279
rect 8861 8245 8895 8279
rect 11161 8245 11195 8279
rect 12449 8245 12483 8279
rect 19717 8245 19751 8279
rect 21925 8245 21959 8279
rect 24133 8245 24167 8279
rect 25421 8245 25455 8279
rect 2421 8041 2455 8075
rect 4813 8041 4847 8075
rect 6285 8041 6319 8075
rect 7573 8041 7607 8075
rect 8493 8041 8527 8075
rect 9413 8041 9447 8075
rect 10425 8041 10459 8075
rect 10793 8041 10827 8075
rect 13185 8041 13219 8075
rect 14565 8041 14599 8075
rect 15025 8041 15059 8075
rect 16129 8041 16163 8075
rect 16773 8041 16807 8075
rect 18153 8041 18187 8075
rect 19717 8041 19751 8075
rect 20637 8041 20671 8075
rect 21557 8041 21591 8075
rect 23213 8041 23247 8075
rect 24041 8041 24075 8075
rect 25421 8041 25455 8075
rect 25789 8041 25823 8075
rect 26157 8041 26191 8075
rect 2789 7973 2823 8007
rect 4445 7973 4479 8007
rect 8401 7973 8435 8007
rect 11244 7973 11278 8007
rect 13553 7973 13587 8007
rect 16681 7973 16715 8007
rect 17141 7973 17175 8007
rect 22100 7973 22134 8007
rect 24501 7973 24535 8007
rect 25053 7973 25087 8007
rect 2881 7905 2915 7939
rect 5172 7905 5206 7939
rect 6929 7905 6963 7939
rect 7297 7905 7331 7939
rect 9873 7905 9907 7939
rect 10977 7905 11011 7939
rect 15301 7905 15335 7939
rect 17233 7905 17267 7939
rect 18593 7905 18627 7939
rect 24409 7905 24443 7939
rect 3065 7837 3099 7871
rect 4905 7837 4939 7871
rect 8677 7837 8711 7871
rect 13645 7837 13679 7871
rect 13737 7837 13771 7871
rect 15485 7837 15519 7871
rect 17325 7837 17359 7871
rect 18337 7837 18371 7871
rect 21833 7837 21867 7871
rect 23765 7837 23799 7871
rect 24593 7837 24627 7871
rect 7113 7769 7147 7803
rect 10057 7769 10091 7803
rect 14197 7769 14231 7803
rect 1685 7701 1719 7735
rect 2145 7701 2179 7735
rect 3709 7701 3743 7735
rect 8033 7701 8067 7735
rect 9045 7701 9079 7735
rect 12357 7701 12391 7735
rect 12633 7701 12667 7735
rect 13001 7701 13035 7735
rect 19993 7701 20027 7735
rect 21097 7701 21131 7735
rect 2053 7497 2087 7531
rect 7941 7497 7975 7531
rect 9597 7497 9631 7531
rect 9873 7497 9907 7531
rect 10793 7497 10827 7531
rect 11805 7497 11839 7531
rect 12265 7497 12299 7531
rect 12449 7497 12483 7531
rect 16037 7497 16071 7531
rect 16405 7497 16439 7531
rect 20821 7497 20855 7531
rect 22201 7497 22235 7531
rect 23673 7497 23707 7531
rect 25053 7497 25087 7531
rect 26157 7497 26191 7531
rect 6285 7429 6319 7463
rect 13461 7429 13495 7463
rect 20729 7429 20763 7463
rect 2697 7361 2731 7395
rect 4261 7361 4295 7395
rect 5825 7361 5859 7395
rect 7297 7361 7331 7395
rect 7389 7361 7423 7395
rect 8401 7361 8435 7395
rect 8953 7361 8987 7395
rect 9045 7361 9079 7395
rect 10333 7361 10367 7395
rect 11437 7361 11471 7395
rect 12909 7361 12943 7395
rect 13001 7361 13035 7395
rect 18521 7361 18555 7395
rect 21281 7361 21315 7395
rect 21465 7361 21499 7395
rect 21833 7361 21867 7395
rect 24133 7361 24167 7395
rect 24317 7361 24351 7395
rect 24777 7361 24811 7395
rect 1961 7293 1995 7327
rect 2513 7293 2547 7327
rect 3525 7293 3559 7327
rect 4077 7293 4111 7327
rect 5089 7293 5123 7327
rect 5641 7293 5675 7327
rect 8861 7293 8895 7327
rect 11253 7293 11287 7327
rect 12817 7293 12851 7327
rect 14289 7293 14323 7327
rect 16497 7293 16531 7327
rect 18613 7293 18647 7327
rect 18880 7293 18914 7327
rect 22477 7293 22511 7327
rect 23029 7293 23063 7327
rect 25237 7293 25271 7327
rect 25789 7293 25823 7327
rect 4721 7225 4755 7259
rect 5549 7225 5583 7259
rect 6561 7225 6595 7259
rect 7205 7225 7239 7259
rect 10609 7225 10643 7259
rect 11161 7225 11195 7259
rect 14197 7225 14231 7259
rect 14556 7225 14590 7259
rect 16773 7225 16807 7259
rect 17325 7225 17359 7259
rect 17877 7225 17911 7259
rect 24041 7225 24075 7259
rect 2421 7157 2455 7191
rect 3157 7157 3191 7191
rect 3617 7157 3651 7191
rect 3985 7157 4019 7191
rect 5181 7157 5215 7191
rect 6837 7157 6871 7191
rect 8493 7157 8527 7191
rect 15669 7157 15703 7191
rect 19993 7157 20027 7191
rect 20361 7157 20395 7191
rect 21189 7157 21223 7191
rect 22661 7157 22695 7191
rect 23489 7157 23523 7191
rect 25421 7157 25455 7191
rect 1777 6953 1811 6987
rect 3249 6953 3283 6987
rect 3709 6953 3743 6987
rect 4997 6953 5031 6987
rect 9045 6953 9079 6987
rect 10057 6953 10091 6987
rect 11161 6953 11195 6987
rect 11345 6953 11379 6987
rect 11713 6953 11747 6987
rect 14749 6953 14783 6987
rect 15117 6953 15151 6987
rect 15669 6953 15703 6987
rect 16865 6953 16899 6987
rect 17785 6953 17819 6987
rect 23765 6953 23799 6987
rect 25881 6953 25915 6987
rect 26157 6953 26191 6987
rect 8401 6885 8435 6919
rect 13277 6885 13311 6919
rect 14933 6885 14967 6919
rect 19441 6885 19475 6919
rect 2605 6817 2639 6851
rect 4629 6817 4663 6851
rect 5641 6817 5675 6851
rect 6837 6817 6871 6851
rect 6929 6817 6963 6851
rect 10793 6817 10827 6851
rect 11805 6817 11839 6851
rect 13369 6817 13403 6851
rect 14289 6817 14323 6851
rect 14841 6817 14875 6851
rect 2697 6749 2731 6783
rect 2789 6749 2823 6783
rect 5733 6749 5767 6783
rect 5917 6749 5951 6783
rect 6469 6749 6503 6783
rect 8493 6749 8527 6783
rect 8677 6749 8711 6783
rect 9505 6749 9539 6783
rect 10149 6749 10183 6783
rect 10333 6749 10367 6783
rect 11897 6749 11931 6783
rect 12817 6749 12851 6783
rect 13461 6749 13495 6783
rect 2237 6681 2271 6715
rect 7573 6681 7607 6715
rect 7941 6681 7975 6715
rect 2053 6613 2087 6647
rect 5273 6613 5307 6647
rect 7113 6613 7147 6647
rect 8033 6613 8067 6647
rect 9689 6613 9723 6647
rect 12449 6613 12483 6647
rect 12909 6613 12943 6647
rect 14013 6613 14047 6647
rect 14841 6613 14875 6647
rect 15761 6817 15795 6851
rect 17233 6817 17267 6851
rect 17877 6817 17911 6851
rect 21281 6817 21315 6851
rect 22845 6817 22879 6851
rect 24409 6817 24443 6851
rect 24501 6817 24535 6851
rect 15853 6749 15887 6783
rect 18061 6749 18095 6783
rect 19533 6749 19567 6783
rect 19717 6749 19751 6783
rect 21373 6749 21407 6783
rect 21557 6749 21591 6783
rect 22937 6749 22971 6783
rect 23029 6749 23063 6783
rect 24593 6749 24627 6783
rect 15301 6681 15335 6715
rect 19073 6681 19107 6715
rect 22293 6681 22327 6715
rect 22477 6681 22511 6715
rect 24041 6681 24075 6715
rect 25053 6681 25087 6715
rect 14933 6613 14967 6647
rect 16313 6613 16347 6647
rect 17417 6613 17451 6647
rect 18521 6613 18555 6647
rect 18797 6613 18831 6647
rect 20085 6613 20119 6647
rect 20545 6613 20579 6647
rect 20913 6613 20947 6647
rect 21925 6613 21959 6647
rect 25421 6613 25455 6647
rect 1961 6409 1995 6443
rect 4445 6409 4479 6443
rect 6653 6409 6687 6443
rect 9689 6409 9723 6443
rect 11529 6409 11563 6443
rect 11897 6409 11931 6443
rect 13369 6409 13403 6443
rect 13829 6409 13863 6443
rect 16129 6409 16163 6443
rect 17509 6409 17543 6443
rect 19165 6409 19199 6443
rect 21373 6409 21407 6443
rect 21741 6409 21775 6443
rect 23673 6409 23707 6443
rect 26157 6409 26191 6443
rect 2329 6341 2363 6375
rect 2697 6341 2731 6375
rect 11253 6341 11287 6375
rect 15669 6341 15703 6375
rect 18061 6341 18095 6375
rect 24777 6341 24811 6375
rect 5457 6273 5491 6307
rect 5641 6273 5675 6307
rect 8585 6273 8619 6307
rect 8677 6273 8711 6307
rect 16681 6273 16715 6307
rect 18705 6273 18739 6307
rect 22293 6273 22327 6307
rect 22477 6273 22511 6307
rect 24225 6273 24259 6307
rect 25053 6273 25087 6307
rect 2789 6205 2823 6239
rect 5365 6205 5399 6239
rect 7021 6205 7055 6239
rect 8493 6205 8527 6239
rect 9873 6205 9907 6239
rect 12633 6205 12667 6239
rect 13921 6205 13955 6239
rect 14188 6205 14222 6239
rect 16589 6205 16623 6239
rect 19625 6205 19659 6239
rect 24041 6205 24075 6239
rect 25237 6205 25271 6239
rect 25789 6205 25823 6239
rect 3034 6137 3068 6171
rect 9413 6137 9447 6171
rect 10118 6137 10152 6171
rect 12909 6137 12943 6171
rect 18521 6137 18555 6171
rect 19870 6137 19904 6171
rect 22201 6137 22235 6171
rect 23489 6137 23523 6171
rect 24133 6137 24167 6171
rect 4169 6069 4203 6103
rect 4813 6069 4847 6103
rect 4997 6069 5031 6103
rect 6009 6069 6043 6103
rect 7205 6069 7239 6103
rect 7665 6069 7699 6103
rect 7941 6069 7975 6103
rect 8125 6069 8159 6103
rect 15301 6069 15335 6103
rect 15945 6069 15979 6103
rect 16497 6069 16531 6103
rect 17877 6069 17911 6103
rect 18429 6069 18463 6103
rect 19533 6069 19567 6103
rect 21005 6069 21039 6103
rect 21833 6069 21867 6103
rect 22937 6069 22971 6103
rect 25421 6069 25455 6103
rect 1685 5865 1719 5899
rect 3157 5865 3191 5899
rect 4537 5865 4571 5899
rect 6377 5865 6411 5899
rect 6837 5865 6871 5899
rect 7941 5865 7975 5899
rect 11069 5865 11103 5899
rect 11345 5865 11379 5899
rect 14657 5865 14691 5899
rect 15025 5865 15059 5899
rect 16681 5865 16715 5899
rect 17141 5865 17175 5899
rect 17509 5865 17543 5899
rect 19533 5865 19567 5899
rect 20913 5865 20947 5899
rect 21741 5865 21775 5899
rect 23305 5865 23339 5899
rect 23673 5865 23707 5899
rect 24133 5865 24167 5899
rect 24409 5865 24443 5899
rect 25513 5865 25547 5899
rect 7573 5797 7607 5831
rect 9045 5797 9079 5831
rect 9934 5797 9968 5831
rect 11713 5797 11747 5831
rect 12265 5797 12299 5831
rect 14105 5797 14139 5831
rect 15568 5797 15602 5831
rect 18052 5797 18086 5831
rect 20729 5797 20763 5831
rect 25881 5797 25915 5831
rect 26157 5797 26191 5831
rect 1777 5729 1811 5763
rect 2044 5729 2078 5763
rect 3525 5729 3559 5763
rect 3893 5729 3927 5763
rect 4629 5729 4663 5763
rect 4896 5729 4930 5763
rect 6929 5729 6963 5763
rect 8401 5729 8435 5763
rect 9689 5729 9723 5763
rect 12624 5729 12658 5763
rect 15301 5729 15335 5763
rect 17785 5729 17819 5763
rect 21465 5729 21499 5763
rect 22192 5729 22226 5763
rect 24777 5729 24811 5763
rect 8493 5661 8527 5695
rect 8677 5661 8711 5695
rect 12357 5661 12391 5695
rect 21925 5661 21959 5695
rect 24869 5661 24903 5695
rect 24961 5661 24995 5695
rect 7113 5593 7147 5627
rect 8033 5593 8067 5627
rect 19901 5593 19935 5627
rect 6009 5525 6043 5559
rect 9505 5525 9539 5559
rect 13737 5525 13771 5559
rect 19165 5525 19199 5559
rect 20361 5525 20395 5559
rect 2513 5321 2547 5355
rect 4261 5321 4295 5355
rect 4997 5321 5031 5355
rect 7297 5321 7331 5355
rect 11437 5321 11471 5355
rect 12173 5321 12207 5355
rect 13461 5321 13495 5355
rect 15025 5321 15059 5355
rect 16497 5321 16531 5355
rect 16865 5321 16899 5355
rect 17877 5321 17911 5355
rect 20729 5321 20763 5355
rect 22201 5321 22235 5355
rect 23489 5321 23523 5355
rect 26157 5321 26191 5355
rect 1869 5185 1903 5219
rect 22477 5253 22511 5287
rect 4629 5185 4663 5219
rect 5641 5185 5675 5219
rect 10517 5185 10551 5219
rect 14013 5185 14047 5219
rect 14197 5185 14231 5219
rect 15117 5185 15151 5219
rect 24225 5185 24259 5219
rect 24777 5185 24811 5219
rect 2881 5117 2915 5151
rect 5549 5117 5583 5151
rect 7757 5117 7791 5151
rect 10333 5117 10367 5151
rect 12449 5117 12483 5151
rect 18245 5117 18279 5151
rect 20821 5117 20855 5151
rect 21077 5117 21111 5151
rect 24041 5117 24075 5151
rect 25237 5117 25271 5151
rect 25789 5117 25823 5151
rect 3126 5049 3160 5083
rect 7665 5049 7699 5083
rect 8024 5049 8058 5083
rect 13921 5049 13955 5083
rect 14657 5049 14691 5083
rect 15362 5049 15396 5083
rect 17509 5049 17543 5083
rect 18512 5049 18546 5083
rect 24133 5049 24167 5083
rect 25145 5049 25179 5083
rect 1777 4981 1811 5015
rect 2329 4981 2363 5015
rect 2513 4981 2547 5015
rect 2697 4981 2731 5015
rect 5089 4981 5123 5015
rect 5457 4981 5491 5015
rect 6193 4981 6227 5015
rect 6653 4981 6687 5015
rect 9137 4981 9171 5015
rect 9413 4981 9447 5015
rect 9781 4981 9815 5015
rect 9965 4981 9999 5015
rect 10425 4981 10459 5015
rect 10977 4981 11011 5015
rect 11805 4981 11839 5015
rect 12633 4981 12667 5015
rect 13001 4981 13035 5015
rect 13553 4981 13587 5015
rect 19625 4981 19659 5015
rect 19993 4981 20027 5015
rect 20269 4981 20303 5015
rect 23029 4981 23063 5015
rect 23673 4981 23707 5015
rect 25421 4981 25455 5015
rect 1593 4777 1627 4811
rect 2881 4777 2915 4811
rect 7297 4777 7331 4811
rect 7757 4777 7791 4811
rect 8125 4777 8159 4811
rect 9689 4777 9723 4811
rect 10701 4777 10735 4811
rect 13093 4777 13127 4811
rect 14013 4777 14047 4811
rect 15025 4777 15059 4811
rect 15669 4777 15703 4811
rect 17509 4777 17543 4811
rect 19073 4777 19107 4811
rect 19533 4777 19567 4811
rect 20361 4777 20395 4811
rect 20913 4777 20947 4811
rect 21373 4777 21407 4811
rect 22017 4777 22051 4811
rect 22937 4777 22971 4811
rect 24041 4777 24075 4811
rect 24409 4777 24443 4811
rect 25145 4777 25179 4811
rect 26249 4777 26283 4811
rect 1961 4709 1995 4743
rect 3893 4709 3927 4743
rect 4537 4709 4571 4743
rect 11704 4709 11738 4743
rect 15761 4709 15795 4743
rect 17877 4709 17911 4743
rect 22845 4709 22879 4743
rect 2789 4641 2823 4675
rect 3525 4641 3559 4675
rect 4445 4641 4479 4675
rect 5917 4641 5951 4675
rect 6173 4641 6207 4675
rect 8493 4641 8527 4675
rect 9137 4641 9171 4675
rect 10057 4641 10091 4675
rect 11437 4641 11471 4675
rect 16589 4641 16623 4675
rect 19441 4641 19475 4675
rect 21281 4641 21315 4675
rect 24501 4641 24535 4675
rect 25789 4641 25823 4675
rect 3065 4573 3099 4607
rect 4629 4573 4663 4607
rect 10149 4573 10183 4607
rect 10241 4573 10275 4607
rect 13553 4573 13587 4607
rect 14105 4573 14139 4607
rect 14197 4573 14231 4607
rect 15945 4573 15979 4607
rect 17969 4573 18003 4607
rect 18061 4573 18095 4607
rect 18981 4573 19015 4607
rect 19717 4573 19751 4607
rect 20729 4573 20763 4607
rect 21465 4573 21499 4607
rect 23029 4573 23063 4607
rect 24685 4573 24719 4607
rect 2421 4505 2455 4539
rect 4077 4505 4111 4539
rect 8677 4505 8711 4539
rect 13645 4505 13679 4539
rect 14749 4505 14783 4539
rect 15301 4505 15335 4539
rect 17325 4505 17359 4539
rect 5089 4437 5123 4471
rect 5457 4437 5491 4471
rect 9413 4437 9447 4471
rect 11345 4437 11379 4471
rect 12817 4437 12851 4471
rect 17049 4437 17083 4471
rect 18521 4437 18555 4471
rect 22385 4437 22419 4471
rect 22477 4437 22511 4471
rect 23673 4437 23707 4471
rect 25421 4437 25455 4471
rect 2053 4233 2087 4267
rect 4445 4233 4479 4267
rect 9873 4233 9907 4267
rect 11529 4233 11563 4267
rect 13737 4233 13771 4267
rect 17417 4233 17451 4267
rect 22569 4233 22603 4267
rect 24685 4233 24719 4267
rect 25145 4233 25179 4267
rect 2421 4165 2455 4199
rect 9229 4165 9263 4199
rect 10057 4165 10091 4199
rect 15577 4165 15611 4199
rect 15945 4165 15979 4199
rect 16313 4165 16347 4199
rect 21005 4165 21039 4199
rect 3341 4097 3375 4131
rect 3433 4097 3467 4131
rect 5089 4097 5123 4131
rect 5549 4097 5583 4131
rect 6837 4097 6871 4131
rect 10609 4097 10643 4131
rect 13093 4097 13127 4131
rect 16865 4097 16899 4131
rect 16957 4097 16991 4131
rect 18981 4097 19015 4131
rect 19809 4097 19843 4131
rect 20545 4097 20579 4131
rect 21925 4097 21959 4131
rect 22109 4097 22143 4131
rect 22937 4097 22971 4131
rect 24225 4097 24259 4131
rect 2789 4029 2823 4063
rect 3249 4029 3283 4063
rect 7849 4029 7883 4063
rect 10425 4029 10459 4063
rect 11805 4029 11839 4063
rect 12817 4029 12851 4063
rect 14197 4029 14231 4063
rect 18797 4029 18831 4063
rect 20269 4029 20303 4063
rect 20361 4029 20395 4063
rect 24133 4029 24167 4063
rect 25237 4029 25271 4063
rect 25973 4029 26007 4063
rect 26341 4029 26375 4063
rect 3893 3961 3927 3995
rect 4813 3961 4847 3995
rect 5917 3961 5951 3995
rect 8094 3961 8128 3995
rect 9505 3961 9539 3995
rect 10517 3961 10551 3995
rect 11069 3961 11103 3995
rect 14105 3961 14139 3995
rect 14442 3961 14476 3995
rect 19441 3961 19475 3995
rect 21833 3961 21867 3995
rect 24041 3961 24075 3995
rect 25513 3961 25547 3995
rect 1685 3893 1719 3927
rect 2881 3893 2915 3927
rect 4261 3893 4295 3927
rect 4905 3893 4939 3927
rect 6377 3893 6411 3927
rect 7389 3893 7423 3927
rect 7665 3893 7699 3927
rect 12173 3893 12207 3927
rect 12449 3893 12483 3927
rect 12909 3893 12943 3927
rect 16405 3893 16439 3927
rect 16773 3893 16807 3927
rect 17785 3893 17819 3927
rect 18337 3893 18371 3927
rect 18705 3893 18739 3927
rect 19901 3893 19935 3927
rect 21281 3893 21315 3927
rect 21465 3893 21499 3927
rect 23489 3893 23523 3927
rect 23673 3893 23707 3927
rect 1409 3689 1443 3723
rect 2973 3689 3007 3723
rect 3801 3689 3835 3723
rect 4077 3689 4111 3723
rect 4445 3689 4479 3723
rect 5549 3689 5583 3723
rect 7573 3689 7607 3723
rect 8217 3689 8251 3723
rect 9045 3689 9079 3723
rect 9505 3689 9539 3723
rect 10149 3689 10183 3723
rect 12817 3689 12851 3723
rect 13185 3689 13219 3723
rect 14657 3689 14691 3723
rect 15117 3689 15151 3723
rect 19073 3689 19107 3723
rect 19533 3689 19567 3723
rect 20913 3689 20947 3723
rect 21373 3689 21407 3723
rect 22017 3689 22051 3723
rect 22385 3689 22419 3723
rect 22477 3689 22511 3723
rect 25421 3689 25455 3723
rect 25789 3689 25823 3723
rect 26157 3689 26191 3723
rect 1777 3621 1811 3655
rect 5089 3621 5123 3655
rect 6162 3621 6196 3655
rect 8585 3621 8619 3655
rect 11713 3621 11747 3655
rect 13277 3621 13311 3655
rect 15568 3621 15602 3655
rect 17325 3621 17359 3655
rect 18613 3621 18647 3655
rect 20269 3621 20303 3655
rect 22937 3621 22971 3655
rect 24501 3621 24535 3655
rect 1869 3553 1903 3587
rect 4537 3553 4571 3587
rect 5917 3553 5951 3587
rect 8309 3553 8343 3587
rect 10057 3553 10091 3587
rect 10793 3553 10827 3587
rect 11621 3553 11655 3587
rect 15301 3553 15335 3587
rect 17877 3553 17911 3587
rect 19441 3553 19475 3587
rect 21281 3553 21315 3587
rect 22845 3553 22879 3587
rect 24409 3553 24443 3587
rect 2053 3485 2087 3519
rect 3249 3485 3283 3519
rect 4721 3485 4755 3519
rect 10241 3485 10275 3519
rect 11805 3485 11839 3519
rect 13461 3485 13495 3519
rect 13829 3485 13863 3519
rect 16957 3485 16991 3519
rect 17969 3485 18003 3519
rect 18061 3485 18095 3519
rect 19625 3485 19659 3519
rect 20729 3485 20763 3519
rect 21557 3485 21591 3519
rect 23029 3485 23063 3519
rect 24685 3485 24719 3519
rect 2421 3417 2455 3451
rect 7297 3417 7331 3451
rect 9689 3417 9723 3451
rect 11253 3417 11287 3451
rect 12541 3417 12575 3451
rect 17509 3417 17543 3451
rect 18889 3417 18923 3451
rect 25053 3417 25087 3451
rect 11069 3349 11103 3383
rect 14381 3349 14415 3383
rect 16681 3349 16715 3383
rect 23765 3349 23799 3383
rect 24041 3349 24075 3383
rect 1409 3145 1443 3179
rect 2881 3145 2915 3179
rect 3433 3145 3467 3179
rect 5273 3145 5307 3179
rect 5641 3145 5675 3179
rect 6929 3145 6963 3179
rect 9873 3145 9907 3179
rect 12449 3145 12483 3179
rect 14841 3145 14875 3179
rect 15945 3145 15979 3179
rect 18061 3145 18095 3179
rect 19533 3145 19567 3179
rect 20637 3145 20671 3179
rect 21189 3145 21223 3179
rect 25053 3145 25087 3179
rect 26341 3145 26375 3179
rect 2421 3077 2455 3111
rect 8309 3077 8343 3111
rect 10701 3077 10735 3111
rect 11713 3077 11747 3111
rect 19073 3077 19107 3111
rect 19625 3077 19659 3111
rect 1869 3009 1903 3043
rect 2053 3009 2087 3043
rect 6285 3009 6319 3043
rect 7481 3009 7515 3043
rect 10609 3009 10643 3043
rect 11161 3009 11195 3043
rect 11253 3009 11287 3043
rect 13093 3009 13127 3043
rect 14197 3009 14231 3043
rect 15577 3009 15611 3043
rect 16405 3009 16439 3043
rect 16681 3009 16715 3043
rect 18613 3009 18647 3043
rect 20177 3009 20211 3043
rect 21005 3009 21039 3043
rect 21649 3009 21683 3043
rect 21741 3009 21775 3043
rect 22477 3009 22511 3043
rect 24225 3009 24259 3043
rect 24685 3009 24719 3043
rect 1777 2941 1811 2975
rect 3525 2941 3559 2975
rect 3792 2941 3826 2975
rect 7297 2941 7331 2975
rect 8033 2941 8067 2975
rect 8493 2941 8527 2975
rect 8749 2941 8783 2975
rect 10149 2941 10183 2975
rect 12817 2941 12851 2975
rect 12909 2941 12943 2975
rect 13829 2941 13863 2975
rect 15301 2941 15335 2975
rect 15393 2941 15427 2975
rect 16497 2941 16531 2975
rect 18521 2941 18555 2975
rect 20085 2941 20119 2975
rect 21557 2941 21591 2975
rect 24041 2941 24075 2975
rect 25237 2941 25271 2975
rect 25973 2941 26007 2975
rect 5733 2873 5767 2907
rect 6653 2873 6687 2907
rect 7389 2873 7423 2907
rect 12265 2873 12299 2907
rect 23489 2873 23523 2907
rect 24133 2873 24167 2907
rect 25513 2873 25547 2907
rect 4905 2805 4939 2839
rect 11069 2805 11103 2839
rect 13461 2805 13495 2839
rect 14933 2805 14967 2839
rect 17509 2805 17543 2839
rect 18429 2805 18463 2839
rect 19993 2805 20027 2839
rect 23029 2805 23063 2839
rect 23673 2805 23707 2839
rect 1409 2601 1443 2635
rect 3617 2601 3651 2635
rect 6101 2601 6135 2635
rect 7205 2601 7239 2635
rect 8861 2601 8895 2635
rect 9505 2601 9539 2635
rect 11713 2601 11747 2635
rect 14013 2601 14047 2635
rect 16497 2601 16531 2635
rect 18153 2601 18187 2635
rect 18705 2601 18739 2635
rect 19717 2601 19751 2635
rect 21189 2601 21223 2635
rect 21649 2601 21683 2635
rect 22753 2601 22787 2635
rect 24041 2601 24075 2635
rect 25421 2601 25455 2635
rect 26433 2601 26467 2635
rect 1777 2533 1811 2567
rect 2881 2533 2915 2567
rect 5733 2533 5767 2567
rect 9229 2533 9263 2567
rect 11989 2533 12023 2567
rect 14565 2533 14599 2567
rect 20913 2533 20947 2567
rect 21557 2533 21591 2567
rect 26065 2533 26099 2567
rect 1869 2465 1903 2499
rect 2421 2465 2455 2499
rect 4077 2465 4111 2499
rect 4344 2465 4378 2499
rect 7481 2465 7515 2499
rect 7748 2465 7782 2499
rect 10241 2465 10275 2499
rect 10600 2465 10634 2499
rect 12900 2465 12934 2499
rect 15853 2465 15887 2499
rect 17049 2465 17083 2499
rect 18797 2465 18831 2499
rect 19993 2465 20027 2499
rect 20545 2465 20579 2499
rect 22845 2465 22879 2499
rect 24409 2465 24443 2499
rect 2053 2397 2087 2431
rect 2973 2397 3007 2431
rect 6745 2397 6779 2431
rect 10333 2397 10367 2431
rect 12449 2397 12483 2431
rect 12633 2397 12667 2431
rect 14841 2397 14875 2431
rect 15945 2397 15979 2431
rect 16129 2397 16163 2431
rect 16957 2397 16991 2431
rect 18981 2397 19015 2431
rect 21741 2397 21775 2431
rect 22201 2397 22235 2431
rect 23765 2397 23799 2431
rect 24501 2397 24535 2431
rect 24685 2397 24719 2431
rect 25053 2397 25087 2431
rect 25605 2397 25639 2431
rect 15485 2329 15519 2363
rect 5457 2261 5491 2295
rect 15301 2261 15335 2295
rect 17233 2261 17267 2295
rect 17601 2261 17635 2295
rect 18337 2261 18371 2295
rect 20177 2261 20211 2295
rect 23029 2261 23063 2295
rect 23489 2261 23523 2295
<< metal1 >>
rect 3510 27548 3516 27600
rect 3568 27588 3574 27600
rect 9122 27588 9128 27600
rect 3568 27560 9128 27588
rect 3568 27548 3574 27560
rect 9122 27548 9128 27560
rect 9180 27548 9186 27600
rect 12069 26571 12127 26577
rect 12069 26537 12081 26571
rect 12115 26568 12127 26571
rect 17405 26571 17463 26577
rect 17405 26568 17417 26571
rect 12115 26540 17417 26568
rect 12115 26537 12127 26540
rect 12069 26531 12127 26537
rect 17405 26537 17417 26540
rect 17451 26537 17463 26571
rect 17405 26531 17463 26537
rect 12529 26503 12587 26509
rect 12529 26469 12541 26503
rect 12575 26500 12587 26503
rect 17313 26503 17371 26509
rect 17313 26500 17325 26503
rect 12575 26472 17325 26500
rect 12575 26469 12587 26472
rect 12529 26463 12587 26469
rect 17313 26469 17325 26472
rect 17359 26469 17371 26503
rect 17313 26463 17371 26469
rect 13357 26367 13415 26373
rect 13357 26333 13369 26367
rect 13403 26364 13415 26367
rect 16577 26367 16635 26373
rect 16577 26364 16589 26367
rect 13403 26336 16589 26364
rect 13403 26333 13415 26336
rect 13357 26327 13415 26333
rect 16577 26333 16589 26336
rect 16623 26333 16635 26367
rect 16577 26327 16635 26333
rect 11146 26296 11152 26308
rect 10704 26268 11152 26296
rect 3326 26188 3332 26240
rect 3384 26228 3390 26240
rect 10704 26228 10732 26268
rect 11146 26256 11152 26268
rect 11204 26256 11210 26308
rect 13909 26299 13967 26305
rect 13909 26296 13921 26299
rect 12084 26268 13921 26296
rect 3384 26200 10732 26228
rect 3384 26188 3390 26200
rect 10778 26188 10784 26240
rect 10836 26228 10842 26240
rect 12084 26228 12112 26268
rect 13909 26265 13921 26268
rect 13955 26265 13967 26299
rect 13909 26259 13967 26265
rect 14458 26256 14464 26308
rect 14516 26296 14522 26308
rect 16114 26296 16120 26308
rect 14516 26268 16120 26296
rect 14516 26256 14522 26268
rect 16114 26256 16120 26268
rect 16172 26256 16178 26308
rect 10836 26200 12112 26228
rect 10836 26188 10842 26200
rect 12342 26188 12348 26240
rect 12400 26228 12406 26240
rect 19518 26228 19524 26240
rect 12400 26200 19524 26228
rect 12400 26188 12406 26200
rect 19518 26188 19524 26200
rect 19576 26188 19582 26240
rect 5534 26120 5540 26172
rect 5592 26160 5598 26172
rect 12069 26163 12127 26169
rect 12069 26160 12081 26163
rect 5592 26132 12081 26160
rect 5592 26120 5598 26132
rect 12069 26129 12081 26132
rect 12115 26129 12127 26163
rect 12069 26123 12127 26129
rect 12253 26163 12311 26169
rect 12253 26129 12265 26163
rect 12299 26160 12311 26163
rect 12529 26163 12587 26169
rect 12529 26160 12541 26163
rect 12299 26132 12541 26160
rect 12299 26129 12311 26132
rect 12253 26123 12311 26129
rect 12529 26129 12541 26132
rect 12575 26129 12587 26163
rect 12529 26123 12587 26129
rect 16577 26163 16635 26169
rect 16577 26129 16589 26163
rect 16623 26160 16635 26163
rect 18138 26160 18144 26172
rect 16623 26132 18144 26160
rect 16623 26129 16635 26132
rect 16577 26123 16635 26129
rect 18138 26120 18144 26132
rect 18196 26120 18202 26172
rect 6730 26052 6736 26104
rect 6788 26092 6794 26104
rect 11793 26095 11851 26101
rect 11793 26092 11805 26095
rect 6788 26064 11805 26092
rect 6788 26052 6794 26064
rect 11793 26061 11805 26064
rect 11839 26061 11851 26095
rect 11793 26055 11851 26061
rect 11882 26052 11888 26104
rect 11940 26092 11946 26104
rect 13357 26095 13415 26101
rect 13357 26092 13369 26095
rect 11940 26064 13369 26092
rect 11940 26052 11946 26064
rect 13357 26061 13369 26064
rect 13403 26061 13415 26095
rect 13357 26055 13415 26061
rect 13446 26052 13452 26104
rect 13504 26092 13510 26104
rect 18874 26092 18880 26104
rect 13504 26064 18880 26092
rect 13504 26052 13510 26064
rect 18874 26052 18880 26064
rect 18932 26052 18938 26104
rect 9214 25984 9220 26036
rect 9272 26024 9278 26036
rect 16574 26024 16580 26036
rect 9272 25996 16580 26024
rect 9272 25984 9278 25996
rect 16574 25984 16580 25996
rect 16632 25984 16638 26036
rect 4614 25916 4620 25968
rect 4672 25956 4678 25968
rect 11790 25956 11796 25968
rect 4672 25928 11796 25956
rect 4672 25916 4678 25928
rect 11790 25916 11796 25928
rect 11848 25916 11854 25968
rect 11882 25916 11888 25968
rect 11940 25956 11946 25968
rect 25130 25956 25136 25968
rect 11940 25928 25136 25956
rect 11940 25916 11946 25928
rect 25130 25916 25136 25928
rect 25188 25916 25194 25968
rect 9950 25848 9956 25900
rect 10008 25888 10014 25900
rect 12158 25888 12164 25900
rect 10008 25860 12164 25888
rect 10008 25848 10014 25860
rect 12158 25848 12164 25860
rect 12216 25848 12222 25900
rect 13538 25848 13544 25900
rect 13596 25888 13602 25900
rect 21266 25888 21272 25900
rect 13596 25860 21272 25888
rect 13596 25848 13602 25860
rect 21266 25848 21272 25860
rect 21324 25848 21330 25900
rect 8018 25780 8024 25832
rect 8076 25820 8082 25832
rect 17126 25820 17132 25832
rect 8076 25792 17132 25820
rect 8076 25780 8082 25792
rect 17126 25780 17132 25792
rect 17184 25780 17190 25832
rect 17313 25823 17371 25829
rect 17313 25789 17325 25823
rect 17359 25820 17371 25823
rect 19518 25820 19524 25832
rect 17359 25792 19524 25820
rect 17359 25789 17371 25792
rect 17313 25783 17371 25789
rect 19518 25780 19524 25792
rect 19576 25780 19582 25832
rect 8938 25712 8944 25764
rect 8996 25752 9002 25764
rect 13814 25752 13820 25764
rect 8996 25724 13820 25752
rect 8996 25712 9002 25724
rect 13814 25712 13820 25724
rect 13872 25712 13878 25764
rect 13909 25755 13967 25761
rect 13909 25721 13921 25755
rect 13955 25752 13967 25755
rect 17218 25752 17224 25764
rect 13955 25724 17224 25752
rect 13955 25721 13967 25724
rect 13909 25715 13967 25721
rect 17218 25712 17224 25724
rect 17276 25712 17282 25764
rect 17405 25755 17463 25761
rect 17405 25721 17417 25755
rect 17451 25752 17463 25755
rect 19150 25752 19156 25764
rect 17451 25724 19156 25752
rect 17451 25721 17463 25724
rect 17405 25715 17463 25721
rect 19150 25712 19156 25724
rect 19208 25712 19214 25764
rect 10686 25644 10692 25696
rect 10744 25684 10750 25696
rect 18322 25684 18328 25696
rect 10744 25656 18328 25684
rect 10744 25644 10750 25656
rect 18322 25644 18328 25656
rect 18380 25644 18386 25696
rect 21910 25644 21916 25696
rect 21968 25684 21974 25696
rect 26510 25684 26516 25696
rect 21968 25656 26516 25684
rect 21968 25644 21974 25656
rect 26510 25644 26516 25656
rect 26568 25644 26574 25696
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 2222 25440 2228 25492
rect 2280 25480 2286 25492
rect 10505 25483 10563 25489
rect 2280 25452 7604 25480
rect 2280 25440 2286 25452
rect 7576 25412 7604 25452
rect 10505 25449 10517 25483
rect 10551 25480 10563 25483
rect 10686 25480 10692 25492
rect 10551 25452 10692 25480
rect 10551 25449 10563 25452
rect 10505 25443 10563 25449
rect 10686 25440 10692 25452
rect 10744 25440 10750 25492
rect 11609 25483 11667 25489
rect 11609 25449 11621 25483
rect 11655 25480 11667 25483
rect 12250 25480 12256 25492
rect 11655 25452 12256 25480
rect 11655 25449 11667 25452
rect 11609 25443 11667 25449
rect 12250 25440 12256 25452
rect 12308 25440 12314 25492
rect 12342 25440 12348 25492
rect 12400 25480 12406 25492
rect 13722 25480 13728 25492
rect 12400 25452 13728 25480
rect 12400 25440 12406 25452
rect 13722 25440 13728 25452
rect 13780 25440 13786 25492
rect 13814 25440 13820 25492
rect 13872 25480 13878 25492
rect 13909 25483 13967 25489
rect 13909 25480 13921 25483
rect 13872 25452 13921 25480
rect 13872 25440 13878 25452
rect 13909 25449 13921 25452
rect 13955 25449 13967 25483
rect 13909 25443 13967 25449
rect 7576 25384 13860 25412
rect 10321 25347 10379 25353
rect 10321 25313 10333 25347
rect 10367 25344 10379 25347
rect 10870 25344 10876 25356
rect 10367 25316 10876 25344
rect 10367 25313 10379 25316
rect 10321 25307 10379 25313
rect 10870 25304 10876 25316
rect 10928 25304 10934 25356
rect 11425 25347 11483 25353
rect 11425 25313 11437 25347
rect 11471 25344 11483 25347
rect 11606 25344 11612 25356
rect 11471 25316 11612 25344
rect 11471 25313 11483 25316
rect 11425 25307 11483 25313
rect 11606 25304 11612 25316
rect 11664 25304 11670 25356
rect 12710 25304 12716 25356
rect 12768 25344 12774 25356
rect 12805 25347 12863 25353
rect 12805 25344 12817 25347
rect 12768 25316 12817 25344
rect 12768 25304 12774 25316
rect 12805 25313 12817 25316
rect 12851 25344 12863 25347
rect 13541 25347 13599 25353
rect 13541 25344 13553 25347
rect 12851 25316 13553 25344
rect 12851 25313 12863 25316
rect 12805 25307 12863 25313
rect 13541 25313 13553 25316
rect 13587 25313 13599 25347
rect 13541 25307 13599 25313
rect 9858 25236 9864 25288
rect 9916 25276 9922 25288
rect 12989 25279 13047 25285
rect 12989 25276 13001 25279
rect 9916 25248 13001 25276
rect 9916 25236 9922 25248
rect 12989 25245 13001 25248
rect 13035 25245 13047 25279
rect 13832 25276 13860 25384
rect 13924 25344 13952 25443
rect 14090 25440 14096 25492
rect 14148 25480 14154 25492
rect 15197 25483 15255 25489
rect 15197 25480 15209 25483
rect 14148 25452 15209 25480
rect 14148 25440 14154 25452
rect 15197 25449 15209 25452
rect 15243 25449 15255 25483
rect 15197 25443 15255 25449
rect 15473 25483 15531 25489
rect 15473 25449 15485 25483
rect 15519 25449 15531 25483
rect 15473 25443 15531 25449
rect 15933 25483 15991 25489
rect 15933 25449 15945 25483
rect 15979 25480 15991 25483
rect 16206 25480 16212 25492
rect 15979 25452 16212 25480
rect 15979 25449 15991 25452
rect 15933 25443 15991 25449
rect 15488 25412 15516 25443
rect 16206 25440 16212 25452
rect 16264 25440 16270 25492
rect 16393 25483 16451 25489
rect 16393 25449 16405 25483
rect 16439 25480 16451 25483
rect 16853 25483 16911 25489
rect 16853 25480 16865 25483
rect 16439 25452 16865 25480
rect 16439 25449 16451 25452
rect 16393 25443 16451 25449
rect 16853 25449 16865 25452
rect 16899 25480 16911 25483
rect 17037 25483 17095 25489
rect 17037 25480 17049 25483
rect 16899 25452 17049 25480
rect 16899 25449 16911 25452
rect 16853 25443 16911 25449
rect 17037 25449 17049 25452
rect 17083 25449 17095 25483
rect 17037 25443 17095 25449
rect 17313 25483 17371 25489
rect 17313 25449 17325 25483
rect 17359 25449 17371 25483
rect 17313 25443 17371 25449
rect 17497 25483 17555 25489
rect 17497 25449 17509 25483
rect 17543 25480 17555 25483
rect 21358 25480 21364 25492
rect 17543 25452 21364 25480
rect 17543 25449 17555 25452
rect 17497 25443 17555 25449
rect 16574 25412 16580 25424
rect 15488 25384 16580 25412
rect 16574 25372 16580 25384
rect 16632 25372 16638 25424
rect 17328 25412 17356 25443
rect 21358 25440 21364 25452
rect 21416 25440 21422 25492
rect 21910 25480 21916 25492
rect 21871 25452 21916 25480
rect 21910 25440 21916 25452
rect 21968 25440 21974 25492
rect 22922 25440 22928 25492
rect 22980 25480 22986 25492
rect 25866 25480 25872 25492
rect 22980 25452 25872 25480
rect 22980 25440 22986 25452
rect 25866 25440 25872 25452
rect 25924 25440 25930 25492
rect 23014 25412 23020 25424
rect 17328 25384 23020 25412
rect 23014 25372 23020 25384
rect 23072 25372 23078 25424
rect 24762 25412 24768 25424
rect 23124 25384 24768 25412
rect 14093 25347 14151 25353
rect 14093 25344 14105 25347
rect 13924 25316 14105 25344
rect 14093 25313 14105 25316
rect 14139 25313 14151 25347
rect 15286 25344 15292 25356
rect 14093 25307 14151 25313
rect 14200 25316 15292 25344
rect 14200 25276 14228 25316
rect 15286 25304 15292 25316
rect 15344 25304 15350 25356
rect 15841 25347 15899 25353
rect 15841 25313 15853 25347
rect 15887 25344 15899 25347
rect 16114 25344 16120 25356
rect 15887 25316 16120 25344
rect 15887 25313 15899 25316
rect 15841 25307 15899 25313
rect 16114 25304 16120 25316
rect 16172 25304 16178 25356
rect 16298 25304 16304 25356
rect 16356 25344 16362 25356
rect 17129 25347 17187 25353
rect 16356 25316 16620 25344
rect 16356 25304 16362 25316
rect 14366 25276 14372 25288
rect 13832 25248 14228 25276
rect 14327 25248 14372 25276
rect 12989 25239 13047 25245
rect 14366 25236 14372 25248
rect 14424 25236 14430 25288
rect 14642 25236 14648 25288
rect 14700 25276 14706 25288
rect 16025 25279 16083 25285
rect 16025 25276 16037 25279
rect 14700 25248 16037 25276
rect 14700 25236 14706 25248
rect 16025 25245 16037 25248
rect 16071 25276 16083 25279
rect 16482 25276 16488 25288
rect 16071 25248 16488 25276
rect 16071 25245 16083 25248
rect 16025 25239 16083 25245
rect 16482 25236 16488 25248
rect 16540 25236 16546 25288
rect 16592 25276 16620 25316
rect 17129 25313 17141 25347
rect 17175 25344 17187 25347
rect 17310 25344 17316 25356
rect 17175 25316 17316 25344
rect 17175 25313 17187 25316
rect 17129 25307 17187 25313
rect 17310 25304 17316 25316
rect 17368 25304 17374 25356
rect 18877 25347 18935 25353
rect 18877 25313 18889 25347
rect 18923 25344 18935 25347
rect 19058 25344 19064 25356
rect 18923 25316 19064 25344
rect 18923 25313 18935 25316
rect 18877 25307 18935 25313
rect 19058 25304 19064 25316
rect 19116 25304 19122 25356
rect 19978 25344 19984 25356
rect 19939 25316 19984 25344
rect 19978 25304 19984 25316
rect 20036 25304 20042 25356
rect 21729 25347 21787 25353
rect 21729 25313 21741 25347
rect 21775 25344 21787 25347
rect 22002 25344 22008 25356
rect 21775 25316 22008 25344
rect 21775 25313 21787 25316
rect 21729 25307 21787 25313
rect 22002 25304 22008 25316
rect 22060 25304 22066 25356
rect 22738 25304 22744 25356
rect 22796 25344 22802 25356
rect 22833 25347 22891 25353
rect 22833 25344 22845 25347
rect 22796 25316 22845 25344
rect 22796 25304 22802 25316
rect 22833 25313 22845 25316
rect 22879 25313 22891 25347
rect 23124 25344 23152 25384
rect 24762 25372 24768 25384
rect 24820 25372 24826 25424
rect 22833 25307 22891 25313
rect 22940 25316 23152 25344
rect 17497 25279 17555 25285
rect 17497 25276 17509 25279
rect 16592 25248 17509 25276
rect 17497 25245 17509 25248
rect 17543 25245 17555 25279
rect 22940 25276 22968 25316
rect 24026 25304 24032 25356
rect 24084 25344 24090 25356
rect 24489 25347 24547 25353
rect 24489 25344 24501 25347
rect 24084 25316 24501 25344
rect 24084 25304 24090 25316
rect 24489 25313 24501 25316
rect 24535 25313 24547 25347
rect 24489 25307 24547 25313
rect 24581 25347 24639 25353
rect 24581 25313 24593 25347
rect 24627 25344 24639 25347
rect 24627 25316 24808 25344
rect 24627 25313 24639 25316
rect 24581 25307 24639 25313
rect 24780 25288 24808 25316
rect 17497 25239 17555 25245
rect 19076 25248 22968 25276
rect 10229 25211 10287 25217
rect 10229 25177 10241 25211
rect 10275 25208 10287 25211
rect 11241 25211 11299 25217
rect 11241 25208 11253 25211
rect 10275 25180 11253 25208
rect 10275 25177 10287 25180
rect 10229 25171 10287 25177
rect 11241 25177 11253 25180
rect 11287 25208 11299 25211
rect 11977 25211 12035 25217
rect 11977 25208 11989 25211
rect 11287 25180 11989 25208
rect 11287 25177 11299 25180
rect 11241 25171 11299 25177
rect 11977 25177 11989 25180
rect 12023 25208 12035 25211
rect 14550 25208 14556 25220
rect 12023 25180 14556 25208
rect 12023 25177 12035 25180
rect 11977 25171 12035 25177
rect 14550 25168 14556 25180
rect 14608 25208 14614 25220
rect 14608 25180 15240 25208
rect 14608 25168 14614 25180
rect 8846 25100 8852 25152
rect 8904 25140 8910 25152
rect 9401 25143 9459 25149
rect 9401 25140 9413 25143
rect 8904 25112 9413 25140
rect 8904 25100 8910 25112
rect 9401 25109 9413 25112
rect 9447 25140 9459 25143
rect 10873 25143 10931 25149
rect 10873 25140 10885 25143
rect 9447 25112 10885 25140
rect 9447 25109 9459 25112
rect 9401 25103 9459 25109
rect 10873 25109 10885 25112
rect 10919 25109 10931 25143
rect 10873 25103 10931 25109
rect 12437 25143 12495 25149
rect 12437 25109 12449 25143
rect 12483 25140 12495 25143
rect 13354 25140 13360 25152
rect 12483 25112 13360 25140
rect 12483 25109 12495 25112
rect 12437 25103 12495 25109
rect 13354 25100 13360 25112
rect 13412 25100 13418 25152
rect 14734 25100 14740 25152
rect 14792 25140 14798 25152
rect 14829 25143 14887 25149
rect 14829 25140 14841 25143
rect 14792 25112 14841 25140
rect 14792 25100 14798 25112
rect 14829 25109 14841 25112
rect 14875 25109 14887 25143
rect 15212 25140 15240 25180
rect 15286 25168 15292 25220
rect 15344 25208 15350 25220
rect 18414 25208 18420 25220
rect 15344 25180 18420 25208
rect 15344 25168 15350 25180
rect 18414 25168 18420 25180
rect 18472 25168 18478 25220
rect 19076 25217 19104 25248
rect 23842 25236 23848 25288
rect 23900 25276 23906 25288
rect 24673 25279 24731 25285
rect 24673 25276 24685 25279
rect 23900 25248 24685 25276
rect 23900 25236 23906 25248
rect 24673 25245 24685 25248
rect 24719 25245 24731 25279
rect 24673 25239 24731 25245
rect 24762 25236 24768 25288
rect 24820 25236 24826 25288
rect 19061 25211 19119 25217
rect 19061 25177 19073 25211
rect 19107 25177 19119 25211
rect 19061 25171 19119 25177
rect 20165 25211 20223 25217
rect 20165 25177 20177 25211
rect 20211 25208 20223 25211
rect 22922 25208 22928 25220
rect 20211 25180 22928 25208
rect 20211 25177 20223 25180
rect 20165 25171 20223 25177
rect 22922 25168 22928 25180
rect 22980 25168 22986 25220
rect 23017 25211 23075 25217
rect 23017 25177 23029 25211
rect 23063 25208 23075 25211
rect 27062 25208 27068 25220
rect 23063 25180 27068 25208
rect 23063 25177 23075 25180
rect 23017 25171 23075 25177
rect 27062 25168 27068 25180
rect 27120 25168 27126 25220
rect 16393 25143 16451 25149
rect 16393 25140 16405 25143
rect 15212 25112 16405 25140
rect 14829 25103 14887 25109
rect 16393 25109 16405 25112
rect 16439 25109 16451 25143
rect 16393 25103 16451 25109
rect 16577 25143 16635 25149
rect 16577 25109 16589 25143
rect 16623 25140 16635 25143
rect 16758 25140 16764 25152
rect 16623 25112 16764 25140
rect 16623 25109 16635 25112
rect 16577 25103 16635 25109
rect 16758 25100 16764 25112
rect 16816 25100 16822 25152
rect 17037 25143 17095 25149
rect 17037 25109 17049 25143
rect 17083 25140 17095 25143
rect 17681 25143 17739 25149
rect 17681 25140 17693 25143
rect 17083 25112 17693 25140
rect 17083 25109 17095 25112
rect 17037 25103 17095 25109
rect 17681 25109 17693 25112
rect 17727 25109 17739 25143
rect 17681 25103 17739 25109
rect 17862 25100 17868 25152
rect 17920 25140 17926 25152
rect 23290 25140 23296 25152
rect 17920 25112 23296 25140
rect 17920 25100 17926 25112
rect 23290 25100 23296 25112
rect 23348 25100 23354 25152
rect 23842 25140 23848 25152
rect 23803 25112 23848 25140
rect 23842 25100 23848 25112
rect 23900 25100 23906 25152
rect 24121 25143 24179 25149
rect 24121 25109 24133 25143
rect 24167 25140 24179 25143
rect 24210 25140 24216 25152
rect 24167 25112 24216 25140
rect 24167 25109 24179 25112
rect 24121 25103 24179 25109
rect 24210 25100 24216 25112
rect 24268 25100 24274 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1578 24936 1584 24948
rect 1539 24908 1584 24936
rect 1578 24896 1584 24908
rect 1636 24896 1642 24948
rect 9214 24936 9220 24948
rect 9175 24908 9220 24936
rect 9214 24896 9220 24908
rect 9272 24896 9278 24948
rect 9306 24896 9312 24948
rect 9364 24936 9370 24948
rect 14366 24936 14372 24948
rect 9364 24908 14372 24936
rect 9364 24896 9370 24908
rect 14366 24896 14372 24908
rect 14424 24896 14430 24948
rect 14642 24936 14648 24948
rect 14603 24908 14648 24936
rect 14642 24896 14648 24908
rect 14700 24896 14706 24948
rect 14734 24896 14740 24948
rect 14792 24936 14798 24948
rect 14792 24908 15148 24936
rect 14792 24896 14798 24908
rect 15120 24880 15148 24908
rect 15286 24896 15292 24948
rect 15344 24936 15350 24948
rect 20349 24939 20407 24945
rect 15344 24908 20300 24936
rect 15344 24896 15350 24908
rect 9677 24871 9735 24877
rect 9677 24837 9689 24871
rect 9723 24868 9735 24871
rect 9858 24868 9864 24880
rect 9723 24840 9864 24868
rect 9723 24837 9735 24840
rect 9677 24831 9735 24837
rect 1397 24735 1455 24741
rect 1397 24701 1409 24735
rect 1443 24732 1455 24735
rect 9033 24735 9091 24741
rect 1443 24704 2084 24732
rect 1443 24701 1455 24704
rect 1397 24695 1455 24701
rect 2056 24605 2084 24704
rect 9033 24701 9045 24735
rect 9079 24732 9091 24735
rect 9692 24732 9720 24831
rect 9858 24828 9864 24840
rect 9916 24828 9922 24880
rect 10321 24871 10379 24877
rect 10321 24837 10333 24871
rect 10367 24868 10379 24871
rect 13446 24868 13452 24880
rect 10367 24840 13452 24868
rect 10367 24837 10379 24840
rect 10321 24831 10379 24837
rect 13446 24828 13452 24840
rect 13504 24828 13510 24880
rect 13722 24828 13728 24880
rect 13780 24868 13786 24880
rect 13780 24840 15056 24868
rect 13780 24828 13786 24840
rect 12253 24803 12311 24809
rect 12253 24769 12265 24803
rect 12299 24800 12311 24803
rect 13633 24803 13691 24809
rect 13633 24800 13645 24803
rect 12299 24772 13645 24800
rect 12299 24769 12311 24772
rect 12253 24763 12311 24769
rect 13633 24769 13645 24772
rect 13679 24800 13691 24803
rect 13998 24800 14004 24812
rect 13679 24772 14004 24800
rect 13679 24769 13691 24772
rect 13633 24763 13691 24769
rect 13998 24760 14004 24772
rect 14056 24760 14062 24812
rect 14274 24760 14280 24812
rect 14332 24800 14338 24812
rect 14826 24800 14832 24812
rect 14332 24772 14832 24800
rect 14332 24760 14338 24772
rect 14826 24760 14832 24772
rect 14884 24760 14890 24812
rect 15028 24800 15056 24840
rect 15102 24828 15108 24880
rect 15160 24828 15166 24880
rect 20272 24868 20300 24908
rect 20349 24905 20361 24939
rect 20395 24936 20407 24939
rect 24670 24936 24676 24948
rect 20395 24908 24676 24936
rect 20395 24905 20407 24908
rect 20349 24899 20407 24905
rect 24670 24896 24676 24908
rect 24728 24896 24734 24948
rect 25590 24936 25596 24948
rect 25551 24908 25596 24936
rect 25590 24896 25596 24908
rect 25648 24896 25654 24948
rect 20714 24868 20720 24880
rect 15212 24840 18552 24868
rect 20272 24840 20720 24868
rect 15212 24800 15240 24840
rect 15028 24772 15240 24800
rect 15381 24803 15439 24809
rect 15381 24769 15393 24803
rect 15427 24800 15439 24803
rect 15470 24800 15476 24812
rect 15427 24772 15476 24800
rect 15427 24769 15439 24772
rect 15381 24763 15439 24769
rect 15470 24760 15476 24772
rect 15528 24800 15534 24812
rect 16390 24800 16396 24812
rect 15528 24772 16396 24800
rect 15528 24760 15534 24772
rect 16390 24760 16396 24772
rect 16448 24800 16454 24812
rect 18524 24809 18552 24840
rect 20714 24828 20720 24840
rect 20772 24828 20778 24880
rect 22649 24871 22707 24877
rect 22649 24837 22661 24871
rect 22695 24837 22707 24871
rect 22649 24831 22707 24837
rect 16853 24803 16911 24809
rect 16853 24800 16865 24803
rect 16448 24772 16865 24800
rect 16448 24760 16454 24772
rect 16853 24769 16865 24772
rect 16899 24769 16911 24803
rect 16853 24763 16911 24769
rect 18509 24803 18567 24809
rect 18509 24769 18521 24803
rect 18555 24769 18567 24803
rect 22664 24800 22692 24831
rect 23842 24828 23848 24880
rect 23900 24868 23906 24880
rect 23900 24840 24532 24868
rect 23900 24828 23906 24840
rect 23382 24800 23388 24812
rect 22664 24772 23388 24800
rect 18509 24763 18567 24769
rect 23382 24760 23388 24772
rect 23440 24760 23446 24812
rect 24504 24809 24532 24840
rect 24489 24803 24547 24809
rect 24489 24769 24501 24803
rect 24535 24800 24547 24803
rect 25041 24803 25099 24809
rect 25041 24800 25053 24803
rect 24535 24772 25053 24800
rect 24535 24769 24547 24772
rect 24489 24763 24547 24769
rect 25041 24769 25053 24772
rect 25087 24769 25099 24803
rect 25041 24763 25099 24769
rect 10137 24735 10195 24741
rect 10137 24732 10149 24735
rect 9079 24704 9720 24732
rect 10060 24704 10149 24732
rect 9079 24701 9091 24704
rect 9033 24695 9091 24701
rect 10060 24608 10088 24704
rect 10137 24701 10149 24704
rect 10183 24701 10195 24735
rect 10137 24695 10195 24701
rect 11241 24735 11299 24741
rect 11241 24701 11253 24735
rect 11287 24701 11299 24735
rect 11241 24695 11299 24701
rect 11256 24608 11284 24695
rect 14458 24692 14464 24744
rect 14516 24732 14522 24744
rect 16298 24732 16304 24744
rect 14516 24704 16304 24732
rect 14516 24692 14522 24704
rect 16298 24692 16304 24704
rect 16356 24692 16362 24744
rect 16574 24692 16580 24744
rect 16632 24732 16638 24744
rect 17586 24732 17592 24744
rect 16632 24704 17592 24732
rect 16632 24692 16638 24704
rect 17586 24692 17592 24704
rect 17644 24692 17650 24744
rect 18325 24735 18383 24741
rect 18325 24732 18337 24735
rect 17788 24704 18337 24732
rect 12897 24667 12955 24673
rect 12897 24633 12909 24667
rect 12943 24664 12955 24667
rect 13170 24664 13176 24676
rect 12943 24636 13176 24664
rect 12943 24633 12955 24636
rect 12897 24627 12955 24633
rect 13170 24624 13176 24636
rect 13228 24664 13234 24676
rect 13449 24667 13507 24673
rect 13449 24664 13461 24667
rect 13228 24636 13461 24664
rect 13228 24624 13234 24636
rect 13449 24633 13461 24636
rect 13495 24633 13507 24667
rect 13449 24627 13507 24633
rect 14277 24667 14335 24673
rect 14277 24633 14289 24667
rect 14323 24664 14335 24667
rect 14826 24664 14832 24676
rect 14323 24636 14832 24664
rect 14323 24633 14335 24636
rect 14277 24627 14335 24633
rect 14826 24624 14832 24636
rect 14884 24664 14890 24676
rect 15197 24667 15255 24673
rect 15197 24664 15209 24667
rect 14884 24636 15209 24664
rect 14884 24624 14890 24636
rect 15197 24633 15209 24636
rect 15243 24633 15255 24667
rect 15197 24627 15255 24633
rect 15841 24667 15899 24673
rect 15841 24633 15853 24667
rect 15887 24664 15899 24667
rect 16206 24664 16212 24676
rect 15887 24636 16212 24664
rect 15887 24633 15899 24636
rect 15841 24627 15899 24633
rect 16206 24624 16212 24636
rect 16264 24624 16270 24676
rect 16666 24664 16672 24676
rect 16627 24636 16672 24664
rect 16666 24624 16672 24636
rect 16724 24624 16730 24676
rect 17788 24608 17816 24704
rect 18325 24701 18337 24704
rect 18371 24701 18383 24735
rect 20162 24732 20168 24744
rect 20075 24704 20168 24732
rect 18325 24695 18383 24701
rect 20162 24692 20168 24704
rect 20220 24732 20226 24744
rect 20717 24735 20775 24741
rect 20717 24732 20729 24735
rect 20220 24704 20729 24732
rect 20220 24692 20226 24704
rect 20717 24701 20729 24704
rect 20763 24701 20775 24735
rect 21269 24735 21327 24741
rect 21269 24732 21281 24735
rect 20717 24695 20775 24701
rect 21100 24704 21281 24732
rect 21100 24608 21128 24704
rect 21269 24701 21281 24704
rect 21315 24701 21327 24735
rect 21269 24695 21327 24701
rect 22465 24735 22523 24741
rect 22465 24701 22477 24735
rect 22511 24732 22523 24735
rect 24213 24735 24271 24741
rect 24213 24732 24225 24735
rect 22511 24704 22876 24732
rect 22511 24701 22523 24704
rect 22465 24695 22523 24701
rect 22848 24608 22876 24704
rect 23492 24704 24225 24732
rect 23492 24608 23520 24704
rect 24213 24701 24225 24704
rect 24259 24701 24271 24735
rect 25409 24735 25467 24741
rect 25409 24732 25421 24735
rect 24213 24695 24271 24701
rect 24872 24704 25421 24732
rect 24118 24624 24124 24676
rect 24176 24664 24182 24676
rect 24305 24667 24363 24673
rect 24305 24664 24317 24667
rect 24176 24636 24317 24664
rect 24176 24624 24182 24636
rect 24305 24633 24317 24636
rect 24351 24633 24363 24667
rect 24305 24627 24363 24633
rect 24872 24608 24900 24704
rect 25409 24701 25421 24704
rect 25455 24732 25467 24735
rect 25961 24735 26019 24741
rect 25961 24732 25973 24735
rect 25455 24704 25973 24732
rect 25455 24701 25467 24704
rect 25409 24695 25467 24701
rect 25961 24701 25973 24704
rect 26007 24701 26019 24735
rect 25961 24695 26019 24701
rect 2041 24599 2099 24605
rect 2041 24565 2053 24599
rect 2087 24596 2099 24599
rect 2222 24596 2228 24608
rect 2087 24568 2228 24596
rect 2087 24565 2099 24568
rect 2041 24559 2099 24565
rect 2222 24556 2228 24568
rect 2280 24556 2286 24608
rect 8665 24599 8723 24605
rect 8665 24565 8677 24599
rect 8711 24596 8723 24599
rect 8846 24596 8852 24608
rect 8711 24568 8852 24596
rect 8711 24565 8723 24568
rect 8665 24559 8723 24565
rect 8846 24556 8852 24568
rect 8904 24556 8910 24608
rect 10042 24596 10048 24608
rect 10003 24568 10048 24596
rect 10042 24556 10048 24568
rect 10100 24556 10106 24608
rect 10781 24599 10839 24605
rect 10781 24565 10793 24599
rect 10827 24596 10839 24599
rect 10870 24596 10876 24608
rect 10827 24568 10876 24596
rect 10827 24565 10839 24568
rect 10781 24559 10839 24565
rect 10870 24556 10876 24568
rect 10928 24556 10934 24608
rect 11149 24599 11207 24605
rect 11149 24565 11161 24599
rect 11195 24596 11207 24599
rect 11238 24596 11244 24608
rect 11195 24568 11244 24596
rect 11195 24565 11207 24568
rect 11149 24559 11207 24565
rect 11238 24556 11244 24568
rect 11296 24556 11302 24608
rect 11422 24596 11428 24608
rect 11383 24568 11428 24596
rect 11422 24556 11428 24568
rect 11480 24556 11486 24608
rect 11606 24556 11612 24608
rect 11664 24596 11670 24608
rect 11885 24599 11943 24605
rect 11885 24596 11897 24599
rect 11664 24568 11897 24596
rect 11664 24556 11670 24568
rect 11885 24565 11897 24568
rect 11931 24596 11943 24599
rect 12250 24596 12256 24608
rect 11931 24568 12256 24596
rect 11931 24565 11943 24568
rect 11885 24559 11943 24565
rect 12250 24556 12256 24568
rect 12308 24556 12314 24608
rect 12986 24596 12992 24608
rect 12947 24568 12992 24596
rect 12986 24556 12992 24568
rect 13044 24556 13050 24608
rect 13354 24596 13360 24608
rect 13315 24568 13360 24596
rect 13354 24556 13360 24568
rect 13412 24556 13418 24608
rect 14737 24599 14795 24605
rect 14737 24565 14749 24599
rect 14783 24596 14795 24599
rect 14918 24596 14924 24608
rect 14783 24568 14924 24596
rect 14783 24565 14795 24568
rect 14737 24559 14795 24565
rect 14918 24556 14924 24568
rect 14976 24556 14982 24608
rect 15102 24596 15108 24608
rect 15063 24568 15108 24596
rect 15102 24556 15108 24568
rect 15160 24556 15166 24608
rect 16114 24596 16120 24608
rect 16075 24568 16120 24596
rect 16114 24556 16120 24568
rect 16172 24556 16178 24608
rect 16298 24596 16304 24608
rect 16259 24568 16304 24596
rect 16298 24556 16304 24568
rect 16356 24556 16362 24608
rect 16758 24596 16764 24608
rect 16719 24568 16764 24596
rect 16758 24556 16764 24568
rect 16816 24556 16822 24608
rect 17310 24596 17316 24608
rect 17271 24568 17316 24596
rect 17310 24556 17316 24568
rect 17368 24556 17374 24608
rect 17770 24596 17776 24608
rect 17731 24568 17776 24596
rect 17770 24556 17776 24568
rect 17828 24556 17834 24608
rect 19058 24596 19064 24608
rect 19019 24568 19064 24596
rect 19058 24556 19064 24568
rect 19116 24556 19122 24608
rect 19978 24596 19984 24608
rect 19939 24568 19984 24596
rect 19978 24556 19984 24568
rect 20036 24556 20042 24608
rect 21082 24596 21088 24608
rect 21043 24568 21088 24596
rect 21082 24556 21088 24568
rect 21140 24556 21146 24608
rect 21453 24599 21511 24605
rect 21453 24565 21465 24599
rect 21499 24596 21511 24599
rect 21726 24596 21732 24608
rect 21499 24568 21732 24596
rect 21499 24565 21511 24568
rect 21453 24559 21511 24565
rect 21726 24556 21732 24568
rect 21784 24556 21790 24608
rect 21913 24599 21971 24605
rect 21913 24565 21925 24599
rect 21959 24596 21971 24599
rect 22002 24596 22008 24608
rect 21959 24568 22008 24596
rect 21959 24565 21971 24568
rect 21913 24559 21971 24565
rect 22002 24556 22008 24568
rect 22060 24556 22066 24608
rect 22830 24556 22836 24608
rect 22888 24596 22894 24608
rect 23017 24599 23075 24605
rect 23017 24596 23029 24599
rect 22888 24568 23029 24596
rect 22888 24556 22894 24568
rect 23017 24565 23029 24568
rect 23063 24565 23075 24599
rect 23474 24596 23480 24608
rect 23435 24568 23480 24596
rect 23017 24559 23075 24565
rect 23474 24556 23480 24568
rect 23532 24556 23538 24608
rect 23750 24556 23756 24608
rect 23808 24596 23814 24608
rect 23845 24599 23903 24605
rect 23845 24596 23857 24599
rect 23808 24568 23857 24596
rect 23808 24556 23814 24568
rect 23845 24565 23857 24568
rect 23891 24565 23903 24599
rect 24854 24596 24860 24608
rect 24815 24568 24860 24596
rect 23845 24559 23903 24565
rect 24854 24556 24860 24568
rect 24912 24556 24918 24608
rect 25041 24599 25099 24605
rect 25041 24565 25053 24599
rect 25087 24596 25099 24599
rect 25314 24596 25320 24608
rect 25087 24568 25320 24596
rect 25087 24565 25099 24568
rect 25041 24559 25099 24565
rect 25314 24556 25320 24568
rect 25372 24556 25378 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1486 24352 1492 24404
rect 1544 24392 1550 24404
rect 1581 24395 1639 24401
rect 1581 24392 1593 24395
rect 1544 24364 1593 24392
rect 1544 24352 1550 24364
rect 1581 24361 1593 24364
rect 1627 24361 1639 24395
rect 1581 24355 1639 24361
rect 7561 24395 7619 24401
rect 7561 24361 7573 24395
rect 7607 24392 7619 24395
rect 7926 24392 7932 24404
rect 7607 24364 7932 24392
rect 7607 24361 7619 24364
rect 7561 24355 7619 24361
rect 7926 24352 7932 24364
rect 7984 24352 7990 24404
rect 8662 24392 8668 24404
rect 8623 24364 8668 24392
rect 8662 24352 8668 24364
rect 8720 24352 8726 24404
rect 11333 24395 11391 24401
rect 11333 24361 11345 24395
rect 11379 24392 11391 24395
rect 11514 24392 11520 24404
rect 11379 24364 11520 24392
rect 11379 24361 11391 24364
rect 11333 24355 11391 24361
rect 11514 24352 11520 24364
rect 11572 24352 11578 24404
rect 13446 24392 13452 24404
rect 13407 24364 13452 24392
rect 13446 24352 13452 24364
rect 13504 24352 13510 24404
rect 13814 24392 13820 24404
rect 13727 24364 13820 24392
rect 13814 24352 13820 24364
rect 13872 24392 13878 24404
rect 14090 24392 14096 24404
rect 13872 24364 14096 24392
rect 13872 24352 13878 24364
rect 14090 24352 14096 24364
rect 14148 24352 14154 24404
rect 14829 24395 14887 24401
rect 14829 24361 14841 24395
rect 14875 24392 14887 24395
rect 15470 24392 15476 24404
rect 14875 24364 15476 24392
rect 14875 24361 14887 24364
rect 14829 24355 14887 24361
rect 15470 24352 15476 24364
rect 15528 24352 15534 24404
rect 15562 24352 15568 24404
rect 15620 24392 15626 24404
rect 15749 24395 15807 24401
rect 15749 24392 15761 24395
rect 15620 24364 15761 24392
rect 15620 24352 15626 24364
rect 15749 24361 15761 24364
rect 15795 24392 15807 24395
rect 15838 24392 15844 24404
rect 15795 24364 15844 24392
rect 15795 24361 15807 24364
rect 15749 24355 15807 24361
rect 15838 24352 15844 24364
rect 15896 24352 15902 24404
rect 16850 24392 16856 24404
rect 16811 24364 16856 24392
rect 16850 24352 16856 24364
rect 16908 24352 16914 24404
rect 18046 24392 18052 24404
rect 18007 24364 18052 24392
rect 18046 24352 18052 24364
rect 18104 24392 18110 24404
rect 18506 24392 18512 24404
rect 18104 24364 18512 24392
rect 18104 24352 18110 24364
rect 18506 24352 18512 24364
rect 18564 24352 18570 24404
rect 19150 24352 19156 24404
rect 19208 24392 19214 24404
rect 19334 24392 19340 24404
rect 19208 24364 19340 24392
rect 19208 24352 19214 24364
rect 19334 24352 19340 24364
rect 19392 24392 19398 24404
rect 21358 24392 21364 24404
rect 19392 24364 20760 24392
rect 21319 24364 21364 24392
rect 19392 24352 19398 24364
rect 15286 24324 15292 24336
rect 10244 24296 15292 24324
rect 10244 24268 10272 24296
rect 15286 24284 15292 24296
rect 15344 24284 15350 24336
rect 17313 24327 17371 24333
rect 17313 24324 17325 24327
rect 15672 24296 17325 24324
rect 1397 24259 1455 24265
rect 1397 24225 1409 24259
rect 1443 24256 1455 24259
rect 2038 24256 2044 24268
rect 1443 24228 2044 24256
rect 1443 24225 1455 24228
rect 1397 24219 1455 24225
rect 2038 24216 2044 24228
rect 2096 24216 2102 24268
rect 7377 24259 7435 24265
rect 7377 24225 7389 24259
rect 7423 24256 7435 24259
rect 7558 24256 7564 24268
rect 7423 24228 7564 24256
rect 7423 24225 7435 24228
rect 7377 24219 7435 24225
rect 7558 24216 7564 24228
rect 7616 24216 7622 24268
rect 8294 24216 8300 24268
rect 8352 24256 8358 24268
rect 8481 24259 8539 24265
rect 8481 24256 8493 24259
rect 8352 24228 8493 24256
rect 8352 24216 8358 24228
rect 8481 24225 8493 24228
rect 8527 24225 8539 24259
rect 10226 24256 10232 24268
rect 10139 24228 10232 24256
rect 8481 24219 8539 24225
rect 10226 24216 10232 24228
rect 10284 24216 10290 24268
rect 11606 24216 11612 24268
rect 11664 24256 11670 24268
rect 11701 24259 11759 24265
rect 11701 24256 11713 24259
rect 11664 24228 11713 24256
rect 11664 24216 11670 24228
rect 11701 24225 11713 24228
rect 11747 24225 11759 24259
rect 11701 24219 11759 24225
rect 11793 24259 11851 24265
rect 11793 24225 11805 24259
rect 11839 24256 11851 24259
rect 12342 24256 12348 24268
rect 11839 24228 12348 24256
rect 11839 24225 11851 24228
rect 11793 24219 11851 24225
rect 12342 24216 12348 24228
rect 12400 24216 12406 24268
rect 14642 24216 14648 24268
rect 14700 24256 14706 24268
rect 15672 24265 15700 24296
rect 17313 24293 17325 24296
rect 17359 24324 17371 24327
rect 17402 24324 17408 24336
rect 17359 24296 17408 24324
rect 17359 24293 17371 24296
rect 17313 24287 17371 24293
rect 17402 24284 17408 24296
rect 17460 24284 17466 24336
rect 20732 24324 20760 24364
rect 21358 24352 21364 24364
rect 21416 24352 21422 24404
rect 21174 24324 21180 24336
rect 20732 24296 21180 24324
rect 21174 24284 21180 24296
rect 21232 24324 21238 24336
rect 21453 24327 21511 24333
rect 21453 24324 21465 24327
rect 21232 24296 21465 24324
rect 21232 24284 21238 24296
rect 21453 24293 21465 24296
rect 21499 24293 21511 24327
rect 21453 24287 21511 24293
rect 15657 24259 15715 24265
rect 15657 24256 15669 24259
rect 14700 24228 15669 24256
rect 14700 24216 14706 24228
rect 15657 24225 15669 24228
rect 15703 24225 15715 24259
rect 15657 24219 15715 24225
rect 16942 24216 16948 24268
rect 17000 24256 17006 24268
rect 17221 24259 17279 24265
rect 17221 24256 17233 24259
rect 17000 24228 17233 24256
rect 17000 24216 17006 24228
rect 17221 24225 17233 24228
rect 17267 24225 17279 24259
rect 17221 24219 17279 24225
rect 18877 24259 18935 24265
rect 18877 24225 18889 24259
rect 18923 24256 18935 24259
rect 19150 24256 19156 24268
rect 18923 24228 19156 24256
rect 18923 24225 18935 24228
rect 18877 24219 18935 24225
rect 19150 24216 19156 24228
rect 19208 24216 19214 24268
rect 22189 24259 22247 24265
rect 22189 24225 22201 24259
rect 22235 24256 22247 24259
rect 23477 24259 23535 24265
rect 23477 24256 23489 24259
rect 22235 24228 23489 24256
rect 22235 24225 22247 24228
rect 22189 24219 22247 24225
rect 23477 24225 23489 24228
rect 23523 24256 23535 24259
rect 23842 24256 23848 24268
rect 23523 24228 23848 24256
rect 23523 24225 23535 24228
rect 23477 24219 23535 24225
rect 23842 24216 23848 24228
rect 23900 24216 23906 24268
rect 25038 24256 25044 24268
rect 24999 24228 25044 24256
rect 25038 24216 25044 24228
rect 25096 24216 25102 24268
rect 11885 24191 11943 24197
rect 11885 24157 11897 24191
rect 11931 24157 11943 24191
rect 13906 24188 13912 24200
rect 13867 24160 13912 24188
rect 11885 24151 11943 24157
rect 10410 24120 10416 24132
rect 10371 24092 10416 24120
rect 10410 24080 10416 24092
rect 10468 24080 10474 24132
rect 11241 24123 11299 24129
rect 11241 24089 11253 24123
rect 11287 24120 11299 24123
rect 11698 24120 11704 24132
rect 11287 24092 11704 24120
rect 11287 24089 11299 24092
rect 11241 24083 11299 24089
rect 11698 24080 11704 24092
rect 11756 24080 11762 24132
rect 11790 24080 11796 24132
rect 11848 24120 11854 24132
rect 11900 24120 11928 24151
rect 13906 24148 13912 24160
rect 13964 24148 13970 24200
rect 14090 24188 14096 24200
rect 14051 24160 14096 24188
rect 14090 24148 14096 24160
rect 14148 24148 14154 24200
rect 15286 24148 15292 24200
rect 15344 24148 15350 24200
rect 15841 24191 15899 24197
rect 15841 24157 15853 24191
rect 15887 24157 15899 24191
rect 15841 24151 15899 24157
rect 11848 24092 11928 24120
rect 15304 24120 15332 24148
rect 15856 24120 15884 24151
rect 16482 24148 16488 24200
rect 16540 24188 16546 24200
rect 17405 24191 17463 24197
rect 17405 24188 17417 24191
rect 16540 24160 17417 24188
rect 16540 24148 16546 24160
rect 17405 24157 17417 24160
rect 17451 24188 17463 24191
rect 18417 24191 18475 24197
rect 18417 24188 18429 24191
rect 17451 24160 18429 24188
rect 17451 24157 17463 24160
rect 17405 24151 17463 24157
rect 18417 24157 18429 24160
rect 18463 24188 18475 24191
rect 18598 24188 18604 24200
rect 18463 24160 18604 24188
rect 18463 24157 18475 24160
rect 18417 24151 18475 24157
rect 18598 24148 18604 24160
rect 18656 24148 18662 24200
rect 19058 24188 19064 24200
rect 19019 24160 19064 24188
rect 19058 24148 19064 24160
rect 19116 24148 19122 24200
rect 21542 24188 21548 24200
rect 21503 24160 21548 24188
rect 21542 24148 21548 24160
rect 21600 24148 21606 24200
rect 22557 24191 22615 24197
rect 22557 24157 22569 24191
rect 22603 24188 22615 24191
rect 23106 24188 23112 24200
rect 22603 24160 23112 24188
rect 22603 24157 22615 24160
rect 22557 24151 22615 24157
rect 23106 24148 23112 24160
rect 23164 24188 23170 24200
rect 23569 24191 23627 24197
rect 23569 24188 23581 24191
rect 23164 24160 23581 24188
rect 23164 24148 23170 24160
rect 23569 24157 23581 24160
rect 23615 24157 23627 24191
rect 23569 24151 23627 24157
rect 23661 24191 23719 24197
rect 23661 24157 23673 24191
rect 23707 24157 23719 24191
rect 23661 24151 23719 24157
rect 15304 24092 15884 24120
rect 11848 24080 11854 24092
rect 15764 24064 15792 24092
rect 23474 24080 23480 24132
rect 23532 24120 23538 24132
rect 23676 24120 23704 24151
rect 24946 24148 24952 24200
rect 25004 24188 25010 24200
rect 25133 24191 25191 24197
rect 25133 24188 25145 24191
rect 25004 24160 25145 24188
rect 25004 24148 25010 24160
rect 25133 24157 25145 24160
rect 25179 24157 25191 24191
rect 25133 24151 25191 24157
rect 25225 24191 25283 24197
rect 25225 24157 25237 24191
rect 25271 24188 25283 24191
rect 25314 24188 25320 24200
rect 25271 24160 25320 24188
rect 25271 24157 25283 24160
rect 25225 24151 25283 24157
rect 24026 24120 24032 24132
rect 23532 24092 23704 24120
rect 23939 24092 24032 24120
rect 23532 24080 23538 24092
rect 8389 24055 8447 24061
rect 8389 24021 8401 24055
rect 8435 24052 8447 24055
rect 8846 24052 8852 24064
rect 8435 24024 8852 24052
rect 8435 24021 8447 24024
rect 8389 24015 8447 24021
rect 8846 24012 8852 24024
rect 8904 24052 8910 24064
rect 9033 24055 9091 24061
rect 9033 24052 9045 24055
rect 8904 24024 9045 24052
rect 8904 24012 8910 24024
rect 9033 24021 9045 24024
rect 9079 24052 9091 24055
rect 9401 24055 9459 24061
rect 9401 24052 9413 24055
rect 9079 24024 9413 24052
rect 9079 24021 9091 24024
rect 9033 24015 9091 24021
rect 9401 24021 9413 24024
rect 9447 24052 9459 24055
rect 9861 24055 9919 24061
rect 9861 24052 9873 24055
rect 9447 24024 9873 24052
rect 9447 24021 9459 24024
rect 9401 24015 9459 24021
rect 9861 24021 9873 24024
rect 9907 24021 9919 24055
rect 10778 24052 10784 24064
rect 10739 24024 10784 24052
rect 9861 24015 9919 24021
rect 10778 24012 10784 24024
rect 10836 24012 10842 24064
rect 12713 24055 12771 24061
rect 12713 24021 12725 24055
rect 12759 24052 12771 24055
rect 12802 24052 12808 24064
rect 12759 24024 12808 24052
rect 12759 24021 12771 24024
rect 12713 24015 12771 24021
rect 12802 24012 12808 24024
rect 12860 24012 12866 24064
rect 13081 24055 13139 24061
rect 13081 24021 13093 24055
rect 13127 24052 13139 24055
rect 13354 24052 13360 24064
rect 13127 24024 13360 24052
rect 13127 24021 13139 24024
rect 13081 24015 13139 24021
rect 13354 24012 13360 24024
rect 13412 24012 13418 24064
rect 15289 24055 15347 24061
rect 15289 24021 15301 24055
rect 15335 24052 15347 24055
rect 15654 24052 15660 24064
rect 15335 24024 15660 24052
rect 15335 24021 15347 24024
rect 15289 24015 15347 24021
rect 15654 24012 15660 24024
rect 15712 24012 15718 24064
rect 15746 24012 15752 24064
rect 15804 24012 15810 24064
rect 16022 24012 16028 24064
rect 16080 24052 16086 24064
rect 16301 24055 16359 24061
rect 16301 24052 16313 24055
rect 16080 24024 16313 24052
rect 16080 24012 16086 24024
rect 16301 24021 16313 24024
rect 16347 24052 16359 24055
rect 16390 24052 16396 24064
rect 16347 24024 16396 24052
rect 16347 24021 16359 24024
rect 16301 24015 16359 24021
rect 16390 24012 16396 24024
rect 16448 24012 16454 24064
rect 16666 24012 16672 24064
rect 16724 24052 16730 24064
rect 16761 24055 16819 24061
rect 16761 24052 16773 24055
rect 16724 24024 16773 24052
rect 16724 24012 16730 24024
rect 16761 24021 16773 24024
rect 16807 24052 16819 24055
rect 16850 24052 16856 24064
rect 16807 24024 16856 24052
rect 16807 24021 16819 24024
rect 16761 24015 16819 24021
rect 16850 24012 16856 24024
rect 16908 24012 16914 24064
rect 19610 24052 19616 24064
rect 19571 24024 19616 24052
rect 19610 24012 19616 24024
rect 19668 24012 19674 24064
rect 20993 24055 21051 24061
rect 20993 24021 21005 24055
rect 21039 24052 21051 24055
rect 22554 24052 22560 24064
rect 21039 24024 22560 24052
rect 21039 24021 21051 24024
rect 20993 24015 21051 24021
rect 22554 24012 22560 24024
rect 22612 24012 22618 24064
rect 22738 24012 22744 24064
rect 22796 24052 22802 24064
rect 22833 24055 22891 24061
rect 22833 24052 22845 24055
rect 22796 24024 22845 24052
rect 22796 24012 22802 24024
rect 22833 24021 22845 24024
rect 22879 24021 22891 24055
rect 22833 24015 22891 24021
rect 23109 24055 23167 24061
rect 23109 24021 23121 24055
rect 23155 24052 23167 24055
rect 23290 24052 23296 24064
rect 23155 24024 23296 24052
rect 23155 24021 23167 24024
rect 23109 24015 23167 24021
rect 23290 24012 23296 24024
rect 23348 24012 23354 24064
rect 23566 24012 23572 24064
rect 23624 24052 23630 24064
rect 23952 24052 23980 24092
rect 24026 24080 24032 24092
rect 24084 24120 24090 24132
rect 24489 24123 24547 24129
rect 24489 24120 24501 24123
rect 24084 24092 24501 24120
rect 24084 24080 24090 24092
rect 24489 24089 24501 24092
rect 24535 24089 24547 24123
rect 24489 24083 24547 24089
rect 24854 24080 24860 24132
rect 24912 24120 24918 24132
rect 25240 24120 25268 24151
rect 25314 24148 25320 24160
rect 25372 24148 25378 24200
rect 24912 24092 25268 24120
rect 24912 24080 24918 24092
rect 24118 24052 24124 24064
rect 23624 24024 23980 24052
rect 24079 24024 24124 24052
rect 23624 24012 23630 24024
rect 24118 24012 24124 24024
rect 24176 24012 24182 24064
rect 24670 24052 24676 24064
rect 24631 24024 24676 24052
rect 24670 24012 24676 24024
rect 24728 24012 24734 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1581 23851 1639 23857
rect 1581 23817 1593 23851
rect 1627 23848 1639 23851
rect 1670 23848 1676 23860
rect 1627 23820 1676 23848
rect 1627 23817 1639 23820
rect 1581 23811 1639 23817
rect 1670 23808 1676 23820
rect 1728 23808 1734 23860
rect 2682 23848 2688 23860
rect 2643 23820 2688 23848
rect 2682 23808 2688 23820
rect 2740 23808 2746 23860
rect 8018 23848 8024 23860
rect 7979 23820 8024 23848
rect 8018 23808 8024 23820
rect 8076 23808 8082 23860
rect 9122 23848 9128 23860
rect 9083 23820 9128 23848
rect 9122 23808 9128 23820
rect 9180 23808 9186 23860
rect 9490 23848 9496 23860
rect 9451 23820 9496 23848
rect 9490 23808 9496 23820
rect 9548 23808 9554 23860
rect 10226 23848 10232 23860
rect 10187 23820 10232 23848
rect 10226 23808 10232 23820
rect 10284 23808 10290 23860
rect 10686 23808 10692 23860
rect 10744 23848 10750 23860
rect 10781 23851 10839 23857
rect 10781 23848 10793 23851
rect 10744 23820 10793 23848
rect 10744 23808 10750 23820
rect 10781 23817 10793 23820
rect 10827 23817 10839 23851
rect 10781 23811 10839 23817
rect 13265 23851 13323 23857
rect 13265 23817 13277 23851
rect 13311 23848 13323 23851
rect 13814 23848 13820 23860
rect 13311 23820 13820 23848
rect 13311 23817 13323 23820
rect 13265 23811 13323 23817
rect 13814 23808 13820 23820
rect 13872 23808 13878 23860
rect 15197 23851 15255 23857
rect 15197 23817 15209 23851
rect 15243 23848 15255 23851
rect 15470 23848 15476 23860
rect 15243 23820 15476 23848
rect 15243 23817 15255 23820
rect 15197 23811 15255 23817
rect 15470 23808 15476 23820
rect 15528 23808 15534 23860
rect 15838 23808 15844 23860
rect 15896 23848 15902 23860
rect 16209 23851 16267 23857
rect 16209 23848 16221 23851
rect 15896 23820 16221 23848
rect 15896 23808 15902 23820
rect 16209 23817 16221 23820
rect 16255 23817 16267 23851
rect 16209 23811 16267 23817
rect 16758 23808 16764 23860
rect 16816 23848 16822 23860
rect 18049 23851 18107 23857
rect 18049 23848 18061 23851
rect 16816 23820 18061 23848
rect 16816 23808 16822 23820
rect 18049 23817 18061 23820
rect 18095 23817 18107 23851
rect 20346 23848 20352 23860
rect 20307 23820 20352 23848
rect 18049 23811 18107 23817
rect 20346 23808 20352 23820
rect 20404 23808 20410 23860
rect 20714 23848 20720 23860
rect 20675 23820 20720 23848
rect 20714 23808 20720 23820
rect 20772 23848 20778 23860
rect 20772 23820 21404 23848
rect 20772 23808 20778 23820
rect 7282 23740 7288 23792
rect 7340 23780 7346 23792
rect 7834 23780 7840 23792
rect 7340 23752 7840 23780
rect 7340 23740 7346 23752
rect 7834 23740 7840 23752
rect 7892 23740 7898 23792
rect 8481 23783 8539 23789
rect 8481 23749 8493 23783
rect 8527 23780 8539 23783
rect 9306 23780 9312 23792
rect 8527 23752 9312 23780
rect 8527 23749 8539 23752
rect 8481 23743 8539 23749
rect 1397 23647 1455 23653
rect 1397 23613 1409 23647
rect 1443 23644 1455 23647
rect 1670 23644 1676 23656
rect 1443 23616 1676 23644
rect 1443 23613 1455 23616
rect 1397 23607 1455 23613
rect 1670 23604 1676 23616
rect 1728 23604 1734 23656
rect 2314 23604 2320 23656
rect 2372 23644 2378 23656
rect 2501 23647 2559 23653
rect 2501 23644 2513 23647
rect 2372 23616 2513 23644
rect 2372 23604 2378 23616
rect 2501 23613 2513 23616
rect 2547 23644 2559 23647
rect 3053 23647 3111 23653
rect 3053 23644 3065 23647
rect 2547 23616 3065 23644
rect 2547 23613 2559 23616
rect 2501 23607 2559 23613
rect 3053 23613 3065 23616
rect 3099 23613 3111 23647
rect 3053 23607 3111 23613
rect 7837 23647 7895 23653
rect 7837 23613 7849 23647
rect 7883 23644 7895 23647
rect 8496 23644 8524 23743
rect 9306 23740 9312 23752
rect 9364 23740 9370 23792
rect 17034 23780 17040 23792
rect 14844 23752 16712 23780
rect 16995 23752 17040 23780
rect 11425 23715 11483 23721
rect 11425 23681 11437 23715
rect 11471 23712 11483 23715
rect 11698 23712 11704 23724
rect 11471 23684 11704 23712
rect 11471 23681 11483 23684
rect 11425 23675 11483 23681
rect 11698 23672 11704 23684
rect 11756 23672 11762 23724
rect 12805 23715 12863 23721
rect 12805 23681 12817 23715
rect 12851 23712 12863 23715
rect 13722 23712 13728 23724
rect 12851 23684 13728 23712
rect 12851 23681 12863 23684
rect 12805 23675 12863 23681
rect 13722 23672 13728 23684
rect 13780 23712 13786 23724
rect 13817 23715 13875 23721
rect 13817 23712 13829 23715
rect 13780 23684 13829 23712
rect 13780 23672 13786 23684
rect 13817 23681 13829 23684
rect 13863 23681 13875 23715
rect 14844 23712 14872 23752
rect 13817 23675 13875 23681
rect 14292 23684 14872 23712
rect 7883 23616 8524 23644
rect 8941 23647 8999 23653
rect 7883 23613 7895 23616
rect 7837 23607 7895 23613
rect 8941 23613 8953 23647
rect 8987 23644 8999 23647
rect 9490 23644 9496 23656
rect 8987 23616 9496 23644
rect 8987 23613 8999 23616
rect 8941 23607 8999 23613
rect 9490 23604 9496 23616
rect 9548 23604 9554 23656
rect 10778 23604 10784 23656
rect 10836 23644 10842 23656
rect 11149 23647 11207 23653
rect 11149 23644 11161 23647
rect 10836 23616 11161 23644
rect 10836 23604 10842 23616
rect 11149 23613 11161 23616
rect 11195 23613 11207 23647
rect 11149 23607 11207 23613
rect 13538 23604 13544 23656
rect 13596 23644 13602 23656
rect 13633 23647 13691 23653
rect 13633 23644 13645 23647
rect 13596 23616 13645 23644
rect 13596 23604 13602 23616
rect 13633 23613 13645 23616
rect 13679 23613 13691 23647
rect 13633 23607 13691 23613
rect 8294 23536 8300 23588
rect 8352 23576 8358 23588
rect 8757 23579 8815 23585
rect 8757 23576 8769 23579
rect 8352 23548 8769 23576
rect 8352 23536 8358 23548
rect 8757 23545 8769 23548
rect 8803 23545 8815 23579
rect 8757 23539 8815 23545
rect 10689 23579 10747 23585
rect 10689 23545 10701 23579
rect 10735 23576 10747 23579
rect 11241 23579 11299 23585
rect 11241 23576 11253 23579
rect 10735 23548 11253 23576
rect 10735 23545 10747 23548
rect 10689 23539 10747 23545
rect 11241 23545 11253 23548
rect 11287 23576 11299 23579
rect 11974 23576 11980 23588
rect 11287 23548 11980 23576
rect 11287 23545 11299 23548
rect 11241 23539 11299 23545
rect 11974 23536 11980 23548
rect 12032 23536 12038 23588
rect 13173 23579 13231 23585
rect 13173 23545 13185 23579
rect 13219 23576 13231 23579
rect 14090 23576 14096 23588
rect 13219 23548 14096 23576
rect 13219 23545 13231 23548
rect 13173 23539 13231 23545
rect 14090 23536 14096 23548
rect 14148 23536 14154 23588
rect 2038 23508 2044 23520
rect 1999 23480 2044 23508
rect 2038 23468 2044 23480
rect 2096 23468 2102 23520
rect 4430 23468 4436 23520
rect 4488 23508 4494 23520
rect 4890 23508 4896 23520
rect 4488 23480 4896 23508
rect 4488 23468 4494 23480
rect 4890 23468 4896 23480
rect 4948 23468 4954 23520
rect 7469 23511 7527 23517
rect 7469 23477 7481 23511
rect 7515 23508 7527 23511
rect 7558 23508 7564 23520
rect 7515 23480 7564 23508
rect 7515 23477 7527 23480
rect 7469 23471 7527 23477
rect 7558 23468 7564 23480
rect 7616 23468 7622 23520
rect 8938 23468 8944 23520
rect 8996 23508 9002 23520
rect 9861 23511 9919 23517
rect 9861 23508 9873 23511
rect 8996 23480 9873 23508
rect 8996 23468 9002 23480
rect 9861 23477 9873 23480
rect 9907 23477 9919 23511
rect 9861 23471 9919 23477
rect 11606 23468 11612 23520
rect 11664 23508 11670 23520
rect 11793 23511 11851 23517
rect 11793 23508 11805 23511
rect 11664 23480 11805 23508
rect 11664 23468 11670 23480
rect 11793 23477 11805 23480
rect 11839 23477 11851 23511
rect 11793 23471 11851 23477
rect 12253 23511 12311 23517
rect 12253 23477 12265 23511
rect 12299 23508 12311 23511
rect 12342 23508 12348 23520
rect 12299 23480 12348 23508
rect 12299 23477 12311 23480
rect 12253 23471 12311 23477
rect 12342 23468 12348 23480
rect 12400 23468 12406 23520
rect 12802 23468 12808 23520
rect 12860 23508 12866 23520
rect 13725 23511 13783 23517
rect 13725 23508 13737 23511
rect 12860 23480 13737 23508
rect 12860 23468 12866 23480
rect 13725 23477 13737 23480
rect 13771 23508 13783 23511
rect 14292 23508 14320 23684
rect 15194 23672 15200 23724
rect 15252 23712 15258 23724
rect 15841 23715 15899 23721
rect 15841 23712 15853 23715
rect 15252 23684 15853 23712
rect 15252 23672 15258 23684
rect 15841 23681 15853 23684
rect 15887 23712 15899 23715
rect 16482 23712 16488 23724
rect 15887 23684 16488 23712
rect 15887 23681 15899 23684
rect 15841 23675 15899 23681
rect 16482 23672 16488 23684
rect 16540 23672 16546 23724
rect 16684 23712 16712 23752
rect 17034 23740 17040 23752
rect 17092 23740 17098 23792
rect 17402 23780 17408 23792
rect 17363 23752 17408 23780
rect 17402 23740 17408 23752
rect 17460 23740 17466 23792
rect 17586 23740 17592 23792
rect 17644 23780 17650 23792
rect 18322 23780 18328 23792
rect 17644 23752 18328 23780
rect 17644 23740 17650 23752
rect 18322 23740 18328 23752
rect 18380 23780 18386 23792
rect 19061 23783 19119 23789
rect 19061 23780 19073 23783
rect 18380 23752 19073 23780
rect 18380 23740 18386 23752
rect 19061 23749 19073 23752
rect 19107 23749 19119 23783
rect 19061 23743 19119 23749
rect 17954 23712 17960 23724
rect 16684 23684 17960 23712
rect 17954 23672 17960 23684
rect 18012 23672 18018 23724
rect 18598 23712 18604 23724
rect 18559 23684 18604 23712
rect 18598 23672 18604 23684
rect 18656 23672 18662 23724
rect 19889 23715 19947 23721
rect 19889 23681 19901 23715
rect 19935 23712 19947 23715
rect 20162 23712 20168 23724
rect 19935 23684 20168 23712
rect 19935 23681 19947 23684
rect 19889 23675 19947 23681
rect 20162 23672 20168 23684
rect 20220 23672 20226 23724
rect 21376 23721 21404 23820
rect 21450 23808 21456 23860
rect 21508 23848 21514 23860
rect 21913 23851 21971 23857
rect 21913 23848 21925 23851
rect 21508 23820 21925 23848
rect 21508 23808 21514 23820
rect 21913 23817 21925 23820
rect 21959 23817 21971 23851
rect 21913 23811 21971 23817
rect 22649 23851 22707 23857
rect 22649 23817 22661 23851
rect 22695 23848 22707 23851
rect 23198 23848 23204 23860
rect 22695 23820 23204 23848
rect 22695 23817 22707 23820
rect 22649 23811 22707 23817
rect 23198 23808 23204 23820
rect 23256 23808 23262 23860
rect 24210 23808 24216 23860
rect 24268 23848 24274 23860
rect 24854 23848 24860 23860
rect 24268 23820 24860 23848
rect 24268 23808 24274 23820
rect 24854 23808 24860 23820
rect 24912 23808 24918 23860
rect 25406 23848 25412 23860
rect 25367 23820 25412 23848
rect 25406 23808 25412 23820
rect 25464 23808 25470 23860
rect 22922 23740 22928 23792
rect 22980 23780 22986 23792
rect 24673 23783 24731 23789
rect 24673 23780 24685 23783
rect 22980 23752 24685 23780
rect 22980 23740 22986 23752
rect 24673 23749 24685 23752
rect 24719 23780 24731 23783
rect 24946 23780 24952 23792
rect 24719 23752 24952 23780
rect 24719 23749 24731 23752
rect 24673 23743 24731 23749
rect 24946 23740 24952 23752
rect 25004 23740 25010 23792
rect 21361 23715 21419 23721
rect 21361 23681 21373 23715
rect 21407 23681 21419 23715
rect 21361 23675 21419 23681
rect 21545 23715 21603 23721
rect 21545 23681 21557 23715
rect 21591 23712 21603 23715
rect 23477 23715 23535 23721
rect 21591 23684 22416 23712
rect 21591 23681 21603 23684
rect 21545 23675 21603 23681
rect 14369 23647 14427 23653
rect 14369 23613 14381 23647
rect 14415 23644 14427 23647
rect 15657 23647 15715 23653
rect 15657 23644 15669 23647
rect 14415 23616 15669 23644
rect 14415 23613 14427 23616
rect 14369 23607 14427 23613
rect 15657 23613 15669 23616
rect 15703 23644 15715 23647
rect 15930 23644 15936 23656
rect 15703 23616 15936 23644
rect 15703 23613 15715 23616
rect 15657 23607 15715 23613
rect 15930 23604 15936 23616
rect 15988 23604 15994 23656
rect 16206 23604 16212 23656
rect 16264 23644 16270 23656
rect 16390 23644 16396 23656
rect 16264 23616 16396 23644
rect 16264 23604 16270 23616
rect 16390 23604 16396 23616
rect 16448 23604 16454 23656
rect 16853 23647 16911 23653
rect 16853 23613 16865 23647
rect 16899 23644 16911 23647
rect 17126 23644 17132 23656
rect 16899 23616 17132 23644
rect 16899 23613 16911 23616
rect 16853 23607 16911 23613
rect 17126 23604 17132 23616
rect 17184 23644 17190 23656
rect 17773 23647 17831 23653
rect 17773 23644 17785 23647
rect 17184 23616 17785 23644
rect 17184 23604 17190 23616
rect 17773 23613 17785 23616
rect 17819 23613 17831 23647
rect 17773 23607 17831 23613
rect 18138 23604 18144 23656
rect 18196 23644 18202 23656
rect 18417 23647 18475 23653
rect 18417 23644 18429 23647
rect 18196 23616 18429 23644
rect 18196 23604 18202 23616
rect 18417 23613 18429 23616
rect 18463 23613 18475 23647
rect 18417 23607 18475 23613
rect 18506 23604 18512 23656
rect 18564 23644 18570 23656
rect 18564 23616 18609 23644
rect 18564 23604 18570 23616
rect 18782 23604 18788 23656
rect 18840 23644 18846 23656
rect 19610 23644 19616 23656
rect 18840 23616 19616 23644
rect 18840 23604 18846 23616
rect 19610 23604 19616 23616
rect 19668 23604 19674 23656
rect 20346 23604 20352 23656
rect 20404 23644 20410 23656
rect 21269 23647 21327 23653
rect 21269 23644 21281 23647
rect 20404 23616 21281 23644
rect 20404 23604 20410 23616
rect 21269 23613 21281 23616
rect 21315 23613 21327 23647
rect 21269 23607 21327 23613
rect 14737 23579 14795 23585
rect 14737 23545 14749 23579
rect 14783 23576 14795 23579
rect 15565 23579 15623 23585
rect 15565 23576 15577 23579
rect 14783 23548 15577 23576
rect 14783 23545 14795 23548
rect 14737 23539 14795 23545
rect 15565 23545 15577 23548
rect 15611 23576 15623 23579
rect 16298 23576 16304 23588
rect 15611 23548 16304 23576
rect 15611 23545 15623 23548
rect 15565 23539 15623 23545
rect 16298 23536 16304 23548
rect 16356 23536 16362 23588
rect 13771 23480 14320 23508
rect 13771 23477 13783 23480
rect 13725 23471 13783 23477
rect 14642 23468 14648 23520
rect 14700 23508 14706 23520
rect 15013 23511 15071 23517
rect 15013 23508 15025 23511
rect 14700 23480 15025 23508
rect 14700 23468 14706 23480
rect 15013 23477 15025 23480
rect 15059 23477 15071 23511
rect 15013 23471 15071 23477
rect 16761 23511 16819 23517
rect 16761 23477 16773 23511
rect 16807 23508 16819 23511
rect 16942 23508 16948 23520
rect 16807 23480 16948 23508
rect 16807 23477 16819 23480
rect 16761 23471 16819 23477
rect 16942 23468 16948 23480
rect 17000 23468 17006 23520
rect 19150 23468 19156 23520
rect 19208 23508 19214 23520
rect 19521 23511 19579 23517
rect 19521 23508 19533 23511
rect 19208 23480 19533 23508
rect 19208 23468 19214 23480
rect 19521 23477 19533 23480
rect 19567 23508 19579 23511
rect 20162 23508 20168 23520
rect 19567 23480 20168 23508
rect 19567 23477 19579 23480
rect 19521 23471 19579 23477
rect 20162 23468 20168 23480
rect 20220 23468 20226 23520
rect 20901 23511 20959 23517
rect 20901 23477 20913 23511
rect 20947 23508 20959 23511
rect 21358 23508 21364 23520
rect 20947 23480 21364 23508
rect 20947 23477 20959 23480
rect 20901 23471 20959 23477
rect 21358 23468 21364 23480
rect 21416 23468 21422 23520
rect 22388 23517 22416 23684
rect 23477 23681 23489 23715
rect 23523 23712 23535 23715
rect 24302 23712 24308 23724
rect 23523 23684 24308 23712
rect 23523 23681 23535 23684
rect 23477 23675 23535 23681
rect 24302 23672 24308 23684
rect 24360 23672 24366 23724
rect 25038 23672 25044 23724
rect 25096 23712 25102 23724
rect 25133 23715 25191 23721
rect 25133 23712 25145 23715
rect 25096 23684 25145 23712
rect 25096 23672 25102 23684
rect 25133 23681 25145 23684
rect 25179 23712 25191 23715
rect 25866 23712 25872 23724
rect 25179 23684 25872 23712
rect 25179 23681 25191 23684
rect 25133 23675 25191 23681
rect 25866 23672 25872 23684
rect 25924 23672 25930 23724
rect 22465 23647 22523 23653
rect 22465 23613 22477 23647
rect 22511 23644 22523 23647
rect 25225 23647 25283 23653
rect 22511 23616 23060 23644
rect 22511 23613 22523 23616
rect 22465 23607 22523 23613
rect 23032 23520 23060 23616
rect 25225 23613 25237 23647
rect 25271 23644 25283 23647
rect 25593 23647 25651 23653
rect 25593 23644 25605 23647
rect 25271 23616 25605 23644
rect 25271 23613 25283 23616
rect 25225 23607 25283 23613
rect 25593 23613 25605 23616
rect 25639 23613 25651 23647
rect 25593 23607 25651 23613
rect 24118 23576 24124 23588
rect 24031 23548 24124 23576
rect 24118 23536 24124 23548
rect 24176 23576 24182 23588
rect 26237 23579 26295 23585
rect 26237 23576 26249 23579
rect 24176 23548 26249 23576
rect 24176 23536 24182 23548
rect 26237 23545 26249 23548
rect 26283 23545 26295 23579
rect 26237 23539 26295 23545
rect 22373 23511 22431 23517
rect 22373 23477 22385 23511
rect 22419 23508 22431 23511
rect 22462 23508 22468 23520
rect 22419 23480 22468 23508
rect 22419 23477 22431 23480
rect 22373 23471 22431 23477
rect 22462 23468 22468 23480
rect 22520 23468 22526 23520
rect 23014 23508 23020 23520
rect 22975 23480 23020 23508
rect 23014 23468 23020 23480
rect 23072 23468 23078 23520
rect 23658 23508 23664 23520
rect 23619 23480 23664 23508
rect 23658 23468 23664 23480
rect 23716 23468 23722 23520
rect 24029 23511 24087 23517
rect 24029 23477 24041 23511
rect 24075 23508 24087 23511
rect 24302 23508 24308 23520
rect 24075 23480 24308 23508
rect 24075 23477 24087 23480
rect 24029 23471 24087 23477
rect 24302 23468 24308 23480
rect 24360 23468 24366 23520
rect 25593 23511 25651 23517
rect 25593 23477 25605 23511
rect 25639 23508 25651 23511
rect 25869 23511 25927 23517
rect 25869 23508 25881 23511
rect 25639 23480 25881 23508
rect 25639 23477 25651 23480
rect 25593 23471 25651 23477
rect 25869 23477 25881 23480
rect 25915 23508 25927 23511
rect 26142 23508 26148 23520
rect 25915 23480 26148 23508
rect 25915 23477 25927 23480
rect 25869 23471 25927 23477
rect 26142 23468 26148 23480
rect 26200 23468 26206 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 7190 23304 7196 23316
rect 7151 23276 7196 23304
rect 7190 23264 7196 23276
rect 7248 23264 7254 23316
rect 11609 23307 11667 23313
rect 11609 23273 11621 23307
rect 11655 23304 11667 23307
rect 11882 23304 11888 23316
rect 11655 23276 11888 23304
rect 11655 23273 11667 23276
rect 11609 23267 11667 23273
rect 11882 23264 11888 23276
rect 11940 23264 11946 23316
rect 15102 23304 15108 23316
rect 15063 23276 15108 23304
rect 15102 23264 15108 23276
rect 15160 23264 15166 23316
rect 16574 23264 16580 23316
rect 16632 23304 16638 23316
rect 16669 23307 16727 23313
rect 16669 23304 16681 23307
rect 16632 23276 16681 23304
rect 16632 23264 16638 23276
rect 16669 23273 16681 23276
rect 16715 23273 16727 23307
rect 16669 23267 16727 23273
rect 17218 23264 17224 23316
rect 17276 23304 17282 23316
rect 17313 23307 17371 23313
rect 17313 23304 17325 23307
rect 17276 23276 17325 23304
rect 17276 23264 17282 23276
rect 17313 23273 17325 23276
rect 17359 23273 17371 23307
rect 18138 23304 18144 23316
rect 18099 23276 18144 23304
rect 17313 23267 17371 23273
rect 18138 23264 18144 23276
rect 18196 23264 18202 23316
rect 18414 23304 18420 23316
rect 18375 23276 18420 23304
rect 18414 23264 18420 23276
rect 18472 23264 18478 23316
rect 18690 23264 18696 23316
rect 18748 23264 18754 23316
rect 21174 23304 21180 23316
rect 21135 23276 21180 23304
rect 21174 23264 21180 23276
rect 21232 23264 21238 23316
rect 23477 23307 23535 23313
rect 23477 23273 23489 23307
rect 23523 23273 23535 23307
rect 25222 23304 25228 23316
rect 25183 23276 25228 23304
rect 23477 23267 23535 23273
rect 7837 23239 7895 23245
rect 7837 23205 7849 23239
rect 7883 23236 7895 23239
rect 8202 23236 8208 23248
rect 7883 23208 8208 23236
rect 7883 23205 7895 23208
rect 7837 23199 7895 23205
rect 8202 23196 8208 23208
rect 8260 23196 8266 23248
rect 11146 23196 11152 23248
rect 11204 23236 11210 23248
rect 14737 23239 14795 23245
rect 11204 23208 14688 23236
rect 11204 23196 11210 23208
rect 2133 23171 2191 23177
rect 2133 23137 2145 23171
rect 2179 23168 2191 23171
rect 2406 23168 2412 23180
rect 2179 23140 2412 23168
rect 2179 23137 2191 23140
rect 2133 23131 2191 23137
rect 2406 23128 2412 23140
rect 2464 23128 2470 23180
rect 7466 23128 7472 23180
rect 7524 23168 7530 23180
rect 7561 23171 7619 23177
rect 7561 23168 7573 23171
rect 7524 23140 7573 23168
rect 7524 23128 7530 23140
rect 7561 23137 7573 23140
rect 7607 23137 7619 23171
rect 7561 23131 7619 23137
rect 9306 23128 9312 23180
rect 9364 23168 9370 23180
rect 9493 23171 9551 23177
rect 9493 23168 9505 23171
rect 9364 23140 9505 23168
rect 9364 23128 9370 23140
rect 9493 23137 9505 23140
rect 9539 23168 9551 23171
rect 10413 23171 10471 23177
rect 10413 23168 10425 23171
rect 9539 23140 10425 23168
rect 9539 23137 9551 23140
rect 9493 23131 9551 23137
rect 10413 23137 10425 23140
rect 10459 23137 10471 23171
rect 10413 23131 10471 23137
rect 10505 23171 10563 23177
rect 10505 23137 10517 23171
rect 10551 23168 10563 23171
rect 10686 23168 10692 23180
rect 10551 23140 10692 23168
rect 10551 23137 10563 23140
rect 10505 23131 10563 23137
rect 10686 23128 10692 23140
rect 10744 23128 10750 23180
rect 11882 23128 11888 23180
rect 11940 23168 11946 23180
rect 11977 23171 12035 23177
rect 11977 23168 11989 23171
rect 11940 23140 11989 23168
rect 11940 23128 11946 23140
rect 11977 23137 11989 23140
rect 12023 23137 12035 23171
rect 11977 23131 12035 23137
rect 13262 23128 13268 23180
rect 13320 23168 13326 23180
rect 13541 23171 13599 23177
rect 13541 23168 13553 23171
rect 13320 23140 13553 23168
rect 13320 23128 13326 23140
rect 13541 23137 13553 23140
rect 13587 23168 13599 23171
rect 14185 23171 14243 23177
rect 14185 23168 14197 23171
rect 13587 23140 14197 23168
rect 13587 23137 13599 23140
rect 13541 23131 13599 23137
rect 14185 23137 14197 23140
rect 14231 23137 14243 23171
rect 14660 23168 14688 23208
rect 14737 23205 14749 23239
rect 14783 23236 14795 23239
rect 15010 23236 15016 23248
rect 14783 23208 15016 23236
rect 14783 23205 14795 23208
rect 14737 23199 14795 23205
rect 15010 23196 15016 23208
rect 15068 23196 15074 23248
rect 15657 23239 15715 23245
rect 15657 23205 15669 23239
rect 15703 23236 15715 23239
rect 15838 23236 15844 23248
rect 15703 23208 15844 23236
rect 15703 23205 15715 23208
rect 15657 23199 15715 23205
rect 15838 23196 15844 23208
rect 15896 23196 15902 23248
rect 17862 23196 17868 23248
rect 17920 23236 17926 23248
rect 18708 23236 18736 23264
rect 23492 23236 23520 23267
rect 25222 23264 25228 23276
rect 25280 23264 25286 23316
rect 24302 23236 24308 23248
rect 17920 23208 18920 23236
rect 23492 23208 24308 23236
rect 17920 23196 17926 23208
rect 15749 23171 15807 23177
rect 15749 23168 15761 23171
rect 14660 23140 15761 23168
rect 14185 23131 14243 23137
rect 15672 23112 15700 23140
rect 15749 23137 15761 23140
rect 15795 23137 15807 23171
rect 15749 23131 15807 23137
rect 17126 23128 17132 23180
rect 17184 23168 17190 23180
rect 17221 23171 17279 23177
rect 17221 23168 17233 23171
rect 17184 23140 17233 23168
rect 17184 23128 17190 23140
rect 17221 23137 17233 23140
rect 17267 23137 17279 23171
rect 17221 23131 17279 23137
rect 18690 23128 18696 23180
rect 18748 23168 18754 23180
rect 18785 23171 18843 23177
rect 18785 23168 18797 23171
rect 18748 23140 18797 23168
rect 18748 23128 18754 23140
rect 18785 23137 18797 23140
rect 18831 23137 18843 23171
rect 18892 23168 18920 23208
rect 24302 23196 24308 23208
rect 24360 23236 24366 23248
rect 25593 23239 25651 23245
rect 25593 23236 25605 23239
rect 24360 23208 25605 23236
rect 24360 23196 24366 23208
rect 25593 23205 25605 23208
rect 25639 23205 25651 23239
rect 25593 23199 25651 23205
rect 19613 23171 19671 23177
rect 19613 23168 19625 23171
rect 18892 23140 19625 23168
rect 18785 23131 18843 23137
rect 1670 23100 1676 23112
rect 1631 23072 1676 23100
rect 1670 23060 1676 23072
rect 1728 23060 1734 23112
rect 2314 23100 2320 23112
rect 2275 23072 2320 23100
rect 2314 23060 2320 23072
rect 2372 23060 2378 23112
rect 10594 23060 10600 23112
rect 10652 23100 10658 23112
rect 12066 23100 12072 23112
rect 10652 23072 10697 23100
rect 12027 23072 12072 23100
rect 10652 23060 10658 23072
rect 12066 23060 12072 23072
rect 12124 23060 12130 23112
rect 12161 23103 12219 23109
rect 12161 23069 12173 23103
rect 12207 23069 12219 23103
rect 12161 23063 12219 23069
rect 12713 23103 12771 23109
rect 12713 23069 12725 23103
rect 12759 23100 12771 23103
rect 13446 23100 13452 23112
rect 12759 23072 13452 23100
rect 12759 23069 12771 23072
rect 12713 23063 12771 23069
rect 9125 23035 9183 23041
rect 9125 23001 9137 23035
rect 9171 23032 9183 23035
rect 9490 23032 9496 23044
rect 9171 23004 9496 23032
rect 9171 23001 9183 23004
rect 9125 22995 9183 23001
rect 9490 22992 9496 23004
rect 9548 23032 9554 23044
rect 10045 23035 10103 23041
rect 10045 23032 10057 23035
rect 9548 23004 10057 23032
rect 9548 22992 9554 23004
rect 10045 23001 10057 23004
rect 10091 23001 10103 23035
rect 10045 22995 10103 23001
rect 11425 23035 11483 23041
rect 11425 23001 11437 23035
rect 11471 23032 11483 23035
rect 11790 23032 11796 23044
rect 11471 23004 11796 23032
rect 11471 23001 11483 23004
rect 11425 22995 11483 23001
rect 11790 22992 11796 23004
rect 11848 23032 11854 23044
rect 12176 23032 12204 23063
rect 13446 23060 13452 23072
rect 13504 23100 13510 23112
rect 13633 23103 13691 23109
rect 13633 23100 13645 23103
rect 13504 23072 13645 23100
rect 13504 23060 13510 23072
rect 13633 23069 13645 23072
rect 13679 23069 13691 23103
rect 13633 23063 13691 23069
rect 13722 23060 13728 23112
rect 13780 23100 13786 23112
rect 13780 23072 13825 23100
rect 13780 23060 13786 23072
rect 15654 23060 15660 23112
rect 15712 23060 15718 23112
rect 15930 23100 15936 23112
rect 15891 23072 15936 23100
rect 15930 23060 15936 23072
rect 15988 23060 15994 23112
rect 16393 23103 16451 23109
rect 16393 23069 16405 23103
rect 16439 23100 16451 23103
rect 17402 23100 17408 23112
rect 16439 23072 17408 23100
rect 16439 23069 16451 23072
rect 16393 23063 16451 23069
rect 11848 23004 12204 23032
rect 11848 22992 11854 23004
rect 13354 22992 13360 23044
rect 13412 23032 13418 23044
rect 13538 23032 13544 23044
rect 13412 23004 13544 23032
rect 13412 22992 13418 23004
rect 13538 22992 13544 23004
rect 13596 22992 13602 23044
rect 13998 22992 14004 23044
rect 14056 23032 14062 23044
rect 16408 23032 16436 23063
rect 17402 23060 17408 23072
rect 17460 23060 17466 23112
rect 18874 23100 18880 23112
rect 18835 23072 18880 23100
rect 18874 23060 18880 23072
rect 18932 23060 18938 23112
rect 18984 23109 19012 23140
rect 19613 23137 19625 23140
rect 19659 23168 19671 23171
rect 20070 23168 20076 23180
rect 19659 23140 20076 23168
rect 19659 23137 19671 23140
rect 19613 23131 19671 23137
rect 20070 23128 20076 23140
rect 20128 23128 20134 23180
rect 21174 23128 21180 23180
rect 21232 23168 21238 23180
rect 22281 23171 22339 23177
rect 22281 23168 22293 23171
rect 21232 23140 22293 23168
rect 21232 23128 21238 23140
rect 22281 23137 22293 23140
rect 22327 23137 22339 23171
rect 23842 23168 23848 23180
rect 23803 23140 23848 23168
rect 22281 23131 22339 23137
rect 23842 23128 23848 23140
rect 23900 23128 23906 23180
rect 25038 23168 25044 23180
rect 24999 23140 25044 23168
rect 25038 23128 25044 23140
rect 25096 23128 25102 23180
rect 18969 23103 19027 23109
rect 18969 23069 18981 23103
rect 19015 23069 19027 23103
rect 18969 23063 19027 23069
rect 21542 23060 21548 23112
rect 21600 23100 21606 23112
rect 22373 23103 22431 23109
rect 22373 23100 22385 23103
rect 21600 23072 22385 23100
rect 21600 23060 21606 23072
rect 22373 23069 22385 23072
rect 22419 23069 22431 23103
rect 22373 23063 22431 23069
rect 22462 23060 22468 23112
rect 22520 23100 22526 23112
rect 23934 23100 23940 23112
rect 22520 23072 22565 23100
rect 23895 23072 23940 23100
rect 22520 23060 22526 23072
rect 23934 23060 23940 23072
rect 23992 23060 23998 23112
rect 24118 23100 24124 23112
rect 24079 23072 24124 23100
rect 24118 23060 24124 23072
rect 24176 23060 24182 23112
rect 14056 23004 16436 23032
rect 22480 23032 22508 23060
rect 24673 23035 24731 23041
rect 24673 23032 24685 23035
rect 22480 23004 24685 23032
rect 14056 22992 14062 23004
rect 24673 23001 24685 23004
rect 24719 23032 24731 23035
rect 24762 23032 24768 23044
rect 24719 23004 24768 23032
rect 24719 23001 24731 23004
rect 24673 22995 24731 23001
rect 24762 22992 24768 23004
rect 24820 22992 24826 23044
rect 6917 22967 6975 22973
rect 6917 22933 6929 22967
rect 6963 22964 6975 22967
rect 7006 22964 7012 22976
rect 6963 22936 7012 22964
rect 6963 22933 6975 22936
rect 6917 22927 6975 22933
rect 7006 22924 7012 22936
rect 7064 22924 7070 22976
rect 8665 22967 8723 22973
rect 8665 22933 8677 22967
rect 8711 22964 8723 22967
rect 8938 22964 8944 22976
rect 8711 22936 8944 22964
rect 8711 22933 8723 22936
rect 8665 22927 8723 22933
rect 8938 22924 8944 22936
rect 8996 22924 9002 22976
rect 9953 22967 10011 22973
rect 9953 22933 9965 22967
rect 9999 22964 10011 22967
rect 10962 22964 10968 22976
rect 9999 22936 10968 22964
rect 9999 22933 10011 22936
rect 9953 22927 10011 22933
rect 10962 22924 10968 22936
rect 11020 22924 11026 22976
rect 12894 22924 12900 22976
rect 12952 22964 12958 22976
rect 12989 22967 13047 22973
rect 12989 22964 13001 22967
rect 12952 22936 13001 22964
rect 12952 22924 12958 22936
rect 12989 22933 13001 22936
rect 13035 22933 13047 22967
rect 12989 22927 13047 22933
rect 13173 22967 13231 22973
rect 13173 22933 13185 22967
rect 13219 22964 13231 22967
rect 13906 22964 13912 22976
rect 13219 22936 13912 22964
rect 13219 22933 13231 22936
rect 13173 22927 13231 22933
rect 13906 22924 13912 22936
rect 13964 22924 13970 22976
rect 15289 22967 15347 22973
rect 15289 22933 15301 22967
rect 15335 22964 15347 22967
rect 16206 22964 16212 22976
rect 15335 22936 16212 22964
rect 15335 22933 15347 22936
rect 15289 22927 15347 22933
rect 16206 22924 16212 22936
rect 16264 22924 16270 22976
rect 16853 22967 16911 22973
rect 16853 22933 16865 22967
rect 16899 22964 16911 22967
rect 17586 22964 17592 22976
rect 16899 22936 17592 22964
rect 16899 22933 16911 22936
rect 16853 22927 16911 22933
rect 17586 22924 17592 22936
rect 17644 22924 17650 22976
rect 20346 22964 20352 22976
rect 20307 22936 20352 22964
rect 20346 22924 20352 22936
rect 20404 22924 20410 22976
rect 20714 22964 20720 22976
rect 20675 22936 20720 22964
rect 20714 22924 20720 22936
rect 20772 22924 20778 22976
rect 21450 22964 21456 22976
rect 21411 22936 21456 22964
rect 21450 22924 21456 22936
rect 21508 22924 21514 22976
rect 21910 22964 21916 22976
rect 21871 22936 21916 22964
rect 21910 22924 21916 22936
rect 21968 22924 21974 22976
rect 23201 22967 23259 22973
rect 23201 22933 23213 22967
rect 23247 22964 23259 22967
rect 23382 22964 23388 22976
rect 23247 22936 23388 22964
rect 23247 22933 23259 22936
rect 23201 22927 23259 22933
rect 23382 22924 23388 22936
rect 23440 22924 23446 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1578 22760 1584 22772
rect 1539 22732 1584 22760
rect 1578 22720 1584 22732
rect 1636 22720 1642 22772
rect 4062 22720 4068 22772
rect 4120 22760 4126 22772
rect 4617 22763 4675 22769
rect 4617 22760 4629 22763
rect 4120 22732 4629 22760
rect 4120 22720 4126 22732
rect 4617 22729 4629 22732
rect 4663 22729 4675 22763
rect 9030 22760 9036 22772
rect 8991 22732 9036 22760
rect 4617 22723 4675 22729
rect 9030 22720 9036 22732
rect 9088 22720 9094 22772
rect 10042 22720 10048 22772
rect 10100 22760 10106 22772
rect 10137 22763 10195 22769
rect 10137 22760 10149 22763
rect 10100 22732 10149 22760
rect 10100 22720 10106 22732
rect 10137 22729 10149 22732
rect 10183 22760 10195 22763
rect 10594 22760 10600 22772
rect 10183 22732 10600 22760
rect 10183 22729 10195 22732
rect 10137 22723 10195 22729
rect 10594 22720 10600 22732
rect 10652 22720 10658 22772
rect 11606 22720 11612 22772
rect 11664 22760 11670 22772
rect 11701 22763 11759 22769
rect 11701 22760 11713 22763
rect 11664 22732 11713 22760
rect 11664 22720 11670 22732
rect 11701 22729 11713 22732
rect 11747 22760 11759 22763
rect 12066 22760 12072 22772
rect 11747 22732 12072 22760
rect 11747 22729 11759 22732
rect 11701 22723 11759 22729
rect 12066 22720 12072 22732
rect 12124 22720 12130 22772
rect 13262 22760 13268 22772
rect 13223 22732 13268 22760
rect 13262 22720 13268 22732
rect 13320 22720 13326 22772
rect 15473 22763 15531 22769
rect 15473 22729 15485 22763
rect 15519 22760 15531 22763
rect 15654 22760 15660 22772
rect 15519 22732 15660 22760
rect 15519 22729 15531 22732
rect 15473 22723 15531 22729
rect 15654 22720 15660 22732
rect 15712 22720 15718 22772
rect 17218 22720 17224 22772
rect 17276 22760 17282 22772
rect 17405 22763 17463 22769
rect 17405 22760 17417 22763
rect 17276 22732 17417 22760
rect 17276 22720 17282 22732
rect 17405 22729 17417 22732
rect 17451 22760 17463 22763
rect 17678 22760 17684 22772
rect 17451 22732 17684 22760
rect 17451 22729 17463 22732
rect 17405 22723 17463 22729
rect 17678 22720 17684 22732
rect 17736 22720 17742 22772
rect 19610 22760 19616 22772
rect 19571 22732 19616 22760
rect 19610 22720 19616 22732
rect 19668 22720 19674 22772
rect 21818 22760 21824 22772
rect 21779 22732 21824 22760
rect 21818 22720 21824 22732
rect 21876 22720 21882 22772
rect 25038 22760 25044 22772
rect 24999 22732 25044 22760
rect 25038 22720 25044 22732
rect 25096 22720 25102 22772
rect 25590 22760 25596 22772
rect 25551 22732 25596 22760
rect 25590 22720 25596 22732
rect 25648 22720 25654 22772
rect 8941 22695 8999 22701
rect 8941 22661 8953 22695
rect 8987 22692 8999 22695
rect 9398 22692 9404 22704
rect 8987 22664 9404 22692
rect 8987 22661 8999 22664
rect 8941 22655 8999 22661
rect 9398 22652 9404 22664
rect 9456 22692 9462 22704
rect 9456 22664 9628 22692
rect 9456 22652 9462 22664
rect 6638 22584 6644 22636
rect 6696 22624 6702 22636
rect 7745 22627 7803 22633
rect 7745 22624 7757 22627
rect 6696 22596 7757 22624
rect 6696 22584 6702 22596
rect 7745 22593 7757 22596
rect 7791 22624 7803 22627
rect 8110 22624 8116 22636
rect 7791 22596 8116 22624
rect 7791 22593 7803 22596
rect 7745 22587 7803 22593
rect 8110 22584 8116 22596
rect 8168 22584 8174 22636
rect 9490 22624 9496 22636
rect 9451 22596 9496 22624
rect 9490 22584 9496 22596
rect 9548 22584 9554 22636
rect 9600 22633 9628 22664
rect 18138 22652 18144 22704
rect 18196 22692 18202 22704
rect 20717 22695 20775 22701
rect 20717 22692 20729 22695
rect 18196 22664 20729 22692
rect 18196 22652 18202 22664
rect 9585 22627 9643 22633
rect 9585 22593 9597 22627
rect 9631 22593 9643 22627
rect 11149 22627 11207 22633
rect 11149 22624 11161 22627
rect 9585 22587 9643 22593
rect 10428 22596 11161 22624
rect 1397 22559 1455 22565
rect 1397 22525 1409 22559
rect 1443 22556 1455 22559
rect 4433 22559 4491 22565
rect 1443 22528 2084 22556
rect 1443 22525 1455 22528
rect 1397 22519 1455 22525
rect 2056 22429 2084 22528
rect 4433 22525 4445 22559
rect 4479 22556 4491 22559
rect 4985 22559 5043 22565
rect 4985 22556 4997 22559
rect 4479 22528 4997 22556
rect 4479 22525 4491 22528
rect 4433 22519 4491 22525
rect 4985 22525 4997 22528
rect 5031 22556 5043 22559
rect 5350 22556 5356 22568
rect 5031 22528 5356 22556
rect 5031 22525 5043 22528
rect 4985 22519 5043 22525
rect 5350 22516 5356 22528
rect 5408 22516 5414 22568
rect 7098 22556 7104 22568
rect 7011 22528 7104 22556
rect 7098 22516 7104 22528
rect 7156 22556 7162 22568
rect 7650 22556 7656 22568
rect 7156 22528 7656 22556
rect 7156 22516 7162 22528
rect 7650 22516 7656 22528
rect 7708 22516 7714 22568
rect 9030 22516 9036 22568
rect 9088 22556 9094 22568
rect 9401 22559 9459 22565
rect 9401 22556 9413 22559
rect 9088 22528 9413 22556
rect 9088 22516 9094 22528
rect 9401 22525 9413 22528
rect 9447 22525 9459 22559
rect 9401 22519 9459 22525
rect 4798 22448 4804 22500
rect 4856 22488 4862 22500
rect 5537 22491 5595 22497
rect 5537 22488 5549 22491
rect 4856 22460 5549 22488
rect 4856 22448 4862 22460
rect 5537 22457 5549 22460
rect 5583 22488 5595 22491
rect 5905 22491 5963 22497
rect 5905 22488 5917 22491
rect 5583 22460 5917 22488
rect 5583 22457 5595 22460
rect 5537 22451 5595 22457
rect 5905 22457 5917 22460
rect 5951 22488 5963 22491
rect 6273 22491 6331 22497
rect 6273 22488 6285 22491
rect 5951 22460 6285 22488
rect 5951 22457 5963 22460
rect 5905 22451 5963 22457
rect 6273 22457 6285 22460
rect 6319 22488 6331 22491
rect 7006 22488 7012 22500
rect 6319 22460 7012 22488
rect 6319 22457 6331 22460
rect 6273 22451 6331 22457
rect 7006 22448 7012 22460
rect 7064 22448 7070 22500
rect 7282 22448 7288 22500
rect 7340 22488 7346 22500
rect 7561 22491 7619 22497
rect 7561 22488 7573 22491
rect 7340 22460 7573 22488
rect 7340 22448 7346 22460
rect 7561 22457 7573 22460
rect 7607 22457 7619 22491
rect 7561 22451 7619 22457
rect 2041 22423 2099 22429
rect 2041 22389 2053 22423
rect 2087 22420 2099 22423
rect 2130 22420 2136 22432
rect 2087 22392 2136 22420
rect 2087 22389 2099 22392
rect 2041 22383 2099 22389
rect 2130 22380 2136 22392
rect 2188 22380 2194 22432
rect 2406 22420 2412 22432
rect 2367 22392 2412 22420
rect 2406 22380 2412 22392
rect 2464 22380 2470 22432
rect 6638 22420 6644 22432
rect 6599 22392 6644 22420
rect 6638 22380 6644 22392
rect 6696 22380 6702 22432
rect 7190 22420 7196 22432
rect 7151 22392 7196 22420
rect 7190 22380 7196 22392
rect 7248 22380 7254 22432
rect 8202 22420 8208 22432
rect 8163 22392 8208 22420
rect 8202 22380 8208 22392
rect 8260 22380 8266 22432
rect 9950 22380 9956 22432
rect 10008 22420 10014 22432
rect 10428 22429 10456 22596
rect 11149 22593 11161 22596
rect 11195 22593 11207 22627
rect 11149 22587 11207 22593
rect 12894 22584 12900 22636
rect 12952 22624 12958 22636
rect 13725 22627 13783 22633
rect 13725 22624 13737 22627
rect 12952 22596 13737 22624
rect 12952 22584 12958 22596
rect 13725 22593 13737 22596
rect 13771 22593 13783 22627
rect 13725 22587 13783 22593
rect 13909 22627 13967 22633
rect 13909 22593 13921 22627
rect 13955 22593 13967 22627
rect 13909 22587 13967 22593
rect 10962 22516 10968 22568
rect 11020 22556 11026 22568
rect 11057 22559 11115 22565
rect 11057 22556 11069 22559
rect 11020 22528 11069 22556
rect 11020 22516 11026 22528
rect 11057 22525 11069 22528
rect 11103 22525 11115 22559
rect 11057 22519 11115 22525
rect 12434 22516 12440 22568
rect 12492 22556 12498 22568
rect 13173 22559 13231 22565
rect 13173 22556 13185 22559
rect 12492 22528 13185 22556
rect 12492 22516 12498 22528
rect 13173 22525 13185 22528
rect 13219 22556 13231 22559
rect 13633 22559 13691 22565
rect 13633 22556 13645 22559
rect 13219 22528 13645 22556
rect 13219 22525 13231 22528
rect 13173 22519 13231 22525
rect 13633 22525 13645 22528
rect 13679 22556 13691 22559
rect 13814 22556 13820 22568
rect 13679 22528 13820 22556
rect 13679 22525 13691 22528
rect 13633 22519 13691 22525
rect 13814 22516 13820 22528
rect 13872 22516 13878 22568
rect 13924 22556 13952 22587
rect 14366 22584 14372 22636
rect 14424 22624 14430 22636
rect 14461 22627 14519 22633
rect 14461 22624 14473 22627
rect 14424 22596 14473 22624
rect 14424 22584 14430 22596
rect 14461 22593 14473 22596
rect 14507 22624 14519 22627
rect 14507 22596 15148 22624
rect 14507 22593 14519 22596
rect 14461 22587 14519 22593
rect 14550 22556 14556 22568
rect 13924 22528 14556 22556
rect 14550 22516 14556 22528
rect 14608 22516 14614 22568
rect 14921 22559 14979 22565
rect 14921 22556 14933 22559
rect 14752 22528 14933 22556
rect 12805 22491 12863 22497
rect 12805 22457 12817 22491
rect 12851 22488 12863 22491
rect 13722 22488 13728 22500
rect 12851 22460 13728 22488
rect 12851 22457 12863 22460
rect 12805 22451 12863 22457
rect 13722 22448 13728 22460
rect 13780 22448 13786 22500
rect 14752 22432 14780 22528
rect 14921 22525 14933 22528
rect 14967 22525 14979 22559
rect 15120 22556 15148 22596
rect 15930 22584 15936 22636
rect 15988 22624 15994 22636
rect 16577 22627 16635 22633
rect 16577 22624 16589 22627
rect 15988 22596 16589 22624
rect 15988 22584 15994 22596
rect 16577 22593 16589 22596
rect 16623 22593 16635 22627
rect 16577 22587 16635 22593
rect 17218 22584 17224 22636
rect 17276 22624 17282 22636
rect 18230 22624 18236 22636
rect 17276 22596 18236 22624
rect 17276 22584 17282 22596
rect 18230 22584 18236 22596
rect 18288 22584 18294 22636
rect 18322 22584 18328 22636
rect 18380 22624 18386 22636
rect 18616 22633 18644 22664
rect 20717 22661 20729 22664
rect 20763 22661 20775 22695
rect 23842 22692 23848 22704
rect 23755 22664 23848 22692
rect 20717 22655 20775 22661
rect 23842 22652 23848 22664
rect 23900 22692 23906 22704
rect 24762 22692 24768 22704
rect 23900 22664 24768 22692
rect 23900 22652 23906 22664
rect 24762 22652 24768 22664
rect 24820 22652 24826 22704
rect 18509 22627 18567 22633
rect 18509 22624 18521 22627
rect 18380 22596 18521 22624
rect 18380 22584 18386 22596
rect 18509 22593 18521 22596
rect 18555 22593 18567 22627
rect 18509 22587 18567 22593
rect 18601 22627 18659 22633
rect 18601 22593 18613 22627
rect 18647 22593 18659 22627
rect 18601 22587 18659 22593
rect 20070 22584 20076 22636
rect 20128 22624 20134 22636
rect 20165 22627 20223 22633
rect 20165 22624 20177 22627
rect 20128 22596 20177 22624
rect 20128 22584 20134 22596
rect 20165 22593 20177 22596
rect 20211 22593 20223 22627
rect 20165 22587 20223 22593
rect 22465 22627 22523 22633
rect 22465 22593 22477 22627
rect 22511 22624 22523 22627
rect 23198 22624 23204 22636
rect 22511 22596 23204 22624
rect 22511 22593 22523 22596
rect 22465 22587 22523 22593
rect 23198 22584 23204 22596
rect 23256 22624 23262 22636
rect 24118 22624 24124 22636
rect 23256 22596 24124 22624
rect 23256 22584 23262 22596
rect 24118 22584 24124 22596
rect 24176 22584 24182 22636
rect 24486 22624 24492 22636
rect 24447 22596 24492 22624
rect 24486 22584 24492 22596
rect 24544 22584 24550 22636
rect 16485 22559 16543 22565
rect 16485 22556 16497 22559
rect 15120 22528 16497 22556
rect 14921 22519 14979 22525
rect 16485 22525 16497 22528
rect 16531 22525 16543 22559
rect 16485 22519 16543 22525
rect 18138 22516 18144 22568
rect 18196 22556 18202 22568
rect 18690 22556 18696 22568
rect 18196 22528 18696 22556
rect 18196 22516 18202 22528
rect 18690 22516 18696 22528
rect 18748 22556 18754 22568
rect 19061 22559 19119 22565
rect 19061 22556 19073 22559
rect 18748 22528 19073 22556
rect 18748 22516 18754 22528
rect 19061 22525 19073 22528
rect 19107 22525 19119 22559
rect 25406 22556 25412 22568
rect 25367 22528 25412 22556
rect 19061 22519 19119 22525
rect 25406 22516 25412 22528
rect 25464 22556 25470 22568
rect 25961 22559 26019 22565
rect 25961 22556 25973 22559
rect 25464 22528 25973 22556
rect 25464 22516 25470 22528
rect 25961 22525 25973 22528
rect 26007 22525 26019 22559
rect 25961 22519 26019 22525
rect 16574 22488 16580 22500
rect 16040 22460 16580 22488
rect 10413 22423 10471 22429
rect 10413 22420 10425 22423
rect 10008 22392 10425 22420
rect 10008 22380 10014 22392
rect 10413 22389 10425 22392
rect 10459 22389 10471 22423
rect 10413 22383 10471 22389
rect 10597 22423 10655 22429
rect 10597 22389 10609 22423
rect 10643 22420 10655 22423
rect 10686 22420 10692 22432
rect 10643 22392 10692 22420
rect 10643 22389 10655 22392
rect 10597 22383 10655 22389
rect 10686 22380 10692 22392
rect 10744 22380 10750 22432
rect 10965 22423 11023 22429
rect 10965 22389 10977 22423
rect 11011 22420 11023 22423
rect 11054 22420 11060 22432
rect 11011 22392 11060 22420
rect 11011 22389 11023 22392
rect 10965 22383 11023 22389
rect 11054 22380 11060 22392
rect 11112 22380 11118 22432
rect 11882 22380 11888 22432
rect 11940 22420 11946 22432
rect 11977 22423 12035 22429
rect 11977 22420 11989 22423
rect 11940 22392 11989 22420
rect 11940 22380 11946 22392
rect 11977 22389 11989 22392
rect 12023 22389 12035 22423
rect 14734 22420 14740 22432
rect 14695 22392 14740 22420
rect 11977 22383 12035 22389
rect 14734 22380 14740 22392
rect 14792 22380 14798 22432
rect 15102 22420 15108 22432
rect 15063 22392 15108 22420
rect 15102 22380 15108 22392
rect 15160 22380 15166 22432
rect 15838 22420 15844 22432
rect 15799 22392 15844 22420
rect 15838 22380 15844 22392
rect 15896 22380 15902 22432
rect 16040 22429 16068 22460
rect 16574 22448 16580 22460
rect 16632 22448 16638 22500
rect 18417 22491 18475 22497
rect 18417 22488 18429 22491
rect 17788 22460 18429 22488
rect 16025 22423 16083 22429
rect 16025 22389 16037 22423
rect 16071 22389 16083 22423
rect 16390 22420 16396 22432
rect 16351 22392 16396 22420
rect 16025 22383 16083 22389
rect 16390 22380 16396 22392
rect 16448 22380 16454 22432
rect 17126 22420 17132 22432
rect 17087 22392 17132 22420
rect 17126 22380 17132 22392
rect 17184 22380 17190 22432
rect 17494 22380 17500 22432
rect 17552 22420 17558 22432
rect 17788 22429 17816 22460
rect 18417 22457 18429 22460
rect 18463 22457 18475 22491
rect 19981 22491 20039 22497
rect 19981 22488 19993 22491
rect 18417 22451 18475 22457
rect 19444 22460 19993 22488
rect 19444 22432 19472 22460
rect 19981 22457 19993 22460
rect 20027 22457 20039 22491
rect 19981 22451 20039 22457
rect 20346 22448 20352 22500
rect 20404 22488 20410 22500
rect 22189 22491 22247 22497
rect 22189 22488 22201 22491
rect 20404 22460 22201 22488
rect 20404 22448 20410 22460
rect 22189 22457 22201 22460
rect 22235 22457 22247 22491
rect 22189 22451 22247 22457
rect 23109 22491 23167 22497
rect 23109 22457 23121 22491
rect 23155 22488 23167 22491
rect 24213 22491 24271 22497
rect 24213 22488 24225 22491
rect 23155 22460 24225 22488
rect 23155 22457 23167 22460
rect 23109 22451 23167 22457
rect 24213 22457 24225 22460
rect 24259 22488 24271 22491
rect 24394 22488 24400 22500
rect 24259 22460 24400 22488
rect 24259 22457 24271 22460
rect 24213 22451 24271 22457
rect 24394 22448 24400 22460
rect 24452 22448 24458 22500
rect 17773 22423 17831 22429
rect 17773 22420 17785 22423
rect 17552 22392 17785 22420
rect 17552 22380 17558 22392
rect 17773 22389 17785 22392
rect 17819 22389 17831 22423
rect 17773 22383 17831 22389
rect 18049 22423 18107 22429
rect 18049 22389 18061 22423
rect 18095 22420 18107 22423
rect 18322 22420 18328 22432
rect 18095 22392 18328 22420
rect 18095 22389 18107 22392
rect 18049 22383 18107 22389
rect 18322 22380 18328 22392
rect 18380 22380 18386 22432
rect 19426 22420 19432 22432
rect 19387 22392 19432 22420
rect 19426 22380 19432 22392
rect 19484 22380 19490 22432
rect 20070 22380 20076 22432
rect 20128 22420 20134 22432
rect 20128 22392 20173 22420
rect 20128 22380 20134 22392
rect 21174 22380 21180 22432
rect 21232 22420 21238 22432
rect 21269 22423 21327 22429
rect 21269 22420 21281 22423
rect 21232 22392 21281 22420
rect 21232 22380 21238 22392
rect 21269 22389 21281 22392
rect 21315 22389 21327 22423
rect 21269 22383 21327 22389
rect 21542 22380 21548 22432
rect 21600 22420 21606 22432
rect 21637 22423 21695 22429
rect 21637 22420 21649 22423
rect 21600 22392 21649 22420
rect 21600 22380 21606 22392
rect 21637 22389 21649 22392
rect 21683 22389 21695 22423
rect 22278 22420 22284 22432
rect 22239 22392 22284 22420
rect 21637 22383 21695 22389
rect 22278 22380 22284 22392
rect 22336 22380 22342 22432
rect 23474 22420 23480 22432
rect 23435 22392 23480 22420
rect 23474 22380 23480 22392
rect 23532 22420 23538 22432
rect 24305 22423 24363 22429
rect 24305 22420 24317 22423
rect 23532 22392 24317 22420
rect 23532 22380 23538 22392
rect 24305 22389 24317 22392
rect 24351 22389 24363 22423
rect 24305 22383 24363 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 4433 22219 4491 22225
rect 4433 22185 4445 22219
rect 4479 22216 4491 22219
rect 4798 22216 4804 22228
rect 4479 22188 4804 22216
rect 4479 22185 4491 22188
rect 4433 22179 4491 22185
rect 4798 22176 4804 22188
rect 4856 22176 4862 22228
rect 13446 22216 13452 22228
rect 13407 22188 13452 22216
rect 13446 22176 13452 22188
rect 13504 22176 13510 22228
rect 13906 22176 13912 22228
rect 13964 22216 13970 22228
rect 14461 22219 14519 22225
rect 14461 22216 14473 22219
rect 13964 22188 14473 22216
rect 13964 22176 13970 22188
rect 14461 22185 14473 22188
rect 14507 22185 14519 22219
rect 14461 22179 14519 22185
rect 15105 22219 15163 22225
rect 15105 22185 15117 22219
rect 15151 22216 15163 22219
rect 16390 22216 16396 22228
rect 15151 22188 16396 22216
rect 15151 22185 15163 22188
rect 15105 22179 15163 22185
rect 16390 22176 16396 22188
rect 16448 22176 16454 22228
rect 20254 22216 20260 22228
rect 16868 22188 20260 22216
rect 5350 22148 5356 22160
rect 5311 22120 5356 22148
rect 5350 22108 5356 22120
rect 5408 22108 5414 22160
rect 9398 22148 9404 22160
rect 8312 22120 9404 22148
rect 1397 22083 1455 22089
rect 1397 22049 1409 22083
rect 1443 22080 1455 22083
rect 2314 22080 2320 22092
rect 1443 22052 2320 22080
rect 1443 22049 1455 22052
rect 1397 22043 1455 22049
rect 2314 22040 2320 22052
rect 2372 22040 2378 22092
rect 4982 22040 4988 22092
rect 5040 22080 5046 22092
rect 7374 22089 7380 22092
rect 5077 22083 5135 22089
rect 5077 22080 5089 22083
rect 5040 22052 5089 22080
rect 5040 22040 5046 22052
rect 5077 22049 5089 22052
rect 5123 22049 5135 22083
rect 7368 22080 7380 22089
rect 7287 22052 7380 22080
rect 5077 22043 5135 22049
rect 7368 22043 7380 22052
rect 7432 22080 7438 22092
rect 8312 22080 8340 22120
rect 9398 22108 9404 22120
rect 9456 22108 9462 22160
rect 10686 22148 10692 22160
rect 9692 22120 10692 22148
rect 7432 22052 8340 22080
rect 9493 22083 9551 22089
rect 7374 22040 7380 22043
rect 7432 22040 7438 22052
rect 9493 22049 9505 22083
rect 9539 22080 9551 22083
rect 9692 22080 9720 22120
rect 10686 22108 10692 22120
rect 10744 22108 10750 22160
rect 11514 22108 11520 22160
rect 11572 22148 11578 22160
rect 12253 22151 12311 22157
rect 12253 22148 12265 22151
rect 11572 22120 12265 22148
rect 11572 22108 11578 22120
rect 12253 22117 12265 22120
rect 12299 22148 12311 22151
rect 13817 22151 13875 22157
rect 13817 22148 13829 22151
rect 12299 22120 12572 22148
rect 13727 22120 13829 22148
rect 12299 22117 12311 22120
rect 12253 22111 12311 22117
rect 9950 22089 9956 22092
rect 9944 22080 9956 22089
rect 9539 22052 9720 22080
rect 9911 22052 9956 22080
rect 9539 22049 9551 22052
rect 9493 22043 9551 22049
rect 9944 22043 9956 22052
rect 9950 22040 9956 22043
rect 10008 22040 10014 22092
rect 11701 22083 11759 22089
rect 11701 22049 11713 22083
rect 11747 22080 11759 22083
rect 11790 22080 11796 22092
rect 11747 22052 11796 22080
rect 11747 22049 11759 22052
rect 11701 22043 11759 22049
rect 11790 22040 11796 22052
rect 11848 22040 11854 22092
rect 12544 22080 12572 22120
rect 13817 22117 13829 22120
rect 13863 22148 13875 22151
rect 13998 22148 14004 22160
rect 13863 22120 14004 22148
rect 13863 22117 13875 22120
rect 13817 22111 13875 22117
rect 12989 22083 13047 22089
rect 12544 22052 12848 22080
rect 12820 22024 12848 22052
rect 12989 22049 13001 22083
rect 13035 22080 13047 22083
rect 13832 22080 13860 22111
rect 13998 22108 14004 22120
rect 14056 22108 14062 22160
rect 15838 22108 15844 22160
rect 15896 22148 15902 22160
rect 16022 22148 16028 22160
rect 15896 22120 16028 22148
rect 15896 22108 15902 22120
rect 16022 22108 16028 22120
rect 16080 22108 16086 22160
rect 16114 22108 16120 22160
rect 16172 22148 16178 22160
rect 16868 22148 16896 22188
rect 20254 22176 20260 22188
rect 20312 22176 20318 22228
rect 20714 22176 20720 22228
rect 20772 22216 20778 22228
rect 21637 22219 21695 22225
rect 21637 22216 21649 22219
rect 20772 22188 21649 22216
rect 20772 22176 20778 22188
rect 21637 22185 21649 22188
rect 21683 22216 21695 22219
rect 22278 22216 22284 22228
rect 21683 22188 22284 22216
rect 21683 22185 21695 22188
rect 21637 22179 21695 22185
rect 22278 22176 22284 22188
rect 22336 22176 22342 22228
rect 23845 22219 23903 22225
rect 23845 22185 23857 22219
rect 23891 22216 23903 22219
rect 23934 22216 23940 22228
rect 23891 22188 23940 22216
rect 23891 22185 23903 22188
rect 23845 22179 23903 22185
rect 23934 22176 23940 22188
rect 23992 22216 23998 22228
rect 23992 22188 24348 22216
rect 23992 22176 23998 22188
rect 16172 22120 16896 22148
rect 17773 22151 17831 22157
rect 16172 22108 16178 22120
rect 17773 22117 17785 22151
rect 17819 22148 17831 22151
rect 17862 22148 17868 22160
rect 17819 22120 17868 22148
rect 17819 22117 17831 22120
rect 17773 22111 17831 22117
rect 13035 22052 13860 22080
rect 13035 22049 13047 22052
rect 12989 22043 13047 22049
rect 14826 22040 14832 22092
rect 14884 22080 14890 22092
rect 16292 22083 16350 22089
rect 14884 22052 16068 22080
rect 14884 22040 14890 22052
rect 7098 22012 7104 22024
rect 7059 21984 7104 22012
rect 7098 21972 7104 21984
rect 7156 21972 7162 22024
rect 8938 21972 8944 22024
rect 8996 22012 9002 22024
rect 9677 22015 9735 22021
rect 9677 22012 9689 22015
rect 8996 21984 9689 22012
rect 8996 21972 9002 21984
rect 9677 21981 9689 21984
rect 9723 21981 9735 22015
rect 12342 22012 12348 22024
rect 12303 21984 12348 22012
rect 9677 21975 9735 21981
rect 12342 21972 12348 21984
rect 12400 21972 12406 22024
rect 12529 22015 12587 22021
rect 12529 21981 12541 22015
rect 12575 22012 12587 22015
rect 12710 22012 12716 22024
rect 12575 21984 12716 22012
rect 12575 21981 12587 21984
rect 12529 21975 12587 21981
rect 12710 21972 12716 21984
rect 12768 21972 12774 22024
rect 12802 21972 12808 22024
rect 12860 21972 12866 22024
rect 13906 22012 13912 22024
rect 13867 21984 13912 22012
rect 13906 21972 13912 21984
rect 13964 21972 13970 22024
rect 14093 22015 14151 22021
rect 14093 21981 14105 22015
rect 14139 22012 14151 22015
rect 14277 22015 14335 22021
rect 14277 22012 14289 22015
rect 14139 21984 14289 22012
rect 14139 21981 14151 21984
rect 14093 21975 14151 21981
rect 14277 21981 14289 21984
rect 14323 22012 14335 22015
rect 14550 22012 14556 22024
rect 14323 21984 14556 22012
rect 14323 21981 14335 21984
rect 14277 21975 14335 21981
rect 14550 21972 14556 21984
rect 14608 21972 14614 22024
rect 15565 22015 15623 22021
rect 15565 21981 15577 22015
rect 15611 22012 15623 22015
rect 15838 22012 15844 22024
rect 15611 21984 15844 22012
rect 15611 21981 15623 21984
rect 15565 21975 15623 21981
rect 15838 21972 15844 21984
rect 15896 21972 15902 22024
rect 16040 22021 16068 22052
rect 16292 22049 16304 22083
rect 16338 22080 16350 22083
rect 16758 22080 16764 22092
rect 16338 22052 16764 22080
rect 16338 22049 16350 22052
rect 16292 22043 16350 22049
rect 16758 22040 16764 22052
rect 16816 22040 16822 22092
rect 16850 22040 16856 22092
rect 16908 22080 16914 22092
rect 17678 22080 17684 22092
rect 16908 22052 17684 22080
rect 16908 22040 16914 22052
rect 17678 22040 17684 22052
rect 17736 22040 17742 22092
rect 16025 22015 16083 22021
rect 16025 21981 16037 22015
rect 16071 21981 16083 22015
rect 16025 21975 16083 21981
rect 1394 21904 1400 21956
rect 1452 21944 1458 21956
rect 1581 21947 1639 21953
rect 1581 21944 1593 21947
rect 1452 21916 1593 21944
rect 1452 21904 1458 21916
rect 1581 21913 1593 21916
rect 1627 21913 1639 21947
rect 1581 21907 1639 21913
rect 8110 21904 8116 21956
rect 8168 21944 8174 21956
rect 8481 21947 8539 21953
rect 8481 21944 8493 21947
rect 8168 21916 8493 21944
rect 8168 21904 8174 21916
rect 8481 21913 8493 21916
rect 8527 21913 8539 21947
rect 8481 21907 8539 21913
rect 11146 21904 11152 21956
rect 11204 21944 11210 21956
rect 11885 21947 11943 21953
rect 11885 21944 11897 21947
rect 11204 21916 11897 21944
rect 11204 21904 11210 21916
rect 11885 21913 11897 21916
rect 11931 21913 11943 21947
rect 11885 21907 11943 21913
rect 12066 21904 12072 21956
rect 12124 21944 12130 21956
rect 14642 21944 14648 21956
rect 12124 21916 14648 21944
rect 12124 21904 12130 21916
rect 14642 21904 14648 21916
rect 14700 21904 14706 21956
rect 17678 21904 17684 21956
rect 17736 21944 17742 21956
rect 17788 21944 17816 22111
rect 17862 22108 17868 22120
rect 17920 22108 17926 22160
rect 18414 22108 18420 22160
rect 18472 22148 18478 22160
rect 18598 22148 18604 22160
rect 18472 22120 18604 22148
rect 18472 22108 18478 22120
rect 18598 22108 18604 22120
rect 18656 22108 18662 22160
rect 21542 22108 21548 22160
rect 21600 22148 21606 22160
rect 21726 22148 21732 22160
rect 21600 22120 21732 22148
rect 21600 22108 21606 22120
rect 21726 22108 21732 22120
rect 21784 22108 21790 22160
rect 21818 22108 21824 22160
rect 21876 22148 21882 22160
rect 22094 22148 22100 22160
rect 21876 22120 22100 22148
rect 21876 22108 21882 22120
rect 22094 22108 22100 22120
rect 22152 22108 22158 22160
rect 23661 22151 23719 22157
rect 23661 22148 23673 22151
rect 22296 22120 23673 22148
rect 17972 22052 18828 22080
rect 17862 21972 17868 22024
rect 17920 22012 17926 22024
rect 17972 22012 18000 22052
rect 18690 22012 18696 22024
rect 17920 21984 18000 22012
rect 18651 21984 18696 22012
rect 17920 21972 17926 21984
rect 18690 21972 18696 21984
rect 18748 21972 18754 22024
rect 18800 22021 18828 22052
rect 19518 22040 19524 22092
rect 19576 22080 19582 22092
rect 20622 22080 20628 22092
rect 19576 22052 20628 22080
rect 19576 22040 19582 22052
rect 20622 22040 20628 22052
rect 20680 22040 20686 22092
rect 20717 22083 20775 22089
rect 20717 22049 20729 22083
rect 20763 22080 20775 22083
rect 22002 22080 22008 22092
rect 20763 22052 22008 22080
rect 20763 22049 20775 22052
rect 20717 22043 20775 22049
rect 22002 22040 22008 22052
rect 22060 22040 22066 22092
rect 22296 22024 22324 22120
rect 23661 22117 23673 22120
rect 23707 22148 23719 22151
rect 24118 22148 24124 22160
rect 23707 22120 24124 22148
rect 23707 22117 23719 22120
rect 23661 22111 23719 22117
rect 24118 22108 24124 22120
rect 24176 22108 24182 22160
rect 22557 22083 22615 22089
rect 22557 22049 22569 22083
rect 22603 22080 22615 22083
rect 23198 22080 23204 22092
rect 22603 22052 23204 22080
rect 22603 22049 22615 22052
rect 22557 22043 22615 22049
rect 23198 22040 23204 22052
rect 23256 22080 23262 22092
rect 23385 22083 23443 22089
rect 23385 22080 23397 22083
rect 23256 22052 23397 22080
rect 23256 22040 23262 22052
rect 23385 22049 23397 22052
rect 23431 22080 23443 22083
rect 23934 22080 23940 22092
rect 23431 22052 23940 22080
rect 23431 22049 23443 22052
rect 23385 22043 23443 22049
rect 23934 22040 23940 22052
rect 23992 22040 23998 22092
rect 24213 22083 24271 22089
rect 24213 22049 24225 22083
rect 24259 22049 24271 22083
rect 24320 22080 24348 22188
rect 24320 22052 24624 22080
rect 24213 22043 24271 22049
rect 18785 22015 18843 22021
rect 18785 21981 18797 22015
rect 18831 21981 18843 22015
rect 18785 21975 18843 21981
rect 19705 22015 19763 22021
rect 19705 21981 19717 22015
rect 19751 22012 19763 22015
rect 20070 22012 20076 22024
rect 19751 21984 20076 22012
rect 19751 21981 19763 21984
rect 19705 21975 19763 21981
rect 20070 21972 20076 21984
rect 20128 22012 20134 22024
rect 20438 22012 20444 22024
rect 20128 21984 20444 22012
rect 20128 21972 20134 21984
rect 20438 21972 20444 21984
rect 20496 21972 20502 22024
rect 20990 21972 20996 22024
rect 21048 22012 21054 22024
rect 21177 22015 21235 22021
rect 21177 22012 21189 22015
rect 21048 21984 21189 22012
rect 21048 21972 21054 21984
rect 21177 21981 21189 21984
rect 21223 22012 21235 22015
rect 22097 22015 22155 22021
rect 22097 22012 22109 22015
rect 21223 21984 22109 22012
rect 21223 21981 21235 21984
rect 21177 21975 21235 21981
rect 22097 21981 22109 21984
rect 22143 21981 22155 22015
rect 22278 22012 22284 22024
rect 22239 21984 22284 22012
rect 22097 21975 22155 21981
rect 22278 21972 22284 21984
rect 22336 21972 22342 22024
rect 23474 21972 23480 22024
rect 23532 22012 23538 22024
rect 24228 22012 24256 22043
rect 23532 21984 24256 22012
rect 24305 22015 24363 22021
rect 23532 21972 23538 21984
rect 24305 21981 24317 22015
rect 24351 21981 24363 22015
rect 24305 21975 24363 21981
rect 18230 21944 18236 21956
rect 17736 21916 17816 21944
rect 18191 21916 18236 21944
rect 17736 21904 17742 21916
rect 18230 21904 18236 21916
rect 18288 21904 18294 21956
rect 18966 21904 18972 21956
rect 19024 21944 19030 21956
rect 21082 21944 21088 21956
rect 19024 21916 21088 21944
rect 19024 21904 19030 21916
rect 21082 21904 21088 21916
rect 21140 21904 21146 21956
rect 21545 21947 21603 21953
rect 21545 21913 21557 21947
rect 21591 21944 21603 21947
rect 22557 21947 22615 21953
rect 22557 21944 22569 21947
rect 21591 21916 22569 21944
rect 21591 21913 21603 21916
rect 21545 21907 21603 21913
rect 22557 21913 22569 21916
rect 22603 21913 22615 21947
rect 22557 21907 22615 21913
rect 23198 21904 23204 21956
rect 23256 21944 23262 21956
rect 24320 21944 24348 21975
rect 24394 21972 24400 22024
rect 24452 22012 24458 22024
rect 24596 22012 24624 22052
rect 24854 22040 24860 22092
rect 24912 22080 24918 22092
rect 25593 22083 25651 22089
rect 25593 22080 25605 22083
rect 24912 22052 25605 22080
rect 24912 22040 24918 22052
rect 25593 22049 25605 22052
rect 25639 22049 25651 22083
rect 25593 22043 25651 22049
rect 25225 22015 25283 22021
rect 25225 22012 25237 22015
rect 24452 21984 24497 22012
rect 24596 21984 25237 22012
rect 24452 21972 24458 21984
rect 25225 21981 25237 21984
rect 25271 21981 25283 22015
rect 25225 21975 25283 21981
rect 23256 21916 24348 21944
rect 23256 21904 23262 21916
rect 5905 21879 5963 21885
rect 5905 21845 5917 21879
rect 5951 21876 5963 21879
rect 6270 21876 6276 21888
rect 5951 21848 6276 21876
rect 5951 21845 5963 21848
rect 5905 21839 5963 21845
rect 6270 21836 6276 21848
rect 6328 21836 6334 21888
rect 6546 21876 6552 21888
rect 6507 21848 6552 21876
rect 6546 21836 6552 21848
rect 6604 21836 6610 21888
rect 6914 21876 6920 21888
rect 6875 21848 6920 21876
rect 6914 21836 6920 21848
rect 6972 21836 6978 21888
rect 9030 21876 9036 21888
rect 8991 21848 9036 21876
rect 9030 21836 9036 21848
rect 9088 21836 9094 21888
rect 9122 21836 9128 21888
rect 9180 21876 9186 21888
rect 9582 21876 9588 21888
rect 9180 21848 9588 21876
rect 9180 21836 9186 21848
rect 9582 21836 9588 21848
rect 9640 21836 9646 21888
rect 10042 21836 10048 21888
rect 10100 21876 10106 21888
rect 11057 21879 11115 21885
rect 11057 21876 11069 21879
rect 10100 21848 11069 21876
rect 10100 21836 10106 21848
rect 11057 21845 11069 21848
rect 11103 21845 11115 21879
rect 13262 21876 13268 21888
rect 13223 21848 13268 21876
rect 11057 21839 11115 21845
rect 13262 21836 13268 21848
rect 13320 21876 13326 21888
rect 14277 21879 14335 21885
rect 14277 21876 14289 21879
rect 13320 21848 14289 21876
rect 13320 21836 13326 21848
rect 14277 21845 14289 21848
rect 14323 21845 14335 21879
rect 15930 21876 15936 21888
rect 15843 21848 15936 21876
rect 14277 21839 14335 21845
rect 15930 21836 15936 21848
rect 15988 21876 15994 21888
rect 17405 21879 17463 21885
rect 17405 21876 17417 21879
rect 15988 21848 17417 21876
rect 15988 21836 15994 21848
rect 17405 21845 17417 21848
rect 17451 21845 17463 21879
rect 17405 21839 17463 21845
rect 18046 21836 18052 21888
rect 18104 21876 18110 21888
rect 18141 21879 18199 21885
rect 18141 21876 18153 21879
rect 18104 21848 18153 21876
rect 18104 21836 18110 21848
rect 18141 21845 18153 21848
rect 18187 21876 18199 21879
rect 18414 21876 18420 21888
rect 18187 21848 18420 21876
rect 18187 21845 18199 21848
rect 18141 21839 18199 21845
rect 18414 21836 18420 21848
rect 18472 21836 18478 21888
rect 18874 21836 18880 21888
rect 18932 21876 18938 21888
rect 19242 21876 19248 21888
rect 18932 21848 19248 21876
rect 18932 21836 18938 21848
rect 19242 21836 19248 21848
rect 19300 21836 19306 21888
rect 20349 21879 20407 21885
rect 20349 21845 20361 21879
rect 20395 21876 20407 21879
rect 20898 21876 20904 21888
rect 20395 21848 20904 21876
rect 20395 21845 20407 21848
rect 20349 21839 20407 21845
rect 20898 21836 20904 21848
rect 20956 21836 20962 21888
rect 22462 21836 22468 21888
rect 22520 21876 22526 21888
rect 22649 21879 22707 21885
rect 22649 21876 22661 21879
rect 22520 21848 22661 21876
rect 22520 21836 22526 21848
rect 22649 21845 22661 21848
rect 22695 21845 22707 21879
rect 22649 21839 22707 21845
rect 24210 21836 24216 21888
rect 24268 21876 24274 21888
rect 24670 21876 24676 21888
rect 24268 21848 24676 21876
rect 24268 21836 24274 21848
rect 24670 21836 24676 21848
rect 24728 21876 24734 21888
rect 24857 21879 24915 21885
rect 24857 21876 24869 21879
rect 24728 21848 24869 21876
rect 24728 21836 24734 21848
rect 24857 21845 24869 21848
rect 24903 21845 24915 21879
rect 24857 21839 24915 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1486 21632 1492 21684
rect 1544 21672 1550 21684
rect 1581 21675 1639 21681
rect 1581 21672 1593 21675
rect 1544 21644 1593 21672
rect 1544 21632 1550 21644
rect 1581 21641 1593 21644
rect 1627 21641 1639 21675
rect 1581 21635 1639 21641
rect 3510 21632 3516 21684
rect 3568 21672 3574 21684
rect 3973 21675 4031 21681
rect 3973 21672 3985 21675
rect 3568 21644 3985 21672
rect 3568 21632 3574 21644
rect 3973 21641 3985 21644
rect 4019 21672 4031 21675
rect 4798 21672 4804 21684
rect 4019 21644 4804 21672
rect 4019 21641 4031 21644
rect 3973 21635 4031 21641
rect 4798 21632 4804 21644
rect 4856 21632 4862 21684
rect 4890 21632 4896 21684
rect 4948 21672 4954 21684
rect 4985 21675 5043 21681
rect 4985 21672 4997 21675
rect 4948 21644 4997 21672
rect 4948 21632 4954 21644
rect 4985 21641 4997 21644
rect 5031 21641 5043 21675
rect 6638 21672 6644 21684
rect 6599 21644 6644 21672
rect 4985 21635 5043 21641
rect 6638 21632 6644 21644
rect 6696 21632 6702 21684
rect 7101 21675 7159 21681
rect 7101 21641 7113 21675
rect 7147 21672 7159 21675
rect 7374 21672 7380 21684
rect 7147 21644 7380 21672
rect 7147 21641 7159 21644
rect 7101 21635 7159 21641
rect 7374 21632 7380 21644
rect 7432 21632 7438 21684
rect 10686 21632 10692 21684
rect 10744 21672 10750 21684
rect 10781 21675 10839 21681
rect 10781 21672 10793 21675
rect 10744 21644 10793 21672
rect 10744 21632 10750 21644
rect 10781 21641 10793 21644
rect 10827 21641 10839 21675
rect 10781 21635 10839 21641
rect 12713 21675 12771 21681
rect 12713 21641 12725 21675
rect 12759 21672 12771 21675
rect 12802 21672 12808 21684
rect 12759 21644 12808 21672
rect 12759 21641 12771 21644
rect 12713 21635 12771 21641
rect 12802 21632 12808 21644
rect 12860 21632 12866 21684
rect 14090 21632 14096 21684
rect 14148 21672 14154 21684
rect 14737 21675 14795 21681
rect 14737 21672 14749 21675
rect 14148 21644 14749 21672
rect 14148 21632 14154 21644
rect 14737 21641 14749 21644
rect 14783 21672 14795 21675
rect 15381 21675 15439 21681
rect 15381 21672 15393 21675
rect 14783 21644 15393 21672
rect 14783 21641 14795 21644
rect 14737 21635 14795 21641
rect 15381 21641 15393 21644
rect 15427 21641 15439 21675
rect 15381 21635 15439 21641
rect 3786 21564 3792 21616
rect 3844 21604 3850 21616
rect 4617 21607 4675 21613
rect 4617 21604 4629 21607
rect 3844 21576 4629 21604
rect 3844 21564 3850 21576
rect 4617 21573 4629 21576
rect 4663 21604 4675 21607
rect 5534 21604 5540 21616
rect 4663 21576 5540 21604
rect 4663 21573 4675 21576
rect 4617 21567 4675 21573
rect 5534 21564 5540 21576
rect 5592 21564 5598 21616
rect 2038 21536 2044 21548
rect 1412 21508 2044 21536
rect 1412 21477 1440 21508
rect 2038 21496 2044 21508
rect 2096 21496 2102 21548
rect 4341 21539 4399 21545
rect 4341 21505 4353 21539
rect 4387 21536 4399 21539
rect 5810 21536 5816 21548
rect 4387 21508 5816 21536
rect 4387 21505 4399 21508
rect 4341 21499 4399 21505
rect 5810 21496 5816 21508
rect 5868 21536 5874 21548
rect 6656 21536 6684 21632
rect 5868 21508 6316 21536
rect 6656 21508 7328 21536
rect 5868 21496 5874 21508
rect 1397 21471 1455 21477
rect 1397 21437 1409 21471
rect 1443 21437 1455 21471
rect 1397 21431 1455 21437
rect 2501 21471 2559 21477
rect 2501 21437 2513 21471
rect 2547 21468 2559 21471
rect 3050 21468 3056 21480
rect 2547 21440 3056 21468
rect 2547 21437 2559 21440
rect 2501 21431 2559 21437
rect 3050 21428 3056 21440
rect 3108 21428 3114 21480
rect 4982 21428 4988 21480
rect 5040 21468 5046 21480
rect 6181 21471 6239 21477
rect 6181 21468 6193 21471
rect 5040 21440 6193 21468
rect 5040 21428 5046 21440
rect 6181 21437 6193 21440
rect 6227 21437 6239 21471
rect 6288 21468 6316 21508
rect 6288 21440 6960 21468
rect 6181 21431 6239 21437
rect 4890 21360 4896 21412
rect 4948 21400 4954 21412
rect 5629 21403 5687 21409
rect 5629 21400 5641 21403
rect 4948 21372 5641 21400
rect 4948 21360 4954 21372
rect 5629 21369 5641 21372
rect 5675 21400 5687 21403
rect 6822 21400 6828 21412
rect 5675 21372 6828 21400
rect 5675 21369 5687 21372
rect 5629 21363 5687 21369
rect 6822 21360 6828 21372
rect 6880 21360 6886 21412
rect 2314 21332 2320 21344
rect 2275 21304 2320 21332
rect 2314 21292 2320 21304
rect 2372 21292 2378 21344
rect 2685 21335 2743 21341
rect 2685 21301 2697 21335
rect 2731 21332 2743 21335
rect 2774 21332 2780 21344
rect 2731 21304 2780 21332
rect 2731 21301 2743 21304
rect 2685 21295 2743 21301
rect 2774 21292 2780 21304
rect 2832 21292 2838 21344
rect 5166 21332 5172 21344
rect 5127 21304 5172 21332
rect 5166 21292 5172 21304
rect 5224 21292 5230 21344
rect 5534 21332 5540 21344
rect 5495 21304 5540 21332
rect 5534 21292 5540 21304
rect 5592 21292 5598 21344
rect 6932 21332 6960 21440
rect 7098 21428 7104 21480
rect 7156 21468 7162 21480
rect 7193 21471 7251 21477
rect 7193 21468 7205 21471
rect 7156 21440 7205 21468
rect 7156 21428 7162 21440
rect 7193 21437 7205 21440
rect 7239 21437 7251 21471
rect 7300 21468 7328 21508
rect 8938 21496 8944 21548
rect 8996 21496 9002 21548
rect 11977 21539 12035 21545
rect 11977 21505 11989 21539
rect 12023 21536 12035 21539
rect 12342 21536 12348 21548
rect 12023 21508 12348 21536
rect 12023 21505 12035 21508
rect 11977 21499 12035 21505
rect 12342 21496 12348 21508
rect 12400 21496 12406 21548
rect 15396 21536 15424 21635
rect 18598 21632 18604 21684
rect 18656 21672 18662 21684
rect 19061 21675 19119 21681
rect 19061 21672 19073 21675
rect 18656 21644 19073 21672
rect 18656 21632 18662 21644
rect 19061 21641 19073 21644
rect 19107 21641 19119 21675
rect 19061 21635 19119 21641
rect 20070 21632 20076 21684
rect 20128 21672 20134 21684
rect 20257 21675 20315 21681
rect 20257 21672 20269 21675
rect 20128 21644 20269 21672
rect 20128 21632 20134 21644
rect 20257 21641 20269 21644
rect 20303 21641 20315 21675
rect 20257 21635 20315 21641
rect 16758 21564 16764 21616
rect 16816 21604 16822 21616
rect 16945 21607 17003 21613
rect 16945 21604 16957 21607
rect 16816 21576 16957 21604
rect 16816 21564 16822 21576
rect 16945 21573 16957 21576
rect 16991 21573 17003 21607
rect 16945 21567 17003 21573
rect 16960 21536 16988 21567
rect 17126 21564 17132 21616
rect 17184 21604 17190 21616
rect 17681 21607 17739 21613
rect 17681 21604 17693 21607
rect 17184 21576 17693 21604
rect 17184 21564 17190 21576
rect 17681 21573 17693 21576
rect 17727 21604 17739 21607
rect 17773 21607 17831 21613
rect 17773 21604 17785 21607
rect 17727 21576 17785 21604
rect 17727 21573 17739 21576
rect 17681 21567 17739 21573
rect 17773 21573 17785 21576
rect 17819 21573 17831 21607
rect 17773 21567 17831 21573
rect 18690 21564 18696 21616
rect 18748 21604 18754 21616
rect 19797 21607 19855 21613
rect 19797 21604 19809 21607
rect 18748 21576 19809 21604
rect 18748 21564 18754 21576
rect 19797 21573 19809 21576
rect 19843 21573 19855 21607
rect 19797 21567 19855 21573
rect 18601 21539 18659 21545
rect 18601 21536 18613 21539
rect 15396 21508 15700 21536
rect 16960 21508 18613 21536
rect 7449 21471 7507 21477
rect 7449 21468 7461 21471
rect 7300 21440 7461 21468
rect 7193 21431 7251 21437
rect 7449 21437 7461 21440
rect 7495 21437 7507 21471
rect 7449 21431 7507 21437
rect 7208 21400 7236 21431
rect 8202 21428 8208 21480
rect 8260 21468 8266 21480
rect 8956 21468 8984 21496
rect 9401 21471 9459 21477
rect 9401 21468 9413 21471
rect 8260 21440 9413 21468
rect 8260 21428 8266 21440
rect 9401 21437 9413 21440
rect 9447 21468 9459 21471
rect 10686 21468 10692 21480
rect 9447 21440 10692 21468
rect 9447 21437 9459 21440
rect 9401 21431 9459 21437
rect 10686 21428 10692 21440
rect 10744 21428 10750 21480
rect 12986 21428 12992 21480
rect 13044 21468 13050 21480
rect 13357 21471 13415 21477
rect 13357 21468 13369 21471
rect 13044 21440 13369 21468
rect 13044 21428 13050 21440
rect 13357 21437 13369 21440
rect 13403 21468 13415 21471
rect 14826 21468 14832 21480
rect 13403 21440 14832 21468
rect 13403 21437 13415 21440
rect 13357 21431 13415 21437
rect 14826 21428 14832 21440
rect 14884 21468 14890 21480
rect 15565 21471 15623 21477
rect 15565 21468 15577 21471
rect 14884 21440 15577 21468
rect 14884 21428 14890 21440
rect 15565 21437 15577 21440
rect 15611 21437 15623 21471
rect 15672 21468 15700 21508
rect 18601 21505 18613 21508
rect 18647 21536 18659 21539
rect 18874 21536 18880 21548
rect 18647 21508 18880 21536
rect 18647 21505 18659 21508
rect 18601 21499 18659 21505
rect 18874 21496 18880 21508
rect 18932 21536 18938 21548
rect 19429 21539 19487 21545
rect 19429 21536 19441 21539
rect 18932 21508 19441 21536
rect 18932 21496 18938 21508
rect 19429 21505 19441 21508
rect 19475 21505 19487 21539
rect 19429 21499 19487 21505
rect 15821 21471 15879 21477
rect 15821 21468 15833 21471
rect 15672 21440 15833 21468
rect 15565 21431 15623 21437
rect 15821 21437 15833 21440
rect 15867 21437 15879 21471
rect 15821 21431 15879 21437
rect 17681 21471 17739 21477
rect 17681 21437 17693 21471
rect 17727 21468 17739 21471
rect 18509 21471 18567 21477
rect 18509 21468 18521 21471
rect 17727 21440 18521 21468
rect 17727 21437 17739 21440
rect 17681 21431 17739 21437
rect 18509 21437 18521 21440
rect 18555 21468 18567 21471
rect 19058 21468 19064 21480
rect 18555 21440 19064 21468
rect 18555 21437 18567 21440
rect 18509 21431 18567 21437
rect 19058 21428 19064 21440
rect 19116 21428 19122 21480
rect 20272 21468 20300 21635
rect 20346 21632 20352 21684
rect 20404 21672 20410 21684
rect 20441 21675 20499 21681
rect 20441 21672 20453 21675
rect 20404 21644 20453 21672
rect 20404 21632 20410 21644
rect 20441 21641 20453 21644
rect 20487 21641 20499 21675
rect 20441 21635 20499 21641
rect 21634 21632 21640 21684
rect 21692 21672 21698 21684
rect 21821 21675 21879 21681
rect 21821 21672 21833 21675
rect 21692 21644 21833 21672
rect 21692 21632 21698 21644
rect 21821 21641 21833 21644
rect 21867 21641 21879 21675
rect 22002 21672 22008 21684
rect 21963 21644 22008 21672
rect 21821 21635 21879 21641
rect 22002 21632 22008 21644
rect 22060 21632 22066 21684
rect 22094 21632 22100 21684
rect 22152 21672 22158 21684
rect 23017 21675 23075 21681
rect 23017 21672 23029 21675
rect 22152 21644 23029 21672
rect 22152 21632 22158 21644
rect 23017 21641 23029 21644
rect 23063 21672 23075 21675
rect 23198 21672 23204 21684
rect 23063 21644 23204 21672
rect 23063 21641 23075 21644
rect 23017 21635 23075 21641
rect 23198 21632 23204 21644
rect 23256 21632 23262 21684
rect 23750 21632 23756 21684
rect 23808 21672 23814 21684
rect 24670 21672 24676 21684
rect 23808 21644 24676 21672
rect 23808 21632 23814 21644
rect 24670 21632 24676 21644
rect 24728 21632 24734 21684
rect 25593 21675 25651 21681
rect 25593 21641 25605 21675
rect 25639 21672 25651 21675
rect 25682 21672 25688 21684
rect 25639 21644 25688 21672
rect 25639 21641 25651 21644
rect 25593 21635 25651 21641
rect 25682 21632 25688 21644
rect 25740 21632 25746 21684
rect 22278 21604 22284 21616
rect 21100 21576 22284 21604
rect 20898 21536 20904 21548
rect 20859 21508 20904 21536
rect 20898 21496 20904 21508
rect 20956 21496 20962 21548
rect 21100 21545 21128 21576
rect 22278 21564 22284 21576
rect 22336 21564 22342 21616
rect 21085 21539 21143 21545
rect 21085 21505 21097 21539
rect 21131 21505 21143 21539
rect 21085 21499 21143 21505
rect 21545 21539 21603 21545
rect 21545 21505 21557 21539
rect 21591 21536 21603 21539
rect 22370 21536 22376 21548
rect 21591 21508 22376 21536
rect 21591 21505 21603 21508
rect 21545 21499 21603 21505
rect 22370 21496 22376 21508
rect 22428 21536 22434 21548
rect 22557 21539 22615 21545
rect 22557 21536 22569 21539
rect 22428 21508 22569 21536
rect 22428 21496 22434 21508
rect 22557 21505 22569 21508
rect 22603 21505 22615 21539
rect 22557 21499 22615 21505
rect 23382 21496 23388 21548
rect 23440 21536 23446 21548
rect 24489 21539 24547 21545
rect 24489 21536 24501 21539
rect 23440 21508 24501 21536
rect 23440 21496 23446 21508
rect 24489 21505 24501 21508
rect 24535 21536 24547 21539
rect 25038 21536 25044 21548
rect 24535 21508 25044 21536
rect 24535 21505 24547 21508
rect 24489 21499 24547 21505
rect 25038 21496 25044 21508
rect 25096 21496 25102 21548
rect 20809 21471 20867 21477
rect 20809 21468 20821 21471
rect 20272 21440 20821 21468
rect 20809 21437 20821 21440
rect 20855 21437 20867 21471
rect 20916 21468 20944 21496
rect 22002 21468 22008 21480
rect 20916 21440 22008 21468
rect 20809 21431 20867 21437
rect 22002 21428 22008 21440
rect 22060 21428 22066 21480
rect 22094 21428 22100 21480
rect 22152 21468 22158 21480
rect 22465 21471 22523 21477
rect 22465 21468 22477 21471
rect 22152 21440 22477 21468
rect 22152 21428 22158 21440
rect 22465 21437 22477 21440
rect 22511 21437 22523 21471
rect 24210 21468 24216 21480
rect 24171 21440 24216 21468
rect 22465 21431 22523 21437
rect 24210 21428 24216 21440
rect 24268 21428 24274 21480
rect 25222 21428 25228 21480
rect 25280 21468 25286 21480
rect 25409 21471 25467 21477
rect 25409 21468 25421 21471
rect 25280 21440 25421 21468
rect 25280 21428 25286 21440
rect 25409 21437 25421 21440
rect 25455 21468 25467 21471
rect 25961 21471 26019 21477
rect 25961 21468 25973 21471
rect 25455 21440 25973 21468
rect 25455 21437 25467 21440
rect 25409 21431 25467 21437
rect 25961 21437 25973 21440
rect 26007 21437 26019 21471
rect 25961 21431 26019 21437
rect 7208 21372 8892 21400
rect 8864 21344 8892 21372
rect 9490 21360 9496 21412
rect 9548 21400 9554 21412
rect 9646 21403 9704 21409
rect 9646 21400 9658 21403
rect 9548 21372 9658 21400
rect 9548 21360 9554 21372
rect 9646 21369 9658 21372
rect 9692 21400 9704 21403
rect 10042 21400 10048 21412
rect 9692 21372 10048 21400
rect 9692 21369 9704 21372
rect 9646 21363 9704 21369
rect 10042 21360 10048 21372
rect 10100 21360 10106 21412
rect 13624 21403 13682 21409
rect 13624 21369 13636 21403
rect 13670 21400 13682 21403
rect 13722 21400 13728 21412
rect 13670 21372 13728 21400
rect 13670 21369 13682 21372
rect 13624 21363 13682 21369
rect 13722 21360 13728 21372
rect 13780 21360 13786 21412
rect 13906 21360 13912 21412
rect 13964 21400 13970 21412
rect 15013 21403 15071 21409
rect 15013 21400 15025 21403
rect 13964 21372 15025 21400
rect 13964 21360 13970 21372
rect 15013 21369 15025 21372
rect 15059 21369 15071 21403
rect 15013 21363 15071 21369
rect 16758 21360 16764 21412
rect 16816 21400 16822 21412
rect 17494 21400 17500 21412
rect 16816 21372 17500 21400
rect 16816 21360 16822 21372
rect 17494 21360 17500 21372
rect 17552 21360 17558 21412
rect 24305 21403 24363 21409
rect 24305 21369 24317 21403
rect 24351 21400 24363 21403
rect 24351 21372 25360 21400
rect 24351 21369 24363 21372
rect 24305 21363 24363 21369
rect 7650 21332 7656 21344
rect 6932 21304 7656 21332
rect 7650 21292 7656 21304
rect 7708 21332 7714 21344
rect 8573 21335 8631 21341
rect 8573 21332 8585 21335
rect 7708 21304 8585 21332
rect 7708 21292 7714 21304
rect 8573 21301 8585 21304
rect 8619 21301 8631 21335
rect 8846 21332 8852 21344
rect 8807 21304 8852 21332
rect 8573 21295 8631 21301
rect 8846 21292 8852 21304
rect 8904 21292 8910 21344
rect 9309 21335 9367 21341
rect 9309 21301 9321 21335
rect 9355 21332 9367 21335
rect 9398 21332 9404 21344
rect 9355 21304 9404 21332
rect 9355 21301 9367 21304
rect 9309 21295 9367 21301
rect 9398 21292 9404 21304
rect 9456 21332 9462 21344
rect 9950 21332 9956 21344
rect 9456 21304 9956 21332
rect 9456 21292 9462 21304
rect 9950 21292 9956 21304
rect 10008 21292 10014 21344
rect 11054 21332 11060 21344
rect 11015 21304 11060 21332
rect 11054 21292 11060 21304
rect 11112 21292 11118 21344
rect 11238 21292 11244 21344
rect 11296 21332 11302 21344
rect 11517 21335 11575 21341
rect 11517 21332 11529 21335
rect 11296 21304 11529 21332
rect 11296 21292 11302 21304
rect 11517 21301 11529 21304
rect 11563 21301 11575 21335
rect 13262 21332 13268 21344
rect 13223 21304 13268 21332
rect 11517 21295 11575 21301
rect 13262 21292 13268 21304
rect 13320 21292 13326 21344
rect 14274 21292 14280 21344
rect 14332 21332 14338 21344
rect 14550 21332 14556 21344
rect 14332 21304 14556 21332
rect 14332 21292 14338 21304
rect 14550 21292 14556 21304
rect 14608 21292 14614 21344
rect 16666 21292 16672 21344
rect 16724 21332 16730 21344
rect 17126 21332 17132 21344
rect 16724 21304 17132 21332
rect 16724 21292 16730 21304
rect 17126 21292 17132 21304
rect 17184 21332 17190 21344
rect 17405 21335 17463 21341
rect 17405 21332 17417 21335
rect 17184 21304 17417 21332
rect 17184 21292 17190 21304
rect 17405 21301 17417 21304
rect 17451 21332 17463 21335
rect 17862 21332 17868 21344
rect 17451 21304 17868 21332
rect 17451 21301 17463 21304
rect 17405 21295 17463 21301
rect 17862 21292 17868 21304
rect 17920 21292 17926 21344
rect 18046 21332 18052 21344
rect 18007 21304 18052 21332
rect 18046 21292 18052 21304
rect 18104 21292 18110 21344
rect 18414 21332 18420 21344
rect 18375 21304 18420 21332
rect 18414 21292 18420 21304
rect 18472 21292 18478 21344
rect 22373 21335 22431 21341
rect 22373 21301 22385 21335
rect 22419 21332 22431 21335
rect 22738 21332 22744 21344
rect 22419 21304 22744 21332
rect 22419 21301 22431 21304
rect 22373 21295 22431 21301
rect 22738 21292 22744 21304
rect 22796 21292 22802 21344
rect 23474 21332 23480 21344
rect 23435 21304 23480 21332
rect 23474 21292 23480 21304
rect 23532 21292 23538 21344
rect 23845 21335 23903 21341
rect 23845 21301 23857 21335
rect 23891 21332 23903 21335
rect 23934 21332 23940 21344
rect 23891 21304 23940 21332
rect 23891 21301 23903 21304
rect 23845 21295 23903 21301
rect 23934 21292 23940 21304
rect 23992 21292 23998 21344
rect 24949 21335 25007 21341
rect 24949 21301 24961 21335
rect 24995 21332 25007 21335
rect 25038 21332 25044 21344
rect 24995 21304 25044 21332
rect 24995 21301 25007 21304
rect 24949 21295 25007 21301
rect 25038 21292 25044 21304
rect 25096 21292 25102 21344
rect 25332 21341 25360 21372
rect 25317 21335 25375 21341
rect 25317 21301 25329 21335
rect 25363 21332 25375 21335
rect 25682 21332 25688 21344
rect 25363 21304 25688 21332
rect 25363 21301 25375 21304
rect 25317 21295 25375 21301
rect 25682 21292 25688 21304
rect 25740 21292 25746 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1578 21128 1584 21140
rect 1539 21100 1584 21128
rect 1578 21088 1584 21100
rect 1636 21088 1642 21140
rect 2590 21088 2596 21140
rect 2648 21128 2654 21140
rect 2685 21131 2743 21137
rect 2685 21128 2697 21131
rect 2648 21100 2697 21128
rect 2648 21088 2654 21100
rect 2685 21097 2697 21100
rect 2731 21097 2743 21131
rect 2685 21091 2743 21097
rect 3145 21131 3203 21137
rect 3145 21097 3157 21131
rect 3191 21128 3203 21131
rect 3510 21128 3516 21140
rect 3191 21100 3516 21128
rect 3191 21097 3203 21100
rect 3145 21091 3203 21097
rect 2225 21063 2283 21069
rect 2225 21029 2237 21063
rect 2271 21060 2283 21063
rect 3160 21060 3188 21091
rect 3510 21088 3516 21100
rect 3568 21088 3574 21140
rect 4890 21128 4896 21140
rect 4851 21100 4896 21128
rect 4890 21088 4896 21100
rect 4948 21088 4954 21140
rect 5534 21088 5540 21140
rect 5592 21128 5598 21140
rect 6273 21131 6331 21137
rect 6273 21128 6285 21131
rect 5592 21100 6285 21128
rect 5592 21088 5598 21100
rect 6273 21097 6285 21100
rect 6319 21097 6331 21131
rect 6273 21091 6331 21097
rect 2271 21032 3188 21060
rect 4433 21063 4491 21069
rect 2271 21029 2283 21032
rect 2225 21023 2283 21029
rect 4433 21029 4445 21063
rect 4479 21060 4491 21063
rect 5442 21060 5448 21072
rect 4479 21032 5448 21060
rect 4479 21029 4491 21032
rect 4433 21023 4491 21029
rect 5442 21020 5448 21032
rect 5500 21020 5506 21072
rect 6288 21060 6316 21091
rect 6546 21088 6552 21140
rect 6604 21128 6610 21140
rect 6917 21131 6975 21137
rect 6917 21128 6929 21131
rect 6604 21100 6929 21128
rect 6604 21088 6610 21100
rect 6917 21097 6929 21100
rect 6963 21097 6975 21131
rect 6917 21091 6975 21097
rect 8021 21131 8079 21137
rect 8021 21097 8033 21131
rect 8067 21128 8079 21131
rect 9030 21128 9036 21140
rect 8067 21100 9036 21128
rect 8067 21097 8079 21100
rect 8021 21091 8079 21097
rect 9030 21088 9036 21100
rect 9088 21088 9094 21140
rect 9674 21088 9680 21140
rect 9732 21128 9738 21140
rect 9861 21131 9919 21137
rect 9861 21128 9873 21131
rect 9732 21100 9873 21128
rect 9732 21088 9738 21100
rect 9861 21097 9873 21100
rect 9907 21097 9919 21131
rect 9861 21091 9919 21097
rect 10134 21088 10140 21140
rect 10192 21128 10198 21140
rect 11146 21128 11152 21140
rect 10192 21100 11152 21128
rect 10192 21088 10198 21100
rect 11146 21088 11152 21100
rect 11204 21088 11210 21140
rect 13633 21131 13691 21137
rect 13633 21097 13645 21131
rect 13679 21128 13691 21131
rect 16390 21128 16396 21140
rect 13679 21100 16396 21128
rect 13679 21097 13691 21100
rect 13633 21091 13691 21097
rect 16390 21088 16396 21100
rect 16448 21088 16454 21140
rect 16577 21131 16635 21137
rect 16577 21097 16589 21131
rect 16623 21128 16635 21131
rect 17770 21128 17776 21140
rect 16623 21100 17776 21128
rect 16623 21097 16635 21100
rect 16577 21091 16635 21097
rect 17770 21088 17776 21100
rect 17828 21088 17834 21140
rect 18138 21128 18144 21140
rect 18099 21100 18144 21128
rect 18138 21088 18144 21100
rect 18196 21088 18202 21140
rect 19518 21128 19524 21140
rect 19479 21100 19524 21128
rect 19518 21088 19524 21100
rect 19576 21088 19582 21140
rect 20990 21128 20996 21140
rect 20951 21100 20996 21128
rect 20990 21088 20996 21100
rect 21048 21088 21054 21140
rect 23382 21128 23388 21140
rect 23343 21100 23388 21128
rect 23382 21088 23388 21100
rect 23440 21088 23446 21140
rect 24854 21088 24860 21140
rect 24912 21128 24918 21140
rect 25133 21131 25191 21137
rect 25133 21128 25145 21131
rect 24912 21100 25145 21128
rect 24912 21088 24918 21100
rect 25133 21097 25145 21100
rect 25179 21097 25191 21131
rect 25133 21091 25191 21097
rect 6825 21063 6883 21069
rect 6825 21060 6837 21063
rect 6288 21032 6837 21060
rect 6825 21029 6837 21032
rect 6871 21029 6883 21063
rect 6825 21023 6883 21029
rect 8662 21020 8668 21072
rect 8720 21060 8726 21072
rect 10594 21060 10600 21072
rect 8720 21032 10600 21060
rect 8720 21020 8726 21032
rect 10594 21020 10600 21032
rect 10652 21020 10658 21072
rect 11048 21063 11106 21069
rect 11048 21029 11060 21063
rect 11094 21060 11106 21063
rect 11238 21060 11244 21072
rect 11094 21032 11244 21060
rect 11094 21029 11106 21032
rect 11048 21023 11106 21029
rect 11238 21020 11244 21032
rect 11296 21060 11302 21072
rect 12437 21063 12495 21069
rect 12437 21060 12449 21063
rect 11296 21032 12449 21060
rect 11296 21020 11302 21032
rect 12437 21029 12449 21032
rect 12483 21060 12495 21063
rect 12710 21060 12716 21072
rect 12483 21032 12716 21060
rect 12483 21029 12495 21032
rect 12437 21023 12495 21029
rect 12710 21020 12716 21032
rect 12768 21020 12774 21072
rect 13081 21063 13139 21069
rect 13081 21029 13093 21063
rect 13127 21060 13139 21063
rect 14090 21060 14096 21072
rect 13127 21032 14096 21060
rect 13127 21029 13139 21032
rect 13081 21023 13139 21029
rect 14090 21020 14096 21032
rect 14148 21020 14154 21072
rect 14274 21020 14280 21072
rect 14332 21020 14338 21072
rect 15120 21032 15424 21060
rect 1397 20995 1455 21001
rect 1397 20961 1409 20995
rect 1443 20992 1455 20995
rect 2038 20992 2044 21004
rect 1443 20964 2044 20992
rect 1443 20961 1455 20964
rect 1397 20955 1455 20961
rect 2038 20952 2044 20964
rect 2096 20952 2102 21004
rect 2501 20995 2559 21001
rect 2501 20961 2513 20995
rect 2547 20992 2559 20995
rect 3142 20992 3148 21004
rect 2547 20964 3148 20992
rect 2547 20961 2559 20964
rect 2501 20955 2559 20961
rect 3142 20952 3148 20964
rect 3200 20952 3206 21004
rect 5261 20995 5319 21001
rect 5261 20992 5273 20995
rect 5000 20964 5273 20992
rect 5000 20936 5028 20964
rect 5261 20961 5273 20964
rect 5307 20961 5319 20995
rect 5261 20955 5319 20961
rect 5353 20995 5411 21001
rect 5353 20961 5365 20995
rect 5399 20992 5411 20995
rect 5534 20992 5540 21004
rect 5399 20964 5540 20992
rect 5399 20961 5411 20964
rect 5353 20955 5411 20961
rect 5534 20952 5540 20964
rect 5592 20952 5598 21004
rect 7561 20995 7619 21001
rect 7561 20961 7573 20995
rect 7607 20992 7619 20995
rect 8018 20992 8024 21004
rect 7607 20964 8024 20992
rect 7607 20961 7619 20964
rect 7561 20955 7619 20961
rect 8018 20952 8024 20964
rect 8076 20992 8082 21004
rect 8389 20995 8447 21001
rect 8389 20992 8401 20995
rect 8076 20964 8401 20992
rect 8076 20952 8082 20964
rect 8389 20961 8401 20964
rect 8435 20961 8447 20995
rect 8389 20955 8447 20961
rect 8481 20995 8539 21001
rect 8481 20961 8493 20995
rect 8527 20992 8539 20995
rect 9582 20992 9588 21004
rect 8527 20964 9588 20992
rect 8527 20961 8539 20964
rect 8481 20955 8539 20961
rect 4982 20884 4988 20936
rect 5040 20884 5046 20936
rect 5074 20884 5080 20936
rect 5132 20924 5138 20936
rect 5445 20927 5503 20933
rect 5445 20924 5457 20927
rect 5132 20896 5457 20924
rect 5132 20884 5138 20896
rect 5445 20893 5457 20896
rect 5491 20924 5503 20927
rect 5810 20924 5816 20936
rect 5491 20896 5816 20924
rect 5491 20893 5503 20896
rect 5445 20887 5503 20893
rect 5810 20884 5816 20896
rect 5868 20884 5874 20936
rect 5994 20884 6000 20936
rect 6052 20924 6058 20936
rect 7009 20927 7067 20933
rect 7009 20924 7021 20927
rect 6052 20896 7021 20924
rect 6052 20884 6058 20896
rect 7009 20893 7021 20896
rect 7055 20893 7067 20927
rect 7009 20887 7067 20893
rect 7929 20927 7987 20933
rect 7929 20893 7941 20927
rect 7975 20924 7987 20927
rect 8496 20924 8524 20955
rect 9582 20952 9588 20964
rect 9640 20952 9646 21004
rect 9677 20995 9735 21001
rect 9677 20961 9689 20995
rect 9723 20992 9735 20995
rect 9858 20992 9864 21004
rect 9723 20964 9864 20992
rect 9723 20961 9735 20964
rect 9677 20955 9735 20961
rect 9858 20952 9864 20964
rect 9916 20952 9922 21004
rect 10686 20952 10692 21004
rect 10744 20992 10750 21004
rect 10781 20995 10839 21001
rect 10781 20992 10793 20995
rect 10744 20964 10793 20992
rect 10744 20952 10750 20964
rect 10781 20961 10793 20964
rect 10827 20961 10839 20995
rect 10781 20955 10839 20961
rect 13814 20952 13820 21004
rect 13872 20992 13878 21004
rect 14001 20995 14059 21001
rect 14001 20992 14013 20995
rect 13872 20964 14013 20992
rect 13872 20952 13878 20964
rect 14001 20961 14013 20964
rect 14047 20992 14059 20995
rect 14292 20992 14320 21020
rect 15120 20992 15148 21032
rect 15286 20992 15292 21004
rect 14047 20964 15148 20992
rect 15247 20964 15292 20992
rect 14047 20961 14059 20964
rect 14001 20955 14059 20961
rect 15286 20952 15292 20964
rect 15344 20952 15350 21004
rect 15396 20992 15424 21032
rect 15470 21020 15476 21072
rect 15528 21060 15534 21072
rect 15565 21063 15623 21069
rect 15565 21060 15577 21063
rect 15528 21032 15577 21060
rect 15528 21020 15534 21032
rect 15565 21029 15577 21032
rect 15611 21029 15623 21063
rect 22278 21060 22284 21072
rect 15565 21023 15623 21029
rect 15764 21032 22284 21060
rect 15764 20992 15792 21032
rect 22278 21020 22284 21032
rect 22336 21020 22342 21072
rect 23658 21020 23664 21072
rect 23716 21060 23722 21072
rect 23716 21032 25084 21060
rect 23716 21020 23722 21032
rect 15396 20964 15792 20992
rect 16574 20952 16580 21004
rect 16632 20992 16638 21004
rect 16945 20995 17003 21001
rect 16945 20992 16957 20995
rect 16632 20964 16957 20992
rect 16632 20952 16638 20964
rect 16945 20961 16957 20964
rect 16991 20961 17003 20995
rect 16945 20955 17003 20961
rect 18509 20995 18567 21001
rect 18509 20961 18521 20995
rect 18555 20992 18567 20995
rect 18690 20992 18696 21004
rect 18555 20964 18696 20992
rect 18555 20961 18567 20964
rect 18509 20955 18567 20961
rect 18690 20952 18696 20964
rect 18748 20992 18754 21004
rect 19242 20992 19248 21004
rect 18748 20964 19248 20992
rect 18748 20952 18754 20964
rect 19242 20952 19248 20964
rect 19300 20952 19306 21004
rect 19702 20992 19708 21004
rect 19663 20964 19708 20992
rect 19702 20952 19708 20964
rect 19760 20952 19766 21004
rect 20714 20952 20720 21004
rect 20772 20992 20778 21004
rect 21361 20995 21419 21001
rect 21361 20992 21373 20995
rect 20772 20964 21373 20992
rect 20772 20952 20778 20964
rect 21361 20961 21373 20964
rect 21407 20961 21419 20995
rect 23750 20992 23756 21004
rect 23711 20964 23756 20992
rect 21361 20955 21419 20961
rect 23750 20952 23756 20964
rect 23808 20952 23814 21004
rect 23845 20995 23903 21001
rect 23845 20961 23857 20995
rect 23891 20992 23903 20995
rect 24026 20992 24032 21004
rect 23891 20964 24032 20992
rect 23891 20961 23903 20964
rect 23845 20955 23903 20961
rect 24026 20952 24032 20964
rect 24084 20992 24090 21004
rect 24765 20995 24823 21001
rect 24765 20992 24777 20995
rect 24084 20964 24777 20992
rect 24084 20952 24090 20964
rect 24765 20961 24777 20964
rect 24811 20961 24823 20995
rect 24946 20992 24952 21004
rect 24907 20964 24952 20992
rect 24765 20955 24823 20961
rect 24946 20952 24952 20964
rect 25004 20952 25010 21004
rect 25056 20992 25084 21032
rect 25130 20992 25136 21004
rect 25056 20964 25136 20992
rect 25130 20952 25136 20964
rect 25188 20952 25194 21004
rect 7975 20896 8524 20924
rect 8573 20927 8631 20933
rect 7975 20893 7987 20896
rect 7929 20887 7987 20893
rect 8573 20893 8585 20927
rect 8619 20924 8631 20927
rect 9401 20927 9459 20933
rect 9401 20924 9413 20927
rect 8619 20896 9413 20924
rect 8619 20893 8631 20896
rect 8573 20887 8631 20893
rect 9401 20893 9413 20896
rect 9447 20924 9459 20927
rect 9490 20924 9496 20936
rect 9447 20896 9496 20924
rect 9447 20893 9459 20896
rect 9401 20887 9459 20893
rect 4801 20859 4859 20865
rect 4801 20825 4813 20859
rect 4847 20856 4859 20859
rect 5534 20856 5540 20868
rect 4847 20828 5540 20856
rect 4847 20825 4859 20828
rect 4801 20819 4859 20825
rect 5534 20816 5540 20828
rect 5592 20856 5598 20868
rect 6457 20859 6515 20865
rect 6457 20856 6469 20859
rect 5592 20828 6469 20856
rect 5592 20816 5598 20828
rect 6457 20825 6469 20828
rect 6503 20825 6515 20859
rect 6457 20819 6515 20825
rect 8294 20816 8300 20868
rect 8352 20856 8358 20868
rect 8588 20856 8616 20887
rect 9490 20884 9496 20896
rect 9548 20884 9554 20936
rect 14277 20927 14335 20933
rect 14277 20893 14289 20927
rect 14323 20924 14335 20927
rect 15930 20924 15936 20936
rect 14323 20896 15936 20924
rect 14323 20893 14335 20896
rect 14277 20887 14335 20893
rect 15930 20884 15936 20896
rect 15988 20884 15994 20936
rect 17034 20924 17040 20936
rect 16995 20896 17040 20924
rect 17034 20884 17040 20896
rect 17092 20884 17098 20936
rect 17221 20927 17279 20933
rect 17221 20893 17233 20927
rect 17267 20924 17279 20927
rect 17402 20924 17408 20936
rect 17267 20896 17408 20924
rect 17267 20893 17279 20896
rect 17221 20887 17279 20893
rect 17402 20884 17408 20896
rect 17460 20884 17466 20936
rect 18138 20884 18144 20936
rect 18196 20924 18202 20936
rect 18601 20927 18659 20933
rect 18601 20924 18613 20927
rect 18196 20896 18613 20924
rect 18196 20884 18202 20896
rect 18601 20893 18613 20896
rect 18647 20893 18659 20927
rect 18601 20887 18659 20893
rect 18785 20927 18843 20933
rect 18785 20893 18797 20927
rect 18831 20924 18843 20927
rect 18874 20924 18880 20936
rect 18831 20896 18880 20924
rect 18831 20893 18843 20896
rect 18785 20887 18843 20893
rect 8352 20828 8616 20856
rect 8352 20816 8358 20828
rect 8846 20816 8852 20868
rect 8904 20856 8910 20868
rect 9950 20856 9956 20868
rect 8904 20828 9956 20856
rect 8904 20816 8910 20828
rect 9950 20816 9956 20828
rect 10008 20856 10014 20868
rect 10597 20859 10655 20865
rect 10597 20856 10609 20859
rect 10008 20828 10609 20856
rect 10008 20816 10014 20828
rect 10597 20825 10609 20828
rect 10643 20825 10655 20859
rect 10597 20819 10655 20825
rect 13449 20859 13507 20865
rect 13449 20825 13461 20859
rect 13495 20856 13507 20859
rect 13722 20856 13728 20868
rect 13495 20828 13728 20856
rect 13495 20825 13507 20828
rect 13449 20819 13507 20825
rect 13722 20816 13728 20828
rect 13780 20816 13786 20868
rect 14737 20859 14795 20865
rect 14737 20825 14749 20859
rect 14783 20856 14795 20859
rect 14826 20856 14832 20868
rect 14783 20828 14832 20856
rect 14783 20825 14795 20828
rect 14737 20819 14795 20825
rect 14826 20816 14832 20828
rect 14884 20856 14890 20868
rect 16117 20859 16175 20865
rect 16117 20856 16129 20859
rect 14884 20828 16129 20856
rect 14884 20816 14890 20828
rect 16117 20825 16129 20828
rect 16163 20856 16175 20859
rect 18049 20859 18107 20865
rect 18049 20856 18061 20859
rect 16163 20828 18061 20856
rect 16163 20825 16175 20828
rect 16117 20819 16175 20825
rect 18049 20825 18061 20828
rect 18095 20856 18107 20859
rect 18800 20856 18828 20887
rect 18874 20884 18880 20896
rect 18932 20884 18938 20936
rect 20990 20884 20996 20936
rect 21048 20924 21054 20936
rect 21453 20927 21511 20933
rect 21453 20924 21465 20927
rect 21048 20896 21465 20924
rect 21048 20884 21054 20896
rect 21453 20893 21465 20896
rect 21499 20893 21511 20927
rect 21453 20887 21511 20893
rect 21637 20927 21695 20933
rect 21637 20893 21649 20927
rect 21683 20924 21695 20927
rect 22370 20924 22376 20936
rect 21683 20896 22376 20924
rect 21683 20893 21695 20896
rect 21637 20887 21695 20893
rect 22370 20884 22376 20896
rect 22428 20884 22434 20936
rect 22925 20927 22983 20933
rect 22925 20893 22937 20927
rect 22971 20924 22983 20927
rect 23658 20924 23664 20936
rect 22971 20896 23664 20924
rect 22971 20893 22983 20896
rect 22925 20887 22983 20893
rect 23658 20884 23664 20896
rect 23716 20884 23722 20936
rect 23937 20927 23995 20933
rect 23937 20893 23949 20927
rect 23983 20924 23995 20927
rect 24854 20924 24860 20936
rect 23983 20896 24860 20924
rect 23983 20893 23995 20896
rect 23937 20887 23995 20893
rect 24854 20884 24860 20896
rect 24912 20884 24918 20936
rect 19886 20856 19892 20868
rect 18095 20828 18828 20856
rect 19847 20828 19892 20856
rect 18095 20825 18107 20828
rect 18049 20819 18107 20825
rect 19886 20816 19892 20828
rect 19944 20816 19950 20868
rect 22097 20859 22155 20865
rect 22097 20825 22109 20859
rect 22143 20856 22155 20859
rect 22738 20856 22744 20868
rect 22143 20828 22744 20856
rect 22143 20825 22155 20828
rect 22097 20819 22155 20825
rect 22738 20816 22744 20828
rect 22796 20816 22802 20868
rect 23293 20859 23351 20865
rect 23293 20825 23305 20859
rect 23339 20856 23351 20859
rect 24118 20856 24124 20868
rect 23339 20828 24124 20856
rect 23339 20825 23351 20828
rect 23293 20819 23351 20825
rect 24118 20816 24124 20828
rect 24176 20816 24182 20868
rect 3881 20791 3939 20797
rect 3881 20757 3893 20791
rect 3927 20788 3939 20791
rect 5166 20788 5172 20800
rect 3927 20760 5172 20788
rect 3927 20757 3939 20760
rect 3881 20751 3939 20757
rect 5166 20748 5172 20760
rect 5224 20748 5230 20800
rect 5997 20791 6055 20797
rect 5997 20757 6009 20791
rect 6043 20788 6055 20791
rect 6178 20788 6184 20800
rect 6043 20760 6184 20788
rect 6043 20757 6055 20760
rect 5997 20751 6055 20757
rect 6178 20748 6184 20760
rect 6236 20748 6242 20800
rect 9125 20791 9183 20797
rect 9125 20757 9137 20791
rect 9171 20788 9183 20791
rect 9490 20788 9496 20800
rect 9171 20760 9496 20788
rect 9171 20757 9183 20760
rect 9125 20751 9183 20757
rect 9490 20748 9496 20760
rect 9548 20748 9554 20800
rect 10318 20788 10324 20800
rect 10279 20760 10324 20788
rect 10318 20748 10324 20760
rect 10376 20748 10382 20800
rect 10686 20748 10692 20800
rect 10744 20788 10750 20800
rect 12161 20791 12219 20797
rect 12161 20788 12173 20791
rect 10744 20760 12173 20788
rect 10744 20748 10750 20760
rect 12161 20757 12173 20760
rect 12207 20757 12219 20791
rect 12161 20751 12219 20757
rect 15105 20791 15163 20797
rect 15105 20757 15117 20791
rect 15151 20788 15163 20791
rect 15378 20788 15384 20800
rect 15151 20760 15384 20788
rect 15151 20757 15163 20760
rect 15105 20751 15163 20757
rect 15378 20748 15384 20760
rect 15436 20748 15442 20800
rect 17310 20748 17316 20800
rect 17368 20788 17374 20800
rect 17589 20791 17647 20797
rect 17589 20788 17601 20791
rect 17368 20760 17601 20788
rect 17368 20748 17374 20760
rect 17589 20757 17601 20760
rect 17635 20757 17647 20791
rect 17589 20751 17647 20757
rect 19058 20748 19064 20800
rect 19116 20788 19122 20800
rect 19153 20791 19211 20797
rect 19153 20788 19165 20791
rect 19116 20760 19165 20788
rect 19116 20748 19122 20760
rect 19153 20757 19165 20760
rect 19199 20757 19211 20791
rect 19153 20751 19211 20757
rect 20533 20791 20591 20797
rect 20533 20757 20545 20791
rect 20579 20788 20591 20791
rect 22278 20788 22284 20800
rect 20579 20760 22284 20788
rect 20579 20757 20591 20760
rect 20533 20751 20591 20757
rect 22278 20748 22284 20760
rect 22336 20788 22342 20800
rect 22373 20791 22431 20797
rect 22373 20788 22385 20791
rect 22336 20760 22385 20788
rect 22336 20748 22342 20760
rect 22373 20757 22385 20760
rect 22419 20788 22431 20791
rect 24397 20791 24455 20797
rect 24397 20788 24409 20791
rect 22419 20760 24409 20788
rect 22419 20757 22431 20760
rect 22373 20751 22431 20757
rect 24397 20757 24409 20760
rect 24443 20757 24455 20791
rect 24397 20751 24455 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 2682 20584 2688 20596
rect 2643 20556 2688 20584
rect 2682 20544 2688 20556
rect 2740 20544 2746 20596
rect 5169 20587 5227 20593
rect 5169 20553 5181 20587
rect 5215 20584 5227 20587
rect 5258 20584 5264 20596
rect 5215 20556 5264 20584
rect 5215 20553 5227 20556
rect 5169 20547 5227 20553
rect 5258 20544 5264 20556
rect 5316 20544 5322 20596
rect 6546 20544 6552 20596
rect 6604 20584 6610 20596
rect 6825 20587 6883 20593
rect 6825 20584 6837 20587
rect 6604 20556 6837 20584
rect 6604 20544 6610 20556
rect 6825 20553 6837 20556
rect 6871 20553 6883 20587
rect 6825 20547 6883 20553
rect 8113 20587 8171 20593
rect 8113 20553 8125 20587
rect 8159 20584 8171 20587
rect 8294 20584 8300 20596
rect 8159 20556 8300 20584
rect 8159 20553 8171 20556
rect 8113 20547 8171 20553
rect 8294 20544 8300 20556
rect 8352 20544 8358 20596
rect 8573 20587 8631 20593
rect 8573 20553 8585 20587
rect 8619 20584 8631 20587
rect 9306 20584 9312 20596
rect 8619 20556 9312 20584
rect 8619 20553 8631 20556
rect 8573 20547 8631 20553
rect 9306 20544 9312 20556
rect 9364 20544 9370 20596
rect 9674 20544 9680 20596
rect 9732 20584 9738 20596
rect 10137 20587 10195 20593
rect 10137 20584 10149 20587
rect 9732 20556 10149 20584
rect 9732 20544 9738 20556
rect 10137 20553 10149 20556
rect 10183 20553 10195 20587
rect 10137 20547 10195 20553
rect 13725 20587 13783 20593
rect 13725 20553 13737 20587
rect 13771 20584 13783 20587
rect 13814 20584 13820 20596
rect 13771 20556 13820 20584
rect 13771 20553 13783 20556
rect 13725 20547 13783 20553
rect 13814 20544 13820 20556
rect 13872 20544 13878 20596
rect 14182 20584 14188 20596
rect 14143 20556 14188 20584
rect 14182 20544 14188 20556
rect 14240 20544 14246 20596
rect 14366 20584 14372 20596
rect 14327 20556 14372 20584
rect 14366 20544 14372 20556
rect 14424 20544 14430 20596
rect 15378 20544 15384 20596
rect 15436 20584 15442 20596
rect 16393 20587 16451 20593
rect 16393 20584 16405 20587
rect 15436 20556 16405 20584
rect 15436 20544 15442 20556
rect 16393 20553 16405 20556
rect 16439 20584 16451 20587
rect 16482 20584 16488 20596
rect 16439 20556 16488 20584
rect 16439 20553 16451 20556
rect 16393 20547 16451 20553
rect 16482 20544 16488 20556
rect 16540 20544 16546 20596
rect 20990 20584 20996 20596
rect 20951 20556 20996 20584
rect 20990 20544 20996 20556
rect 21048 20544 21054 20596
rect 21818 20544 21824 20596
rect 21876 20584 21882 20596
rect 24946 20584 24952 20596
rect 21876 20556 24952 20584
rect 21876 20544 21882 20556
rect 24946 20544 24952 20556
rect 25004 20544 25010 20596
rect 25406 20584 25412 20596
rect 25367 20556 25412 20584
rect 25406 20544 25412 20556
rect 25464 20544 25470 20596
rect 2038 20516 2044 20528
rect 1999 20488 2044 20516
rect 2038 20476 2044 20488
rect 2096 20476 2102 20528
rect 3878 20476 3884 20528
rect 3936 20516 3942 20528
rect 8386 20516 8392 20528
rect 3936 20488 8392 20516
rect 3936 20476 3942 20488
rect 8386 20476 8392 20488
rect 8444 20476 8450 20528
rect 9585 20519 9643 20525
rect 9585 20485 9597 20519
rect 9631 20516 9643 20519
rect 9631 20488 10732 20516
rect 9631 20485 9643 20488
rect 9585 20479 9643 20485
rect 5534 20408 5540 20460
rect 5592 20408 5598 20460
rect 5718 20448 5724 20460
rect 5679 20420 5724 20448
rect 5718 20408 5724 20420
rect 5776 20408 5782 20460
rect 6914 20408 6920 20460
rect 6972 20448 6978 20460
rect 7285 20451 7343 20457
rect 7285 20448 7297 20451
rect 6972 20420 7297 20448
rect 6972 20408 6978 20420
rect 7285 20417 7297 20420
rect 7331 20417 7343 20451
rect 7285 20411 7343 20417
rect 7377 20451 7435 20457
rect 7377 20417 7389 20451
rect 7423 20417 7435 20451
rect 7377 20411 7435 20417
rect 8481 20451 8539 20457
rect 8481 20417 8493 20451
rect 8527 20448 8539 20451
rect 8662 20448 8668 20460
rect 8527 20420 8668 20448
rect 8527 20417 8539 20420
rect 8481 20411 8539 20417
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20380 1455 20383
rect 1443 20352 2452 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 2424 20256 2452 20352
rect 2498 20340 2504 20392
rect 2556 20380 2562 20392
rect 3421 20383 3479 20389
rect 3421 20380 3433 20383
rect 2556 20352 3433 20380
rect 2556 20340 2562 20352
rect 3421 20349 3433 20352
rect 3467 20349 3479 20383
rect 3602 20380 3608 20392
rect 3515 20352 3608 20380
rect 3421 20343 3479 20349
rect 3602 20340 3608 20352
rect 3660 20380 3666 20392
rect 4157 20383 4215 20389
rect 4157 20380 4169 20383
rect 3660 20352 4169 20380
rect 3660 20340 3666 20352
rect 4157 20349 4169 20352
rect 4203 20349 4215 20383
rect 5552 20380 5580 20408
rect 5629 20383 5687 20389
rect 5629 20380 5641 20383
rect 5552 20352 5641 20380
rect 4157 20343 4215 20349
rect 5629 20349 5641 20352
rect 5675 20349 5687 20383
rect 6638 20380 6644 20392
rect 6551 20352 6644 20380
rect 5629 20343 5687 20349
rect 6638 20340 6644 20352
rect 6696 20380 6702 20392
rect 7392 20380 7420 20411
rect 8662 20408 8668 20420
rect 8720 20448 8726 20460
rect 9217 20451 9275 20457
rect 9217 20448 9229 20451
rect 8720 20420 9229 20448
rect 8720 20408 8726 20420
rect 9217 20417 9229 20420
rect 9263 20448 9275 20451
rect 9398 20448 9404 20460
rect 9263 20420 9404 20448
rect 9263 20417 9275 20420
rect 9217 20411 9275 20417
rect 9398 20408 9404 20420
rect 9456 20448 9462 20460
rect 9600 20448 9628 20479
rect 10704 20460 10732 20488
rect 10686 20448 10692 20460
rect 9456 20420 9628 20448
rect 10647 20420 10692 20448
rect 9456 20408 9462 20420
rect 10686 20408 10692 20420
rect 10744 20408 10750 20460
rect 12710 20408 12716 20460
rect 12768 20448 12774 20460
rect 12989 20451 13047 20457
rect 12989 20448 13001 20451
rect 12768 20420 13001 20448
rect 12768 20408 12774 20420
rect 12989 20417 13001 20420
rect 13035 20417 13047 20451
rect 14200 20448 14228 20544
rect 15473 20519 15531 20525
rect 15473 20485 15485 20519
rect 15519 20516 15531 20519
rect 15930 20516 15936 20528
rect 15519 20488 15936 20516
rect 15519 20485 15531 20488
rect 15473 20479 15531 20485
rect 15930 20476 15936 20488
rect 15988 20476 15994 20528
rect 17862 20476 17868 20528
rect 17920 20516 17926 20528
rect 18049 20519 18107 20525
rect 18049 20516 18061 20519
rect 17920 20488 18061 20516
rect 17920 20476 17926 20488
rect 18049 20485 18061 20488
rect 18095 20485 18107 20519
rect 18049 20479 18107 20485
rect 18138 20476 18144 20528
rect 18196 20516 18202 20528
rect 19153 20519 19211 20525
rect 19153 20516 19165 20519
rect 18196 20488 19165 20516
rect 18196 20476 18202 20488
rect 19153 20485 19165 20488
rect 19199 20516 19211 20519
rect 22465 20519 22523 20525
rect 22465 20516 22477 20519
rect 19199 20488 20300 20516
rect 19199 20485 19211 20488
rect 19153 20479 19211 20485
rect 14829 20451 14887 20457
rect 14829 20448 14841 20451
rect 14200 20420 14841 20448
rect 12989 20411 13047 20417
rect 14829 20417 14841 20420
rect 14875 20417 14887 20451
rect 14829 20411 14887 20417
rect 14918 20408 14924 20460
rect 14976 20448 14982 20460
rect 14976 20420 15021 20448
rect 14976 20408 14982 20420
rect 15838 20408 15844 20460
rect 15896 20448 15902 20460
rect 16209 20451 16267 20457
rect 16209 20448 16221 20451
rect 15896 20420 16221 20448
rect 15896 20408 15902 20420
rect 16209 20417 16221 20420
rect 16255 20448 16267 20451
rect 16945 20451 17003 20457
rect 16945 20448 16957 20451
rect 16255 20420 16957 20448
rect 16255 20417 16267 20420
rect 16209 20411 16267 20417
rect 16945 20417 16957 20420
rect 16991 20448 17003 20451
rect 17310 20448 17316 20460
rect 16991 20420 17316 20448
rect 16991 20417 17003 20420
rect 16945 20411 17003 20417
rect 17310 20408 17316 20420
rect 17368 20448 17374 20460
rect 18601 20451 18659 20457
rect 18601 20448 18613 20451
rect 17368 20420 18613 20448
rect 17368 20408 17374 20420
rect 18601 20417 18613 20420
rect 18647 20417 18659 20451
rect 18601 20411 18659 20417
rect 20070 20408 20076 20460
rect 20128 20448 20134 20460
rect 20165 20451 20223 20457
rect 20165 20448 20177 20451
rect 20128 20420 20177 20448
rect 20128 20408 20134 20420
rect 20165 20417 20177 20420
rect 20211 20417 20223 20451
rect 20165 20411 20223 20417
rect 6696 20352 7420 20380
rect 6696 20340 6702 20352
rect 10318 20340 10324 20392
rect 10376 20380 10382 20392
rect 10597 20383 10655 20389
rect 10597 20380 10609 20383
rect 10376 20352 10609 20380
rect 10376 20340 10382 20352
rect 10597 20349 10609 20352
rect 10643 20380 10655 20383
rect 10778 20380 10784 20392
rect 10643 20352 10784 20380
rect 10643 20349 10655 20352
rect 10597 20343 10655 20349
rect 10778 20340 10784 20352
rect 10836 20340 10842 20392
rect 15930 20340 15936 20392
rect 15988 20380 15994 20392
rect 16390 20380 16396 20392
rect 15988 20352 16396 20380
rect 15988 20340 15994 20352
rect 16390 20340 16396 20352
rect 16448 20340 16454 20392
rect 18414 20380 18420 20392
rect 18375 20352 18420 20380
rect 18414 20340 18420 20352
rect 18472 20340 18478 20392
rect 18506 20340 18512 20392
rect 18564 20380 18570 20392
rect 18564 20352 18609 20380
rect 18564 20340 18570 20352
rect 19426 20340 19432 20392
rect 19484 20380 19490 20392
rect 19981 20383 20039 20389
rect 19981 20380 19993 20383
rect 19484 20352 19993 20380
rect 19484 20340 19490 20352
rect 19981 20349 19993 20352
rect 20027 20349 20039 20383
rect 19981 20343 20039 20349
rect 3142 20312 3148 20324
rect 3103 20284 3148 20312
rect 3142 20272 3148 20284
rect 3200 20272 3206 20324
rect 4617 20315 4675 20321
rect 4617 20281 4629 20315
rect 4663 20312 4675 20315
rect 5074 20312 5080 20324
rect 4663 20284 5080 20312
rect 4663 20281 4675 20284
rect 4617 20275 4675 20281
rect 5074 20272 5080 20284
rect 5132 20272 5138 20324
rect 5534 20312 5540 20324
rect 5495 20284 5540 20312
rect 5534 20272 5540 20284
rect 5592 20272 5598 20324
rect 8938 20312 8944 20324
rect 8899 20284 8944 20312
rect 8938 20272 8944 20284
rect 8996 20272 9002 20324
rect 12253 20315 12311 20321
rect 12253 20281 12265 20315
rect 12299 20312 12311 20315
rect 12897 20315 12955 20321
rect 12897 20312 12909 20315
rect 12299 20284 12909 20312
rect 12299 20281 12311 20284
rect 12253 20275 12311 20281
rect 12897 20281 12909 20284
rect 12943 20312 12955 20315
rect 13170 20312 13176 20324
rect 12943 20284 13176 20312
rect 12943 20281 12955 20284
rect 12897 20275 12955 20281
rect 13170 20272 13176 20284
rect 13228 20272 13234 20324
rect 16853 20315 16911 20321
rect 16853 20312 16865 20315
rect 15948 20284 16865 20312
rect 15948 20256 15976 20284
rect 16853 20281 16865 20284
rect 16899 20281 16911 20315
rect 19702 20312 19708 20324
rect 16853 20275 16911 20281
rect 19444 20284 19708 20312
rect 1394 20204 1400 20256
rect 1452 20244 1458 20256
rect 1581 20247 1639 20253
rect 1581 20244 1593 20247
rect 1452 20216 1593 20244
rect 1452 20204 1458 20216
rect 1581 20213 1593 20216
rect 1627 20213 1639 20247
rect 2406 20244 2412 20256
rect 2367 20216 2412 20244
rect 1581 20207 1639 20213
rect 2406 20204 2412 20216
rect 2464 20204 2470 20256
rect 3786 20244 3792 20256
rect 3747 20216 3792 20244
rect 3786 20204 3792 20216
rect 3844 20204 3850 20256
rect 4982 20244 4988 20256
rect 4895 20216 4988 20244
rect 4982 20204 4988 20216
rect 5040 20244 5046 20256
rect 5258 20244 5264 20256
rect 5040 20216 5264 20244
rect 5040 20204 5046 20216
rect 5258 20204 5264 20216
rect 5316 20204 5322 20256
rect 5994 20204 6000 20256
rect 6052 20244 6058 20256
rect 6181 20247 6239 20253
rect 6181 20244 6193 20247
rect 6052 20216 6193 20244
rect 6052 20204 6058 20216
rect 6181 20213 6193 20216
rect 6227 20213 6239 20247
rect 7190 20244 7196 20256
rect 7151 20216 7196 20244
rect 6181 20207 6239 20213
rect 7190 20204 7196 20216
rect 7248 20204 7254 20256
rect 9033 20247 9091 20253
rect 9033 20213 9045 20247
rect 9079 20244 9091 20247
rect 9122 20244 9128 20256
rect 9079 20216 9128 20244
rect 9079 20213 9091 20216
rect 9033 20207 9091 20213
rect 9122 20204 9128 20216
rect 9180 20204 9186 20256
rect 9582 20204 9588 20256
rect 9640 20244 9646 20256
rect 9953 20247 10011 20253
rect 9953 20244 9965 20247
rect 9640 20216 9965 20244
rect 9640 20204 9646 20216
rect 9953 20213 9965 20216
rect 9999 20244 10011 20247
rect 10505 20247 10563 20253
rect 10505 20244 10517 20247
rect 9999 20216 10517 20244
rect 9999 20213 10011 20216
rect 9953 20207 10011 20213
rect 10505 20213 10517 20216
rect 10551 20213 10563 20247
rect 11238 20244 11244 20256
rect 11199 20216 11244 20244
rect 10505 20207 10563 20213
rect 11238 20204 11244 20216
rect 11296 20244 11302 20256
rect 11517 20247 11575 20253
rect 11517 20244 11529 20247
rect 11296 20216 11529 20244
rect 11296 20204 11302 20216
rect 11517 20213 11529 20216
rect 11563 20213 11575 20247
rect 11517 20207 11575 20213
rect 12434 20204 12440 20256
rect 12492 20244 12498 20256
rect 12802 20244 12808 20256
rect 12492 20216 12537 20244
rect 12763 20216 12808 20244
rect 12492 20204 12498 20216
rect 12802 20204 12808 20216
rect 12860 20204 12866 20256
rect 14642 20204 14648 20256
rect 14700 20244 14706 20256
rect 14737 20247 14795 20253
rect 14737 20244 14749 20247
rect 14700 20216 14749 20244
rect 14700 20204 14706 20216
rect 14737 20213 14749 20216
rect 14783 20213 14795 20247
rect 15930 20244 15936 20256
rect 15891 20216 15936 20244
rect 14737 20207 14795 20213
rect 15930 20204 15936 20216
rect 15988 20204 15994 20256
rect 16758 20244 16764 20256
rect 16719 20216 16764 20244
rect 16758 20204 16764 20216
rect 16816 20204 16822 20256
rect 17402 20244 17408 20256
rect 17363 20216 17408 20244
rect 17402 20204 17408 20216
rect 17460 20204 17466 20256
rect 17862 20244 17868 20256
rect 17823 20216 17868 20244
rect 17862 20204 17868 20216
rect 17920 20204 17926 20256
rect 19242 20204 19248 20256
rect 19300 20244 19306 20256
rect 19444 20253 19472 20284
rect 19702 20272 19708 20284
rect 19760 20272 19766 20324
rect 19429 20247 19487 20253
rect 19429 20244 19441 20247
rect 19300 20216 19441 20244
rect 19300 20204 19306 20216
rect 19429 20213 19441 20216
rect 19475 20213 19487 20247
rect 19429 20207 19487 20213
rect 19518 20204 19524 20256
rect 19576 20244 19582 20256
rect 19613 20247 19671 20253
rect 19613 20244 19625 20247
rect 19576 20216 19625 20244
rect 19576 20204 19582 20216
rect 19613 20213 19625 20216
rect 19659 20213 19671 20247
rect 19613 20207 19671 20213
rect 20073 20247 20131 20253
rect 20073 20213 20085 20247
rect 20119 20244 20131 20247
rect 20272 20244 20300 20488
rect 21560 20488 22477 20516
rect 20714 20448 20720 20460
rect 20675 20420 20720 20448
rect 20714 20408 20720 20420
rect 20772 20408 20778 20460
rect 21560 20389 21588 20488
rect 22465 20485 22477 20488
rect 22511 20485 22523 20519
rect 24210 20516 24216 20528
rect 22465 20479 22523 20485
rect 23400 20488 24216 20516
rect 21634 20408 21640 20460
rect 21692 20448 21698 20460
rect 21729 20451 21787 20457
rect 21729 20448 21741 20451
rect 21692 20420 21741 20448
rect 21692 20408 21698 20420
rect 21729 20417 21741 20420
rect 21775 20448 21787 20451
rect 22189 20451 22247 20457
rect 22189 20448 22201 20451
rect 21775 20420 22201 20448
rect 21775 20417 21787 20420
rect 21729 20411 21787 20417
rect 22189 20417 22201 20420
rect 22235 20417 22247 20451
rect 22189 20411 22247 20417
rect 21545 20383 21603 20389
rect 21545 20349 21557 20383
rect 21591 20349 21603 20383
rect 22204 20380 22232 20411
rect 22370 20408 22376 20460
rect 22428 20448 22434 20460
rect 22649 20451 22707 20457
rect 22649 20448 22661 20451
rect 22428 20420 22661 20448
rect 22428 20408 22434 20420
rect 22649 20417 22661 20420
rect 22695 20448 22707 20451
rect 23198 20448 23204 20460
rect 22695 20420 23204 20448
rect 22695 20417 22707 20420
rect 22649 20411 22707 20417
rect 23198 20408 23204 20420
rect 23256 20408 23262 20460
rect 23400 20380 23428 20488
rect 24210 20476 24216 20488
rect 24268 20476 24274 20528
rect 24578 20476 24584 20528
rect 24636 20516 24642 20528
rect 24854 20516 24860 20528
rect 24636 20488 24860 20516
rect 24636 20476 24642 20488
rect 24854 20476 24860 20488
rect 24912 20476 24918 20528
rect 24118 20448 24124 20460
rect 24079 20420 24124 20448
rect 24118 20408 24124 20420
rect 24176 20408 24182 20460
rect 24305 20451 24363 20457
rect 24305 20417 24317 20451
rect 24351 20448 24363 20451
rect 24762 20448 24768 20460
rect 24351 20420 24768 20448
rect 24351 20417 24363 20420
rect 24305 20411 24363 20417
rect 24762 20408 24768 20420
rect 24820 20408 24826 20460
rect 22204 20352 23428 20380
rect 21545 20343 21603 20349
rect 23658 20340 23664 20392
rect 23716 20380 23722 20392
rect 23716 20352 23980 20380
rect 23716 20340 23722 20352
rect 21358 20272 21364 20324
rect 21416 20312 21422 20324
rect 22278 20312 22284 20324
rect 21416 20284 22284 20312
rect 21416 20272 21422 20284
rect 22278 20272 22284 20284
rect 22336 20272 22342 20324
rect 22370 20272 22376 20324
rect 22428 20312 22434 20324
rect 22830 20312 22836 20324
rect 22428 20284 22836 20312
rect 22428 20272 22434 20284
rect 22830 20272 22836 20284
rect 22888 20272 22894 20324
rect 23952 20312 23980 20352
rect 24946 20340 24952 20392
rect 25004 20380 25010 20392
rect 25225 20383 25283 20389
rect 25225 20380 25237 20383
rect 25004 20352 25237 20380
rect 25004 20340 25010 20352
rect 25225 20349 25237 20352
rect 25271 20380 25283 20383
rect 25777 20383 25835 20389
rect 25777 20380 25789 20383
rect 25271 20352 25789 20380
rect 25271 20349 25283 20352
rect 25225 20343 25283 20349
rect 25777 20349 25789 20352
rect 25823 20349 25835 20383
rect 25777 20343 25835 20349
rect 24029 20315 24087 20321
rect 24029 20312 24041 20315
rect 23952 20284 24041 20312
rect 24029 20281 24041 20284
rect 24075 20281 24087 20315
rect 24029 20275 24087 20281
rect 20806 20244 20812 20256
rect 20119 20216 20812 20244
rect 20119 20213 20131 20216
rect 20073 20207 20131 20213
rect 20806 20204 20812 20216
rect 20864 20204 20870 20256
rect 21174 20244 21180 20256
rect 21135 20216 21180 20244
rect 21174 20204 21180 20216
rect 21232 20204 21238 20256
rect 21634 20244 21640 20256
rect 21595 20216 21640 20244
rect 21634 20204 21640 20216
rect 21692 20204 21698 20256
rect 22465 20247 22523 20253
rect 22465 20213 22477 20247
rect 22511 20244 22523 20247
rect 23017 20247 23075 20253
rect 23017 20244 23029 20247
rect 22511 20216 23029 20244
rect 22511 20213 22523 20216
rect 22465 20207 22523 20213
rect 23017 20213 23029 20216
rect 23063 20244 23075 20247
rect 23106 20244 23112 20256
rect 23063 20216 23112 20244
rect 23063 20213 23075 20216
rect 23017 20207 23075 20213
rect 23106 20204 23112 20216
rect 23164 20204 23170 20256
rect 23474 20244 23480 20256
rect 23435 20216 23480 20244
rect 23474 20204 23480 20216
rect 23532 20204 23538 20256
rect 23661 20247 23719 20253
rect 23661 20213 23673 20247
rect 23707 20244 23719 20247
rect 23750 20244 23756 20256
rect 23707 20216 23756 20244
rect 23707 20213 23719 20216
rect 23661 20207 23719 20213
rect 23750 20204 23756 20216
rect 23808 20244 23814 20256
rect 24210 20244 24216 20256
rect 23808 20216 24216 20244
rect 23808 20204 23814 20216
rect 24210 20204 24216 20216
rect 24268 20204 24274 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 4246 20040 4252 20052
rect 4207 20012 4252 20040
rect 4246 20000 4252 20012
rect 4304 20000 4310 20052
rect 4706 20040 4712 20052
rect 4667 20012 4712 20040
rect 4706 20000 4712 20012
rect 4764 20000 4770 20052
rect 5721 20043 5779 20049
rect 5721 20009 5733 20043
rect 5767 20040 5779 20043
rect 6086 20040 6092 20052
rect 5767 20012 6092 20040
rect 5767 20009 5779 20012
rect 5721 20003 5779 20009
rect 6086 20000 6092 20012
rect 6144 20000 6150 20052
rect 7561 20043 7619 20049
rect 7561 20009 7573 20043
rect 7607 20040 7619 20043
rect 7650 20040 7656 20052
rect 7607 20012 7656 20040
rect 7607 20009 7619 20012
rect 7561 20003 7619 20009
rect 7650 20000 7656 20012
rect 7708 20000 7714 20052
rect 8018 20040 8024 20052
rect 7979 20012 8024 20040
rect 8018 20000 8024 20012
rect 8076 20000 8082 20052
rect 9858 20040 9864 20052
rect 9819 20012 9864 20040
rect 9858 20000 9864 20012
rect 9916 20000 9922 20052
rect 11054 20040 11060 20052
rect 11015 20012 11060 20040
rect 11054 20000 11060 20012
rect 11112 20000 11118 20052
rect 11514 20040 11520 20052
rect 11475 20012 11520 20040
rect 11514 20000 11520 20012
rect 11572 20000 11578 20052
rect 12529 20043 12587 20049
rect 12529 20009 12541 20043
rect 12575 20040 12587 20043
rect 12802 20040 12808 20052
rect 12575 20012 12808 20040
rect 12575 20009 12587 20012
rect 12529 20003 12587 20009
rect 12802 20000 12808 20012
rect 12860 20000 12866 20052
rect 13722 20000 13728 20052
rect 13780 20040 13786 20052
rect 14369 20043 14427 20049
rect 14369 20040 14381 20043
rect 13780 20012 14381 20040
rect 13780 20000 13786 20012
rect 14369 20009 14381 20012
rect 14415 20009 14427 20043
rect 15102 20040 15108 20052
rect 15063 20012 15108 20040
rect 14369 20003 14427 20009
rect 15102 20000 15108 20012
rect 15160 20000 15166 20052
rect 15289 20043 15347 20049
rect 15289 20009 15301 20043
rect 15335 20040 15347 20043
rect 16574 20040 16580 20052
rect 15335 20012 16580 20040
rect 15335 20009 15347 20012
rect 15289 20003 15347 20009
rect 16574 20000 16580 20012
rect 16632 20000 16638 20052
rect 18230 20000 18236 20052
rect 18288 20040 18294 20052
rect 18509 20043 18567 20049
rect 18509 20040 18521 20043
rect 18288 20012 18521 20040
rect 18288 20000 18294 20012
rect 18509 20009 18521 20012
rect 18555 20009 18567 20043
rect 18966 20040 18972 20052
rect 18927 20012 18972 20040
rect 18509 20003 18567 20009
rect 18966 20000 18972 20012
rect 19024 20000 19030 20052
rect 20070 20040 20076 20052
rect 20031 20012 20076 20040
rect 20070 20000 20076 20012
rect 20128 20000 20134 20052
rect 22094 20000 22100 20052
rect 22152 20040 22158 20052
rect 22465 20043 22523 20049
rect 22465 20040 22477 20043
rect 22152 20012 22477 20040
rect 22152 20000 22158 20012
rect 22465 20009 22477 20012
rect 22511 20009 22523 20043
rect 24026 20040 24032 20052
rect 23987 20012 24032 20040
rect 22465 20003 22523 20009
rect 24026 20000 24032 20012
rect 24084 20000 24090 20052
rect 24210 20000 24216 20052
rect 24268 20040 24274 20052
rect 25041 20043 25099 20049
rect 25041 20040 25053 20043
rect 24268 20012 25053 20040
rect 24268 20000 24274 20012
rect 25041 20009 25053 20012
rect 25087 20009 25099 20043
rect 25041 20003 25099 20009
rect 1949 19975 2007 19981
rect 1949 19941 1961 19975
rect 1995 19972 2007 19975
rect 2498 19972 2504 19984
rect 1995 19944 2504 19972
rect 1995 19941 2007 19944
rect 1949 19935 2007 19941
rect 2498 19932 2504 19944
rect 2556 19932 2562 19984
rect 2590 19932 2596 19984
rect 2648 19972 2654 19984
rect 2648 19944 4660 19972
rect 2648 19932 2654 19944
rect 4632 19913 4660 19944
rect 4798 19932 4804 19984
rect 4856 19972 4862 19984
rect 6822 19972 6828 19984
rect 4856 19944 6828 19972
rect 4856 19932 4862 19944
rect 1673 19907 1731 19913
rect 1673 19873 1685 19907
rect 1719 19904 1731 19907
rect 4617 19907 4675 19913
rect 1719 19876 3280 19904
rect 1719 19873 1731 19876
rect 1673 19867 1731 19873
rect 2314 19660 2320 19712
rect 2372 19700 2378 19712
rect 2409 19703 2467 19709
rect 2409 19700 2421 19703
rect 2372 19672 2421 19700
rect 2372 19660 2378 19672
rect 2409 19669 2421 19672
rect 2455 19669 2467 19703
rect 2866 19700 2872 19712
rect 2827 19672 2872 19700
rect 2409 19663 2467 19669
rect 2866 19660 2872 19672
rect 2924 19660 2930 19712
rect 3252 19709 3280 19876
rect 4617 19873 4629 19907
rect 4663 19904 4675 19907
rect 4982 19904 4988 19916
rect 4663 19876 4988 19904
rect 4663 19873 4675 19876
rect 4617 19867 4675 19873
rect 4982 19864 4988 19876
rect 5040 19864 5046 19916
rect 5353 19907 5411 19913
rect 5353 19873 5365 19907
rect 5399 19904 5411 19907
rect 5718 19904 5724 19916
rect 5399 19876 5724 19904
rect 5399 19873 5411 19876
rect 5353 19867 5411 19873
rect 5718 19864 5724 19876
rect 5776 19864 5782 19916
rect 5828 19913 5856 19944
rect 6822 19932 6828 19944
rect 6880 19932 6886 19984
rect 7190 19932 7196 19984
rect 7248 19972 7254 19984
rect 9401 19975 9459 19981
rect 9401 19972 9413 19975
rect 7248 19944 9413 19972
rect 7248 19932 7254 19944
rect 9401 19941 9413 19944
rect 9447 19941 9459 19975
rect 9401 19935 9459 19941
rect 11146 19932 11152 19984
rect 11204 19972 11210 19984
rect 11425 19975 11483 19981
rect 11425 19972 11437 19975
rect 11204 19944 11437 19972
rect 11204 19932 11210 19944
rect 11425 19941 11437 19944
rect 11471 19972 11483 19975
rect 12342 19972 12348 19984
rect 11471 19944 12348 19972
rect 11471 19941 11483 19944
rect 11425 19935 11483 19941
rect 12342 19932 12348 19944
rect 12400 19932 12406 19984
rect 12986 19932 12992 19984
rect 13044 19972 13050 19984
rect 14642 19972 14648 19984
rect 13044 19944 14504 19972
rect 14603 19944 14648 19972
rect 13044 19932 13050 19944
rect 6086 19913 6092 19916
rect 5813 19907 5871 19913
rect 5813 19873 5825 19907
rect 5859 19873 5871 19907
rect 6080 19904 6092 19913
rect 5999 19876 6092 19904
rect 5813 19867 5871 19873
rect 6080 19867 6092 19876
rect 6144 19904 6150 19916
rect 6638 19904 6644 19916
rect 6144 19876 6644 19904
rect 6086 19864 6092 19867
rect 6144 19864 6150 19876
rect 6638 19864 6644 19876
rect 6696 19864 6702 19916
rect 8386 19904 8392 19916
rect 8299 19876 8392 19904
rect 8386 19864 8392 19876
rect 8444 19904 8450 19916
rect 10045 19907 10103 19913
rect 10045 19904 10057 19907
rect 8444 19876 10057 19904
rect 8444 19864 8450 19876
rect 10045 19873 10057 19876
rect 10091 19873 10103 19907
rect 11698 19904 11704 19916
rect 10045 19867 10103 19873
rect 10428 19876 11704 19904
rect 3697 19839 3755 19845
rect 3697 19805 3709 19839
rect 3743 19836 3755 19839
rect 4798 19836 4804 19848
rect 3743 19808 4804 19836
rect 3743 19805 3755 19808
rect 3697 19799 3755 19805
rect 4798 19796 4804 19808
rect 4856 19836 4862 19848
rect 4893 19839 4951 19845
rect 4893 19836 4905 19839
rect 4856 19808 4905 19836
rect 4856 19796 4862 19808
rect 4893 19805 4905 19808
rect 4939 19836 4951 19839
rect 5074 19836 5080 19848
rect 4939 19808 5080 19836
rect 4939 19805 4951 19808
rect 4893 19799 4951 19805
rect 5074 19796 5080 19808
rect 5132 19796 5138 19848
rect 8018 19796 8024 19848
rect 8076 19836 8082 19848
rect 8481 19839 8539 19845
rect 8481 19836 8493 19839
rect 8076 19808 8493 19836
rect 8076 19796 8082 19808
rect 8481 19805 8493 19808
rect 8527 19805 8539 19839
rect 8662 19836 8668 19848
rect 8623 19808 8668 19836
rect 8481 19799 8539 19805
rect 8662 19796 8668 19808
rect 8720 19796 8726 19848
rect 9858 19796 9864 19848
rect 9916 19836 9922 19848
rect 10428 19836 10456 19876
rect 11698 19864 11704 19876
rect 11756 19904 11762 19916
rect 12710 19904 12716 19916
rect 11756 19876 12716 19904
rect 11756 19864 11762 19876
rect 12710 19864 12716 19876
rect 12768 19864 12774 19916
rect 13262 19913 13268 19916
rect 12897 19907 12955 19913
rect 12897 19873 12909 19907
rect 12943 19904 12955 19907
rect 13256 19904 13268 19913
rect 12943 19876 13268 19904
rect 12943 19873 12955 19876
rect 12897 19867 12955 19873
rect 13256 19867 13268 19876
rect 13320 19904 13326 19916
rect 13722 19904 13728 19916
rect 13320 19876 13728 19904
rect 13262 19864 13268 19867
rect 13320 19864 13326 19876
rect 13722 19864 13728 19876
rect 13780 19864 13786 19916
rect 14476 19904 14504 19944
rect 14642 19932 14648 19944
rect 14700 19932 14706 19984
rect 16209 19975 16267 19981
rect 16209 19941 16221 19975
rect 16255 19972 16267 19975
rect 16758 19972 16764 19984
rect 16255 19944 16764 19972
rect 16255 19941 16267 19944
rect 16209 19935 16267 19941
rect 16758 19932 16764 19944
rect 16816 19932 16822 19984
rect 21361 19975 21419 19981
rect 21361 19941 21373 19975
rect 21407 19972 21419 19975
rect 21407 19944 22416 19972
rect 21407 19941 21419 19944
rect 21361 19935 21419 19941
rect 15378 19904 15384 19916
rect 14476 19876 15384 19904
rect 15378 19864 15384 19876
rect 15436 19904 15442 19916
rect 16301 19907 16359 19913
rect 16301 19904 16313 19907
rect 15436 19876 16313 19904
rect 15436 19864 15442 19876
rect 16301 19873 16313 19876
rect 16347 19873 16359 19907
rect 16301 19867 16359 19873
rect 16390 19864 16396 19916
rect 16448 19904 16454 19916
rect 16557 19907 16615 19913
rect 16557 19904 16569 19907
rect 16448 19876 16569 19904
rect 16448 19864 16454 19876
rect 16557 19873 16569 19876
rect 16603 19873 16615 19907
rect 16557 19867 16615 19873
rect 18506 19864 18512 19916
rect 18564 19904 18570 19916
rect 18877 19907 18935 19913
rect 18877 19904 18889 19907
rect 18564 19876 18889 19904
rect 18564 19864 18570 19876
rect 18877 19873 18889 19876
rect 18923 19873 18935 19907
rect 18877 19867 18935 19873
rect 21269 19907 21327 19913
rect 21269 19873 21281 19907
rect 21315 19904 21327 19907
rect 22002 19904 22008 19916
rect 21315 19876 22008 19904
rect 21315 19873 21327 19876
rect 21269 19867 21327 19873
rect 22002 19864 22008 19876
rect 22060 19864 22066 19916
rect 9916 19808 10456 19836
rect 9916 19796 9922 19808
rect 11238 19796 11244 19848
rect 11296 19836 11302 19848
rect 11609 19839 11667 19845
rect 11609 19836 11621 19839
rect 11296 19808 11621 19836
rect 11296 19796 11302 19808
rect 11609 19805 11621 19808
rect 11655 19805 11667 19839
rect 12986 19836 12992 19848
rect 12947 19808 12992 19836
rect 11609 19799 11667 19805
rect 12986 19796 12992 19808
rect 13044 19796 13050 19848
rect 19058 19796 19064 19848
rect 19116 19836 19122 19848
rect 21542 19836 21548 19848
rect 19116 19808 19161 19836
rect 21503 19808 21548 19836
rect 19116 19796 19122 19808
rect 21542 19796 21548 19808
rect 21600 19796 21606 19848
rect 7929 19771 7987 19777
rect 7929 19737 7941 19771
rect 7975 19768 7987 19771
rect 8680 19768 8708 19796
rect 7975 19740 8708 19768
rect 7975 19737 7987 19740
rect 7929 19731 7987 19737
rect 9582 19728 9588 19780
rect 9640 19768 9646 19780
rect 12069 19771 12127 19777
rect 12069 19768 12081 19771
rect 9640 19740 12081 19768
rect 9640 19728 9646 19740
rect 12069 19737 12081 19740
rect 12115 19768 12127 19771
rect 12250 19768 12256 19780
rect 12115 19740 12256 19768
rect 12115 19737 12127 19740
rect 12069 19731 12127 19737
rect 12250 19728 12256 19740
rect 12308 19728 12314 19780
rect 22388 19777 22416 19944
rect 23934 19932 23940 19984
rect 23992 19972 23998 19984
rect 24397 19975 24455 19981
rect 24397 19972 24409 19975
rect 23992 19944 24409 19972
rect 23992 19932 23998 19944
rect 24397 19941 24409 19944
rect 24443 19972 24455 19975
rect 24854 19972 24860 19984
rect 24443 19944 24860 19972
rect 24443 19941 24455 19944
rect 24397 19935 24455 19941
rect 24854 19932 24860 19944
rect 24912 19932 24918 19984
rect 22830 19904 22836 19916
rect 22791 19876 22836 19904
rect 22830 19864 22836 19876
rect 22888 19864 22894 19916
rect 23474 19864 23480 19916
rect 23532 19904 23538 19916
rect 24026 19904 24032 19916
rect 23532 19876 24032 19904
rect 23532 19864 23538 19876
rect 24026 19864 24032 19876
rect 24084 19904 24090 19916
rect 24578 19904 24584 19916
rect 24084 19876 24584 19904
rect 24084 19864 24090 19876
rect 24578 19864 24584 19876
rect 24636 19864 24642 19916
rect 25038 19864 25044 19916
rect 25096 19904 25102 19916
rect 25409 19907 25467 19913
rect 25409 19904 25421 19907
rect 25096 19876 25421 19904
rect 25096 19864 25102 19876
rect 25409 19873 25421 19876
rect 25455 19873 25467 19907
rect 25409 19867 25467 19873
rect 22922 19836 22928 19848
rect 22883 19808 22928 19836
rect 22922 19796 22928 19808
rect 22980 19796 22986 19848
rect 23109 19839 23167 19845
rect 23109 19805 23121 19839
rect 23155 19836 23167 19839
rect 23198 19836 23204 19848
rect 23155 19808 23204 19836
rect 23155 19805 23167 19808
rect 23109 19799 23167 19805
rect 23198 19796 23204 19808
rect 23256 19796 23262 19848
rect 23290 19796 23296 19848
rect 23348 19836 23354 19848
rect 24486 19836 24492 19848
rect 23348 19808 24492 19836
rect 23348 19796 23354 19808
rect 24486 19796 24492 19808
rect 24544 19796 24550 19848
rect 24673 19839 24731 19845
rect 24673 19805 24685 19839
rect 24719 19836 24731 19839
rect 24762 19836 24768 19848
rect 24719 19808 24768 19836
rect 24719 19805 24731 19808
rect 24673 19799 24731 19805
rect 22373 19771 22431 19777
rect 22373 19737 22385 19771
rect 22419 19768 22431 19771
rect 23382 19768 23388 19780
rect 22419 19740 23388 19768
rect 22419 19737 22431 19740
rect 22373 19731 22431 19737
rect 23382 19728 23388 19740
rect 23440 19728 23446 19780
rect 24688 19768 24716 19799
rect 24762 19796 24768 19808
rect 24820 19796 24826 19848
rect 24320 19740 24716 19768
rect 3237 19703 3295 19709
rect 3237 19669 3249 19703
rect 3283 19700 3295 19703
rect 4246 19700 4252 19712
rect 3283 19672 4252 19700
rect 3283 19669 3295 19672
rect 3237 19663 3295 19669
rect 4246 19660 4252 19672
rect 4304 19660 4310 19712
rect 7190 19700 7196 19712
rect 7151 19672 7196 19700
rect 7190 19660 7196 19672
rect 7248 19660 7254 19712
rect 9122 19700 9128 19712
rect 9083 19672 9128 19700
rect 9122 19660 9128 19672
rect 9180 19660 9186 19712
rect 10873 19703 10931 19709
rect 10873 19669 10885 19703
rect 10919 19700 10931 19703
rect 11238 19700 11244 19712
rect 10919 19672 11244 19700
rect 10919 19669 10931 19672
rect 10873 19663 10931 19669
rect 11238 19660 11244 19672
rect 11296 19660 11302 19712
rect 15838 19700 15844 19712
rect 15799 19672 15844 19700
rect 15838 19660 15844 19672
rect 15896 19700 15902 19712
rect 17681 19703 17739 19709
rect 17681 19700 17693 19703
rect 15896 19672 17693 19700
rect 15896 19660 15902 19672
rect 17681 19669 17693 19672
rect 17727 19669 17739 19703
rect 18230 19700 18236 19712
rect 18191 19672 18236 19700
rect 17681 19663 17739 19669
rect 18230 19660 18236 19672
rect 18288 19660 18294 19712
rect 19426 19660 19432 19712
rect 19484 19700 19490 19712
rect 19702 19700 19708 19712
rect 19484 19672 19708 19700
rect 19484 19660 19490 19672
rect 19702 19660 19708 19672
rect 19760 19660 19766 19712
rect 20346 19700 20352 19712
rect 20307 19672 20352 19700
rect 20346 19660 20352 19672
rect 20404 19660 20410 19712
rect 20898 19700 20904 19712
rect 20859 19672 20904 19700
rect 20898 19660 20904 19672
rect 20956 19660 20962 19712
rect 21082 19660 21088 19712
rect 21140 19700 21146 19712
rect 21634 19700 21640 19712
rect 21140 19672 21640 19700
rect 21140 19660 21146 19672
rect 21634 19660 21640 19672
rect 21692 19700 21698 19712
rect 21913 19703 21971 19709
rect 21913 19700 21925 19703
rect 21692 19672 21925 19700
rect 21692 19660 21698 19672
rect 21913 19669 21925 19672
rect 21959 19669 21971 19703
rect 21913 19663 21971 19669
rect 23753 19703 23811 19709
rect 23753 19669 23765 19703
rect 23799 19700 23811 19703
rect 24320 19700 24348 19740
rect 23799 19672 24348 19700
rect 23799 19669 23811 19672
rect 23753 19663 23811 19669
rect 25222 19660 25228 19712
rect 25280 19700 25286 19712
rect 25777 19703 25835 19709
rect 25777 19700 25789 19703
rect 25280 19672 25789 19700
rect 25280 19660 25286 19672
rect 25777 19669 25789 19672
rect 25823 19669 25835 19703
rect 25777 19663 25835 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 2038 19456 2044 19508
rect 2096 19496 2102 19508
rect 2222 19496 2228 19508
rect 2096 19468 2228 19496
rect 2096 19456 2102 19468
rect 2222 19456 2228 19468
rect 2280 19456 2286 19508
rect 4706 19496 4712 19508
rect 4667 19468 4712 19496
rect 4706 19456 4712 19468
rect 4764 19456 4770 19508
rect 8386 19496 8392 19508
rect 8347 19468 8392 19496
rect 8386 19456 8392 19468
rect 8444 19456 8450 19508
rect 10778 19496 10784 19508
rect 10739 19468 10784 19496
rect 10778 19456 10784 19468
rect 10836 19456 10842 19508
rect 11514 19456 11520 19508
rect 11572 19496 11578 19508
rect 11793 19499 11851 19505
rect 11793 19496 11805 19499
rect 11572 19468 11805 19496
rect 11572 19456 11578 19468
rect 11793 19465 11805 19468
rect 11839 19465 11851 19499
rect 11793 19459 11851 19465
rect 12437 19499 12495 19505
rect 12437 19465 12449 19499
rect 12483 19496 12495 19499
rect 12526 19496 12532 19508
rect 12483 19468 12532 19496
rect 12483 19465 12495 19468
rect 12437 19459 12495 19465
rect 12526 19456 12532 19468
rect 12584 19456 12590 19508
rect 12894 19456 12900 19508
rect 12952 19496 12958 19508
rect 12952 19468 13216 19496
rect 12952 19456 12958 19468
rect 4798 19428 4804 19440
rect 4264 19400 4804 19428
rect 4264 19369 4292 19400
rect 4798 19388 4804 19400
rect 4856 19388 4862 19440
rect 6454 19388 6460 19440
rect 6512 19428 6518 19440
rect 7098 19428 7104 19440
rect 6512 19400 7104 19428
rect 6512 19388 6518 19400
rect 7098 19388 7104 19400
rect 7156 19388 7162 19440
rect 12250 19388 12256 19440
rect 12308 19428 12314 19440
rect 13188 19428 13216 19468
rect 14182 19456 14188 19508
rect 14240 19496 14246 19508
rect 14550 19496 14556 19508
rect 14240 19468 14556 19496
rect 14240 19456 14246 19468
rect 14550 19456 14556 19468
rect 14608 19456 14614 19508
rect 15657 19499 15715 19505
rect 15657 19465 15669 19499
rect 15703 19496 15715 19499
rect 16390 19496 16396 19508
rect 15703 19468 16396 19496
rect 15703 19465 15715 19468
rect 15657 19459 15715 19465
rect 16390 19456 16396 19468
rect 16448 19496 16454 19508
rect 16448 19468 16712 19496
rect 16448 19456 16454 19468
rect 15194 19428 15200 19440
rect 12308 19400 13124 19428
rect 13188 19400 15200 19428
rect 12308 19388 12314 19400
rect 2593 19363 2651 19369
rect 2593 19329 2605 19363
rect 2639 19329 2651 19363
rect 2593 19323 2651 19329
rect 4249 19363 4307 19369
rect 4249 19329 4261 19363
rect 4295 19329 4307 19363
rect 4249 19323 4307 19329
rect 5813 19363 5871 19369
rect 5813 19329 5825 19363
rect 5859 19360 5871 19363
rect 6086 19360 6092 19372
rect 5859 19332 6092 19360
rect 5859 19329 5871 19332
rect 5813 19323 5871 19329
rect 2608 19292 2636 19323
rect 6086 19320 6092 19332
rect 6144 19320 6150 19372
rect 7469 19363 7527 19369
rect 7469 19329 7481 19363
rect 7515 19360 7527 19363
rect 7650 19360 7656 19372
rect 7515 19332 7656 19360
rect 7515 19329 7527 19332
rect 7469 19323 7527 19329
rect 7650 19320 7656 19332
rect 7708 19320 7714 19372
rect 11146 19360 11152 19372
rect 10704 19332 11152 19360
rect 1872 19264 2636 19292
rect 3513 19295 3571 19301
rect 1872 19165 1900 19264
rect 3513 19261 3525 19295
rect 3559 19292 3571 19295
rect 3602 19292 3608 19304
rect 3559 19264 3608 19292
rect 3559 19261 3571 19264
rect 3513 19255 3571 19261
rect 3602 19252 3608 19264
rect 3660 19292 3666 19304
rect 3970 19292 3976 19304
rect 3660 19264 3976 19292
rect 3660 19252 3666 19264
rect 3970 19252 3976 19264
rect 4028 19252 4034 19304
rect 4065 19295 4123 19301
rect 4065 19261 4077 19295
rect 4111 19292 4123 19295
rect 4338 19292 4344 19304
rect 4111 19264 4344 19292
rect 4111 19261 4123 19264
rect 4065 19255 4123 19261
rect 4338 19252 4344 19264
rect 4396 19252 4402 19304
rect 5166 19252 5172 19304
rect 5224 19292 5230 19304
rect 5629 19295 5687 19301
rect 5629 19292 5641 19295
rect 5224 19264 5641 19292
rect 5224 19252 5230 19264
rect 5629 19261 5641 19264
rect 5675 19261 5687 19295
rect 5629 19255 5687 19261
rect 6641 19295 6699 19301
rect 6641 19261 6653 19295
rect 6687 19292 6699 19295
rect 7006 19292 7012 19304
rect 6687 19264 7012 19292
rect 6687 19261 6699 19264
rect 6641 19255 6699 19261
rect 7006 19252 7012 19264
rect 7064 19292 7070 19304
rect 7285 19295 7343 19301
rect 7285 19292 7297 19295
rect 7064 19264 7297 19292
rect 7064 19252 7070 19264
rect 7285 19261 7297 19264
rect 7331 19261 7343 19295
rect 7285 19255 7343 19261
rect 8202 19252 8208 19304
rect 8260 19292 8266 19304
rect 8573 19295 8631 19301
rect 8573 19292 8585 19295
rect 8260 19264 8585 19292
rect 8260 19252 8266 19264
rect 8573 19261 8585 19264
rect 8619 19292 8631 19295
rect 9398 19292 9404 19304
rect 8619 19264 9404 19292
rect 8619 19261 8631 19264
rect 8573 19255 8631 19261
rect 9398 19252 9404 19264
rect 9456 19252 9462 19304
rect 10226 19252 10232 19304
rect 10284 19292 10290 19304
rect 10704 19292 10732 19332
rect 11146 19320 11152 19332
rect 11204 19320 11210 19372
rect 11238 19320 11244 19372
rect 11296 19360 11302 19372
rect 11425 19363 11483 19369
rect 11425 19360 11437 19363
rect 11296 19332 11437 19360
rect 11296 19320 11302 19332
rect 11425 19329 11437 19332
rect 11471 19360 11483 19363
rect 11471 19332 11744 19360
rect 11471 19329 11483 19332
rect 11425 19323 11483 19329
rect 10284 19264 10732 19292
rect 10284 19252 10290 19264
rect 10778 19252 10784 19304
rect 10836 19292 10842 19304
rect 10962 19292 10968 19304
rect 10836 19264 10968 19292
rect 10836 19252 10842 19264
rect 10962 19252 10968 19264
rect 11020 19252 11026 19304
rect 11716 19236 11744 19332
rect 12066 19320 12072 19372
rect 12124 19320 12130 19372
rect 12161 19363 12219 19369
rect 12161 19329 12173 19363
rect 12207 19360 12219 19363
rect 12989 19363 13047 19369
rect 12989 19360 13001 19363
rect 12207 19332 13001 19360
rect 12207 19329 12219 19332
rect 12161 19323 12219 19329
rect 12989 19329 13001 19332
rect 13035 19329 13047 19363
rect 12989 19323 13047 19329
rect 12084 19236 12112 19320
rect 2774 19224 2780 19236
rect 2056 19196 2780 19224
rect 2056 19165 2084 19196
rect 2774 19184 2780 19196
rect 2832 19184 2838 19236
rect 5537 19227 5595 19233
rect 5537 19224 5549 19227
rect 3620 19196 5549 19224
rect 937 19159 995 19165
rect 937 19125 949 19159
rect 983 19156 995 19159
rect 1857 19159 1915 19165
rect 1857 19156 1869 19159
rect 983 19128 1869 19156
rect 983 19125 995 19128
rect 937 19119 995 19125
rect 1857 19125 1869 19128
rect 1903 19125 1915 19159
rect 1857 19119 1915 19125
rect 2041 19159 2099 19165
rect 2041 19125 2053 19159
rect 2087 19125 2099 19159
rect 2041 19119 2099 19125
rect 2314 19116 2320 19168
rect 2372 19156 2378 19168
rect 2409 19159 2467 19165
rect 2409 19156 2421 19159
rect 2372 19128 2421 19156
rect 2372 19116 2378 19128
rect 2409 19125 2421 19128
rect 2455 19125 2467 19159
rect 2409 19119 2467 19125
rect 2501 19159 2559 19165
rect 2501 19125 2513 19159
rect 2547 19156 2559 19159
rect 2866 19156 2872 19168
rect 2547 19128 2872 19156
rect 2547 19125 2559 19128
rect 2501 19119 2559 19125
rect 2866 19116 2872 19128
rect 2924 19116 2930 19168
rect 3050 19156 3056 19168
rect 3011 19128 3056 19156
rect 3050 19116 3056 19128
rect 3108 19116 3114 19168
rect 3620 19165 3648 19196
rect 5537 19193 5549 19196
rect 5583 19224 5595 19227
rect 6270 19224 6276 19236
rect 5583 19196 6276 19224
rect 5583 19193 5595 19196
rect 5537 19187 5595 19193
rect 6270 19184 6276 19196
rect 6328 19184 6334 19236
rect 7193 19227 7251 19233
rect 7193 19224 7205 19227
rect 6380 19196 7205 19224
rect 6380 19168 6408 19196
rect 7193 19193 7205 19196
rect 7239 19193 7251 19227
rect 7193 19187 7251 19193
rect 8294 19184 8300 19236
rect 8352 19224 8358 19236
rect 8818 19227 8876 19233
rect 8818 19224 8830 19227
rect 8352 19196 8830 19224
rect 8352 19184 8358 19196
rect 8818 19193 8830 19196
rect 8864 19193 8876 19227
rect 10689 19227 10747 19233
rect 8818 19187 8876 19193
rect 9968 19196 10640 19224
rect 3605 19159 3663 19165
rect 3605 19125 3617 19159
rect 3651 19125 3663 19159
rect 3970 19156 3976 19168
rect 3931 19128 3976 19156
rect 3605 19119 3663 19125
rect 3970 19116 3976 19128
rect 4028 19116 4034 19168
rect 4982 19156 4988 19168
rect 4943 19128 4988 19156
rect 4982 19116 4988 19128
rect 5040 19116 5046 19168
rect 5169 19159 5227 19165
rect 5169 19125 5181 19159
rect 5215 19156 5227 19159
rect 5350 19156 5356 19168
rect 5215 19128 5356 19156
rect 5215 19125 5227 19128
rect 5169 19119 5227 19125
rect 5350 19116 5356 19128
rect 5408 19116 5414 19168
rect 6181 19159 6239 19165
rect 6181 19125 6193 19159
rect 6227 19156 6239 19159
rect 6362 19156 6368 19168
rect 6227 19128 6368 19156
rect 6227 19125 6239 19128
rect 6181 19119 6239 19125
rect 6362 19116 6368 19128
rect 6420 19116 6426 19168
rect 6638 19116 6644 19168
rect 6696 19156 6702 19168
rect 6825 19159 6883 19165
rect 6825 19156 6837 19159
rect 6696 19128 6837 19156
rect 6696 19116 6702 19128
rect 6825 19125 6837 19128
rect 6871 19125 6883 19159
rect 8018 19156 8024 19168
rect 7979 19128 8024 19156
rect 6825 19119 6883 19125
rect 8018 19116 8024 19128
rect 8076 19116 8082 19168
rect 9968 19165 9996 19196
rect 9953 19159 10011 19165
rect 9953 19125 9965 19159
rect 9999 19125 10011 19159
rect 10612 19156 10640 19196
rect 10689 19193 10701 19227
rect 10735 19224 10747 19227
rect 11149 19227 11207 19233
rect 11149 19224 11161 19227
rect 10735 19196 11161 19224
rect 10735 19193 10747 19196
rect 10689 19187 10747 19193
rect 11149 19193 11161 19196
rect 11195 19193 11207 19227
rect 11149 19187 11207 19193
rect 10962 19156 10968 19168
rect 10612 19128 10968 19156
rect 9953 19119 10011 19125
rect 10962 19116 10968 19128
rect 11020 19116 11026 19168
rect 11164 19156 11192 19187
rect 11238 19184 11244 19236
rect 11296 19224 11302 19236
rect 11296 19196 11341 19224
rect 11296 19184 11302 19196
rect 11698 19184 11704 19236
rect 11756 19184 11762 19236
rect 12066 19184 12072 19236
rect 12124 19184 12130 19236
rect 11790 19156 11796 19168
rect 11164 19128 11796 19156
rect 11790 19116 11796 19128
rect 11848 19116 11854 19168
rect 11974 19116 11980 19168
rect 12032 19156 12038 19168
rect 12176 19156 12204 19323
rect 12897 19295 12955 19301
rect 12897 19261 12909 19295
rect 12943 19292 12955 19295
rect 13096 19292 13124 19400
rect 15194 19388 15200 19400
rect 15252 19388 15258 19440
rect 16684 19428 16712 19468
rect 16758 19456 16764 19508
rect 16816 19496 16822 19508
rect 18049 19499 18107 19505
rect 18049 19496 18061 19499
rect 16816 19468 18061 19496
rect 16816 19456 16822 19468
rect 18049 19465 18061 19468
rect 18095 19465 18107 19499
rect 18049 19459 18107 19465
rect 20622 19456 20628 19508
rect 20680 19496 20686 19508
rect 22465 19499 22523 19505
rect 22465 19496 22477 19499
rect 20680 19468 22477 19496
rect 20680 19456 20686 19468
rect 22465 19465 22477 19468
rect 22511 19496 22523 19499
rect 22830 19496 22836 19508
rect 22511 19468 22836 19496
rect 22511 19465 22523 19468
rect 22465 19459 22523 19465
rect 22830 19456 22836 19468
rect 22888 19456 22894 19508
rect 23658 19496 23664 19508
rect 23619 19468 23664 19496
rect 23658 19456 23664 19468
rect 23716 19456 23722 19508
rect 16684 19400 18644 19428
rect 14550 19360 14556 19372
rect 14511 19332 14556 19360
rect 14550 19320 14556 19332
rect 14608 19320 14614 19372
rect 15378 19320 15384 19372
rect 15436 19360 15442 19372
rect 18616 19369 18644 19400
rect 20070 19388 20076 19440
rect 20128 19428 20134 19440
rect 24578 19428 24584 19440
rect 20128 19400 21772 19428
rect 20128 19388 20134 19400
rect 15749 19363 15807 19369
rect 15749 19360 15761 19363
rect 15436 19332 15761 19360
rect 15436 19320 15442 19332
rect 15749 19329 15761 19332
rect 15795 19329 15807 19363
rect 15749 19323 15807 19329
rect 18601 19363 18659 19369
rect 18601 19329 18613 19363
rect 18647 19329 18659 19363
rect 18601 19323 18659 19329
rect 20165 19363 20223 19369
rect 20165 19329 20177 19363
rect 20211 19360 20223 19363
rect 20346 19360 20352 19372
rect 20211 19332 20352 19360
rect 20211 19329 20223 19332
rect 20165 19323 20223 19329
rect 12943 19264 13124 19292
rect 12943 19261 12955 19264
rect 12897 19255 12955 19261
rect 13446 19252 13452 19304
rect 13504 19292 13510 19304
rect 13814 19292 13820 19304
rect 13504 19264 13820 19292
rect 13504 19252 13510 19264
rect 13814 19252 13820 19264
rect 13872 19252 13878 19304
rect 13909 19295 13967 19301
rect 13909 19261 13921 19295
rect 13955 19292 13967 19295
rect 14090 19292 14096 19304
rect 13955 19264 14096 19292
rect 13955 19261 13967 19264
rect 13909 19255 13967 19261
rect 14090 19252 14096 19264
rect 14148 19292 14154 19304
rect 14461 19295 14519 19301
rect 14461 19292 14473 19295
rect 14148 19264 14473 19292
rect 14148 19252 14154 19264
rect 14461 19261 14473 19264
rect 14507 19261 14519 19295
rect 15286 19292 15292 19304
rect 15247 19264 15292 19292
rect 14461 19255 14519 19261
rect 15286 19252 15292 19264
rect 15344 19252 15350 19304
rect 14369 19227 14427 19233
rect 14369 19224 14381 19227
rect 13464 19196 14381 19224
rect 13464 19168 13492 19196
rect 14369 19193 14381 19196
rect 14415 19193 14427 19227
rect 14369 19187 14427 19193
rect 12032 19128 12204 19156
rect 12032 19116 12038 19128
rect 12618 19116 12624 19168
rect 12676 19156 12682 19168
rect 12805 19159 12863 19165
rect 12805 19156 12817 19159
rect 12676 19128 12817 19156
rect 12676 19116 12682 19128
rect 12805 19125 12817 19128
rect 12851 19125 12863 19159
rect 13446 19156 13452 19168
rect 13407 19128 13452 19156
rect 12805 19119 12863 19125
rect 13446 19116 13452 19128
rect 13504 19116 13510 19168
rect 13906 19116 13912 19168
rect 13964 19156 13970 19168
rect 14001 19159 14059 19165
rect 14001 19156 14013 19159
rect 13964 19128 14013 19156
rect 13964 19116 13970 19128
rect 14001 19125 14013 19128
rect 14047 19125 14059 19159
rect 15764 19156 15792 19323
rect 20346 19320 20352 19332
rect 20404 19320 20410 19372
rect 21744 19369 21772 19400
rect 24320 19400 24584 19428
rect 21729 19363 21787 19369
rect 21729 19329 21741 19363
rect 21775 19360 21787 19363
rect 21818 19360 21824 19372
rect 21775 19332 21824 19360
rect 21775 19329 21787 19332
rect 21729 19323 21787 19329
rect 21818 19320 21824 19332
rect 21876 19320 21882 19372
rect 22278 19320 22284 19372
rect 22336 19360 22342 19372
rect 23934 19360 23940 19372
rect 22336 19332 23940 19360
rect 22336 19320 22342 19332
rect 23934 19320 23940 19332
rect 23992 19320 23998 19372
rect 24320 19369 24348 19400
rect 24578 19388 24584 19400
rect 24636 19388 24642 19440
rect 24305 19363 24363 19369
rect 24305 19329 24317 19363
rect 24351 19329 24363 19363
rect 24305 19323 24363 19329
rect 15838 19252 15844 19304
rect 15896 19292 15902 19304
rect 16005 19295 16063 19301
rect 16005 19292 16017 19295
rect 15896 19264 16017 19292
rect 15896 19252 15902 19264
rect 16005 19261 16017 19264
rect 16051 19261 16063 19295
rect 16005 19255 16063 19261
rect 16574 19252 16580 19304
rect 16632 19292 16638 19304
rect 17405 19295 17463 19301
rect 17405 19292 17417 19295
rect 16632 19264 17417 19292
rect 16632 19252 16638 19264
rect 17405 19261 17417 19264
rect 17451 19292 17463 19295
rect 18417 19295 18475 19301
rect 18417 19292 18429 19295
rect 17451 19264 18429 19292
rect 17451 19261 17463 19264
rect 17405 19255 17463 19261
rect 18417 19261 18429 19264
rect 18463 19261 18475 19295
rect 18417 19255 18475 19261
rect 18966 19252 18972 19304
rect 19024 19292 19030 19304
rect 19061 19295 19119 19301
rect 19061 19292 19073 19295
rect 19024 19264 19073 19292
rect 19024 19252 19030 19264
rect 19061 19261 19073 19264
rect 19107 19261 19119 19295
rect 19061 19255 19119 19261
rect 19334 19252 19340 19304
rect 19392 19252 19398 19304
rect 19521 19295 19579 19301
rect 19521 19261 19533 19295
rect 19567 19292 19579 19295
rect 19981 19295 20039 19301
rect 19981 19292 19993 19295
rect 19567 19264 19993 19292
rect 19567 19261 19579 19264
rect 19521 19255 19579 19261
rect 19981 19261 19993 19264
rect 20027 19292 20039 19295
rect 20254 19292 20260 19304
rect 20027 19264 20260 19292
rect 20027 19261 20039 19264
rect 19981 19255 20039 19261
rect 20254 19252 20260 19264
rect 20312 19252 20318 19304
rect 20622 19252 20628 19304
rect 20680 19292 20686 19304
rect 20993 19295 21051 19301
rect 20993 19292 21005 19295
rect 20680 19264 21005 19292
rect 20680 19252 20686 19264
rect 20993 19261 21005 19264
rect 21039 19292 21051 19295
rect 21545 19295 21603 19301
rect 21545 19292 21557 19295
rect 21039 19264 21557 19292
rect 21039 19261 21051 19264
rect 20993 19255 21051 19261
rect 21545 19261 21557 19264
rect 21591 19261 21603 19295
rect 21545 19255 21603 19261
rect 22738 19252 22744 19304
rect 22796 19292 22802 19304
rect 22922 19292 22928 19304
rect 22796 19264 22928 19292
rect 22796 19252 22802 19264
rect 22922 19252 22928 19264
rect 22980 19252 22986 19304
rect 24121 19295 24179 19301
rect 24121 19261 24133 19295
rect 24167 19292 24179 19295
rect 24670 19292 24676 19304
rect 24167 19264 24676 19292
rect 24167 19261 24179 19264
rect 24121 19255 24179 19261
rect 24670 19252 24676 19264
rect 24728 19252 24734 19304
rect 24854 19252 24860 19304
rect 24912 19292 24918 19304
rect 25041 19295 25099 19301
rect 25041 19292 25053 19295
rect 24912 19264 25053 19292
rect 24912 19252 24918 19264
rect 25041 19261 25053 19264
rect 25087 19261 25099 19295
rect 25041 19255 25099 19261
rect 25225 19295 25283 19301
rect 25225 19261 25237 19295
rect 25271 19292 25283 19295
rect 25498 19292 25504 19304
rect 25271 19264 25504 19292
rect 25271 19261 25283 19264
rect 25225 19255 25283 19261
rect 25498 19252 25504 19264
rect 25556 19292 25562 19304
rect 25777 19295 25835 19301
rect 25777 19292 25789 19295
rect 25556 19264 25789 19292
rect 25556 19252 25562 19264
rect 25777 19261 25789 19264
rect 25823 19261 25835 19295
rect 26234 19292 26240 19304
rect 26195 19264 26240 19292
rect 25777 19255 25835 19261
rect 26234 19252 26240 19264
rect 26292 19252 26298 19304
rect 18230 19184 18236 19236
rect 18288 19224 18294 19236
rect 18984 19224 19012 19252
rect 18288 19196 19012 19224
rect 19352 19224 19380 19252
rect 21637 19227 21695 19233
rect 21637 19224 21649 19227
rect 19352 19196 20116 19224
rect 18288 19184 18294 19196
rect 15838 19156 15844 19168
rect 15764 19128 15844 19156
rect 14001 19119 14059 19125
rect 15838 19116 15844 19128
rect 15896 19116 15902 19168
rect 16850 19116 16856 19168
rect 16908 19156 16914 19168
rect 17129 19159 17187 19165
rect 17129 19156 17141 19159
rect 16908 19128 17141 19156
rect 16908 19116 16914 19128
rect 17129 19125 17141 19128
rect 17175 19156 17187 19159
rect 17402 19156 17408 19168
rect 17175 19128 17408 19156
rect 17175 19125 17187 19128
rect 17129 19119 17187 19125
rect 17402 19116 17408 19128
rect 17460 19116 17466 19168
rect 17678 19116 17684 19168
rect 17736 19156 17742 19168
rect 17773 19159 17831 19165
rect 17773 19156 17785 19159
rect 17736 19128 17785 19156
rect 17736 19116 17742 19128
rect 17773 19125 17785 19128
rect 17819 19156 17831 19159
rect 18509 19159 18567 19165
rect 18509 19156 18521 19159
rect 17819 19128 18521 19156
rect 17819 19125 17831 19128
rect 17773 19119 17831 19125
rect 18509 19125 18521 19128
rect 18555 19156 18567 19159
rect 18598 19156 18604 19168
rect 18555 19128 18604 19156
rect 18555 19125 18567 19128
rect 18509 19119 18567 19125
rect 18598 19116 18604 19128
rect 18656 19116 18662 19168
rect 19334 19116 19340 19168
rect 19392 19156 19398 19168
rect 20088 19165 20116 19196
rect 20732 19196 21649 19224
rect 20732 19168 20760 19196
rect 21637 19193 21649 19196
rect 21683 19193 21695 19227
rect 21637 19187 21695 19193
rect 24029 19227 24087 19233
rect 24029 19193 24041 19227
rect 24075 19224 24087 19227
rect 24075 19196 25084 19224
rect 24075 19193 24087 19196
rect 24029 19187 24087 19193
rect 25056 19168 25084 19196
rect 19613 19159 19671 19165
rect 19613 19156 19625 19159
rect 19392 19128 19625 19156
rect 19392 19116 19398 19128
rect 19613 19125 19625 19128
rect 19659 19125 19671 19159
rect 19613 19119 19671 19125
rect 20073 19159 20131 19165
rect 20073 19125 20085 19159
rect 20119 19156 20131 19159
rect 20254 19156 20260 19168
rect 20119 19128 20260 19156
rect 20119 19125 20131 19128
rect 20073 19119 20131 19125
rect 20254 19116 20260 19128
rect 20312 19116 20318 19168
rect 20714 19156 20720 19168
rect 20675 19128 20720 19156
rect 20714 19116 20720 19128
rect 20772 19116 20778 19168
rect 21174 19156 21180 19168
rect 21135 19128 21180 19156
rect 21174 19116 21180 19128
rect 21232 19116 21238 19168
rect 23290 19116 23296 19168
rect 23348 19156 23354 19168
rect 23385 19159 23443 19165
rect 23385 19156 23397 19159
rect 23348 19128 23397 19156
rect 23348 19116 23354 19128
rect 23385 19125 23397 19128
rect 23431 19125 23443 19159
rect 24762 19156 24768 19168
rect 24723 19128 24768 19156
rect 23385 19119 23443 19125
rect 24762 19116 24768 19128
rect 24820 19116 24826 19168
rect 25038 19116 25044 19168
rect 25096 19116 25102 19168
rect 25409 19159 25467 19165
rect 25409 19125 25421 19159
rect 25455 19156 25467 19159
rect 25590 19156 25596 19168
rect 25455 19128 25596 19156
rect 25455 19125 25467 19128
rect 25409 19119 25467 19125
rect 25590 19116 25596 19128
rect 25648 19116 25654 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1854 18912 1860 18964
rect 1912 18952 1918 18964
rect 2317 18955 2375 18961
rect 2317 18952 2329 18955
rect 1912 18924 2329 18952
rect 1912 18912 1918 18924
rect 2317 18921 2329 18924
rect 2363 18952 2375 18955
rect 2777 18955 2835 18961
rect 2777 18952 2789 18955
rect 2363 18924 2789 18952
rect 2363 18921 2375 18924
rect 2317 18915 2375 18921
rect 2777 18921 2789 18924
rect 2823 18921 2835 18955
rect 2777 18915 2835 18921
rect 2869 18955 2927 18961
rect 2869 18921 2881 18955
rect 2915 18952 2927 18955
rect 2958 18952 2964 18964
rect 2915 18924 2964 18952
rect 2915 18921 2927 18924
rect 2869 18915 2927 18921
rect 2958 18912 2964 18924
rect 3016 18912 3022 18964
rect 3694 18952 3700 18964
rect 3655 18924 3700 18952
rect 3694 18912 3700 18924
rect 3752 18912 3758 18964
rect 4249 18955 4307 18961
rect 4249 18921 4261 18955
rect 4295 18921 4307 18955
rect 4706 18952 4712 18964
rect 4667 18924 4712 18952
rect 4249 18915 4307 18921
rect 1946 18844 1952 18896
rect 2004 18884 2010 18896
rect 4264 18884 4292 18915
rect 4706 18912 4712 18924
rect 4764 18912 4770 18964
rect 5353 18955 5411 18961
rect 5353 18921 5365 18955
rect 5399 18952 5411 18955
rect 5442 18952 5448 18964
rect 5399 18924 5448 18952
rect 5399 18921 5411 18924
rect 5353 18915 5411 18921
rect 5442 18912 5448 18924
rect 5500 18912 5506 18964
rect 5721 18955 5779 18961
rect 5721 18921 5733 18955
rect 5767 18952 5779 18955
rect 6178 18952 6184 18964
rect 5767 18924 6184 18952
rect 5767 18921 5779 18924
rect 5721 18915 5779 18921
rect 2004 18856 4292 18884
rect 2004 18844 2010 18856
rect 5258 18844 5264 18896
rect 5316 18884 5322 18896
rect 5736 18884 5764 18915
rect 6178 18912 6184 18924
rect 6236 18912 6242 18964
rect 7006 18952 7012 18964
rect 6748 18924 7012 18952
rect 5316 18856 5764 18884
rect 5316 18844 5322 18856
rect 6086 18844 6092 18896
rect 6144 18884 6150 18896
rect 6362 18884 6368 18896
rect 6144 18856 6368 18884
rect 6144 18844 6150 18856
rect 6362 18844 6368 18856
rect 6420 18844 6426 18896
rect 4065 18819 4123 18825
rect 4065 18785 4077 18819
rect 4111 18816 4123 18819
rect 4614 18816 4620 18828
rect 4111 18788 4620 18816
rect 4111 18785 4123 18788
rect 4065 18779 4123 18785
rect 4614 18776 4620 18788
rect 4672 18776 4678 18828
rect 5074 18776 5080 18828
rect 5132 18816 5138 18828
rect 5169 18819 5227 18825
rect 5169 18816 5181 18819
rect 5132 18788 5181 18816
rect 5132 18776 5138 18788
rect 5169 18785 5181 18788
rect 5215 18816 5227 18819
rect 6104 18816 6132 18844
rect 5215 18788 6132 18816
rect 5215 18785 5227 18788
rect 5169 18779 5227 18785
rect 3050 18748 3056 18760
rect 3011 18720 3056 18748
rect 3050 18708 3056 18720
rect 3108 18708 3114 18760
rect 5534 18708 5540 18760
rect 5592 18748 5598 18760
rect 5813 18751 5871 18757
rect 5813 18748 5825 18751
rect 5592 18720 5825 18748
rect 5592 18708 5598 18720
rect 5813 18717 5825 18720
rect 5859 18717 5871 18751
rect 5994 18748 6000 18760
rect 5955 18720 6000 18748
rect 5813 18711 5871 18717
rect 5994 18708 6000 18720
rect 6052 18708 6058 18760
rect 1118 18640 1124 18692
rect 1176 18680 1182 18692
rect 6748 18680 6776 18924
rect 7006 18912 7012 18924
rect 7064 18912 7070 18964
rect 8294 18952 8300 18964
rect 8255 18924 8300 18952
rect 8294 18912 8300 18924
rect 8352 18952 8358 18964
rect 8941 18955 8999 18961
rect 8941 18952 8953 18955
rect 8352 18924 8953 18952
rect 8352 18912 8358 18924
rect 8941 18921 8953 18924
rect 8987 18921 8999 18955
rect 8941 18915 8999 18921
rect 11054 18912 11060 18964
rect 11112 18952 11118 18964
rect 11149 18955 11207 18961
rect 11149 18952 11161 18955
rect 11112 18924 11161 18952
rect 11112 18912 11118 18924
rect 11149 18921 11161 18924
rect 11195 18921 11207 18955
rect 11149 18915 11207 18921
rect 13722 18912 13728 18964
rect 13780 18952 13786 18964
rect 14185 18955 14243 18961
rect 14185 18952 14197 18955
rect 13780 18924 14197 18952
rect 13780 18912 13786 18924
rect 14185 18921 14197 18924
rect 14231 18952 14243 18955
rect 15841 18955 15899 18961
rect 14231 18924 14780 18952
rect 14231 18921 14243 18924
rect 14185 18915 14243 18921
rect 8478 18844 8484 18896
rect 8536 18884 8542 18896
rect 8573 18887 8631 18893
rect 8573 18884 8585 18887
rect 8536 18856 8585 18884
rect 8536 18844 8542 18856
rect 8573 18853 8585 18856
rect 8619 18853 8631 18887
rect 8573 18847 8631 18853
rect 9858 18844 9864 18896
rect 9916 18884 9922 18896
rect 11514 18884 11520 18896
rect 9916 18856 11520 18884
rect 9916 18844 9922 18856
rect 11514 18844 11520 18856
rect 11572 18844 11578 18896
rect 11790 18844 11796 18896
rect 11848 18884 11854 18896
rect 11848 18856 12940 18884
rect 11848 18844 11854 18856
rect 6822 18776 6828 18828
rect 6880 18816 6886 18828
rect 7190 18825 7196 18828
rect 6917 18819 6975 18825
rect 6917 18816 6929 18819
rect 6880 18788 6929 18816
rect 6880 18776 6886 18788
rect 6917 18785 6929 18788
rect 6963 18785 6975 18819
rect 7184 18816 7196 18825
rect 7151 18788 7196 18816
rect 6917 18779 6975 18785
rect 7184 18779 7196 18788
rect 7190 18776 7196 18779
rect 7248 18776 7254 18828
rect 9950 18776 9956 18828
rect 10008 18816 10014 18828
rect 10318 18816 10324 18828
rect 10008 18788 10324 18816
rect 10008 18776 10014 18788
rect 10318 18776 10324 18788
rect 10376 18776 10382 18828
rect 10870 18776 10876 18828
rect 10928 18776 10934 18828
rect 11532 18816 11560 18844
rect 12802 18816 12808 18828
rect 11532 18788 11928 18816
rect 12763 18788 12808 18816
rect 10888 18748 10916 18776
rect 11900 18760 11928 18788
rect 12802 18776 12808 18788
rect 12860 18776 12866 18828
rect 12912 18816 12940 18856
rect 12986 18844 12992 18896
rect 13044 18893 13050 18896
rect 13044 18887 13108 18893
rect 13044 18853 13062 18887
rect 13096 18884 13108 18887
rect 14461 18887 14519 18893
rect 14461 18884 14473 18887
rect 13096 18856 14473 18884
rect 13096 18853 13108 18856
rect 13044 18847 13108 18853
rect 14461 18853 14473 18856
rect 14507 18884 14519 18887
rect 14550 18884 14556 18896
rect 14507 18856 14556 18884
rect 14507 18853 14519 18856
rect 14461 18847 14519 18853
rect 13044 18844 13050 18847
rect 14550 18844 14556 18856
rect 14608 18844 14614 18896
rect 14752 18884 14780 18924
rect 15841 18921 15853 18955
rect 15887 18952 15899 18955
rect 16298 18952 16304 18964
rect 15887 18924 16304 18952
rect 15887 18921 15899 18924
rect 15841 18915 15899 18921
rect 16298 18912 16304 18924
rect 16356 18912 16362 18964
rect 16390 18912 16396 18964
rect 16448 18952 16454 18964
rect 16577 18955 16635 18961
rect 16577 18952 16589 18955
rect 16448 18924 16589 18952
rect 16448 18912 16454 18924
rect 16577 18921 16589 18924
rect 16623 18952 16635 18955
rect 16758 18952 16764 18964
rect 16623 18924 16764 18952
rect 16623 18921 16635 18924
rect 16577 18915 16635 18921
rect 16758 18912 16764 18924
rect 16816 18912 16822 18964
rect 17678 18912 17684 18964
rect 17736 18952 17742 18964
rect 20622 18952 20628 18964
rect 17736 18924 20628 18952
rect 17736 18912 17742 18924
rect 20622 18912 20628 18924
rect 20680 18912 20686 18964
rect 21818 18912 21824 18964
rect 21876 18952 21882 18964
rect 21913 18955 21971 18961
rect 21913 18952 21925 18955
rect 21876 18924 21925 18952
rect 21876 18912 21882 18924
rect 21913 18921 21925 18924
rect 21959 18921 21971 18955
rect 21913 18915 21971 18921
rect 22186 18912 22192 18964
rect 22244 18952 22250 18964
rect 22925 18955 22983 18961
rect 22925 18952 22937 18955
rect 22244 18924 22937 18952
rect 22244 18912 22250 18924
rect 22925 18921 22937 18924
rect 22971 18921 22983 18955
rect 22925 18915 22983 18921
rect 23474 18912 23480 18964
rect 23532 18952 23538 18964
rect 23658 18952 23664 18964
rect 23532 18924 23664 18952
rect 23532 18912 23538 18924
rect 23658 18912 23664 18924
rect 23716 18912 23722 18964
rect 24029 18955 24087 18961
rect 24029 18921 24041 18955
rect 24075 18952 24087 18955
rect 24118 18952 24124 18964
rect 24075 18924 24124 18952
rect 24075 18921 24087 18924
rect 24029 18915 24087 18921
rect 24118 18912 24124 18924
rect 24176 18912 24182 18964
rect 24486 18952 24492 18964
rect 24447 18924 24492 18952
rect 24486 18912 24492 18924
rect 24544 18952 24550 18964
rect 25041 18955 25099 18961
rect 25041 18952 25053 18955
rect 24544 18924 25053 18952
rect 24544 18912 24550 18924
rect 25041 18921 25053 18924
rect 25087 18921 25099 18955
rect 25041 18915 25099 18921
rect 19058 18884 19064 18896
rect 14752 18856 19064 18884
rect 19058 18844 19064 18856
rect 19116 18844 19122 18896
rect 19337 18887 19395 18893
rect 19337 18853 19349 18887
rect 19383 18853 19395 18887
rect 19337 18847 19395 18853
rect 22373 18887 22431 18893
rect 22373 18853 22385 18887
rect 22419 18884 22431 18887
rect 23198 18884 23204 18896
rect 22419 18856 23204 18884
rect 22419 18853 22431 18856
rect 22373 18847 22431 18853
rect 15378 18816 15384 18828
rect 12912 18788 15384 18816
rect 15378 18776 15384 18788
rect 15436 18816 15442 18828
rect 15657 18819 15715 18825
rect 15657 18816 15669 18819
rect 15436 18788 15669 18816
rect 15436 18776 15442 18788
rect 15657 18785 15669 18788
rect 15703 18785 15715 18819
rect 15657 18779 15715 18785
rect 15838 18776 15844 18828
rect 15896 18816 15902 18828
rect 16761 18819 16819 18825
rect 16761 18816 16773 18819
rect 15896 18788 16773 18816
rect 15896 18776 15902 18788
rect 16761 18785 16773 18788
rect 16807 18785 16819 18819
rect 16761 18779 16819 18785
rect 11146 18748 11152 18760
rect 10888 18720 11152 18748
rect 11146 18708 11152 18720
rect 11204 18708 11210 18760
rect 11514 18708 11520 18760
rect 11572 18748 11578 18760
rect 11609 18751 11667 18757
rect 11609 18748 11621 18751
rect 11572 18720 11621 18748
rect 11572 18708 11578 18720
rect 11609 18717 11621 18720
rect 11655 18717 11667 18751
rect 11609 18711 11667 18717
rect 11698 18708 11704 18760
rect 11756 18748 11762 18760
rect 11756 18720 11801 18748
rect 11756 18708 11762 18720
rect 11882 18708 11888 18760
rect 11940 18708 11946 18760
rect 12526 18708 12532 18760
rect 12584 18708 12590 18760
rect 16482 18748 16488 18760
rect 15488 18720 16488 18748
rect 12544 18680 12572 18708
rect 1176 18652 6776 18680
rect 11624 18652 12572 18680
rect 1176 18640 1182 18652
rect 11624 18624 11652 18652
rect 13814 18640 13820 18692
rect 13872 18680 13878 18692
rect 15488 18689 15516 18720
rect 16482 18708 16488 18720
rect 16540 18708 16546 18760
rect 15473 18683 15531 18689
rect 15473 18680 15485 18683
rect 13872 18652 15485 18680
rect 13872 18640 13878 18652
rect 15473 18649 15485 18652
rect 15519 18649 15531 18683
rect 15473 18643 15531 18649
rect 1946 18612 1952 18624
rect 1907 18584 1952 18612
rect 1946 18572 1952 18584
rect 2004 18572 2010 18624
rect 2409 18615 2467 18621
rect 2409 18581 2421 18615
rect 2455 18612 2467 18615
rect 2498 18612 2504 18624
rect 2455 18584 2504 18612
rect 2455 18581 2467 18584
rect 2409 18575 2467 18581
rect 2498 18572 2504 18584
rect 2556 18572 2562 18624
rect 6822 18612 6828 18624
rect 6783 18584 6828 18612
rect 6822 18572 6828 18584
rect 6880 18572 6886 18624
rect 7558 18572 7564 18624
rect 7616 18612 7622 18624
rect 9309 18615 9367 18621
rect 9309 18612 9321 18615
rect 7616 18584 9321 18612
rect 7616 18572 7622 18584
rect 9309 18581 9321 18584
rect 9355 18581 9367 18615
rect 9858 18612 9864 18624
rect 9819 18584 9864 18612
rect 9309 18575 9367 18581
rect 9858 18572 9864 18584
rect 9916 18572 9922 18624
rect 10318 18612 10324 18624
rect 10279 18584 10324 18612
rect 10318 18572 10324 18584
rect 10376 18572 10382 18624
rect 10873 18615 10931 18621
rect 10873 18581 10885 18615
rect 10919 18612 10931 18615
rect 10962 18612 10968 18624
rect 10919 18584 10968 18612
rect 10919 18581 10931 18584
rect 10873 18575 10931 18581
rect 10962 18572 10968 18584
rect 11020 18612 11026 18624
rect 11606 18612 11612 18624
rect 11020 18584 11612 18612
rect 11020 18572 11026 18584
rect 11606 18572 11612 18584
rect 11664 18572 11670 18624
rect 12526 18612 12532 18624
rect 12487 18584 12532 18612
rect 12526 18572 12532 18584
rect 12584 18572 12590 18624
rect 14826 18612 14832 18624
rect 14787 18584 14832 18612
rect 14826 18572 14832 18584
rect 14884 18572 14890 18624
rect 16298 18612 16304 18624
rect 16259 18584 16304 18612
rect 16298 18572 16304 18584
rect 16356 18572 16362 18624
rect 16776 18612 16804 18779
rect 16850 18776 16856 18828
rect 16908 18816 16914 18828
rect 17017 18819 17075 18825
rect 17017 18816 17029 18819
rect 16908 18788 17029 18816
rect 16908 18776 16914 18788
rect 17017 18785 17029 18788
rect 17063 18785 17075 18819
rect 17017 18779 17075 18785
rect 19352 18680 19380 18847
rect 23198 18844 23204 18856
rect 23256 18844 23262 18896
rect 23934 18844 23940 18896
rect 23992 18884 23998 18896
rect 24397 18887 24455 18893
rect 24397 18884 24409 18887
rect 23992 18856 24409 18884
rect 23992 18844 23998 18856
rect 24397 18853 24409 18856
rect 24443 18853 24455 18887
rect 24397 18847 24455 18853
rect 19426 18776 19432 18828
rect 19484 18816 19490 18828
rect 21269 18819 21327 18825
rect 19484 18788 19529 18816
rect 19484 18776 19490 18788
rect 21269 18785 21281 18819
rect 21315 18816 21327 18819
rect 21818 18816 21824 18828
rect 21315 18788 21824 18816
rect 21315 18785 21327 18788
rect 21269 18779 21327 18785
rect 21818 18776 21824 18788
rect 21876 18776 21882 18828
rect 22094 18776 22100 18828
rect 22152 18816 22158 18828
rect 22833 18819 22891 18825
rect 22152 18788 22508 18816
rect 22152 18776 22158 18788
rect 19518 18748 19524 18760
rect 19479 18720 19524 18748
rect 19518 18708 19524 18720
rect 19576 18708 19582 18760
rect 21358 18748 21364 18760
rect 21319 18720 21364 18748
rect 21358 18708 21364 18720
rect 21416 18708 21422 18760
rect 21545 18751 21603 18757
rect 21545 18717 21557 18751
rect 21591 18748 21603 18751
rect 21634 18748 21640 18760
rect 21591 18720 21640 18748
rect 21591 18717 21603 18720
rect 21545 18711 21603 18717
rect 21634 18708 21640 18720
rect 21692 18708 21698 18760
rect 19426 18680 19432 18692
rect 19352 18652 19432 18680
rect 19426 18640 19432 18652
rect 19484 18640 19490 18692
rect 20901 18683 20959 18689
rect 20901 18649 20913 18683
rect 20947 18680 20959 18683
rect 21910 18680 21916 18692
rect 20947 18652 21916 18680
rect 20947 18649 20959 18652
rect 20901 18643 20959 18649
rect 21910 18640 21916 18652
rect 21968 18640 21974 18692
rect 22480 18689 22508 18788
rect 22833 18785 22845 18819
rect 22879 18816 22891 18819
rect 23474 18816 23480 18828
rect 22879 18788 23480 18816
rect 22879 18785 22891 18788
rect 22833 18779 22891 18785
rect 23474 18776 23480 18788
rect 23532 18776 23538 18828
rect 24412 18816 24440 18847
rect 24670 18844 24676 18896
rect 24728 18884 24734 18896
rect 25409 18887 25467 18893
rect 25409 18884 25421 18887
rect 24728 18856 25421 18884
rect 24728 18844 24734 18856
rect 25409 18853 25421 18856
rect 25455 18853 25467 18887
rect 25409 18847 25467 18853
rect 25038 18816 25044 18828
rect 24412 18788 25044 18816
rect 25038 18776 25044 18788
rect 25096 18776 25102 18828
rect 23106 18748 23112 18760
rect 23067 18720 23112 18748
rect 23106 18708 23112 18720
rect 23164 18708 23170 18760
rect 23290 18708 23296 18760
rect 23348 18748 23354 18760
rect 24581 18751 24639 18757
rect 24581 18748 24593 18751
rect 23348 18720 24593 18748
rect 23348 18708 23354 18720
rect 24581 18717 24593 18720
rect 24627 18748 24639 18751
rect 24670 18748 24676 18760
rect 24627 18720 24676 18748
rect 24627 18717 24639 18720
rect 24581 18711 24639 18717
rect 24670 18708 24676 18720
rect 24728 18708 24734 18760
rect 22465 18683 22523 18689
rect 22465 18649 22477 18683
rect 22511 18649 22523 18683
rect 22465 18643 22523 18649
rect 17402 18612 17408 18624
rect 16776 18584 17408 18612
rect 17402 18572 17408 18584
rect 17460 18572 17466 18624
rect 18138 18612 18144 18624
rect 18099 18584 18144 18612
rect 18138 18572 18144 18584
rect 18196 18572 18202 18624
rect 18506 18612 18512 18624
rect 18467 18584 18512 18612
rect 18506 18572 18512 18584
rect 18564 18572 18570 18624
rect 18966 18612 18972 18624
rect 18927 18584 18972 18612
rect 18966 18572 18972 18584
rect 19024 18572 19030 18624
rect 20073 18615 20131 18621
rect 20073 18581 20085 18615
rect 20119 18612 20131 18615
rect 20254 18612 20260 18624
rect 20119 18584 20260 18612
rect 20119 18581 20131 18584
rect 20073 18575 20131 18581
rect 20254 18572 20260 18584
rect 20312 18572 20318 18624
rect 20717 18615 20775 18621
rect 20717 18581 20729 18615
rect 20763 18612 20775 18615
rect 20806 18612 20812 18624
rect 20763 18584 20812 18612
rect 20763 18581 20775 18584
rect 20717 18575 20775 18581
rect 20806 18572 20812 18584
rect 20864 18612 20870 18624
rect 21542 18612 21548 18624
rect 20864 18584 21548 18612
rect 20864 18572 20870 18584
rect 21542 18572 21548 18584
rect 21600 18572 21606 18624
rect 22278 18572 22284 18624
rect 22336 18612 22342 18624
rect 24946 18612 24952 18624
rect 22336 18584 24952 18612
rect 22336 18572 22342 18584
rect 24946 18572 24952 18584
rect 25004 18572 25010 18624
rect 25222 18572 25228 18624
rect 25280 18612 25286 18624
rect 25869 18615 25927 18621
rect 25869 18612 25881 18615
rect 25280 18584 25881 18612
rect 25280 18572 25286 18584
rect 25869 18581 25881 18584
rect 25915 18612 25927 18615
rect 26234 18612 26240 18624
rect 25915 18584 26240 18612
rect 25915 18581 25927 18584
rect 25869 18575 25927 18581
rect 26234 18572 26240 18584
rect 26292 18572 26298 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 2958 18368 2964 18420
rect 3016 18408 3022 18420
rect 3053 18411 3111 18417
rect 3053 18408 3065 18411
rect 3016 18380 3065 18408
rect 3016 18368 3022 18380
rect 3053 18377 3065 18380
rect 3099 18377 3111 18411
rect 4614 18408 4620 18420
rect 4575 18380 4620 18408
rect 3053 18371 3111 18377
rect 4614 18368 4620 18380
rect 4672 18368 4678 18420
rect 5074 18408 5080 18420
rect 5035 18380 5080 18408
rect 5074 18368 5080 18380
rect 5132 18368 5138 18420
rect 5994 18368 6000 18420
rect 6052 18408 6058 18420
rect 6273 18411 6331 18417
rect 6273 18408 6285 18411
rect 6052 18380 6285 18408
rect 6052 18368 6058 18380
rect 6273 18377 6285 18380
rect 6319 18408 6331 18411
rect 7190 18408 7196 18420
rect 6319 18380 7196 18408
rect 6319 18377 6331 18380
rect 6273 18371 6331 18377
rect 7190 18368 7196 18380
rect 7248 18368 7254 18420
rect 9306 18368 9312 18420
rect 9364 18408 9370 18420
rect 9364 18380 11091 18408
rect 9364 18368 9370 18380
rect 842 18300 848 18352
rect 900 18340 906 18352
rect 3421 18343 3479 18349
rect 3421 18340 3433 18343
rect 900 18312 3433 18340
rect 900 18300 906 18312
rect 3421 18309 3433 18312
rect 3467 18309 3479 18343
rect 3421 18303 3479 18309
rect 1946 18232 1952 18284
rect 2004 18272 2010 18284
rect 2590 18272 2596 18284
rect 2004 18244 2596 18272
rect 2004 18232 2010 18244
rect 2590 18232 2596 18244
rect 2648 18232 2654 18284
rect 1578 18164 1584 18216
rect 1636 18204 1642 18216
rect 3436 18204 3464 18303
rect 4249 18275 4307 18281
rect 4249 18241 4261 18275
rect 4295 18272 4307 18275
rect 4338 18272 4344 18284
rect 4295 18244 4344 18272
rect 4295 18241 4307 18244
rect 4249 18235 4307 18241
rect 4338 18232 4344 18244
rect 4396 18272 4402 18284
rect 4706 18272 4712 18284
rect 4396 18244 4712 18272
rect 4396 18232 4402 18244
rect 4706 18232 4712 18244
rect 4764 18232 4770 18284
rect 5092 18272 5120 18368
rect 7006 18340 7012 18352
rect 6967 18312 7012 18340
rect 7006 18300 7012 18312
rect 7064 18300 7070 18352
rect 7926 18300 7932 18352
rect 7984 18340 7990 18352
rect 8294 18340 8300 18352
rect 7984 18312 8300 18340
rect 7984 18300 7990 18312
rect 8294 18300 8300 18312
rect 8352 18340 8358 18352
rect 11063 18340 11091 18380
rect 12986 18368 12992 18420
rect 13044 18408 13050 18420
rect 13446 18408 13452 18420
rect 13044 18380 13452 18408
rect 13044 18368 13050 18380
rect 13446 18368 13452 18380
rect 13504 18368 13510 18420
rect 13998 18408 14004 18420
rect 13959 18380 14004 18408
rect 13998 18368 14004 18380
rect 14056 18368 14062 18420
rect 15378 18368 15384 18420
rect 15436 18408 15442 18420
rect 15657 18411 15715 18417
rect 15657 18408 15669 18411
rect 15436 18380 15669 18408
rect 15436 18368 15442 18380
rect 15657 18377 15669 18380
rect 15703 18408 15715 18411
rect 15841 18411 15899 18417
rect 15841 18408 15853 18411
rect 15703 18380 15853 18408
rect 15703 18377 15715 18380
rect 15657 18371 15715 18377
rect 15841 18377 15853 18380
rect 15887 18377 15899 18411
rect 15841 18371 15899 18377
rect 15930 18368 15936 18420
rect 15988 18408 15994 18420
rect 16209 18411 16267 18417
rect 16209 18408 16221 18411
rect 15988 18380 16221 18408
rect 15988 18368 15994 18380
rect 16209 18377 16221 18380
rect 16255 18377 16267 18411
rect 17678 18408 17684 18420
rect 16209 18371 16267 18377
rect 16316 18380 17684 18408
rect 12250 18340 12256 18352
rect 8352 18312 9168 18340
rect 11063 18312 12256 18340
rect 8352 18300 8358 18312
rect 5721 18275 5779 18281
rect 5721 18272 5733 18275
rect 5092 18244 5733 18272
rect 5721 18241 5733 18244
rect 5767 18241 5779 18275
rect 5721 18235 5779 18241
rect 6822 18232 6828 18284
rect 6880 18272 6886 18284
rect 7466 18272 7472 18284
rect 6880 18244 7472 18272
rect 6880 18232 6886 18244
rect 7466 18232 7472 18244
rect 7524 18232 7530 18284
rect 7561 18275 7619 18281
rect 7561 18241 7573 18275
rect 7607 18241 7619 18275
rect 7561 18235 7619 18241
rect 8481 18275 8539 18281
rect 8481 18241 8493 18275
rect 8527 18272 8539 18275
rect 9030 18272 9036 18284
rect 8527 18244 9036 18272
rect 8527 18241 8539 18244
rect 8481 18235 8539 18241
rect 3878 18204 3884 18216
rect 1636 18176 2544 18204
rect 3436 18176 3884 18204
rect 1636 18164 1642 18176
rect 2409 18139 2467 18145
rect 2409 18136 2421 18139
rect 1872 18108 2421 18136
rect 1486 18028 1492 18080
rect 1544 18068 1550 18080
rect 1872 18077 1900 18108
rect 2409 18105 2421 18108
rect 2455 18105 2467 18139
rect 2516 18136 2544 18176
rect 3878 18164 3884 18176
rect 3936 18204 3942 18216
rect 3973 18207 4031 18213
rect 3973 18204 3985 18207
rect 3936 18176 3985 18204
rect 3936 18164 3942 18176
rect 3973 18173 3985 18176
rect 4019 18173 4031 18207
rect 3973 18167 4031 18173
rect 4062 18164 4068 18216
rect 4120 18204 4126 18216
rect 4522 18204 4528 18216
rect 4120 18176 4528 18204
rect 4120 18164 4126 18176
rect 4522 18164 4528 18176
rect 4580 18164 4586 18216
rect 6641 18207 6699 18213
rect 6641 18173 6653 18207
rect 6687 18204 6699 18207
rect 7576 18204 7604 18235
rect 9030 18232 9036 18244
rect 9088 18232 9094 18284
rect 9140 18281 9168 18312
rect 12250 18300 12256 18312
rect 12308 18300 12314 18352
rect 13722 18300 13728 18352
rect 13780 18340 13786 18352
rect 16316 18340 16344 18380
rect 17678 18368 17684 18380
rect 17736 18368 17742 18420
rect 17954 18368 17960 18420
rect 18012 18408 18018 18420
rect 18049 18411 18107 18417
rect 18049 18408 18061 18411
rect 18012 18380 18061 18408
rect 18012 18368 18018 18380
rect 18049 18377 18061 18380
rect 18095 18377 18107 18411
rect 18049 18371 18107 18377
rect 19613 18411 19671 18417
rect 19613 18377 19625 18411
rect 19659 18408 19671 18411
rect 21358 18408 21364 18420
rect 19659 18380 21364 18408
rect 19659 18377 19671 18380
rect 19613 18371 19671 18377
rect 21358 18368 21364 18380
rect 21416 18368 21422 18420
rect 23382 18368 23388 18420
rect 23440 18408 23446 18420
rect 23661 18411 23719 18417
rect 23661 18408 23673 18411
rect 23440 18380 23673 18408
rect 23440 18368 23446 18380
rect 23661 18377 23673 18380
rect 23707 18377 23719 18411
rect 23661 18371 23719 18377
rect 23750 18368 23756 18420
rect 23808 18408 23814 18420
rect 24946 18408 24952 18420
rect 23808 18380 24952 18408
rect 23808 18368 23814 18380
rect 24946 18368 24952 18380
rect 25004 18368 25010 18420
rect 13780 18312 16344 18340
rect 13780 18300 13786 18312
rect 16574 18300 16580 18352
rect 16632 18340 16638 18352
rect 22094 18340 22100 18352
rect 16632 18312 22100 18340
rect 16632 18300 16638 18312
rect 22094 18300 22100 18312
rect 22152 18340 22158 18352
rect 22278 18340 22284 18352
rect 22152 18312 22284 18340
rect 22152 18300 22158 18312
rect 22278 18300 22284 18312
rect 22336 18300 22342 18352
rect 23106 18300 23112 18352
rect 23164 18340 23170 18352
rect 24670 18340 24676 18352
rect 23164 18312 24256 18340
rect 24631 18312 24676 18340
rect 23164 18300 23170 18312
rect 9125 18275 9183 18281
rect 9125 18241 9137 18275
rect 9171 18241 9183 18275
rect 9861 18275 9919 18281
rect 9861 18272 9873 18275
rect 9125 18235 9183 18241
rect 9324 18244 9873 18272
rect 8202 18204 8208 18216
rect 6687 18176 8208 18204
rect 6687 18173 6699 18176
rect 6641 18167 6699 18173
rect 8202 18164 8208 18176
rect 8260 18164 8266 18216
rect 8570 18164 8576 18216
rect 8628 18204 8634 18216
rect 8941 18207 8999 18213
rect 8941 18204 8953 18207
rect 8628 18176 8953 18204
rect 8628 18164 8634 18176
rect 8941 18173 8953 18176
rect 8987 18204 8999 18207
rect 9324 18204 9352 18244
rect 9861 18241 9873 18244
rect 9907 18241 9919 18275
rect 9861 18235 9919 18241
rect 10045 18275 10103 18281
rect 10045 18241 10057 18275
rect 10091 18272 10103 18275
rect 10091 18244 10272 18272
rect 10091 18241 10103 18244
rect 10045 18235 10103 18241
rect 8987 18176 9352 18204
rect 8987 18173 8999 18176
rect 8941 18167 8999 18173
rect 9398 18164 9404 18216
rect 9456 18204 9462 18216
rect 10137 18207 10195 18213
rect 10137 18204 10149 18207
rect 9456 18176 10149 18204
rect 9456 18164 9462 18176
rect 10137 18173 10149 18176
rect 10183 18173 10195 18207
rect 10244 18204 10272 18244
rect 12802 18232 12808 18284
rect 12860 18272 12866 18284
rect 12989 18275 13047 18281
rect 12989 18272 13001 18275
rect 12860 18244 13001 18272
rect 12860 18232 12866 18244
rect 12989 18241 13001 18244
rect 13035 18241 13047 18275
rect 14550 18272 14556 18284
rect 14511 18244 14556 18272
rect 12989 18235 13047 18241
rect 14550 18232 14556 18244
rect 14608 18232 14614 18284
rect 16758 18272 16764 18284
rect 16719 18244 16764 18272
rect 16758 18232 16764 18244
rect 16816 18232 16822 18284
rect 18693 18275 18751 18281
rect 18693 18241 18705 18275
rect 18739 18272 18751 18275
rect 19058 18272 19064 18284
rect 18739 18244 19064 18272
rect 18739 18241 18751 18244
rect 18693 18235 18751 18241
rect 19058 18232 19064 18244
rect 19116 18272 19122 18284
rect 19337 18275 19395 18281
rect 19337 18272 19349 18275
rect 19116 18244 19349 18272
rect 19116 18232 19122 18244
rect 19337 18241 19349 18244
rect 19383 18241 19395 18275
rect 19337 18235 19395 18241
rect 19521 18275 19579 18281
rect 19521 18241 19533 18275
rect 19567 18272 19579 18275
rect 19610 18272 19616 18284
rect 19567 18244 19616 18272
rect 19567 18241 19579 18244
rect 19521 18235 19579 18241
rect 19610 18232 19616 18244
rect 19668 18232 19674 18284
rect 20257 18275 20315 18281
rect 20257 18241 20269 18275
rect 20303 18272 20315 18275
rect 20346 18272 20352 18284
rect 20303 18244 20352 18272
rect 20303 18241 20315 18244
rect 20257 18235 20315 18241
rect 20346 18232 20352 18244
rect 20404 18272 20410 18284
rect 21821 18275 21879 18281
rect 21821 18272 21833 18275
rect 20404 18244 21833 18272
rect 20404 18232 20410 18244
rect 21821 18241 21833 18244
rect 21867 18272 21879 18275
rect 21867 18244 22968 18272
rect 21867 18241 21879 18244
rect 21821 18235 21879 18241
rect 10404 18207 10462 18213
rect 10404 18204 10416 18207
rect 10244 18176 10416 18204
rect 10137 18167 10195 18173
rect 10404 18173 10416 18176
rect 10450 18204 10462 18207
rect 11238 18204 11244 18216
rect 10450 18176 11244 18204
rect 10450 18173 10462 18176
rect 10404 18167 10462 18173
rect 11238 18164 11244 18176
rect 11296 18164 11302 18216
rect 11514 18164 11520 18216
rect 11572 18204 11578 18216
rect 11793 18207 11851 18213
rect 11793 18204 11805 18207
rect 11572 18176 11805 18204
rect 11572 18164 11578 18176
rect 11793 18173 11805 18176
rect 11839 18173 11851 18207
rect 11793 18167 11851 18173
rect 13906 18164 13912 18216
rect 13964 18204 13970 18216
rect 14461 18207 14519 18213
rect 14461 18204 14473 18207
rect 13964 18176 14473 18204
rect 13964 18164 13970 18176
rect 14461 18173 14473 18176
rect 14507 18173 14519 18207
rect 19242 18204 19248 18216
rect 14461 18167 14519 18173
rect 18524 18176 19248 18204
rect 5537 18139 5595 18145
rect 5537 18136 5549 18139
rect 2516 18108 5549 18136
rect 2409 18099 2467 18105
rect 5537 18105 5549 18108
rect 5583 18136 5595 18139
rect 7377 18139 7435 18145
rect 5583 18108 5856 18136
rect 5583 18105 5595 18108
rect 5537 18099 5595 18105
rect 1857 18071 1915 18077
rect 1857 18068 1869 18071
rect 1544 18040 1869 18068
rect 1544 18028 1550 18040
rect 1857 18037 1869 18040
rect 1903 18037 1915 18071
rect 2038 18068 2044 18080
rect 1999 18040 2044 18068
rect 1857 18031 1915 18037
rect 2038 18028 2044 18040
rect 2096 18028 2102 18080
rect 2222 18028 2228 18080
rect 2280 18068 2286 18080
rect 2501 18071 2559 18077
rect 2501 18068 2513 18071
rect 2280 18040 2513 18068
rect 2280 18028 2286 18040
rect 2501 18037 2513 18040
rect 2547 18068 2559 18071
rect 2682 18068 2688 18080
rect 2547 18040 2688 18068
rect 2547 18037 2559 18040
rect 2501 18031 2559 18037
rect 2682 18028 2688 18040
rect 2740 18028 2746 18080
rect 3605 18071 3663 18077
rect 3605 18037 3617 18071
rect 3651 18068 3663 18071
rect 3878 18068 3884 18080
rect 3651 18040 3884 18068
rect 3651 18037 3663 18040
rect 3605 18031 3663 18037
rect 3878 18028 3884 18040
rect 3936 18028 3942 18080
rect 5169 18071 5227 18077
rect 5169 18037 5181 18071
rect 5215 18068 5227 18071
rect 5442 18068 5448 18080
rect 5215 18040 5448 18068
rect 5215 18037 5227 18040
rect 5169 18031 5227 18037
rect 5442 18028 5448 18040
rect 5500 18028 5506 18080
rect 5626 18028 5632 18080
rect 5684 18068 5690 18080
rect 5828 18068 5856 18108
rect 7377 18105 7389 18139
rect 7423 18136 7435 18139
rect 7423 18108 9720 18136
rect 7423 18105 7435 18108
rect 7377 18099 7435 18105
rect 7558 18068 7564 18080
rect 5684 18040 5729 18068
rect 5828 18040 7564 18068
rect 5684 18028 5690 18040
rect 7558 18028 7564 18040
rect 7616 18028 7622 18080
rect 7926 18028 7932 18080
rect 7984 18068 7990 18080
rect 8021 18071 8079 18077
rect 8021 18068 8033 18071
rect 7984 18040 8033 18068
rect 7984 18028 7990 18040
rect 8021 18037 8033 18040
rect 8067 18037 8079 18071
rect 8570 18068 8576 18080
rect 8531 18040 8576 18068
rect 8021 18031 8079 18037
rect 8570 18028 8576 18040
rect 8628 18028 8634 18080
rect 9692 18077 9720 18108
rect 10686 18096 10692 18148
rect 10744 18136 10750 18148
rect 10778 18136 10784 18148
rect 10744 18108 10784 18136
rect 10744 18096 10750 18108
rect 10778 18096 10784 18108
rect 10836 18096 10842 18148
rect 11054 18136 11060 18148
rect 10888 18108 11060 18136
rect 9677 18071 9735 18077
rect 9677 18037 9689 18071
rect 9723 18068 9735 18071
rect 9766 18068 9772 18080
rect 9723 18040 9772 18068
rect 9723 18037 9735 18040
rect 9677 18031 9735 18037
rect 9766 18028 9772 18040
rect 9824 18028 9830 18080
rect 9861 18071 9919 18077
rect 9861 18037 9873 18071
rect 9907 18068 9919 18071
rect 10888 18068 10916 18108
rect 11054 18096 11060 18108
rect 11112 18096 11118 18148
rect 12897 18139 12955 18145
rect 12176 18108 12848 18136
rect 12176 18080 12204 18108
rect 9907 18040 10916 18068
rect 9907 18037 9919 18040
rect 9861 18031 9919 18037
rect 10962 18028 10968 18080
rect 11020 18068 11026 18080
rect 11517 18071 11575 18077
rect 11517 18068 11529 18071
rect 11020 18040 11529 18068
rect 11020 18028 11026 18040
rect 11517 18037 11529 18040
rect 11563 18068 11575 18071
rect 11698 18068 11704 18080
rect 11563 18040 11704 18068
rect 11563 18037 11575 18040
rect 11517 18031 11575 18037
rect 11698 18028 11704 18040
rect 11756 18028 11762 18080
rect 12158 18068 12164 18080
rect 12119 18040 12164 18068
rect 12158 18028 12164 18040
rect 12216 18028 12222 18080
rect 12434 18068 12440 18080
rect 12395 18040 12440 18068
rect 12434 18028 12440 18040
rect 12492 18028 12498 18080
rect 12820 18077 12848 18108
rect 12897 18105 12909 18139
rect 12943 18136 12955 18139
rect 12943 18108 15148 18136
rect 12943 18105 12955 18108
rect 12897 18099 12955 18105
rect 15120 18080 15148 18108
rect 15378 18096 15384 18148
rect 15436 18136 15442 18148
rect 16025 18139 16083 18145
rect 16025 18136 16037 18139
rect 15436 18108 16037 18136
rect 15436 18096 15442 18108
rect 16025 18105 16037 18108
rect 16071 18136 16083 18139
rect 16669 18139 16727 18145
rect 16669 18136 16681 18139
rect 16071 18108 16681 18136
rect 16071 18105 16083 18108
rect 16025 18099 16083 18105
rect 16669 18105 16681 18108
rect 16715 18105 16727 18139
rect 16669 18099 16727 18105
rect 17310 18096 17316 18148
rect 17368 18136 17374 18148
rect 17773 18139 17831 18145
rect 17773 18136 17785 18139
rect 17368 18108 17785 18136
rect 17368 18096 17374 18108
rect 17773 18105 17785 18108
rect 17819 18136 17831 18139
rect 18417 18139 18475 18145
rect 18417 18136 18429 18139
rect 17819 18108 18429 18136
rect 17819 18105 17831 18108
rect 17773 18099 17831 18105
rect 18417 18105 18429 18108
rect 18463 18105 18475 18139
rect 18417 18099 18475 18105
rect 12805 18071 12863 18077
rect 12805 18037 12817 18071
rect 12851 18068 12863 18071
rect 13170 18068 13176 18080
rect 12851 18040 13176 18068
rect 12851 18037 12863 18040
rect 12805 18031 12863 18037
rect 13170 18028 13176 18040
rect 13228 18028 13234 18080
rect 13909 18071 13967 18077
rect 13909 18037 13921 18071
rect 13955 18068 13967 18071
rect 14366 18068 14372 18080
rect 13955 18040 14372 18068
rect 13955 18037 13967 18040
rect 13909 18031 13967 18037
rect 14366 18028 14372 18040
rect 14424 18028 14430 18080
rect 15102 18068 15108 18080
rect 15063 18040 15108 18068
rect 15102 18028 15108 18040
rect 15160 18028 15166 18080
rect 15838 18068 15844 18080
rect 15799 18040 15844 18068
rect 15838 18028 15844 18040
rect 15896 18028 15902 18080
rect 16574 18068 16580 18080
rect 16535 18040 16580 18068
rect 16574 18028 16580 18040
rect 16632 18028 16638 18080
rect 17126 18028 17132 18080
rect 17184 18068 17190 18080
rect 18524 18077 18552 18176
rect 19242 18164 19248 18176
rect 19300 18164 19306 18216
rect 19628 18204 19656 18232
rect 19628 18176 20116 18204
rect 20088 18145 20116 18176
rect 20898 18164 20904 18216
rect 20956 18204 20962 18216
rect 21637 18207 21695 18213
rect 21637 18204 21649 18207
rect 20956 18176 21649 18204
rect 20956 18164 20962 18176
rect 21637 18173 21649 18176
rect 21683 18173 21695 18207
rect 21637 18167 21695 18173
rect 19981 18139 20039 18145
rect 19981 18136 19993 18139
rect 19076 18108 19993 18136
rect 19076 18080 19104 18108
rect 19981 18105 19993 18108
rect 20027 18105 20039 18139
rect 19981 18099 20039 18105
rect 20073 18139 20131 18145
rect 20073 18105 20085 18139
rect 20119 18105 20131 18139
rect 20714 18136 20720 18148
rect 20675 18108 20720 18136
rect 20073 18099 20131 18105
rect 20714 18096 20720 18108
rect 20772 18136 20778 18148
rect 22940 18145 22968 18244
rect 23658 18232 23664 18284
rect 23716 18272 23722 18284
rect 24228 18281 24256 18312
rect 24670 18300 24676 18312
rect 24728 18300 24734 18352
rect 24121 18275 24179 18281
rect 24121 18272 24133 18275
rect 23716 18244 24133 18272
rect 23716 18232 23722 18244
rect 24121 18241 24133 18244
rect 24167 18241 24179 18275
rect 24121 18235 24179 18241
rect 24213 18275 24271 18281
rect 24213 18241 24225 18275
rect 24259 18241 24271 18275
rect 25498 18272 25504 18284
rect 25459 18244 25504 18272
rect 24213 18235 24271 18241
rect 25498 18232 25504 18244
rect 25556 18232 25562 18284
rect 26326 18272 26332 18284
rect 26287 18244 26332 18272
rect 26326 18232 26332 18244
rect 26384 18232 26390 18284
rect 23842 18164 23848 18216
rect 23900 18204 23906 18216
rect 24029 18207 24087 18213
rect 24029 18204 24041 18207
rect 23900 18176 24041 18204
rect 23900 18164 23906 18176
rect 24029 18173 24041 18176
rect 24075 18173 24087 18207
rect 25222 18204 25228 18216
rect 25183 18176 25228 18204
rect 24029 18167 24087 18173
rect 25222 18164 25228 18176
rect 25280 18204 25286 18216
rect 25961 18207 26019 18213
rect 25961 18204 25973 18207
rect 25280 18176 25973 18204
rect 25280 18164 25286 18176
rect 25961 18173 25973 18176
rect 26007 18173 26019 18207
rect 25961 18167 26019 18173
rect 21545 18139 21603 18145
rect 21545 18136 21557 18139
rect 20772 18108 21557 18136
rect 20772 18096 20778 18108
rect 21545 18105 21557 18108
rect 21591 18105 21603 18139
rect 21545 18099 21603 18105
rect 22925 18139 22983 18145
rect 22925 18105 22937 18139
rect 22971 18136 22983 18139
rect 23750 18136 23756 18148
rect 22971 18108 23756 18136
rect 22971 18105 22983 18108
rect 22925 18099 22983 18105
rect 23750 18096 23756 18108
rect 23808 18096 23814 18148
rect 17405 18071 17463 18077
rect 17405 18068 17417 18071
rect 17184 18040 17417 18068
rect 17184 18028 17190 18040
rect 17405 18037 17417 18040
rect 17451 18068 17463 18071
rect 18509 18071 18567 18077
rect 18509 18068 18521 18071
rect 17451 18040 18521 18068
rect 17451 18037 17463 18040
rect 17405 18031 17463 18037
rect 18509 18037 18521 18040
rect 18555 18037 18567 18071
rect 19058 18068 19064 18080
rect 19019 18040 19064 18068
rect 18509 18031 18567 18037
rect 19058 18028 19064 18040
rect 19116 18028 19122 18080
rect 19242 18068 19248 18080
rect 19203 18040 19248 18068
rect 19242 18028 19248 18040
rect 19300 18028 19306 18080
rect 20898 18028 20904 18080
rect 20956 18068 20962 18080
rect 20993 18071 21051 18077
rect 20993 18068 21005 18071
rect 20956 18040 21005 18068
rect 20956 18028 20962 18040
rect 20993 18037 21005 18040
rect 21039 18037 21051 18071
rect 20993 18031 21051 18037
rect 21177 18071 21235 18077
rect 21177 18037 21189 18071
rect 21223 18068 21235 18071
rect 21358 18068 21364 18080
rect 21223 18040 21364 18068
rect 21223 18037 21235 18040
rect 21177 18031 21235 18037
rect 21358 18028 21364 18040
rect 21416 18028 21422 18080
rect 22557 18071 22615 18077
rect 22557 18037 22569 18071
rect 22603 18068 22615 18071
rect 23106 18068 23112 18080
rect 22603 18040 23112 18068
rect 22603 18037 22615 18040
rect 22557 18031 22615 18037
rect 23106 18028 23112 18040
rect 23164 18068 23170 18080
rect 23385 18071 23443 18077
rect 23385 18068 23397 18071
rect 23164 18040 23397 18068
rect 23164 18028 23170 18040
rect 23385 18037 23397 18040
rect 23431 18037 23443 18071
rect 23385 18031 23443 18037
rect 25133 18071 25191 18077
rect 25133 18037 25145 18071
rect 25179 18068 25191 18071
rect 25222 18068 25228 18080
rect 25179 18040 25228 18068
rect 25179 18037 25191 18040
rect 25133 18031 25191 18037
rect 25222 18028 25228 18040
rect 25280 18028 25286 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 2406 17864 2412 17876
rect 2367 17836 2412 17864
rect 2406 17824 2412 17836
rect 2464 17824 2470 17876
rect 4338 17864 4344 17876
rect 4299 17836 4344 17864
rect 4338 17824 4344 17836
rect 4396 17824 4402 17876
rect 4525 17867 4583 17873
rect 4525 17833 4537 17867
rect 4571 17864 4583 17867
rect 5258 17864 5264 17876
rect 4571 17836 5264 17864
rect 4571 17833 4583 17836
rect 4525 17827 4583 17833
rect 5258 17824 5264 17836
rect 5316 17824 5322 17876
rect 5994 17824 6000 17876
rect 6052 17864 6058 17876
rect 6914 17864 6920 17876
rect 6052 17836 6920 17864
rect 6052 17824 6058 17836
rect 6914 17824 6920 17836
rect 6972 17824 6978 17876
rect 7190 17824 7196 17876
rect 7248 17864 7254 17876
rect 7745 17867 7803 17873
rect 7745 17864 7757 17867
rect 7248 17836 7757 17864
rect 7248 17824 7254 17836
rect 7745 17833 7757 17836
rect 7791 17833 7803 17867
rect 8478 17864 8484 17876
rect 8439 17836 8484 17864
rect 7745 17827 7803 17833
rect 8478 17824 8484 17836
rect 8536 17824 8542 17876
rect 8846 17864 8852 17876
rect 8807 17836 8852 17864
rect 8846 17824 8852 17836
rect 8904 17824 8910 17876
rect 10689 17867 10747 17873
rect 10689 17833 10701 17867
rect 10735 17864 10747 17867
rect 13078 17864 13084 17876
rect 10735 17836 13084 17864
rect 10735 17833 10747 17836
rect 10689 17827 10747 17833
rect 13078 17824 13084 17836
rect 13136 17824 13142 17876
rect 13446 17824 13452 17876
rect 13504 17864 13510 17876
rect 13633 17867 13691 17873
rect 13633 17864 13645 17867
rect 13504 17836 13645 17864
rect 13504 17824 13510 17836
rect 13633 17833 13645 17836
rect 13679 17833 13691 17867
rect 14182 17864 14188 17876
rect 14143 17836 14188 17864
rect 13633 17827 13691 17833
rect 14182 17824 14188 17836
rect 14240 17824 14246 17876
rect 15102 17864 15108 17876
rect 15063 17836 15108 17864
rect 15102 17824 15108 17836
rect 15160 17824 15166 17876
rect 15286 17864 15292 17876
rect 15247 17836 15292 17864
rect 15286 17824 15292 17836
rect 15344 17824 15350 17876
rect 15749 17867 15807 17873
rect 15749 17833 15761 17867
rect 15795 17864 15807 17867
rect 15930 17864 15936 17876
rect 15795 17836 15936 17864
rect 15795 17833 15807 17836
rect 15749 17827 15807 17833
rect 15930 17824 15936 17836
rect 15988 17824 15994 17876
rect 16390 17864 16396 17876
rect 16351 17836 16396 17864
rect 16390 17824 16396 17836
rect 16448 17824 16454 17876
rect 16850 17864 16856 17876
rect 16811 17836 16856 17864
rect 16850 17824 16856 17836
rect 16908 17824 16914 17876
rect 17402 17824 17408 17876
rect 17460 17824 17466 17876
rect 17954 17824 17960 17876
rect 18012 17864 18018 17876
rect 19061 17867 19119 17873
rect 19061 17864 19073 17867
rect 18012 17836 19073 17864
rect 18012 17824 18018 17836
rect 19061 17833 19073 17836
rect 19107 17864 19119 17867
rect 19518 17864 19524 17876
rect 19107 17836 19524 17864
rect 19107 17833 19119 17836
rect 19061 17827 19119 17833
rect 19518 17824 19524 17836
rect 19576 17824 19582 17876
rect 19978 17864 19984 17876
rect 19628 17836 19984 17864
rect 1946 17756 1952 17808
rect 2004 17796 2010 17808
rect 2590 17796 2596 17808
rect 2004 17768 2596 17796
rect 2004 17756 2010 17768
rect 2590 17756 2596 17768
rect 2648 17796 2654 17808
rect 2777 17799 2835 17805
rect 2777 17796 2789 17799
rect 2648 17768 2789 17796
rect 2648 17756 2654 17768
rect 2777 17765 2789 17768
rect 2823 17765 2835 17799
rect 2777 17759 2835 17765
rect 4356 17728 4384 17824
rect 4893 17799 4951 17805
rect 4893 17765 4905 17799
rect 4939 17796 4951 17799
rect 6638 17796 6644 17808
rect 4939 17768 6644 17796
rect 4939 17765 4951 17768
rect 4893 17759 4951 17765
rect 6638 17756 6644 17768
rect 6696 17756 6702 17808
rect 9674 17796 9680 17808
rect 9635 17768 9680 17796
rect 9674 17756 9680 17768
rect 9732 17756 9738 17808
rect 10597 17799 10655 17805
rect 10597 17765 10609 17799
rect 10643 17796 10655 17799
rect 10962 17796 10968 17808
rect 10643 17768 10968 17796
rect 10643 17765 10655 17768
rect 10597 17759 10655 17765
rect 10962 17756 10968 17768
rect 11020 17756 11026 17808
rect 11149 17799 11207 17805
rect 11149 17765 11161 17799
rect 11195 17796 11207 17799
rect 11330 17796 11336 17808
rect 11195 17768 11336 17796
rect 11195 17765 11207 17768
rect 11149 17759 11207 17765
rect 6178 17728 6184 17740
rect 3068 17700 6184 17728
rect 2866 17660 2872 17672
rect 2827 17632 2872 17660
rect 2866 17620 2872 17632
rect 2924 17620 2930 17672
rect 3068 17669 3096 17700
rect 6178 17688 6184 17700
rect 6236 17728 6242 17740
rect 6345 17731 6403 17737
rect 6345 17728 6357 17731
rect 6236 17700 6357 17728
rect 6236 17688 6242 17700
rect 6345 17697 6357 17700
rect 6391 17697 6403 17731
rect 6345 17691 6403 17697
rect 7558 17688 7564 17740
rect 7616 17728 7622 17740
rect 8297 17731 8355 17737
rect 8297 17728 8309 17731
rect 7616 17700 8309 17728
rect 7616 17688 7622 17700
rect 8297 17697 8309 17700
rect 8343 17697 8355 17731
rect 8297 17691 8355 17697
rect 8386 17688 8392 17740
rect 8444 17728 8450 17740
rect 9217 17731 9275 17737
rect 9217 17728 9229 17731
rect 8444 17700 9229 17728
rect 8444 17688 8450 17700
rect 9217 17697 9229 17700
rect 9263 17697 9275 17731
rect 11054 17728 11060 17740
rect 11015 17700 11060 17728
rect 9217 17691 9275 17697
rect 11054 17688 11060 17700
rect 11112 17688 11118 17740
rect 3053 17663 3111 17669
rect 3053 17629 3065 17663
rect 3099 17629 3111 17663
rect 3053 17623 3111 17629
rect 3878 17620 3884 17672
rect 3936 17660 3942 17672
rect 4982 17660 4988 17672
rect 3936 17632 4988 17660
rect 3936 17620 3942 17632
rect 4982 17620 4988 17632
rect 5040 17620 5046 17672
rect 5074 17620 5080 17672
rect 5132 17660 5138 17672
rect 5132 17632 5177 17660
rect 5132 17620 5138 17632
rect 5534 17620 5540 17672
rect 5592 17660 5598 17672
rect 5905 17663 5963 17669
rect 5905 17660 5917 17663
rect 5592 17632 5917 17660
rect 5592 17620 5598 17632
rect 5905 17629 5917 17632
rect 5951 17629 5963 17663
rect 5905 17623 5963 17629
rect 5994 17620 6000 17672
rect 6052 17660 6058 17672
rect 6089 17663 6147 17669
rect 6089 17660 6101 17663
rect 6052 17632 6101 17660
rect 6052 17620 6058 17632
rect 6089 17629 6101 17632
rect 6135 17629 6147 17663
rect 6089 17623 6147 17629
rect 10962 17620 10968 17672
rect 11020 17660 11026 17672
rect 11164 17660 11192 17759
rect 11330 17756 11336 17768
rect 11388 17756 11394 17808
rect 11793 17799 11851 17805
rect 11793 17765 11805 17799
rect 11839 17796 11851 17799
rect 11882 17796 11888 17808
rect 11839 17768 11888 17796
rect 11839 17765 11851 17768
rect 11793 17759 11851 17765
rect 11882 17756 11888 17768
rect 11940 17756 11946 17808
rect 12529 17799 12587 17805
rect 12529 17765 12541 17799
rect 12575 17796 12587 17799
rect 12802 17796 12808 17808
rect 12575 17768 12808 17796
rect 12575 17765 12587 17768
rect 12529 17759 12587 17765
rect 12802 17756 12808 17768
rect 12860 17756 12866 17808
rect 14550 17756 14556 17808
rect 14608 17796 14614 17808
rect 17420 17796 17448 17824
rect 18506 17796 18512 17808
rect 14608 17768 15884 17796
rect 14608 17756 14614 17768
rect 12894 17688 12900 17740
rect 12952 17728 12958 17740
rect 12989 17731 13047 17737
rect 12989 17728 13001 17731
rect 12952 17700 13001 17728
rect 12952 17688 12958 17700
rect 12989 17697 13001 17700
rect 13035 17697 13047 17731
rect 12989 17691 13047 17697
rect 14642 17688 14648 17740
rect 14700 17728 14706 17740
rect 15657 17731 15715 17737
rect 15657 17728 15669 17731
rect 14700 17700 15669 17728
rect 14700 17688 14706 17700
rect 15657 17697 15669 17700
rect 15703 17697 15715 17731
rect 15657 17691 15715 17697
rect 11330 17660 11336 17672
rect 11020 17632 11192 17660
rect 11291 17632 11336 17660
rect 11020 17620 11026 17632
rect 11330 17620 11336 17632
rect 11388 17620 11394 17672
rect 13078 17660 13084 17672
rect 13039 17632 13084 17660
rect 13078 17620 13084 17632
rect 13136 17620 13142 17672
rect 13173 17663 13231 17669
rect 13173 17629 13185 17663
rect 13219 17629 13231 17663
rect 13173 17623 13231 17629
rect 12161 17595 12219 17601
rect 12161 17561 12173 17595
rect 12207 17592 12219 17595
rect 13188 17592 13216 17623
rect 14366 17620 14372 17672
rect 14424 17660 14430 17672
rect 14734 17660 14740 17672
rect 14424 17632 14740 17660
rect 14424 17620 14430 17632
rect 14734 17620 14740 17632
rect 14792 17620 14798 17672
rect 13446 17592 13452 17604
rect 12207 17564 13452 17592
rect 12207 17561 12219 17564
rect 12161 17555 12219 17561
rect 13446 17552 13452 17564
rect 13504 17552 13510 17604
rect 14918 17552 14924 17604
rect 14976 17552 14982 17604
rect 15672 17592 15700 17691
rect 15856 17669 15884 17768
rect 17144 17768 18512 17796
rect 17144 17737 17172 17768
rect 18506 17756 18512 17768
rect 18564 17756 18570 17808
rect 19628 17805 19656 17836
rect 19978 17824 19984 17836
rect 20036 17824 20042 17876
rect 20165 17867 20223 17873
rect 20165 17833 20177 17867
rect 20211 17864 20223 17867
rect 20346 17864 20352 17876
rect 20211 17836 20352 17864
rect 20211 17833 20223 17836
rect 20165 17827 20223 17833
rect 19613 17799 19671 17805
rect 19613 17765 19625 17799
rect 19659 17765 19671 17799
rect 19613 17759 19671 17765
rect 20070 17756 20076 17808
rect 20128 17796 20134 17808
rect 20180 17796 20208 17827
rect 20346 17824 20352 17836
rect 20404 17824 20410 17876
rect 20717 17867 20775 17873
rect 20717 17833 20729 17867
rect 20763 17864 20775 17867
rect 22002 17864 22008 17876
rect 20763 17836 22008 17864
rect 20763 17833 20775 17836
rect 20717 17827 20775 17833
rect 22002 17824 22008 17836
rect 22060 17824 22066 17876
rect 22186 17824 22192 17876
rect 22244 17864 22250 17876
rect 22465 17867 22523 17873
rect 22465 17864 22477 17867
rect 22244 17836 22477 17864
rect 22244 17824 22250 17836
rect 22465 17833 22477 17836
rect 22511 17833 22523 17867
rect 23290 17864 23296 17876
rect 23251 17836 23296 17864
rect 22465 17827 22523 17833
rect 23290 17824 23296 17836
rect 23348 17824 23354 17876
rect 23842 17824 23848 17876
rect 23900 17864 23906 17876
rect 24213 17867 24271 17873
rect 24213 17864 24225 17867
rect 23900 17836 24225 17864
rect 23900 17824 23906 17836
rect 24213 17833 24225 17836
rect 24259 17833 24271 17867
rect 24213 17827 24271 17833
rect 24302 17824 24308 17876
rect 24360 17864 24366 17876
rect 24360 17836 24992 17864
rect 24360 17824 24366 17836
rect 20128 17768 20208 17796
rect 21177 17799 21235 17805
rect 20128 17756 20134 17768
rect 21177 17765 21189 17799
rect 21223 17796 21235 17799
rect 21542 17796 21548 17808
rect 21223 17768 21548 17796
rect 21223 17765 21235 17768
rect 21177 17759 21235 17765
rect 21542 17756 21548 17768
rect 21600 17756 21606 17808
rect 21818 17756 21824 17808
rect 21876 17796 21882 17808
rect 24026 17796 24032 17808
rect 21876 17768 24032 17796
rect 21876 17756 21882 17768
rect 24026 17756 24032 17768
rect 24084 17796 24090 17808
rect 24857 17799 24915 17805
rect 24857 17796 24869 17799
rect 24084 17768 24869 17796
rect 24084 17756 24090 17768
rect 24857 17765 24869 17768
rect 24903 17765 24915 17799
rect 24857 17759 24915 17765
rect 17402 17737 17408 17740
rect 17129 17731 17187 17737
rect 17129 17697 17141 17731
rect 17175 17697 17187 17731
rect 17396 17728 17408 17737
rect 17363 17700 17408 17728
rect 17129 17691 17187 17697
rect 17396 17691 17408 17700
rect 17402 17688 17408 17691
rect 17460 17688 17466 17740
rect 19337 17731 19395 17737
rect 19337 17697 19349 17731
rect 19383 17728 19395 17731
rect 19978 17728 19984 17740
rect 19383 17700 19984 17728
rect 19383 17697 19395 17700
rect 19337 17691 19395 17697
rect 19978 17688 19984 17700
rect 20036 17728 20042 17740
rect 20346 17728 20352 17740
rect 20036 17700 20352 17728
rect 20036 17688 20042 17700
rect 20346 17688 20352 17700
rect 20404 17688 20410 17740
rect 21358 17688 21364 17740
rect 21416 17728 21422 17740
rect 21637 17731 21695 17737
rect 21637 17728 21649 17731
rect 21416 17700 21649 17728
rect 21416 17688 21422 17700
rect 21637 17697 21649 17700
rect 21683 17697 21695 17731
rect 21637 17691 21695 17697
rect 22370 17688 22376 17740
rect 22428 17728 22434 17740
rect 23198 17728 23204 17740
rect 22428 17700 23204 17728
rect 22428 17688 22434 17700
rect 23198 17688 23204 17700
rect 23256 17688 23262 17740
rect 24670 17688 24676 17740
rect 24728 17728 24734 17740
rect 24765 17731 24823 17737
rect 24765 17728 24777 17731
rect 24728 17700 24777 17728
rect 24728 17688 24734 17700
rect 24765 17697 24777 17700
rect 24811 17697 24823 17731
rect 24765 17691 24823 17697
rect 15841 17663 15899 17669
rect 15841 17629 15853 17663
rect 15887 17629 15899 17663
rect 15841 17623 15899 17629
rect 20898 17620 20904 17672
rect 20956 17660 20962 17672
rect 21729 17663 21787 17669
rect 21729 17660 21741 17663
rect 20956 17632 21741 17660
rect 20956 17620 20962 17632
rect 21729 17629 21741 17632
rect 21775 17629 21787 17663
rect 21729 17623 21787 17629
rect 21821 17663 21879 17669
rect 21821 17629 21833 17663
rect 21867 17629 21879 17663
rect 23382 17660 23388 17672
rect 23343 17632 23388 17660
rect 21821 17623 21879 17629
rect 16482 17592 16488 17604
rect 15672 17564 16488 17592
rect 16482 17552 16488 17564
rect 16540 17552 16546 17604
rect 21174 17552 21180 17604
rect 21232 17592 21238 17604
rect 21836 17592 21864 17623
rect 23382 17620 23388 17632
rect 23440 17620 23446 17672
rect 23934 17620 23940 17672
rect 23992 17660 23998 17672
rect 24964 17669 24992 17836
rect 25038 17824 25044 17876
rect 25096 17864 25102 17876
rect 25409 17867 25467 17873
rect 25409 17864 25421 17867
rect 25096 17836 25421 17864
rect 25096 17824 25102 17836
rect 25409 17833 25421 17836
rect 25455 17833 25467 17867
rect 25409 17827 25467 17833
rect 24949 17663 25007 17669
rect 23992 17632 24900 17660
rect 23992 17620 23998 17632
rect 21232 17564 21864 17592
rect 21232 17552 21238 17564
rect 22002 17552 22008 17604
rect 22060 17592 22066 17604
rect 22833 17595 22891 17601
rect 22833 17592 22845 17595
rect 22060 17564 22845 17592
rect 22060 17552 22066 17564
rect 22833 17561 22845 17564
rect 22879 17561 22891 17595
rect 22833 17555 22891 17561
rect 23474 17552 23480 17604
rect 23532 17592 23538 17604
rect 24397 17595 24455 17601
rect 24397 17592 24409 17595
rect 23532 17564 24409 17592
rect 23532 17552 23538 17564
rect 24397 17561 24409 17564
rect 24443 17561 24455 17595
rect 24872 17592 24900 17632
rect 24949 17629 24961 17663
rect 24995 17660 25007 17663
rect 25038 17660 25044 17672
rect 24995 17632 25044 17660
rect 24995 17629 25007 17632
rect 24949 17623 25007 17629
rect 25038 17620 25044 17632
rect 25096 17620 25102 17672
rect 25777 17595 25835 17601
rect 25777 17592 25789 17595
rect 24872 17564 25789 17592
rect 24397 17555 24455 17561
rect 25777 17561 25789 17564
rect 25823 17561 25835 17595
rect 25777 17555 25835 17561
rect 1670 17524 1676 17536
rect 1631 17496 1676 17524
rect 1670 17484 1676 17496
rect 1728 17484 1734 17536
rect 2133 17527 2191 17533
rect 2133 17493 2145 17527
rect 2179 17524 2191 17527
rect 2682 17524 2688 17536
rect 2179 17496 2688 17524
rect 2179 17493 2191 17496
rect 2133 17487 2191 17493
rect 2682 17484 2688 17496
rect 2740 17484 2746 17536
rect 3050 17484 3056 17536
rect 3108 17524 3114 17536
rect 3605 17527 3663 17533
rect 3605 17524 3617 17527
rect 3108 17496 3617 17524
rect 3108 17484 3114 17496
rect 3605 17493 3617 17496
rect 3651 17524 3663 17527
rect 4062 17524 4068 17536
rect 3651 17496 4068 17524
rect 3651 17493 3663 17496
rect 3605 17487 3663 17493
rect 4062 17484 4068 17496
rect 4120 17484 4126 17536
rect 5629 17527 5687 17533
rect 5629 17493 5641 17527
rect 5675 17524 5687 17527
rect 5994 17524 6000 17536
rect 5675 17496 6000 17524
rect 5675 17493 5687 17496
rect 5629 17487 5687 17493
rect 5994 17484 6000 17496
rect 6052 17484 6058 17536
rect 6362 17484 6368 17536
rect 6420 17524 6426 17536
rect 7469 17527 7527 17533
rect 7469 17524 7481 17527
rect 6420 17496 7481 17524
rect 6420 17484 6426 17496
rect 7469 17493 7481 17496
rect 7515 17493 7527 17527
rect 8110 17524 8116 17536
rect 8071 17496 8116 17524
rect 7469 17487 7527 17493
rect 8110 17484 8116 17496
rect 8168 17484 8174 17536
rect 9766 17484 9772 17536
rect 9824 17524 9830 17536
rect 10137 17527 10195 17533
rect 10137 17524 10149 17527
rect 9824 17496 10149 17524
rect 9824 17484 9830 17496
rect 10137 17493 10149 17496
rect 10183 17493 10195 17527
rect 10137 17487 10195 17493
rect 12621 17527 12679 17533
rect 12621 17493 12633 17527
rect 12667 17524 12679 17527
rect 13814 17524 13820 17536
rect 12667 17496 13820 17524
rect 12667 17493 12679 17496
rect 12621 17487 12679 17493
rect 13814 17484 13820 17496
rect 13872 17484 13878 17536
rect 13906 17484 13912 17536
rect 13964 17524 13970 17536
rect 14001 17527 14059 17533
rect 14001 17524 14013 17527
rect 13964 17496 14013 17524
rect 13964 17484 13970 17496
rect 14001 17493 14013 17496
rect 14047 17493 14059 17527
rect 14734 17524 14740 17536
rect 14695 17496 14740 17524
rect 14001 17487 14059 17493
rect 14734 17484 14740 17496
rect 14792 17484 14798 17536
rect 14936 17524 14964 17552
rect 16758 17524 16764 17536
rect 14936 17496 16764 17524
rect 16758 17484 16764 17496
rect 16816 17484 16822 17536
rect 18509 17527 18567 17533
rect 18509 17493 18521 17527
rect 18555 17524 18567 17527
rect 18874 17524 18880 17536
rect 18555 17496 18880 17524
rect 18555 17493 18567 17496
rect 18509 17487 18567 17493
rect 18874 17484 18880 17496
rect 18932 17484 18938 17536
rect 21269 17527 21327 17533
rect 21269 17493 21281 17527
rect 21315 17524 21327 17527
rect 21634 17524 21640 17536
rect 21315 17496 21640 17524
rect 21315 17493 21327 17496
rect 21269 17487 21327 17493
rect 21634 17484 21640 17496
rect 21692 17484 21698 17536
rect 23937 17527 23995 17533
rect 23937 17493 23949 17527
rect 23983 17524 23995 17527
rect 24210 17524 24216 17536
rect 23983 17496 24216 17524
rect 23983 17493 23995 17496
rect 23937 17487 23995 17493
rect 24210 17484 24216 17496
rect 24268 17484 24274 17536
rect 24412 17524 24440 17555
rect 25222 17524 25228 17536
rect 24412 17496 25228 17524
rect 25222 17484 25228 17496
rect 25280 17484 25286 17536
rect 26234 17524 26240 17536
rect 26195 17496 26240 17524
rect 26234 17484 26240 17496
rect 26292 17484 26298 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1578 17320 1584 17332
rect 1539 17292 1584 17320
rect 1578 17280 1584 17292
rect 1636 17280 1642 17332
rect 2590 17320 2596 17332
rect 2551 17292 2596 17320
rect 2590 17280 2596 17292
rect 2648 17280 2654 17332
rect 5813 17323 5871 17329
rect 5813 17289 5825 17323
rect 5859 17320 5871 17323
rect 6362 17320 6368 17332
rect 5859 17292 6368 17320
rect 5859 17289 5871 17292
rect 5813 17283 5871 17289
rect 6362 17280 6368 17292
rect 6420 17280 6426 17332
rect 6730 17280 6736 17332
rect 6788 17320 6794 17332
rect 7009 17323 7067 17329
rect 7009 17320 7021 17323
rect 6788 17292 7021 17320
rect 6788 17280 6794 17292
rect 7009 17289 7021 17292
rect 7055 17289 7067 17323
rect 7009 17283 7067 17289
rect 7466 17280 7472 17332
rect 7524 17320 7530 17332
rect 8113 17323 8171 17329
rect 8113 17320 8125 17323
rect 7524 17292 8125 17320
rect 7524 17280 7530 17292
rect 8113 17289 8125 17292
rect 8159 17289 8171 17323
rect 8113 17283 8171 17289
rect 8294 17280 8300 17332
rect 8352 17320 8358 17332
rect 9493 17323 9551 17329
rect 9493 17320 9505 17323
rect 8352 17292 9505 17320
rect 8352 17280 8358 17292
rect 9493 17289 9505 17292
rect 9539 17289 9551 17323
rect 9493 17283 9551 17289
rect 2501 17255 2559 17261
rect 2501 17221 2513 17255
rect 2547 17252 2559 17255
rect 4249 17255 4307 17261
rect 2547 17224 3832 17252
rect 2547 17221 2559 17224
rect 2501 17215 2559 17221
rect 2222 17184 2228 17196
rect 2183 17156 2228 17184
rect 2222 17144 2228 17156
rect 2280 17144 2286 17196
rect 3418 17144 3424 17196
rect 3476 17184 3482 17196
rect 3697 17187 3755 17193
rect 3697 17184 3709 17187
rect 3476 17156 3709 17184
rect 3476 17144 3482 17156
rect 3697 17153 3709 17156
rect 3743 17153 3755 17187
rect 3804 17184 3832 17224
rect 4249 17221 4261 17255
rect 4295 17252 4307 17255
rect 5074 17252 5080 17264
rect 4295 17224 5080 17252
rect 4295 17221 4307 17224
rect 4249 17215 4307 17221
rect 5074 17212 5080 17224
rect 5132 17212 5138 17264
rect 6178 17252 6184 17264
rect 6139 17224 6184 17252
rect 6178 17212 6184 17224
rect 6236 17212 6242 17264
rect 8938 17252 8944 17264
rect 6288 17224 8944 17252
rect 4617 17187 4675 17193
rect 4617 17184 4629 17187
rect 3804 17156 4629 17184
rect 3697 17147 3755 17153
rect 4617 17153 4629 17156
rect 4663 17184 4675 17187
rect 5166 17184 5172 17196
rect 4663 17156 5172 17184
rect 4663 17153 4675 17156
rect 4617 17147 4675 17153
rect 5166 17144 5172 17156
rect 5224 17144 5230 17196
rect 5258 17144 5264 17196
rect 5316 17184 5322 17196
rect 5316 17156 5361 17184
rect 5316 17144 5322 17156
rect 6086 17144 6092 17196
rect 6144 17184 6150 17196
rect 6288 17184 6316 17224
rect 8938 17212 8944 17224
rect 8996 17212 9002 17264
rect 6144 17156 6316 17184
rect 8021 17187 8079 17193
rect 6144 17144 6150 17156
rect 8021 17153 8033 17187
rect 8067 17184 8079 17187
rect 8754 17184 8760 17196
rect 8067 17156 8760 17184
rect 8067 17153 8079 17156
rect 8021 17147 8079 17153
rect 8754 17144 8760 17156
rect 8812 17144 8818 17196
rect 9306 17144 9312 17196
rect 9364 17144 9370 17196
rect 9508 17184 9536 17283
rect 10042 17280 10048 17332
rect 10100 17320 10106 17332
rect 10778 17320 10784 17332
rect 10100 17292 10784 17320
rect 10100 17280 10106 17292
rect 10778 17280 10784 17292
rect 10836 17280 10842 17332
rect 11057 17323 11115 17329
rect 11057 17289 11069 17323
rect 11103 17320 11115 17323
rect 11238 17320 11244 17332
rect 11103 17292 11244 17320
rect 11103 17289 11115 17292
rect 11057 17283 11115 17289
rect 11238 17280 11244 17292
rect 11296 17280 11302 17332
rect 13998 17280 14004 17332
rect 14056 17320 14062 17332
rect 14458 17320 14464 17332
rect 14056 17292 14464 17320
rect 14056 17280 14062 17292
rect 14458 17280 14464 17292
rect 14516 17280 14522 17332
rect 14826 17320 14832 17332
rect 14787 17292 14832 17320
rect 14826 17280 14832 17292
rect 14884 17280 14890 17332
rect 18046 17320 18052 17332
rect 18007 17292 18052 17320
rect 18046 17280 18052 17292
rect 18104 17280 18110 17332
rect 19153 17323 19211 17329
rect 19153 17289 19165 17323
rect 19199 17320 19211 17323
rect 19242 17320 19248 17332
rect 19199 17292 19248 17320
rect 19199 17289 19211 17292
rect 19153 17283 19211 17289
rect 19242 17280 19248 17292
rect 19300 17280 19306 17332
rect 19426 17280 19432 17332
rect 19484 17320 19490 17332
rect 19613 17323 19671 17329
rect 19613 17320 19625 17323
rect 19484 17292 19625 17320
rect 19484 17280 19490 17292
rect 19613 17289 19625 17292
rect 19659 17289 19671 17323
rect 19613 17283 19671 17289
rect 22370 17280 22376 17332
rect 22428 17320 22434 17332
rect 22646 17320 22652 17332
rect 22428 17292 22652 17320
rect 22428 17280 22434 17292
rect 22646 17280 22652 17292
rect 22704 17280 22710 17332
rect 23750 17280 23756 17332
rect 23808 17320 23814 17332
rect 24670 17320 24676 17332
rect 23808 17292 24676 17320
rect 23808 17280 23814 17292
rect 24670 17280 24676 17292
rect 24728 17320 24734 17332
rect 25041 17323 25099 17329
rect 25041 17320 25053 17323
rect 24728 17292 25053 17320
rect 24728 17280 24734 17292
rect 25041 17289 25053 17292
rect 25087 17289 25099 17323
rect 26326 17320 26332 17332
rect 26287 17292 26332 17320
rect 25041 17283 25099 17289
rect 26326 17280 26332 17292
rect 26384 17280 26390 17332
rect 10962 17212 10968 17264
rect 11020 17252 11026 17264
rect 11333 17255 11391 17261
rect 11333 17252 11345 17255
rect 11020 17224 11345 17252
rect 11020 17212 11026 17224
rect 11333 17221 11345 17224
rect 11379 17221 11391 17255
rect 11333 17215 11391 17221
rect 12250 17212 12256 17264
rect 12308 17252 12314 17264
rect 14642 17252 14648 17264
rect 12308 17224 12388 17252
rect 12308 17212 12314 17224
rect 9508 17156 9812 17184
rect 2866 17076 2872 17128
rect 2924 17116 2930 17128
rect 3053 17119 3111 17125
rect 3053 17116 3065 17119
rect 2924 17088 3065 17116
rect 2924 17076 2930 17088
rect 3053 17085 3065 17088
rect 3099 17116 3111 17119
rect 3602 17116 3608 17128
rect 3099 17088 3608 17116
rect 3099 17085 3111 17088
rect 3053 17079 3111 17085
rect 3602 17076 3608 17088
rect 3660 17076 3666 17128
rect 5074 17116 5080 17128
rect 5035 17088 5080 17116
rect 5074 17076 5080 17088
rect 5132 17076 5138 17128
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17116 6883 17119
rect 7098 17116 7104 17128
rect 6871 17088 7104 17116
rect 6871 17085 6883 17088
rect 6825 17079 6883 17085
rect 7098 17076 7104 17088
rect 7156 17116 7162 17128
rect 7377 17119 7435 17125
rect 7377 17116 7389 17119
rect 7156 17088 7389 17116
rect 7156 17076 7162 17088
rect 7377 17085 7389 17088
rect 7423 17085 7435 17119
rect 7377 17079 7435 17085
rect 8481 17119 8539 17125
rect 8481 17085 8493 17119
rect 8527 17116 8539 17119
rect 8570 17116 8576 17128
rect 8527 17088 8576 17116
rect 8527 17085 8539 17088
rect 8481 17079 8539 17085
rect 8570 17076 8576 17088
rect 8628 17076 8634 17128
rect 9324 17116 9352 17144
rect 9582 17116 9588 17128
rect 9324 17088 9588 17116
rect 9582 17076 9588 17088
rect 9640 17116 9646 17128
rect 9677 17119 9735 17125
rect 9677 17116 9689 17119
rect 9640 17088 9689 17116
rect 9640 17076 9646 17088
rect 9677 17085 9689 17088
rect 9723 17085 9735 17119
rect 9784 17116 9812 17156
rect 11054 17144 11060 17196
rect 11112 17184 11118 17196
rect 11701 17187 11759 17193
rect 11701 17184 11713 17187
rect 11112 17156 11713 17184
rect 11112 17144 11118 17156
rect 11701 17153 11713 17156
rect 11747 17153 11759 17187
rect 11701 17147 11759 17153
rect 9933 17119 9991 17125
rect 9933 17116 9945 17119
rect 9784 17088 9945 17116
rect 9677 17079 9735 17085
rect 9933 17085 9945 17088
rect 9979 17116 9991 17119
rect 9979 17088 10088 17116
rect 9979 17085 9991 17088
rect 9933 17079 9991 17085
rect 1670 17008 1676 17060
rect 1728 17048 1734 17060
rect 1949 17051 2007 17057
rect 1949 17048 1961 17051
rect 1728 17020 1961 17048
rect 1728 17008 1734 17020
rect 1949 17017 1961 17020
rect 1995 17048 2007 17051
rect 2501 17051 2559 17057
rect 2501 17048 2513 17051
rect 1995 17020 2513 17048
rect 1995 17017 2007 17020
rect 1949 17011 2007 17017
rect 2501 17017 2513 17020
rect 2547 17017 2559 17051
rect 2501 17011 2559 17017
rect 2682 17008 2688 17060
rect 2740 17048 2746 17060
rect 4982 17048 4988 17060
rect 2740 17020 4988 17048
rect 2740 17008 2746 17020
rect 4982 17008 4988 17020
rect 5040 17008 5046 17060
rect 7558 17008 7564 17060
rect 7616 17048 7622 17060
rect 9125 17051 9183 17057
rect 9125 17048 9137 17051
rect 7616 17020 9137 17048
rect 7616 17008 7622 17020
rect 9125 17017 9137 17020
rect 9171 17048 9183 17051
rect 9306 17048 9312 17060
rect 9171 17020 9312 17048
rect 9171 17017 9183 17020
rect 9125 17011 9183 17017
rect 9306 17008 9312 17020
rect 9364 17008 9370 17060
rect 10060 17048 10088 17088
rect 10134 17048 10140 17060
rect 10060 17020 10140 17048
rect 10134 17008 10140 17020
rect 10192 17008 10198 17060
rect 12253 17051 12311 17057
rect 12253 17017 12265 17051
rect 12299 17048 12311 17051
rect 12360 17048 12388 17224
rect 14476 17224 14648 17252
rect 13541 17187 13599 17193
rect 13541 17153 13553 17187
rect 13587 17184 13599 17187
rect 13587 17156 14044 17184
rect 13587 17153 13599 17156
rect 13541 17147 13599 17153
rect 13170 17116 13176 17128
rect 12636 17088 13176 17116
rect 12636 17048 12664 17088
rect 13170 17076 13176 17088
rect 13228 17116 13234 17128
rect 13357 17119 13415 17125
rect 13357 17116 13369 17119
rect 13228 17088 13369 17116
rect 13228 17076 13234 17088
rect 13357 17085 13369 17088
rect 13403 17085 13415 17119
rect 13357 17079 13415 17085
rect 12299 17020 12664 17048
rect 12299 17017 12311 17020
rect 12253 17011 12311 17017
rect 12710 17008 12716 17060
rect 12768 17048 12774 17060
rect 12805 17051 12863 17057
rect 12805 17048 12817 17051
rect 12768 17020 12817 17048
rect 12768 17008 12774 17020
rect 12805 17017 12817 17020
rect 12851 17048 12863 17051
rect 12851 17020 13308 17048
rect 12851 17017 12863 17020
rect 12805 17011 12863 17017
rect 2041 16983 2099 16989
rect 2041 16949 2053 16983
rect 2087 16980 2099 16983
rect 2406 16980 2412 16992
rect 2087 16952 2412 16980
rect 2087 16949 2099 16952
rect 2041 16943 2099 16949
rect 2406 16940 2412 16952
rect 2464 16940 2470 16992
rect 3142 16980 3148 16992
rect 3103 16952 3148 16980
rect 3142 16940 3148 16952
rect 3200 16940 3206 16992
rect 3510 16980 3516 16992
rect 3471 16952 3516 16980
rect 3510 16940 3516 16952
rect 3568 16940 3574 16992
rect 3605 16983 3663 16989
rect 3605 16949 3617 16983
rect 3651 16980 3663 16983
rect 3970 16980 3976 16992
rect 3651 16952 3976 16980
rect 3651 16949 3663 16952
rect 3605 16943 3663 16949
rect 3970 16940 3976 16952
rect 4028 16940 4034 16992
rect 4706 16980 4712 16992
rect 4667 16952 4712 16980
rect 4706 16940 4712 16952
rect 4764 16940 4770 16992
rect 6454 16940 6460 16992
rect 6512 16980 6518 16992
rect 6549 16983 6607 16989
rect 6549 16980 6561 16983
rect 6512 16952 6561 16980
rect 6512 16940 6518 16952
rect 6549 16949 6561 16952
rect 6595 16949 6607 16983
rect 6549 16943 6607 16949
rect 8110 16940 8116 16992
rect 8168 16980 8174 16992
rect 8573 16983 8631 16989
rect 8573 16980 8585 16983
rect 8168 16952 8585 16980
rect 8168 16940 8174 16952
rect 8573 16949 8585 16952
rect 8619 16949 8631 16983
rect 12894 16980 12900 16992
rect 12855 16952 12900 16980
rect 8573 16943 8631 16949
rect 12894 16940 12900 16952
rect 12952 16940 12958 16992
rect 13280 16989 13308 17020
rect 13265 16983 13323 16989
rect 13265 16949 13277 16983
rect 13311 16980 13323 16983
rect 13630 16980 13636 16992
rect 13311 16952 13636 16980
rect 13311 16949 13323 16952
rect 13265 16943 13323 16949
rect 13630 16940 13636 16952
rect 13688 16940 13694 16992
rect 14016 16989 14044 17156
rect 14476 17128 14504 17224
rect 14642 17212 14648 17224
rect 14700 17212 14706 17264
rect 17129 17255 17187 17261
rect 17129 17221 17141 17255
rect 17175 17221 17187 17255
rect 17129 17215 17187 17221
rect 17144 17184 17172 17215
rect 24026 17212 24032 17264
rect 24084 17252 24090 17264
rect 24765 17255 24823 17261
rect 24765 17252 24777 17255
rect 24084 17224 24777 17252
rect 24084 17212 24090 17224
rect 24765 17221 24777 17224
rect 24811 17221 24823 17255
rect 24765 17215 24823 17221
rect 25314 17212 25320 17264
rect 25372 17252 25378 17264
rect 25866 17252 25872 17264
rect 25372 17224 25872 17252
rect 25372 17212 25378 17224
rect 25866 17212 25872 17224
rect 25924 17212 25930 17264
rect 17402 17184 17408 17196
rect 17144 17156 17408 17184
rect 17402 17144 17408 17156
rect 17460 17184 17466 17196
rect 17865 17187 17923 17193
rect 17865 17184 17877 17187
rect 17460 17156 17877 17184
rect 17460 17144 17466 17156
rect 17865 17153 17877 17156
rect 17911 17184 17923 17187
rect 18690 17184 18696 17196
rect 17911 17156 18696 17184
rect 17911 17153 17923 17156
rect 17865 17147 17923 17153
rect 18690 17144 18696 17156
rect 18748 17144 18754 17196
rect 19426 17144 19432 17196
rect 19484 17184 19490 17196
rect 19521 17187 19579 17193
rect 19521 17184 19533 17187
rect 19484 17156 19533 17184
rect 19484 17144 19490 17156
rect 19521 17153 19533 17156
rect 19567 17184 19579 17187
rect 20165 17187 20223 17193
rect 20165 17184 20177 17187
rect 19567 17156 20177 17184
rect 19567 17153 19579 17156
rect 19521 17147 19579 17153
rect 20165 17153 20177 17156
rect 20211 17153 20223 17187
rect 20165 17147 20223 17153
rect 21542 17144 21548 17196
rect 21600 17184 21606 17196
rect 22373 17187 22431 17193
rect 22373 17184 22385 17187
rect 21600 17156 22385 17184
rect 21600 17144 21606 17156
rect 22373 17153 22385 17156
rect 22419 17153 22431 17187
rect 22373 17147 22431 17153
rect 23106 17144 23112 17196
rect 23164 17184 23170 17196
rect 23658 17184 23664 17196
rect 23164 17156 23664 17184
rect 23164 17144 23170 17156
rect 23658 17144 23664 17156
rect 23716 17144 23722 17196
rect 24210 17144 24216 17196
rect 24268 17184 24274 17196
rect 24305 17187 24363 17193
rect 24305 17184 24317 17187
rect 24268 17156 24317 17184
rect 24268 17144 24274 17156
rect 24305 17153 24317 17156
rect 24351 17153 24363 17187
rect 25406 17184 25412 17196
rect 25367 17156 25412 17184
rect 24305 17147 24363 17153
rect 14458 17116 14464 17128
rect 14419 17088 14464 17116
rect 14458 17076 14464 17088
rect 14516 17076 14522 17128
rect 14642 17116 14648 17128
rect 14603 17088 14648 17116
rect 14642 17076 14648 17088
rect 14700 17076 14706 17128
rect 15194 17076 15200 17128
rect 15252 17116 15258 17128
rect 15749 17119 15807 17125
rect 15749 17116 15761 17119
rect 15252 17088 15761 17116
rect 15252 17076 15258 17088
rect 15749 17085 15761 17088
rect 15795 17116 15807 17119
rect 18046 17116 18052 17128
rect 15795 17088 18052 17116
rect 15795 17085 15807 17088
rect 15749 17079 15807 17085
rect 18046 17076 18052 17088
rect 18104 17076 18110 17128
rect 18506 17116 18512 17128
rect 18419 17088 18512 17116
rect 18506 17076 18512 17088
rect 18564 17116 18570 17128
rect 19242 17116 19248 17128
rect 18564 17088 19248 17116
rect 18564 17076 18570 17088
rect 19242 17076 19248 17088
rect 19300 17076 19306 17128
rect 21818 17076 21824 17128
rect 21876 17116 21882 17128
rect 23017 17119 23075 17125
rect 23017 17116 23029 17119
rect 21876 17088 23029 17116
rect 21876 17076 21882 17088
rect 23017 17085 23029 17088
rect 23063 17116 23075 17119
rect 24121 17119 24179 17125
rect 24121 17116 24133 17119
rect 23063 17088 24133 17116
rect 23063 17085 23075 17088
rect 23017 17079 23075 17085
rect 24121 17085 24133 17088
rect 24167 17085 24179 17119
rect 24320 17116 24348 17147
rect 25406 17144 25412 17156
rect 25464 17144 25470 17196
rect 24762 17116 24768 17128
rect 24320 17088 24768 17116
rect 24121 17079 24179 17085
rect 24762 17076 24768 17088
rect 24820 17076 24826 17128
rect 24946 17076 24952 17128
rect 25004 17116 25010 17128
rect 25225 17119 25283 17125
rect 25225 17116 25237 17119
rect 25004 17088 25237 17116
rect 25004 17076 25010 17088
rect 25225 17085 25237 17088
rect 25271 17116 25283 17119
rect 25961 17119 26019 17125
rect 25961 17116 25973 17119
rect 25271 17088 25973 17116
rect 25271 17085 25283 17088
rect 25225 17079 25283 17085
rect 25961 17085 25973 17088
rect 26007 17085 26019 17119
rect 25961 17079 26019 17085
rect 16016 17051 16074 17057
rect 16016 17017 16028 17051
rect 16062 17048 16074 17051
rect 16574 17048 16580 17060
rect 16062 17020 16580 17048
rect 16062 17017 16074 17020
rect 16016 17011 16074 17017
rect 16574 17008 16580 17020
rect 16632 17048 16638 17060
rect 17405 17051 17463 17057
rect 17405 17048 17417 17051
rect 16632 17020 17417 17048
rect 16632 17008 16638 17020
rect 17405 17017 17417 17020
rect 17451 17048 17463 17051
rect 17678 17048 17684 17060
rect 17451 17020 17684 17048
rect 17451 17017 17463 17020
rect 17405 17011 17463 17017
rect 17678 17008 17684 17020
rect 17736 17008 17742 17060
rect 18417 17051 18475 17057
rect 18417 17017 18429 17051
rect 18463 17048 18475 17051
rect 18598 17048 18604 17060
rect 18463 17020 18604 17048
rect 18463 17017 18475 17020
rect 18417 17011 18475 17017
rect 18598 17008 18604 17020
rect 18656 17008 18662 17060
rect 19981 17051 20039 17057
rect 19981 17048 19993 17051
rect 19352 17020 19993 17048
rect 19352 16992 19380 17020
rect 19981 17017 19993 17020
rect 20027 17017 20039 17051
rect 19981 17011 20039 17017
rect 20346 17008 20352 17060
rect 20404 17048 20410 17060
rect 23474 17048 23480 17060
rect 20404 17020 23480 17048
rect 20404 17008 20410 17020
rect 14001 16983 14059 16989
rect 14001 16949 14013 16983
rect 14047 16980 14059 16983
rect 14090 16980 14096 16992
rect 14047 16952 14096 16980
rect 14047 16949 14059 16952
rect 14001 16943 14059 16949
rect 14090 16940 14096 16952
rect 14148 16940 14154 16992
rect 15102 16940 15108 16992
rect 15160 16980 15166 16992
rect 15289 16983 15347 16989
rect 15289 16980 15301 16983
rect 15160 16952 15301 16980
rect 15160 16940 15166 16952
rect 15289 16949 15301 16952
rect 15335 16980 15347 16983
rect 15930 16980 15936 16992
rect 15335 16952 15936 16980
rect 15335 16949 15347 16952
rect 15289 16943 15347 16949
rect 15930 16940 15936 16952
rect 15988 16940 15994 16992
rect 19334 16940 19340 16992
rect 19392 16940 19398 16992
rect 20070 16980 20076 16992
rect 20031 16952 20076 16980
rect 20070 16940 20076 16952
rect 20128 16940 20134 16992
rect 20898 16980 20904 16992
rect 20859 16952 20904 16980
rect 20898 16940 20904 16952
rect 20956 16940 20962 16992
rect 21174 16940 21180 16992
rect 21232 16980 21238 16992
rect 21269 16983 21327 16989
rect 21269 16980 21281 16983
rect 21232 16952 21281 16980
rect 21232 16940 21238 16952
rect 21269 16949 21281 16952
rect 21315 16949 21327 16983
rect 21269 16943 21327 16949
rect 21542 16940 21548 16992
rect 21600 16980 21606 16992
rect 21637 16983 21695 16989
rect 21637 16980 21649 16983
rect 21600 16952 21649 16980
rect 21600 16940 21606 16952
rect 21637 16949 21649 16952
rect 21683 16949 21695 16983
rect 21637 16943 21695 16949
rect 21821 16983 21879 16989
rect 21821 16949 21833 16983
rect 21867 16980 21879 16983
rect 22002 16980 22008 16992
rect 21867 16952 22008 16980
rect 21867 16949 21879 16952
rect 21821 16943 21879 16949
rect 22002 16940 22008 16952
rect 22060 16940 22066 16992
rect 22204 16989 22232 17020
rect 23474 17008 23480 17020
rect 23532 17008 23538 17060
rect 23584 17020 23888 17048
rect 22189 16983 22247 16989
rect 22189 16949 22201 16983
rect 22235 16949 22247 16983
rect 22189 16943 22247 16949
rect 22281 16983 22339 16989
rect 22281 16949 22293 16983
rect 22327 16980 22339 16983
rect 23290 16980 23296 16992
rect 22327 16952 23296 16980
rect 22327 16949 22339 16952
rect 22281 16943 22339 16949
rect 23290 16940 23296 16952
rect 23348 16940 23354 16992
rect 23385 16983 23443 16989
rect 23385 16949 23397 16983
rect 23431 16980 23443 16983
rect 23584 16980 23612 17020
rect 23431 16952 23612 16980
rect 23661 16983 23719 16989
rect 23431 16949 23443 16952
rect 23385 16943 23443 16949
rect 23661 16949 23673 16983
rect 23707 16980 23719 16983
rect 23750 16980 23756 16992
rect 23707 16952 23756 16980
rect 23707 16949 23719 16952
rect 23661 16943 23719 16949
rect 23750 16940 23756 16952
rect 23808 16940 23814 16992
rect 23860 16980 23888 17020
rect 24026 16980 24032 16992
rect 23860 16952 24032 16980
rect 24026 16940 24032 16952
rect 24084 16940 24090 16992
rect 24210 16940 24216 16992
rect 24268 16980 24274 16992
rect 24670 16980 24676 16992
rect 24268 16952 24676 16980
rect 24268 16940 24274 16952
rect 24670 16940 24676 16952
rect 24728 16940 24734 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 2222 16736 2228 16788
rect 2280 16776 2286 16788
rect 2958 16776 2964 16788
rect 2280 16748 2820 16776
rect 2919 16748 2964 16776
rect 2280 16736 2286 16748
rect 1670 16668 1676 16720
rect 1728 16708 1734 16720
rect 1765 16711 1823 16717
rect 1765 16708 1777 16711
rect 1728 16680 1777 16708
rect 1728 16668 1734 16680
rect 1765 16677 1777 16680
rect 1811 16677 1823 16711
rect 2406 16708 2412 16720
rect 2367 16680 2412 16708
rect 1765 16671 1823 16677
rect 2406 16668 2412 16680
rect 2464 16708 2470 16720
rect 2685 16711 2743 16717
rect 2685 16708 2697 16711
rect 2464 16680 2697 16708
rect 2464 16668 2470 16680
rect 2685 16677 2697 16680
rect 2731 16677 2743 16711
rect 2792 16708 2820 16748
rect 2958 16736 2964 16748
rect 3016 16736 3022 16788
rect 3881 16779 3939 16785
rect 3881 16745 3893 16779
rect 3927 16776 3939 16779
rect 4338 16776 4344 16788
rect 3927 16748 4344 16776
rect 3927 16745 3939 16748
rect 3881 16739 3939 16745
rect 2869 16711 2927 16717
rect 2869 16708 2881 16711
rect 2792 16680 2881 16708
rect 2685 16671 2743 16677
rect 2869 16677 2881 16680
rect 2915 16708 2927 16711
rect 3896 16708 3924 16739
rect 4338 16736 4344 16748
rect 4396 16736 4402 16788
rect 5629 16779 5687 16785
rect 5629 16776 5641 16779
rect 5460 16748 5641 16776
rect 4706 16708 4712 16720
rect 2915 16680 3924 16708
rect 4448 16680 4712 16708
rect 2915 16677 2927 16680
rect 2869 16671 2927 16677
rect 4154 16600 4160 16652
rect 4212 16640 4218 16652
rect 4448 16649 4476 16680
rect 4706 16668 4712 16680
rect 4764 16668 4770 16720
rect 5460 16649 5488 16748
rect 5629 16745 5641 16748
rect 5675 16745 5687 16779
rect 5629 16739 5687 16745
rect 5997 16779 6055 16785
rect 5997 16745 6009 16779
rect 6043 16776 6055 16779
rect 6086 16776 6092 16788
rect 6043 16748 6092 16776
rect 6043 16745 6055 16748
rect 5997 16739 6055 16745
rect 6086 16736 6092 16748
rect 6144 16776 6150 16788
rect 7190 16776 7196 16788
rect 6144 16748 6408 16776
rect 7151 16748 7196 16776
rect 6144 16736 6150 16748
rect 4433 16643 4491 16649
rect 4433 16640 4445 16643
rect 4212 16612 4445 16640
rect 4212 16600 4218 16612
rect 4433 16609 4445 16612
rect 4479 16609 4491 16643
rect 4433 16603 4491 16609
rect 4525 16643 4583 16649
rect 4525 16609 4537 16643
rect 4571 16640 4583 16643
rect 5445 16643 5503 16649
rect 5445 16640 5457 16643
rect 4571 16612 5457 16640
rect 4571 16609 4583 16612
rect 4525 16603 4583 16609
rect 5445 16609 5457 16612
rect 5491 16609 5503 16643
rect 5445 16603 5503 16609
rect 1857 16575 1915 16581
rect 1857 16541 1869 16575
rect 1903 16572 1915 16575
rect 1946 16572 1952 16584
rect 1903 16544 1952 16572
rect 1903 16541 1915 16544
rect 1857 16535 1915 16541
rect 1946 16532 1952 16544
rect 2004 16532 2010 16584
rect 2041 16575 2099 16581
rect 2041 16541 2053 16575
rect 2087 16572 2099 16575
rect 2130 16572 2136 16584
rect 2087 16544 2136 16572
rect 2087 16541 2099 16544
rect 2041 16535 2099 16541
rect 2130 16532 2136 16544
rect 2188 16532 2194 16584
rect 3418 16532 3424 16584
rect 3476 16572 3482 16584
rect 4617 16575 4675 16581
rect 4617 16572 4629 16575
rect 3476 16544 4629 16572
rect 3476 16532 3482 16544
rect 4617 16541 4629 16544
rect 4663 16541 4675 16575
rect 6086 16572 6092 16584
rect 6047 16544 6092 16572
rect 4617 16535 4675 16541
rect 6086 16532 6092 16544
rect 6144 16532 6150 16584
rect 6178 16532 6184 16584
rect 6236 16572 6242 16584
rect 6236 16544 6281 16572
rect 6236 16532 6242 16544
rect 2685 16507 2743 16513
rect 2685 16473 2697 16507
rect 2731 16504 2743 16507
rect 6380 16504 6408 16748
rect 7190 16736 7196 16748
rect 7248 16736 7254 16788
rect 7653 16779 7711 16785
rect 7653 16745 7665 16779
rect 7699 16776 7711 16779
rect 7742 16776 7748 16788
rect 7699 16748 7748 16776
rect 7699 16745 7711 16748
rect 7653 16739 7711 16745
rect 7742 16736 7748 16748
rect 7800 16736 7806 16788
rect 8386 16776 8392 16788
rect 8347 16748 8392 16776
rect 8386 16736 8392 16748
rect 8444 16736 8450 16788
rect 8570 16736 8576 16788
rect 8628 16776 8634 16788
rect 8665 16779 8723 16785
rect 8665 16776 8677 16779
rect 8628 16748 8677 16776
rect 8628 16736 8634 16748
rect 8665 16745 8677 16748
rect 8711 16745 8723 16779
rect 9030 16776 9036 16788
rect 8991 16748 9036 16776
rect 8665 16739 8723 16745
rect 9030 16736 9036 16748
rect 9088 16736 9094 16788
rect 9398 16776 9404 16788
rect 9359 16748 9404 16776
rect 9398 16736 9404 16748
rect 9456 16736 9462 16788
rect 9950 16736 9956 16788
rect 10008 16736 10014 16788
rect 10134 16736 10140 16788
rect 10192 16776 10198 16788
rect 11057 16779 11115 16785
rect 11057 16776 11069 16779
rect 10192 16748 11069 16776
rect 10192 16736 10198 16748
rect 11057 16745 11069 16748
rect 11103 16745 11115 16779
rect 11330 16776 11336 16788
rect 11291 16748 11336 16776
rect 11057 16739 11115 16745
rect 11330 16736 11336 16748
rect 11388 16736 11394 16788
rect 12894 16736 12900 16788
rect 12952 16776 12958 16788
rect 13725 16779 13783 16785
rect 13725 16776 13737 16779
rect 12952 16748 13737 16776
rect 12952 16736 12958 16748
rect 13725 16745 13737 16748
rect 13771 16745 13783 16779
rect 14366 16776 14372 16788
rect 14327 16748 14372 16776
rect 13725 16739 13783 16745
rect 14366 16736 14372 16748
rect 14424 16736 14430 16788
rect 14642 16776 14648 16788
rect 14603 16748 14648 16776
rect 14642 16736 14648 16748
rect 14700 16736 14706 16788
rect 16574 16736 16580 16788
rect 16632 16776 16638 16788
rect 16669 16779 16727 16785
rect 16669 16776 16681 16779
rect 16632 16748 16681 16776
rect 16632 16736 16638 16748
rect 16669 16745 16681 16748
rect 16715 16745 16727 16779
rect 16669 16739 16727 16745
rect 17221 16779 17279 16785
rect 17221 16745 17233 16779
rect 17267 16776 17279 16779
rect 17402 16776 17408 16788
rect 17267 16748 17408 16776
rect 17267 16745 17279 16748
rect 17221 16739 17279 16745
rect 17402 16736 17408 16748
rect 17460 16736 17466 16788
rect 17497 16779 17555 16785
rect 17497 16745 17509 16779
rect 17543 16776 17555 16779
rect 17862 16776 17868 16788
rect 17543 16748 17868 16776
rect 17543 16745 17555 16748
rect 17497 16739 17555 16745
rect 17862 16736 17868 16748
rect 17920 16736 17926 16788
rect 19518 16736 19524 16788
rect 19576 16776 19582 16788
rect 19889 16779 19947 16785
rect 19889 16776 19901 16779
rect 19576 16748 19901 16776
rect 19576 16736 19582 16748
rect 19889 16745 19901 16748
rect 19935 16745 19947 16779
rect 20346 16776 20352 16788
rect 20307 16748 20352 16776
rect 19889 16739 19947 16745
rect 20346 16736 20352 16748
rect 20404 16736 20410 16788
rect 21269 16779 21327 16785
rect 21269 16745 21281 16779
rect 21315 16776 21327 16779
rect 21358 16776 21364 16788
rect 21315 16748 21364 16776
rect 21315 16745 21327 16748
rect 21269 16739 21327 16745
rect 21358 16736 21364 16748
rect 21416 16736 21422 16788
rect 22370 16736 22376 16788
rect 22428 16736 22434 16788
rect 23109 16779 23167 16785
rect 23109 16745 23121 16779
rect 23155 16776 23167 16779
rect 23382 16776 23388 16788
rect 23155 16748 23388 16776
rect 23155 16745 23167 16748
rect 23109 16739 23167 16745
rect 23382 16736 23388 16748
rect 23440 16736 23446 16788
rect 23658 16736 23664 16788
rect 23716 16776 23722 16788
rect 24765 16779 24823 16785
rect 24765 16776 24777 16779
rect 23716 16748 24777 16776
rect 23716 16736 23722 16748
rect 24765 16745 24777 16748
rect 24811 16745 24823 16779
rect 24765 16739 24823 16745
rect 24854 16736 24860 16788
rect 24912 16776 24918 16788
rect 24949 16779 25007 16785
rect 24949 16776 24961 16779
rect 24912 16748 24961 16776
rect 24912 16736 24918 16748
rect 24949 16745 24961 16748
rect 24995 16745 25007 16779
rect 24949 16739 25007 16745
rect 9968 16708 9996 16736
rect 10226 16708 10232 16720
rect 9968 16680 10232 16708
rect 10226 16668 10232 16680
rect 10284 16668 10290 16720
rect 11348 16708 11376 16736
rect 12066 16708 12072 16720
rect 11348 16680 12072 16708
rect 12066 16668 12072 16680
rect 12124 16708 12130 16720
rect 12314 16711 12372 16717
rect 12314 16708 12326 16711
rect 12124 16680 12326 16708
rect 12124 16668 12130 16680
rect 12314 16677 12326 16680
rect 12360 16708 12372 16711
rect 14090 16708 14096 16720
rect 12360 16680 14096 16708
rect 12360 16677 12372 16680
rect 12314 16671 12372 16677
rect 14090 16668 14096 16680
rect 14148 16668 14154 16720
rect 14550 16668 14556 16720
rect 14608 16708 14614 16720
rect 15013 16711 15071 16717
rect 15013 16708 15025 16711
rect 14608 16680 15025 16708
rect 14608 16668 14614 16680
rect 15013 16677 15025 16680
rect 15059 16677 15071 16711
rect 18776 16711 18834 16717
rect 15013 16671 15071 16677
rect 15120 16680 18644 16708
rect 6638 16640 6644 16652
rect 6599 16612 6644 16640
rect 6638 16600 6644 16612
rect 6696 16600 6702 16652
rect 7009 16643 7067 16649
rect 7009 16640 7021 16643
rect 6840 16612 7021 16640
rect 6546 16532 6552 16584
rect 6604 16572 6610 16584
rect 6840 16572 6868 16612
rect 7009 16609 7021 16612
rect 7055 16609 7067 16643
rect 7009 16603 7067 16609
rect 7561 16643 7619 16649
rect 7561 16609 7573 16643
rect 7607 16640 7619 16643
rect 7650 16640 7656 16652
rect 7607 16612 7656 16640
rect 7607 16609 7619 16612
rect 7561 16603 7619 16609
rect 7650 16600 7656 16612
rect 7708 16600 7714 16652
rect 8754 16600 8760 16652
rect 8812 16640 8818 16652
rect 9950 16649 9956 16652
rect 9944 16640 9956 16649
rect 8812 16612 9956 16640
rect 8812 16600 8818 16612
rect 9944 16603 9956 16612
rect 9950 16600 9956 16603
rect 10008 16600 10014 16652
rect 11793 16643 11851 16649
rect 11793 16609 11805 16643
rect 11839 16640 11851 16643
rect 11882 16640 11888 16652
rect 11839 16612 11888 16640
rect 11839 16609 11851 16612
rect 11793 16603 11851 16609
rect 11882 16600 11888 16612
rect 11940 16600 11946 16652
rect 12084 16612 13124 16640
rect 6604 16544 6868 16572
rect 6604 16532 6610 16544
rect 7466 16532 7472 16584
rect 7524 16572 7530 16584
rect 7745 16575 7803 16581
rect 7745 16572 7757 16575
rect 7524 16544 7757 16572
rect 7524 16532 7530 16544
rect 7745 16541 7757 16544
rect 7791 16541 7803 16575
rect 7745 16535 7803 16541
rect 9582 16532 9588 16584
rect 9640 16572 9646 16584
rect 12084 16581 12112 16612
rect 9677 16575 9735 16581
rect 9677 16572 9689 16575
rect 9640 16544 9689 16572
rect 9640 16532 9646 16544
rect 9677 16541 9689 16544
rect 9723 16541 9735 16575
rect 9677 16535 9735 16541
rect 12069 16575 12127 16581
rect 12069 16541 12081 16575
rect 12115 16541 12127 16575
rect 12069 16535 12127 16541
rect 6638 16504 6644 16516
rect 2731 16476 6644 16504
rect 2731 16473 2743 16476
rect 2685 16467 2743 16473
rect 6638 16464 6644 16476
rect 6696 16464 6702 16516
rect 1397 16439 1455 16445
rect 1397 16405 1409 16439
rect 1443 16436 1455 16439
rect 1854 16436 1860 16448
rect 1443 16408 1860 16436
rect 1443 16405 1455 16408
rect 1397 16399 1455 16405
rect 1854 16396 1860 16408
rect 1912 16396 1918 16448
rect 2038 16396 2044 16448
rect 2096 16436 2102 16448
rect 3418 16436 3424 16448
rect 2096 16408 3424 16436
rect 2096 16396 2102 16408
rect 3418 16396 3424 16408
rect 3476 16396 3482 16448
rect 4062 16436 4068 16448
rect 4023 16408 4068 16436
rect 4062 16396 4068 16408
rect 4120 16396 4126 16448
rect 5166 16436 5172 16448
rect 5127 16408 5172 16436
rect 5166 16396 5172 16408
rect 5224 16396 5230 16448
rect 8294 16396 8300 16448
rect 8352 16436 8358 16448
rect 8570 16436 8576 16448
rect 8352 16408 8576 16436
rect 8352 16396 8358 16408
rect 8570 16396 8576 16408
rect 8628 16436 8634 16448
rect 9692 16436 9720 16535
rect 11330 16504 11336 16516
rect 10612 16476 11336 16504
rect 10612 16436 10640 16476
rect 11330 16464 11336 16476
rect 11388 16504 11394 16516
rect 12084 16504 12112 16535
rect 11388 16476 12112 16504
rect 11388 16464 11394 16476
rect 8628 16408 10640 16436
rect 8628 16396 8634 16408
rect 11790 16396 11796 16448
rect 11848 16436 11854 16448
rect 12434 16436 12440 16448
rect 11848 16408 12440 16436
rect 11848 16396 11854 16408
rect 12434 16396 12440 16408
rect 12492 16396 12498 16448
rect 13096 16436 13124 16612
rect 13262 16600 13268 16652
rect 13320 16640 13326 16652
rect 13630 16640 13636 16652
rect 13320 16612 13636 16640
rect 13320 16600 13326 16612
rect 13630 16600 13636 16612
rect 13688 16640 13694 16652
rect 15120 16640 15148 16680
rect 13688 16612 15148 16640
rect 13688 16600 13694 16612
rect 15194 16600 15200 16652
rect 15252 16640 15258 16652
rect 15289 16643 15347 16649
rect 15289 16640 15301 16643
rect 15252 16612 15301 16640
rect 15252 16600 15258 16612
rect 15289 16609 15301 16612
rect 15335 16609 15347 16643
rect 15289 16603 15347 16609
rect 15556 16643 15614 16649
rect 15556 16609 15568 16643
rect 15602 16640 15614 16643
rect 16298 16640 16304 16652
rect 15602 16612 16304 16640
rect 15602 16609 15614 16612
rect 15556 16603 15614 16609
rect 16298 16600 16304 16612
rect 16356 16640 16362 16652
rect 17034 16640 17040 16652
rect 16356 16612 17040 16640
rect 16356 16600 16362 16612
rect 17034 16600 17040 16612
rect 17092 16600 17098 16652
rect 18046 16600 18052 16652
rect 18104 16640 18110 16652
rect 18509 16643 18567 16649
rect 18509 16640 18521 16643
rect 18104 16612 18521 16640
rect 18104 16600 18110 16612
rect 18509 16609 18521 16612
rect 18555 16609 18567 16643
rect 18616 16640 18644 16680
rect 18776 16677 18788 16711
rect 18822 16708 18834 16711
rect 18874 16708 18880 16720
rect 18822 16680 18880 16708
rect 18822 16677 18834 16680
rect 18776 16671 18834 16677
rect 18874 16668 18880 16680
rect 18932 16668 18938 16720
rect 18966 16668 18972 16720
rect 19024 16708 19030 16720
rect 19150 16708 19156 16720
rect 19024 16680 19156 16708
rect 19024 16668 19030 16680
rect 19150 16668 19156 16680
rect 19208 16668 19214 16720
rect 21542 16668 21548 16720
rect 21600 16717 21606 16720
rect 21600 16711 21664 16717
rect 21600 16677 21618 16711
rect 21652 16677 21664 16711
rect 21600 16671 21664 16677
rect 21600 16668 21606 16671
rect 19610 16640 19616 16652
rect 18616 16612 19616 16640
rect 18509 16603 18567 16609
rect 19610 16600 19616 16612
rect 19668 16600 19674 16652
rect 13906 16532 13912 16584
rect 13964 16572 13970 16584
rect 14274 16572 14280 16584
rect 13964 16544 14280 16572
rect 13964 16532 13970 16544
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 14366 16532 14372 16584
rect 14424 16572 14430 16584
rect 15212 16572 15240 16600
rect 22388 16584 22416 16736
rect 24029 16711 24087 16717
rect 24029 16677 24041 16711
rect 24075 16708 24087 16711
rect 24397 16711 24455 16717
rect 24397 16708 24409 16711
rect 24075 16680 24409 16708
rect 24075 16677 24087 16680
rect 24029 16671 24087 16677
rect 24397 16677 24409 16680
rect 24443 16677 24455 16711
rect 24397 16671 24455 16677
rect 24581 16711 24639 16717
rect 24581 16677 24593 16711
rect 24627 16708 24639 16711
rect 25038 16708 25044 16720
rect 24627 16680 25044 16708
rect 24627 16677 24639 16680
rect 24581 16671 24639 16677
rect 25038 16668 25044 16680
rect 25096 16668 25102 16720
rect 26234 16708 26240 16720
rect 25148 16680 26240 16708
rect 25148 16652 25176 16680
rect 26234 16668 26240 16680
rect 26292 16668 26298 16720
rect 22738 16600 22744 16652
rect 22796 16640 22802 16652
rect 23937 16643 23995 16649
rect 23937 16640 23949 16643
rect 22796 16612 23949 16640
rect 22796 16600 22802 16612
rect 23937 16609 23949 16612
rect 23983 16640 23995 16643
rect 24670 16640 24676 16652
rect 23983 16612 24676 16640
rect 23983 16609 23995 16612
rect 23937 16603 23995 16609
rect 24670 16600 24676 16612
rect 24728 16600 24734 16652
rect 25130 16640 25136 16652
rect 25091 16612 25136 16640
rect 25130 16600 25136 16612
rect 25188 16600 25194 16652
rect 25406 16640 25412 16652
rect 25367 16612 25412 16640
rect 25406 16600 25412 16612
rect 25464 16600 25470 16652
rect 25498 16600 25504 16652
rect 25556 16640 25562 16652
rect 25774 16640 25780 16652
rect 25556 16612 25780 16640
rect 25556 16600 25562 16612
rect 25774 16600 25780 16612
rect 25832 16600 25838 16652
rect 14424 16544 15240 16572
rect 14424 16532 14430 16544
rect 20530 16532 20536 16584
rect 20588 16572 20594 16584
rect 21361 16575 21419 16581
rect 21361 16572 21373 16575
rect 20588 16544 21373 16572
rect 20588 16532 20594 16544
rect 21361 16541 21373 16544
rect 21407 16541 21419 16575
rect 21361 16535 21419 16541
rect 22370 16532 22376 16584
rect 22428 16532 22434 16584
rect 23477 16575 23535 16581
rect 23477 16541 23489 16575
rect 23523 16572 23535 16575
rect 23842 16572 23848 16584
rect 23523 16544 23848 16572
rect 23523 16541 23535 16544
rect 23477 16535 23535 16541
rect 23842 16532 23848 16544
rect 23900 16572 23906 16584
rect 24121 16575 24179 16581
rect 24121 16572 24133 16575
rect 23900 16544 24133 16572
rect 23900 16532 23906 16544
rect 24121 16541 24133 16544
rect 24167 16541 24179 16575
rect 24121 16535 24179 16541
rect 24765 16575 24823 16581
rect 24765 16541 24777 16575
rect 24811 16572 24823 16575
rect 25869 16575 25927 16581
rect 25869 16572 25881 16575
rect 24811 16544 25881 16572
rect 24811 16541 24823 16544
rect 24765 16535 24823 16541
rect 25148 16516 25176 16544
rect 25869 16541 25881 16544
rect 25915 16572 25927 16575
rect 26237 16575 26295 16581
rect 26237 16572 26249 16575
rect 25915 16544 26249 16572
rect 25915 16541 25927 16544
rect 25869 16535 25927 16541
rect 26237 16541 26249 16544
rect 26283 16572 26295 16575
rect 26326 16572 26332 16584
rect 26283 16544 26332 16572
rect 26283 16541 26295 16544
rect 26237 16535 26295 16541
rect 26326 16532 26332 16544
rect 26384 16532 26390 16584
rect 13446 16504 13452 16516
rect 13407 16476 13452 16504
rect 13446 16464 13452 16476
rect 13504 16464 13510 16516
rect 13630 16464 13636 16516
rect 13688 16504 13694 16516
rect 15102 16504 15108 16516
rect 13688 16476 15108 16504
rect 13688 16464 13694 16476
rect 15102 16464 15108 16476
rect 15160 16464 15166 16516
rect 23290 16504 23296 16516
rect 22287 16476 23296 16504
rect 16758 16436 16764 16448
rect 13096 16408 16764 16436
rect 16758 16396 16764 16408
rect 16816 16396 16822 16448
rect 18141 16439 18199 16445
rect 18141 16405 18153 16439
rect 18187 16436 18199 16439
rect 18414 16436 18420 16448
rect 18187 16408 18420 16436
rect 18187 16405 18199 16408
rect 18141 16399 18199 16405
rect 18414 16396 18420 16408
rect 18472 16396 18478 16448
rect 20717 16439 20775 16445
rect 20717 16405 20729 16439
rect 20763 16436 20775 16439
rect 22287 16436 22315 16476
rect 23290 16464 23296 16476
rect 23348 16464 23354 16516
rect 23569 16507 23627 16513
rect 23569 16473 23581 16507
rect 23615 16504 23627 16507
rect 23934 16504 23940 16516
rect 23615 16476 23940 16504
rect 23615 16473 23627 16476
rect 23569 16467 23627 16473
rect 23934 16464 23940 16476
rect 23992 16464 23998 16516
rect 25130 16464 25136 16516
rect 25188 16464 25194 16516
rect 20763 16408 22315 16436
rect 20763 16405 20775 16408
rect 20717 16399 20775 16405
rect 22462 16396 22468 16448
rect 22520 16436 22526 16448
rect 22741 16439 22799 16445
rect 22741 16436 22753 16439
rect 22520 16408 22753 16436
rect 22520 16396 22526 16408
rect 22741 16405 22753 16408
rect 22787 16405 22799 16439
rect 22741 16399 22799 16405
rect 23842 16396 23848 16448
rect 23900 16436 23906 16448
rect 24397 16439 24455 16445
rect 24397 16436 24409 16439
rect 23900 16408 24409 16436
rect 23900 16396 23906 16408
rect 24397 16405 24409 16408
rect 24443 16405 24455 16439
rect 24397 16399 24455 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 934 16192 940 16244
rect 992 16232 998 16244
rect 3326 16232 3332 16244
rect 992 16204 3332 16232
rect 992 16192 998 16204
rect 3326 16192 3332 16204
rect 3384 16192 3390 16244
rect 3418 16192 3424 16244
rect 3476 16232 3482 16244
rect 3881 16235 3939 16241
rect 3881 16232 3893 16235
rect 3476 16204 3893 16232
rect 3476 16192 3482 16204
rect 3881 16201 3893 16204
rect 3927 16201 3939 16235
rect 3881 16195 3939 16201
rect 6089 16235 6147 16241
rect 6089 16201 6101 16235
rect 6135 16232 6147 16235
rect 6638 16232 6644 16244
rect 6135 16204 6644 16232
rect 6135 16201 6147 16204
rect 6089 16195 6147 16201
rect 6638 16192 6644 16204
rect 6696 16192 6702 16244
rect 7742 16192 7748 16244
rect 7800 16232 7806 16244
rect 7929 16235 7987 16241
rect 7929 16232 7941 16235
rect 7800 16204 7941 16232
rect 7800 16192 7806 16204
rect 7929 16201 7941 16204
rect 7975 16201 7987 16235
rect 7929 16195 7987 16201
rect 10134 16192 10140 16244
rect 10192 16232 10198 16244
rect 10321 16235 10379 16241
rect 10321 16232 10333 16235
rect 10192 16204 10333 16232
rect 10192 16192 10198 16204
rect 10321 16201 10333 16204
rect 10367 16201 10379 16235
rect 10502 16232 10508 16244
rect 10463 16204 10508 16232
rect 10321 16195 10379 16201
rect 4433 16167 4491 16173
rect 4433 16133 4445 16167
rect 4479 16164 4491 16167
rect 6454 16164 6460 16176
rect 4479 16136 6460 16164
rect 4479 16133 4491 16136
rect 4433 16127 4491 16133
rect 6454 16124 6460 16136
rect 6512 16164 6518 16176
rect 6512 16136 6776 16164
rect 6512 16124 6518 16136
rect 2038 16096 2044 16108
rect 1999 16068 2044 16096
rect 2038 16056 2044 16068
rect 2096 16056 2102 16108
rect 4341 16099 4399 16105
rect 4341 16065 4353 16099
rect 4387 16096 4399 16099
rect 4985 16099 5043 16105
rect 4985 16096 4997 16099
rect 4387 16068 4997 16096
rect 4387 16065 4399 16068
rect 4341 16059 4399 16065
rect 4985 16065 4997 16068
rect 5031 16096 5043 16099
rect 5350 16096 5356 16108
rect 5031 16068 5356 16096
rect 5031 16065 5043 16068
rect 4985 16059 5043 16065
rect 5350 16056 5356 16068
rect 5408 16056 5414 16108
rect 1762 16028 1768 16040
rect 1723 16000 1768 16028
rect 1762 15988 1768 16000
rect 1820 16028 1826 16040
rect 2222 16028 2228 16040
rect 1820 16000 2228 16028
rect 1820 15988 1826 16000
rect 2222 15988 2228 16000
rect 2280 15988 2286 16040
rect 2958 16028 2964 16040
rect 2919 16000 2964 16028
rect 2958 15988 2964 16000
rect 3016 15988 3022 16040
rect 4801 16031 4859 16037
rect 4801 15997 4813 16031
rect 4847 16028 4859 16031
rect 5442 16028 5448 16040
rect 4847 16000 5448 16028
rect 4847 15997 4859 16000
rect 4801 15991 4859 15997
rect 5442 15988 5448 16000
rect 5500 15988 5506 16040
rect 6748 16028 6776 16136
rect 7098 16096 7104 16108
rect 7059 16068 7104 16096
rect 7098 16056 7104 16068
rect 7156 16056 7162 16108
rect 8294 16056 8300 16108
rect 8352 16096 8358 16108
rect 8352 16068 8397 16096
rect 8352 16056 8358 16068
rect 6825 16031 6883 16037
rect 6825 16028 6837 16031
rect 6748 16000 6837 16028
rect 6825 15997 6837 16000
rect 6871 15997 6883 16031
rect 6825 15991 6883 15997
rect 8386 15988 8392 16040
rect 8444 16028 8450 16040
rect 8553 16031 8611 16037
rect 8553 16028 8565 16031
rect 8444 16000 8565 16028
rect 8444 15988 8450 16000
rect 8553 15997 8565 16000
rect 8599 15997 8611 16031
rect 10336 16028 10364 16195
rect 10502 16192 10508 16204
rect 10560 16192 10566 16244
rect 11609 16235 11667 16241
rect 11609 16232 11621 16235
rect 10980 16204 11621 16232
rect 10980 16105 11008 16204
rect 11609 16201 11621 16204
rect 11655 16232 11667 16235
rect 11790 16232 11796 16244
rect 11655 16204 11796 16232
rect 11655 16201 11667 16204
rect 11609 16195 11667 16201
rect 11790 16192 11796 16204
rect 11848 16192 11854 16244
rect 12066 16232 12072 16244
rect 12027 16204 12072 16232
rect 12066 16192 12072 16204
rect 12124 16192 12130 16244
rect 12989 16235 13047 16241
rect 12989 16201 13001 16235
rect 13035 16232 13047 16235
rect 13078 16232 13084 16244
rect 13035 16204 13084 16232
rect 13035 16201 13047 16204
rect 12989 16195 13047 16201
rect 13078 16192 13084 16204
rect 13136 16192 13142 16244
rect 14366 16232 14372 16244
rect 13740 16204 14372 16232
rect 10965 16099 11023 16105
rect 10965 16065 10977 16099
rect 11011 16065 11023 16099
rect 10965 16059 11023 16065
rect 11057 16099 11115 16105
rect 11057 16065 11069 16099
rect 11103 16065 11115 16099
rect 11057 16059 11115 16065
rect 11072 16028 11100 16059
rect 11606 16056 11612 16108
rect 11664 16096 11670 16108
rect 11790 16096 11796 16108
rect 11664 16068 11796 16096
rect 11664 16056 11670 16068
rect 11790 16056 11796 16068
rect 11848 16056 11854 16108
rect 13630 16056 13636 16108
rect 13688 16096 13694 16108
rect 13740 16105 13768 16204
rect 14366 16192 14372 16204
rect 14424 16192 14430 16244
rect 15654 16192 15660 16244
rect 15712 16232 15718 16244
rect 15749 16235 15807 16241
rect 15749 16232 15761 16235
rect 15712 16204 15761 16232
rect 15712 16192 15718 16204
rect 15749 16201 15761 16204
rect 15795 16232 15807 16235
rect 16298 16232 16304 16244
rect 15795 16204 16304 16232
rect 15795 16201 15807 16204
rect 15749 16195 15807 16201
rect 16298 16192 16304 16204
rect 16356 16232 16362 16244
rect 17034 16232 17040 16244
rect 16356 16204 16436 16232
rect 16947 16204 17040 16232
rect 16356 16192 16362 16204
rect 15105 16167 15163 16173
rect 15105 16133 15117 16167
rect 15151 16164 15163 16167
rect 16206 16164 16212 16176
rect 15151 16136 16212 16164
rect 15151 16133 15163 16136
rect 15105 16127 15163 16133
rect 16206 16124 16212 16136
rect 16264 16124 16270 16176
rect 16408 16105 16436 16204
rect 17034 16192 17040 16204
rect 17092 16232 17098 16244
rect 17862 16232 17868 16244
rect 17092 16204 17868 16232
rect 17092 16192 17098 16204
rect 17862 16192 17868 16204
rect 17920 16192 17926 16244
rect 18874 16192 18880 16244
rect 18932 16232 18938 16244
rect 19061 16235 19119 16241
rect 19061 16232 19073 16235
rect 18932 16204 19073 16232
rect 18932 16192 18938 16204
rect 19061 16201 19073 16204
rect 19107 16201 19119 16235
rect 20530 16232 20536 16244
rect 19061 16195 19119 16201
rect 19628 16204 20536 16232
rect 17497 16167 17555 16173
rect 17497 16133 17509 16167
rect 17543 16164 17555 16167
rect 18046 16164 18052 16176
rect 17543 16136 18052 16164
rect 17543 16133 17555 16136
rect 17497 16127 17555 16133
rect 18046 16124 18052 16136
rect 18104 16124 18110 16176
rect 18598 16124 18604 16176
rect 18656 16164 18662 16176
rect 19628 16164 19656 16204
rect 20530 16192 20536 16204
rect 20588 16192 20594 16244
rect 21821 16235 21879 16241
rect 21821 16201 21833 16235
rect 21867 16232 21879 16235
rect 21910 16232 21916 16244
rect 21867 16204 21916 16232
rect 21867 16201 21879 16204
rect 21821 16195 21879 16201
rect 21910 16192 21916 16204
rect 21968 16192 21974 16244
rect 22094 16192 22100 16244
rect 22152 16232 22158 16244
rect 23382 16232 23388 16244
rect 22152 16204 23244 16232
rect 23343 16204 23388 16232
rect 22152 16192 22158 16204
rect 18656 16136 19656 16164
rect 18656 16124 18662 16136
rect 13725 16099 13783 16105
rect 13725 16096 13737 16099
rect 13688 16068 13737 16096
rect 13688 16056 13694 16068
rect 13725 16065 13737 16068
rect 13771 16065 13783 16099
rect 13725 16059 13783 16065
rect 16393 16099 16451 16105
rect 16393 16065 16405 16099
rect 16439 16065 16451 16099
rect 16393 16059 16451 16065
rect 16485 16099 16543 16105
rect 16485 16065 16497 16099
rect 16531 16065 16543 16099
rect 18690 16096 18696 16108
rect 18651 16068 18696 16096
rect 16485 16059 16543 16065
rect 15381 16031 15439 16037
rect 15381 16028 15393 16031
rect 10336 16000 11100 16028
rect 13832 16000 15393 16028
rect 8553 15991 8611 15997
rect 1670 15920 1676 15972
rect 1728 15960 1734 15972
rect 3234 15960 3240 15972
rect 1728 15932 2912 15960
rect 3195 15932 3240 15960
rect 1728 15920 1734 15932
rect 1394 15892 1400 15904
rect 1355 15864 1400 15892
rect 1394 15852 1400 15864
rect 1452 15852 1458 15904
rect 1854 15892 1860 15904
rect 1815 15864 1860 15892
rect 1854 15852 1860 15864
rect 1912 15852 1918 15904
rect 1946 15852 1952 15904
rect 2004 15892 2010 15904
rect 2501 15895 2559 15901
rect 2501 15892 2513 15895
rect 2004 15864 2513 15892
rect 2004 15852 2010 15864
rect 2501 15861 2513 15864
rect 2547 15892 2559 15895
rect 2682 15892 2688 15904
rect 2547 15864 2688 15892
rect 2547 15861 2559 15864
rect 2501 15855 2559 15861
rect 2682 15852 2688 15864
rect 2740 15852 2746 15904
rect 2884 15901 2912 15932
rect 3234 15920 3240 15932
rect 3292 15920 3298 15972
rect 5721 15963 5779 15969
rect 5721 15929 5733 15963
rect 5767 15960 5779 15963
rect 6086 15960 6092 15972
rect 5767 15932 6092 15960
rect 5767 15929 5779 15932
rect 5721 15923 5779 15929
rect 6086 15920 6092 15932
rect 6144 15960 6150 15972
rect 7190 15960 7196 15972
rect 6144 15932 7196 15960
rect 6144 15920 6150 15932
rect 7190 15920 7196 15932
rect 7248 15920 7254 15972
rect 9950 15960 9956 15972
rect 9692 15932 9956 15960
rect 2869 15895 2927 15901
rect 2869 15861 2881 15895
rect 2915 15892 2927 15895
rect 3694 15892 3700 15904
rect 2915 15864 3700 15892
rect 2915 15861 2927 15864
rect 2869 15855 2927 15861
rect 3694 15852 3700 15864
rect 3752 15852 3758 15904
rect 4893 15895 4951 15901
rect 4893 15861 4905 15895
rect 4939 15892 4951 15895
rect 5534 15892 5540 15904
rect 4939 15864 5540 15892
rect 4939 15861 4951 15864
rect 4893 15855 4951 15861
rect 5534 15852 5540 15864
rect 5592 15852 5598 15904
rect 6270 15852 6276 15904
rect 6328 15892 6334 15904
rect 6549 15895 6607 15901
rect 6549 15892 6561 15895
rect 6328 15864 6561 15892
rect 6328 15852 6334 15864
rect 6549 15861 6561 15864
rect 6595 15892 6607 15895
rect 7466 15892 7472 15904
rect 6595 15864 7472 15892
rect 6595 15861 6607 15864
rect 6549 15855 6607 15861
rect 7466 15852 7472 15864
rect 7524 15852 7530 15904
rect 7650 15892 7656 15904
rect 7611 15864 7656 15892
rect 7650 15852 7656 15864
rect 7708 15852 7714 15904
rect 9692 15901 9720 15932
rect 9950 15920 9956 15932
rect 10008 15960 10014 15972
rect 10045 15963 10103 15969
rect 10045 15960 10057 15963
rect 10008 15932 10057 15960
rect 10008 15920 10014 15932
rect 10045 15929 10057 15932
rect 10091 15960 10103 15963
rect 12437 15963 12495 15969
rect 10091 15932 11008 15960
rect 10091 15929 10103 15932
rect 10045 15923 10103 15929
rect 9677 15895 9735 15901
rect 9677 15861 9689 15895
rect 9723 15861 9735 15895
rect 10870 15892 10876 15904
rect 10831 15864 10876 15892
rect 9677 15855 9735 15861
rect 10870 15852 10876 15864
rect 10928 15852 10934 15904
rect 10980 15892 11008 15932
rect 12437 15929 12449 15963
rect 12483 15960 12495 15963
rect 13832 15960 13860 16000
rect 15381 15997 15393 16000
rect 15427 16028 15439 16031
rect 16301 16031 16359 16037
rect 16301 16028 16313 16031
rect 15427 16000 16313 16028
rect 15427 15997 15439 16000
rect 15381 15991 15439 15997
rect 16301 15997 16313 16000
rect 16347 15997 16359 16031
rect 16301 15991 16359 15997
rect 13992 15963 14050 15969
rect 13992 15960 14004 15963
rect 12483 15932 13860 15960
rect 13924 15932 14004 15960
rect 12483 15929 12495 15932
rect 12437 15923 12495 15929
rect 12802 15892 12808 15904
rect 10980 15864 12808 15892
rect 12802 15852 12808 15864
rect 12860 15852 12866 15904
rect 13633 15895 13691 15901
rect 13633 15861 13645 15895
rect 13679 15892 13691 15895
rect 13924 15892 13952 15932
rect 13992 15929 14004 15932
rect 14038 15960 14050 15963
rect 14366 15960 14372 15972
rect 14038 15932 14372 15960
rect 14038 15929 14050 15932
rect 13992 15923 14050 15929
rect 14366 15920 14372 15932
rect 14424 15920 14430 15972
rect 15654 15920 15660 15972
rect 15712 15960 15718 15972
rect 16206 15960 16212 15972
rect 15712 15932 16212 15960
rect 15712 15920 15718 15932
rect 16206 15920 16212 15932
rect 16264 15960 16270 15972
rect 16500 15960 16528 16059
rect 18690 16056 18696 16068
rect 18748 16056 18754 16108
rect 19628 16105 19656 16136
rect 21361 16167 21419 16173
rect 21361 16133 21373 16167
rect 21407 16164 21419 16167
rect 21542 16164 21548 16176
rect 21407 16136 21548 16164
rect 21407 16133 21419 16136
rect 21361 16127 21419 16133
rect 21542 16124 21548 16136
rect 21600 16164 21606 16176
rect 22738 16164 22744 16176
rect 21600 16136 22744 16164
rect 21600 16124 21606 16136
rect 22738 16124 22744 16136
rect 22796 16124 22802 16176
rect 19613 16099 19671 16105
rect 19613 16065 19625 16099
rect 19659 16065 19671 16099
rect 22462 16096 22468 16108
rect 19613 16059 19671 16065
rect 21652 16068 22468 16096
rect 17586 15988 17592 16040
rect 17644 16028 17650 16040
rect 17681 16031 17739 16037
rect 17681 16028 17693 16031
rect 17644 16000 17693 16028
rect 17644 15988 17650 16000
rect 17681 15997 17693 16000
rect 17727 15997 17739 16031
rect 18414 16028 18420 16040
rect 18375 16000 18420 16028
rect 17681 15991 17739 15997
rect 18414 15988 18420 16000
rect 18472 15988 18478 16040
rect 18509 15963 18567 15969
rect 18509 15960 18521 15963
rect 16264 15932 16528 15960
rect 17328 15932 18521 15960
rect 16264 15920 16270 15932
rect 15930 15892 15936 15904
rect 13679 15864 13952 15892
rect 15891 15864 15936 15892
rect 13679 15861 13691 15864
rect 13633 15855 13691 15861
rect 15930 15852 15936 15864
rect 15988 15852 15994 15904
rect 17126 15852 17132 15904
rect 17184 15892 17190 15904
rect 17328 15901 17356 15932
rect 18509 15929 18521 15932
rect 18555 15960 18567 15963
rect 19058 15960 19064 15972
rect 18555 15932 19064 15960
rect 18555 15929 18567 15932
rect 18509 15923 18567 15929
rect 19058 15920 19064 15932
rect 19116 15920 19122 15972
rect 21652 15969 21680 16068
rect 22462 16056 22468 16068
rect 22520 16056 22526 16108
rect 23216 16028 23244 16204
rect 23382 16192 23388 16204
rect 23440 16192 23446 16244
rect 23474 16192 23480 16244
rect 23532 16232 23538 16244
rect 23661 16235 23719 16241
rect 23661 16232 23673 16235
rect 23532 16204 23673 16232
rect 23532 16192 23538 16204
rect 23661 16201 23673 16204
rect 23707 16201 23719 16235
rect 23661 16195 23719 16201
rect 24670 16192 24676 16244
rect 24728 16232 24734 16244
rect 25409 16235 25467 16241
rect 24728 16204 24808 16232
rect 24728 16192 24734 16204
rect 23400 16164 23428 16192
rect 23400 16136 24164 16164
rect 23382 16056 23388 16108
rect 23440 16096 23446 16108
rect 24026 16096 24032 16108
rect 23440 16068 24032 16096
rect 23440 16056 23446 16068
rect 24026 16056 24032 16068
rect 24084 16056 24090 16108
rect 24136 16105 24164 16136
rect 24121 16099 24179 16105
rect 24121 16065 24133 16099
rect 24167 16065 24179 16099
rect 24121 16059 24179 16065
rect 24305 16099 24363 16105
rect 24305 16065 24317 16099
rect 24351 16096 24363 16099
rect 24670 16096 24676 16108
rect 24351 16068 24676 16096
rect 24351 16065 24363 16068
rect 24305 16059 24363 16065
rect 24670 16056 24676 16068
rect 24728 16056 24734 16108
rect 24780 16105 24808 16204
rect 25409 16201 25421 16235
rect 25455 16232 25467 16235
rect 26050 16232 26056 16244
rect 25455 16204 26056 16232
rect 25455 16201 25467 16204
rect 25409 16195 25467 16201
rect 26050 16192 26056 16204
rect 26108 16192 26114 16244
rect 26234 16232 26240 16244
rect 26195 16204 26240 16232
rect 26234 16192 26240 16204
rect 26292 16192 26298 16244
rect 24765 16099 24823 16105
rect 24765 16065 24777 16099
rect 24811 16096 24823 16099
rect 26326 16096 26332 16108
rect 24811 16068 26332 16096
rect 24811 16065 24823 16068
rect 24765 16059 24823 16065
rect 26326 16056 26332 16068
rect 26384 16056 26390 16108
rect 23474 16028 23480 16040
rect 23216 16000 23480 16028
rect 23474 15988 23480 16000
rect 23532 15988 23538 16040
rect 25222 16028 25228 16040
rect 25183 16000 25228 16028
rect 25222 15988 25228 16000
rect 25280 16028 25286 16040
rect 25777 16031 25835 16037
rect 25777 16028 25789 16031
rect 25280 16000 25789 16028
rect 25280 15988 25286 16000
rect 25777 15997 25789 16000
rect 25823 15997 25835 16031
rect 25777 15991 25835 15997
rect 19521 15963 19579 15969
rect 19521 15929 19533 15963
rect 19567 15960 19579 15963
rect 19858 15963 19916 15969
rect 19858 15960 19870 15963
rect 19567 15932 19870 15960
rect 19567 15929 19579 15932
rect 19521 15923 19579 15929
rect 19858 15929 19870 15932
rect 19904 15960 19916 15963
rect 21637 15963 21695 15969
rect 21637 15960 21649 15963
rect 19904 15932 21649 15960
rect 19904 15929 19916 15932
rect 19858 15923 19916 15929
rect 21637 15929 21649 15932
rect 21683 15929 21695 15963
rect 21637 15923 21695 15929
rect 22094 15920 22100 15972
rect 22152 15960 22158 15972
rect 22281 15963 22339 15969
rect 22281 15960 22293 15963
rect 22152 15932 22293 15960
rect 22152 15920 22158 15932
rect 22281 15929 22293 15932
rect 22327 15960 22339 15963
rect 23566 15960 23572 15972
rect 22327 15932 23572 15960
rect 22327 15929 22339 15932
rect 22281 15923 22339 15929
rect 23566 15920 23572 15932
rect 23624 15920 23630 15972
rect 24029 15963 24087 15969
rect 24029 15929 24041 15963
rect 24075 15960 24087 15963
rect 24075 15932 25084 15960
rect 24075 15929 24087 15932
rect 24029 15923 24087 15929
rect 25056 15904 25084 15932
rect 17313 15895 17371 15901
rect 17313 15892 17325 15895
rect 17184 15864 17325 15892
rect 17184 15852 17190 15864
rect 17313 15861 17325 15864
rect 17359 15861 17371 15895
rect 18046 15892 18052 15904
rect 18007 15864 18052 15892
rect 17313 15855 17371 15861
rect 18046 15852 18052 15864
rect 18104 15852 18110 15904
rect 20990 15892 20996 15904
rect 20951 15864 20996 15892
rect 20990 15852 20996 15864
rect 21048 15852 21054 15904
rect 22002 15852 22008 15904
rect 22060 15892 22066 15904
rect 22186 15892 22192 15904
rect 22060 15864 22192 15892
rect 22060 15852 22066 15864
rect 22186 15852 22192 15864
rect 22244 15852 22250 15904
rect 23109 15895 23167 15901
rect 23109 15861 23121 15895
rect 23155 15892 23167 15895
rect 23842 15892 23848 15904
rect 23155 15864 23848 15892
rect 23155 15861 23167 15864
rect 23109 15855 23167 15861
rect 23842 15852 23848 15864
rect 23900 15852 23906 15904
rect 25038 15892 25044 15904
rect 24999 15864 25044 15892
rect 25038 15852 25044 15864
rect 25096 15852 25102 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 2130 15648 2136 15700
rect 2188 15688 2194 15700
rect 5166 15688 5172 15700
rect 2188 15660 5172 15688
rect 2188 15648 2194 15660
rect 5166 15648 5172 15660
rect 5224 15688 5230 15700
rect 5997 15691 6055 15697
rect 5997 15688 6009 15691
rect 5224 15660 6009 15688
rect 5224 15648 5230 15660
rect 5997 15657 6009 15660
rect 6043 15688 6055 15691
rect 6178 15688 6184 15700
rect 6043 15660 6184 15688
rect 6043 15657 6055 15660
rect 5997 15651 6055 15657
rect 6178 15648 6184 15660
rect 6236 15648 6242 15700
rect 6546 15688 6552 15700
rect 6507 15660 6552 15688
rect 6546 15648 6552 15660
rect 6604 15688 6610 15700
rect 6914 15688 6920 15700
rect 6604 15660 6920 15688
rect 6604 15648 6610 15660
rect 6914 15648 6920 15660
rect 6972 15648 6978 15700
rect 9398 15688 9404 15700
rect 9359 15660 9404 15688
rect 9398 15648 9404 15660
rect 9456 15648 9462 15700
rect 9674 15648 9680 15700
rect 9732 15688 9738 15700
rect 9861 15691 9919 15697
rect 9861 15688 9873 15691
rect 9732 15660 9873 15688
rect 9732 15648 9738 15660
rect 9861 15657 9873 15660
rect 9907 15657 9919 15691
rect 9861 15651 9919 15657
rect 10873 15691 10931 15697
rect 10873 15657 10885 15691
rect 10919 15688 10931 15691
rect 12437 15691 12495 15697
rect 12437 15688 12449 15691
rect 10919 15660 12449 15688
rect 10919 15657 10931 15660
rect 10873 15651 10931 15657
rect 12437 15657 12449 15660
rect 12483 15688 12495 15691
rect 12894 15688 12900 15700
rect 12483 15660 12900 15688
rect 12483 15657 12495 15660
rect 12437 15651 12495 15657
rect 12894 15648 12900 15660
rect 12952 15648 12958 15700
rect 14277 15691 14335 15697
rect 14277 15657 14289 15691
rect 14323 15688 14335 15691
rect 14366 15688 14372 15700
rect 14323 15660 14372 15688
rect 14323 15657 14335 15660
rect 14277 15651 14335 15657
rect 14366 15648 14372 15660
rect 14424 15648 14430 15700
rect 14458 15648 14464 15700
rect 14516 15648 14522 15700
rect 15470 15648 15476 15700
rect 15528 15688 15534 15700
rect 15930 15688 15936 15700
rect 15528 15660 15936 15688
rect 15528 15648 15534 15660
rect 15930 15648 15936 15660
rect 15988 15648 15994 15700
rect 16206 15648 16212 15700
rect 16264 15688 16270 15700
rect 16301 15691 16359 15697
rect 16301 15688 16313 15691
rect 16264 15660 16313 15688
rect 16264 15648 16270 15660
rect 16301 15657 16313 15660
rect 16347 15657 16359 15691
rect 16301 15651 16359 15657
rect 21269 15691 21327 15697
rect 21269 15657 21281 15691
rect 21315 15688 21327 15691
rect 22094 15688 22100 15700
rect 21315 15660 22100 15688
rect 21315 15657 21327 15660
rect 21269 15651 21327 15657
rect 22094 15648 22100 15660
rect 22152 15648 22158 15700
rect 22186 15648 22192 15700
rect 22244 15688 22250 15700
rect 23017 15691 23075 15697
rect 23017 15688 23029 15691
rect 22244 15660 23029 15688
rect 22244 15648 22250 15660
rect 23017 15657 23029 15660
rect 23063 15657 23075 15691
rect 23566 15688 23572 15700
rect 23527 15660 23572 15688
rect 23017 15651 23075 15657
rect 23566 15648 23572 15660
rect 23624 15648 23630 15700
rect 24026 15688 24032 15700
rect 23987 15660 24032 15688
rect 24026 15648 24032 15660
rect 24084 15648 24090 15700
rect 25041 15691 25099 15697
rect 25041 15657 25053 15691
rect 25087 15688 25099 15691
rect 25130 15688 25136 15700
rect 25087 15660 25136 15688
rect 25087 15657 25099 15660
rect 25041 15651 25099 15657
rect 25130 15648 25136 15660
rect 25188 15648 25194 15700
rect 25314 15688 25320 15700
rect 25275 15660 25320 15688
rect 25314 15648 25320 15660
rect 25372 15648 25378 15700
rect 4706 15620 4712 15632
rect 1780 15592 4712 15620
rect 1780 15561 1808 15592
rect 4706 15580 4712 15592
rect 4764 15580 4770 15632
rect 5626 15580 5632 15632
rect 5684 15620 5690 15632
rect 6365 15623 6423 15629
rect 6365 15620 6377 15623
rect 5684 15592 6377 15620
rect 5684 15580 5690 15592
rect 6365 15589 6377 15592
rect 6411 15589 6423 15623
rect 6365 15583 6423 15589
rect 8389 15623 8447 15629
rect 8389 15589 8401 15623
rect 8435 15620 8447 15623
rect 8662 15620 8668 15632
rect 8435 15592 8668 15620
rect 8435 15589 8447 15592
rect 8389 15583 8447 15589
rect 8662 15580 8668 15592
rect 8720 15580 8726 15632
rect 845 15555 903 15561
rect 845 15521 857 15555
rect 891 15552 903 15555
rect 1765 15555 1823 15561
rect 1765 15552 1777 15555
rect 891 15524 1777 15552
rect 891 15521 903 15524
rect 845 15515 903 15521
rect 1765 15521 1777 15524
rect 1811 15521 1823 15555
rect 1765 15515 1823 15521
rect 3510 15512 3516 15564
rect 3568 15512 3574 15564
rect 4614 15561 4620 15564
rect 4608 15552 4620 15561
rect 4575 15524 4620 15552
rect 4608 15515 4620 15524
rect 4614 15512 4620 15515
rect 4672 15512 4678 15564
rect 6917 15555 6975 15561
rect 6917 15521 6929 15555
rect 6963 15552 6975 15555
rect 7929 15555 7987 15561
rect 7929 15552 7941 15555
rect 6963 15524 7941 15552
rect 6963 15521 6975 15524
rect 6917 15515 6975 15521
rect 7929 15521 7941 15524
rect 7975 15521 7987 15555
rect 8110 15552 8116 15564
rect 8071 15524 8116 15552
rect 7929 15515 7987 15521
rect 1670 15444 1676 15496
rect 1728 15484 1734 15496
rect 1857 15487 1915 15493
rect 1857 15484 1869 15487
rect 1728 15456 1869 15484
rect 1728 15444 1734 15456
rect 1857 15453 1869 15456
rect 1903 15453 1915 15487
rect 1857 15447 1915 15453
rect 2041 15487 2099 15493
rect 2041 15453 2053 15487
rect 2087 15453 2099 15487
rect 2041 15447 2099 15453
rect 1397 15351 1455 15357
rect 1397 15317 1409 15351
rect 1443 15348 1455 15351
rect 1762 15348 1768 15360
rect 1443 15320 1768 15348
rect 1443 15317 1455 15320
rect 1397 15311 1455 15317
rect 1762 15308 1768 15320
rect 1820 15308 1826 15360
rect 1946 15308 1952 15360
rect 2004 15348 2010 15360
rect 2056 15348 2084 15447
rect 3142 15376 3148 15428
rect 3200 15416 3206 15428
rect 3528 15416 3556 15512
rect 4341 15487 4399 15493
rect 4341 15453 4353 15487
rect 4387 15453 4399 15487
rect 4341 15447 4399 15453
rect 7009 15487 7067 15493
rect 7009 15453 7021 15487
rect 7055 15453 7067 15487
rect 7009 15447 7067 15453
rect 3697 15419 3755 15425
rect 3697 15416 3709 15419
rect 3200 15388 3709 15416
rect 3200 15376 3206 15388
rect 3697 15385 3709 15388
rect 3743 15385 3755 15419
rect 3697 15379 3755 15385
rect 2409 15351 2467 15357
rect 2409 15348 2421 15351
rect 2004 15320 2421 15348
rect 2004 15308 2010 15320
rect 2409 15317 2421 15320
rect 2455 15317 2467 15351
rect 2958 15348 2964 15360
rect 2919 15320 2964 15348
rect 2409 15311 2467 15317
rect 2958 15308 2964 15320
rect 3016 15308 3022 15360
rect 3418 15348 3424 15360
rect 3379 15320 3424 15348
rect 3418 15308 3424 15320
rect 3476 15308 3482 15360
rect 4356 15348 4384 15447
rect 5721 15419 5779 15425
rect 5721 15385 5733 15419
rect 5767 15416 5779 15419
rect 6086 15416 6092 15428
rect 5767 15388 6092 15416
rect 5767 15385 5779 15388
rect 5721 15379 5779 15385
rect 6086 15376 6092 15388
rect 6144 15376 6150 15428
rect 7024 15416 7052 15447
rect 7098 15444 7104 15496
rect 7156 15484 7162 15496
rect 7944 15484 7972 15515
rect 8110 15512 8116 15524
rect 8168 15512 8174 15564
rect 9416 15552 9444 15648
rect 10410 15580 10416 15632
rect 10468 15620 10474 15632
rect 11054 15620 11060 15632
rect 10468 15592 11060 15620
rect 10468 15580 10474 15592
rect 11054 15580 11060 15592
rect 11112 15580 11118 15632
rect 13164 15623 13222 15629
rect 13164 15589 13176 15623
rect 13210 15620 13222 15623
rect 13446 15620 13452 15632
rect 13210 15592 13452 15620
rect 13210 15589 13222 15592
rect 13164 15583 13222 15589
rect 13446 15580 13452 15592
rect 13504 15580 13510 15632
rect 14476 15620 14504 15648
rect 15657 15623 15715 15629
rect 15657 15620 15669 15623
rect 14476 15592 15669 15620
rect 15657 15589 15669 15592
rect 15703 15620 15715 15623
rect 15838 15620 15844 15632
rect 15703 15592 15844 15620
rect 15703 15589 15715 15592
rect 15657 15583 15715 15589
rect 15838 15580 15844 15592
rect 15896 15580 15902 15632
rect 16117 15623 16175 15629
rect 16117 15589 16129 15623
rect 16163 15620 16175 15623
rect 18049 15623 18107 15629
rect 18049 15620 18061 15623
rect 16163 15592 18061 15620
rect 16163 15589 16175 15592
rect 16117 15583 16175 15589
rect 9677 15555 9735 15561
rect 9677 15552 9689 15555
rect 9416 15524 9689 15552
rect 9677 15521 9689 15524
rect 9723 15521 9735 15555
rect 11238 15552 11244 15564
rect 11151 15524 11244 15552
rect 9677 15515 9735 15521
rect 11238 15512 11244 15524
rect 11296 15552 11302 15564
rect 11606 15552 11612 15564
rect 11296 15524 11612 15552
rect 11296 15512 11302 15524
rect 11606 15512 11612 15524
rect 11664 15512 11670 15564
rect 12897 15555 12955 15561
rect 12897 15521 12909 15555
rect 12943 15552 12955 15555
rect 13630 15552 13636 15564
rect 12943 15524 13636 15552
rect 12943 15521 12955 15524
rect 12897 15515 12955 15521
rect 13630 15512 13636 15524
rect 13688 15512 13694 15564
rect 15286 15512 15292 15564
rect 15344 15552 15350 15564
rect 15470 15552 15476 15564
rect 15344 15524 15476 15552
rect 15344 15512 15350 15524
rect 15470 15512 15476 15524
rect 15528 15512 15534 15564
rect 15749 15555 15807 15561
rect 15749 15521 15761 15555
rect 15795 15552 15807 15555
rect 16206 15552 16212 15564
rect 15795 15524 16212 15552
rect 15795 15521 15807 15524
rect 15749 15515 15807 15521
rect 16206 15512 16212 15524
rect 16264 15512 16270 15564
rect 16574 15512 16580 15564
rect 16632 15552 16638 15564
rect 17405 15555 17463 15561
rect 17405 15552 17417 15555
rect 16632 15524 17417 15552
rect 16632 15512 16638 15524
rect 17405 15521 17417 15524
rect 17451 15521 17463 15555
rect 17405 15515 17463 15521
rect 17497 15555 17555 15561
rect 17497 15521 17509 15555
rect 17543 15552 17555 15555
rect 17862 15552 17868 15564
rect 17543 15524 17868 15552
rect 17543 15521 17555 15524
rect 17497 15515 17555 15521
rect 17862 15512 17868 15524
rect 17920 15512 17926 15564
rect 8202 15484 8208 15496
rect 7156 15456 7201 15484
rect 7944 15456 8208 15484
rect 7156 15444 7162 15456
rect 8202 15444 8208 15456
rect 8260 15444 8266 15496
rect 11054 15444 11060 15496
rect 11112 15484 11118 15496
rect 11333 15487 11391 15493
rect 11333 15484 11345 15487
rect 11112 15456 11345 15484
rect 11112 15444 11118 15456
rect 11333 15453 11345 15456
rect 11379 15453 11391 15487
rect 11333 15447 11391 15453
rect 11422 15444 11428 15496
rect 11480 15484 11486 15496
rect 11882 15484 11888 15496
rect 11480 15456 11888 15484
rect 11480 15444 11486 15456
rect 11882 15444 11888 15456
rect 11940 15444 11946 15496
rect 13906 15444 13912 15496
rect 13964 15484 13970 15496
rect 15933 15487 15991 15493
rect 13964 15456 15424 15484
rect 13964 15444 13970 15456
rect 7024 15388 7696 15416
rect 7668 15360 7696 15388
rect 14366 15376 14372 15428
rect 14424 15416 14430 15428
rect 14645 15419 14703 15425
rect 14645 15416 14657 15419
rect 14424 15388 14657 15416
rect 14424 15376 14430 15388
rect 14645 15385 14657 15388
rect 14691 15416 14703 15419
rect 15289 15419 15347 15425
rect 15289 15416 15301 15419
rect 14691 15388 15301 15416
rect 14691 15385 14703 15388
rect 14645 15379 14703 15385
rect 15289 15385 15301 15388
rect 15335 15385 15347 15419
rect 15289 15379 15347 15385
rect 4522 15348 4528 15360
rect 4356 15320 4528 15348
rect 4522 15308 4528 15320
rect 4580 15348 4586 15360
rect 6546 15348 6552 15360
rect 4580 15320 6552 15348
rect 4580 15308 4586 15320
rect 6546 15308 6552 15320
rect 6604 15348 6610 15360
rect 6822 15348 6828 15360
rect 6604 15320 6828 15348
rect 6604 15308 6610 15320
rect 6822 15308 6828 15320
rect 6880 15308 6886 15360
rect 7650 15348 7656 15360
rect 7611 15320 7656 15348
rect 7650 15308 7656 15320
rect 7708 15308 7714 15360
rect 8386 15308 8392 15360
rect 8444 15348 8450 15360
rect 8849 15351 8907 15357
rect 8849 15348 8861 15351
rect 8444 15320 8861 15348
rect 8444 15308 8450 15320
rect 8849 15317 8861 15320
rect 8895 15317 8907 15351
rect 10318 15348 10324 15360
rect 10279 15320 10324 15348
rect 8849 15311 8907 15317
rect 10318 15308 10324 15320
rect 10376 15308 10382 15360
rect 10686 15348 10692 15360
rect 10647 15320 10692 15348
rect 10686 15308 10692 15320
rect 10744 15308 10750 15360
rect 11422 15308 11428 15360
rect 11480 15348 11486 15360
rect 11885 15351 11943 15357
rect 11885 15348 11897 15351
rect 11480 15320 11897 15348
rect 11480 15308 11486 15320
rect 11885 15317 11897 15320
rect 11931 15317 11943 15351
rect 11885 15311 11943 15317
rect 14826 15308 14832 15360
rect 14884 15348 14890 15360
rect 15013 15351 15071 15357
rect 15013 15348 15025 15351
rect 14884 15320 15025 15348
rect 14884 15308 14890 15320
rect 15013 15317 15025 15320
rect 15059 15317 15071 15351
rect 15396 15348 15424 15456
rect 15933 15453 15945 15487
rect 15979 15484 15991 15487
rect 16390 15484 16396 15496
rect 15979 15456 16396 15484
rect 15979 15453 15991 15456
rect 15933 15447 15991 15453
rect 15654 15376 15660 15428
rect 15712 15416 15718 15428
rect 15948 15416 15976 15447
rect 16390 15444 16396 15456
rect 16448 15444 16454 15496
rect 17678 15484 17684 15496
rect 17639 15456 17684 15484
rect 17678 15444 17684 15456
rect 17736 15444 17742 15496
rect 15712 15388 15976 15416
rect 16853 15419 16911 15425
rect 15712 15376 15718 15388
rect 16853 15385 16865 15419
rect 16899 15416 16911 15419
rect 17696 15416 17724 15444
rect 17972 15428 18000 15592
rect 18049 15589 18061 15592
rect 18095 15589 18107 15623
rect 18049 15583 18107 15589
rect 23477 15623 23535 15629
rect 23477 15589 23489 15623
rect 23523 15620 23535 15623
rect 24670 15620 24676 15632
rect 23523 15592 24676 15620
rect 23523 15589 23535 15592
rect 23477 15583 23535 15589
rect 24670 15580 24676 15592
rect 24728 15580 24734 15632
rect 25148 15620 25176 15648
rect 25685 15623 25743 15629
rect 25685 15620 25697 15623
rect 25148 15592 25697 15620
rect 25332 15564 25360 15592
rect 25685 15589 25697 15592
rect 25731 15620 25743 15623
rect 26053 15623 26111 15629
rect 26053 15620 26065 15623
rect 25731 15592 26065 15620
rect 25731 15589 25743 15592
rect 25685 15583 25743 15589
rect 26053 15589 26065 15592
rect 26099 15589 26111 15623
rect 26053 15583 26111 15589
rect 18509 15555 18567 15561
rect 18509 15521 18521 15555
rect 18555 15552 18567 15555
rect 18690 15552 18696 15564
rect 18555 15524 18696 15552
rect 18555 15521 18567 15524
rect 18509 15515 18567 15521
rect 18690 15512 18696 15524
rect 18748 15552 18754 15564
rect 18868 15555 18926 15561
rect 18868 15552 18880 15555
rect 18748 15524 18880 15552
rect 18748 15512 18754 15524
rect 18868 15521 18880 15524
rect 18914 15552 18926 15555
rect 19150 15552 19156 15564
rect 18914 15524 19156 15552
rect 18914 15521 18926 15524
rect 18868 15515 18926 15521
rect 19150 15512 19156 15524
rect 19208 15512 19214 15564
rect 20622 15512 20628 15564
rect 20680 15552 20686 15564
rect 20717 15555 20775 15561
rect 20717 15552 20729 15555
rect 20680 15524 20729 15552
rect 20680 15512 20686 15524
rect 20717 15521 20729 15524
rect 20763 15521 20775 15555
rect 20717 15515 20775 15521
rect 21174 15512 21180 15564
rect 21232 15552 21238 15564
rect 21628 15555 21686 15561
rect 21628 15552 21640 15555
rect 21232 15524 21640 15552
rect 21232 15512 21238 15524
rect 21628 15521 21640 15524
rect 21674 15552 21686 15555
rect 22002 15552 22008 15564
rect 21674 15524 22008 15552
rect 21674 15521 21686 15524
rect 21628 15515 21686 15521
rect 22002 15512 22008 15524
rect 22060 15512 22066 15564
rect 23934 15552 23940 15564
rect 23895 15524 23940 15552
rect 23934 15512 23940 15524
rect 23992 15512 23998 15564
rect 25130 15552 25136 15564
rect 25091 15524 25136 15552
rect 25130 15512 25136 15524
rect 25188 15512 25194 15564
rect 25314 15512 25320 15564
rect 25372 15512 25378 15564
rect 18598 15484 18604 15496
rect 18559 15456 18604 15484
rect 18598 15444 18604 15456
rect 18656 15444 18662 15496
rect 19978 15444 19984 15496
rect 20036 15484 20042 15496
rect 20257 15487 20315 15493
rect 20257 15484 20269 15487
rect 20036 15456 20269 15484
rect 20036 15444 20042 15456
rect 20257 15453 20269 15456
rect 20303 15453 20315 15487
rect 20257 15447 20315 15453
rect 20346 15444 20352 15496
rect 20404 15444 20410 15496
rect 20530 15444 20536 15496
rect 20588 15484 20594 15496
rect 21361 15487 21419 15493
rect 21361 15484 21373 15487
rect 20588 15456 21373 15484
rect 20588 15444 20594 15456
rect 21361 15453 21373 15456
rect 21407 15453 21419 15487
rect 21361 15447 21419 15453
rect 24121 15487 24179 15493
rect 24121 15453 24133 15487
rect 24167 15453 24179 15487
rect 24121 15447 24179 15453
rect 16899 15388 17724 15416
rect 16899 15385 16911 15388
rect 16853 15379 16911 15385
rect 17954 15376 17960 15428
rect 18012 15376 18018 15428
rect 20070 15376 20076 15428
rect 20128 15416 20134 15428
rect 20364 15416 20392 15444
rect 22738 15416 22744 15428
rect 20128 15388 20392 15416
rect 22651 15388 22744 15416
rect 20128 15376 20134 15388
rect 22738 15376 22744 15388
rect 22796 15416 22802 15428
rect 24136 15416 24164 15447
rect 22796 15388 24164 15416
rect 22796 15376 22802 15388
rect 16117 15351 16175 15357
rect 16117 15348 16129 15351
rect 15396 15320 16129 15348
rect 15013 15311 15071 15317
rect 16117 15317 16129 15320
rect 16163 15317 16175 15351
rect 16117 15311 16175 15317
rect 16942 15308 16948 15360
rect 17000 15348 17006 15360
rect 17037 15351 17095 15357
rect 17037 15348 17049 15351
rect 17000 15320 17049 15348
rect 17000 15308 17006 15320
rect 17037 15317 17049 15320
rect 17083 15317 17095 15351
rect 17037 15311 17095 15317
rect 19981 15351 20039 15357
rect 19981 15317 19993 15351
rect 20027 15348 20039 15351
rect 20346 15348 20352 15360
rect 20027 15320 20352 15348
rect 20027 15317 20039 15320
rect 19981 15311 20039 15317
rect 20346 15308 20352 15320
rect 20404 15308 20410 15360
rect 22922 15308 22928 15360
rect 22980 15348 22986 15360
rect 24581 15351 24639 15357
rect 24581 15348 24593 15351
rect 22980 15320 24593 15348
rect 22980 15308 22986 15320
rect 24581 15317 24593 15320
rect 24627 15317 24639 15351
rect 24581 15311 24639 15317
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 3697 15147 3755 15153
rect 3697 15113 3709 15147
rect 3743 15144 3755 15147
rect 4154 15144 4160 15156
rect 3743 15116 4160 15144
rect 3743 15113 3755 15116
rect 3697 15107 3755 15113
rect 4154 15104 4160 15116
rect 4212 15104 4218 15156
rect 5534 15104 5540 15156
rect 5592 15144 5598 15156
rect 5994 15144 6000 15156
rect 5592 15116 6000 15144
rect 5592 15104 5598 15116
rect 5994 15104 6000 15116
rect 6052 15144 6058 15156
rect 6825 15147 6883 15153
rect 6825 15144 6837 15147
rect 6052 15116 6837 15144
rect 6052 15104 6058 15116
rect 6825 15113 6837 15116
rect 6871 15113 6883 15147
rect 6825 15107 6883 15113
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 8389 15147 8447 15153
rect 8389 15144 8401 15147
rect 8352 15116 8401 15144
rect 8352 15104 8358 15116
rect 8389 15113 8401 15116
rect 8435 15113 8447 15147
rect 8389 15107 8447 15113
rect 8846 15104 8852 15156
rect 8904 15144 8910 15156
rect 9401 15147 9459 15153
rect 9401 15144 9413 15147
rect 8904 15116 9413 15144
rect 8904 15104 8910 15116
rect 9401 15113 9413 15116
rect 9447 15144 9459 15147
rect 9677 15147 9735 15153
rect 9677 15144 9689 15147
rect 9447 15116 9689 15144
rect 9447 15113 9459 15116
rect 9401 15107 9459 15113
rect 9677 15113 9689 15116
rect 9723 15113 9735 15147
rect 9950 15144 9956 15156
rect 9911 15116 9956 15144
rect 9677 15107 9735 15113
rect 9950 15104 9956 15116
rect 10008 15104 10014 15156
rect 11425 15147 11483 15153
rect 11425 15113 11437 15147
rect 11471 15144 11483 15147
rect 11606 15144 11612 15156
rect 11471 15116 11612 15144
rect 11471 15113 11483 15116
rect 11425 15107 11483 15113
rect 11606 15104 11612 15116
rect 11664 15104 11670 15156
rect 11882 15104 11888 15156
rect 11940 15144 11946 15156
rect 11977 15147 12035 15153
rect 11977 15144 11989 15147
rect 11940 15116 11989 15144
rect 11940 15104 11946 15116
rect 11977 15113 11989 15116
rect 12023 15113 12035 15147
rect 11977 15107 12035 15113
rect 12805 15147 12863 15153
rect 12805 15113 12817 15147
rect 12851 15144 12863 15147
rect 13446 15144 13452 15156
rect 12851 15116 13452 15144
rect 12851 15113 12863 15116
rect 12805 15107 12863 15113
rect 13446 15104 13452 15116
rect 13504 15104 13510 15156
rect 14090 15104 14096 15156
rect 14148 15144 14154 15156
rect 15013 15147 15071 15153
rect 15013 15144 15025 15147
rect 14148 15116 15025 15144
rect 14148 15104 14154 15116
rect 15013 15113 15025 15116
rect 15059 15144 15071 15147
rect 15654 15144 15660 15156
rect 15059 15116 15660 15144
rect 15059 15113 15071 15116
rect 15013 15107 15071 15113
rect 15654 15104 15660 15116
rect 15712 15104 15718 15156
rect 16301 15147 16359 15153
rect 16301 15113 16313 15147
rect 16347 15144 16359 15147
rect 16574 15144 16580 15156
rect 16347 15116 16580 15144
rect 16347 15113 16359 15116
rect 16301 15107 16359 15113
rect 16574 15104 16580 15116
rect 16632 15104 16638 15156
rect 17034 15104 17040 15156
rect 17092 15144 17098 15156
rect 18414 15144 18420 15156
rect 17092 15116 18420 15144
rect 17092 15104 17098 15116
rect 18414 15104 18420 15116
rect 18472 15104 18478 15156
rect 19150 15144 19156 15156
rect 19111 15116 19156 15144
rect 19150 15104 19156 15116
rect 19208 15104 19214 15156
rect 19613 15147 19671 15153
rect 19613 15113 19625 15147
rect 19659 15144 19671 15147
rect 20162 15144 20168 15156
rect 19659 15116 20168 15144
rect 19659 15113 19671 15116
rect 19613 15107 19671 15113
rect 20162 15104 20168 15116
rect 20220 15104 20226 15156
rect 20717 15147 20775 15153
rect 20717 15113 20729 15147
rect 20763 15144 20775 15147
rect 21542 15144 21548 15156
rect 20763 15116 21548 15144
rect 20763 15113 20775 15116
rect 20717 15107 20775 15113
rect 21542 15104 21548 15116
rect 21600 15104 21606 15156
rect 22002 15104 22008 15156
rect 22060 15144 22066 15156
rect 22097 15147 22155 15153
rect 22097 15144 22109 15147
rect 22060 15116 22109 15144
rect 22060 15104 22066 15116
rect 22097 15113 22109 15116
rect 22143 15113 22155 15147
rect 22738 15144 22744 15156
rect 22699 15116 22744 15144
rect 22097 15107 22155 15113
rect 22738 15104 22744 15116
rect 22796 15104 22802 15156
rect 23290 15104 23296 15156
rect 23348 15144 23354 15156
rect 23661 15147 23719 15153
rect 23661 15144 23673 15147
rect 23348 15116 23673 15144
rect 23348 15104 23354 15116
rect 23661 15113 23673 15116
rect 23707 15113 23719 15147
rect 23661 15107 23719 15113
rect 24026 15104 24032 15156
rect 24084 15144 24090 15156
rect 24673 15147 24731 15153
rect 24673 15144 24685 15147
rect 24084 15116 24685 15144
rect 24084 15104 24090 15116
rect 24673 15113 24685 15116
rect 24719 15113 24731 15147
rect 24673 15107 24731 15113
rect 25130 15104 25136 15156
rect 25188 15144 25194 15156
rect 25961 15147 26019 15153
rect 25961 15144 25973 15147
rect 25188 15116 25973 15144
rect 25188 15104 25194 15116
rect 25961 15113 25973 15116
rect 26007 15113 26019 15147
rect 25961 15107 26019 15113
rect 1210 15036 1216 15088
rect 1268 15076 1274 15088
rect 2409 15079 2467 15085
rect 2409 15076 2421 15079
rect 1268 15048 2421 15076
rect 1268 15036 1274 15048
rect 2409 15045 2421 15048
rect 2455 15045 2467 15079
rect 2409 15039 2467 15045
rect 6086 15036 6092 15088
rect 6144 15076 6150 15088
rect 6273 15079 6331 15085
rect 6273 15076 6285 15079
rect 6144 15048 6285 15076
rect 6144 15036 6150 15048
rect 6273 15045 6285 15048
rect 6319 15076 6331 15079
rect 6319 15048 7420 15076
rect 6319 15045 6331 15048
rect 6273 15039 6331 15045
rect 2498 14968 2504 15020
rect 2556 15008 2562 15020
rect 2961 15011 3019 15017
rect 2961 15008 2973 15011
rect 2556 14980 2973 15008
rect 2556 14968 2562 14980
rect 2961 14977 2973 14980
rect 3007 14977 3019 15011
rect 4522 15008 4528 15020
rect 4483 14980 4528 15008
rect 2961 14971 3019 14977
rect 4522 14968 4528 14980
rect 4580 14968 4586 15020
rect 1673 14943 1731 14949
rect 1673 14909 1685 14943
rect 1719 14940 1731 14943
rect 2038 14940 2044 14952
rect 1719 14912 2044 14940
rect 1719 14909 1731 14912
rect 1673 14903 1731 14909
rect 2038 14900 2044 14912
rect 2096 14900 2102 14952
rect 2774 14900 2780 14952
rect 2832 14940 2838 14952
rect 4062 14940 4068 14952
rect 2832 14912 4068 14940
rect 2832 14900 2838 14912
rect 4062 14900 4068 14912
rect 4120 14900 4126 14952
rect 4798 14949 4804 14952
rect 4792 14940 4804 14949
rect 4711 14912 4804 14940
rect 3510 14872 3516 14884
rect 1688 14844 3516 14872
rect 1688 14816 1716 14844
rect 3510 14832 3516 14844
rect 3568 14832 3574 14884
rect 3973 14875 4031 14881
rect 3973 14841 3985 14875
rect 4019 14872 4031 14875
rect 4724 14872 4752 14912
rect 4792 14903 4804 14912
rect 4856 14940 4862 14952
rect 6104 14940 6132 15036
rect 6914 14968 6920 15020
rect 6972 15008 6978 15020
rect 7392 15017 7420 15048
rect 11238 15036 11244 15088
rect 11296 15076 11302 15088
rect 11517 15079 11575 15085
rect 11517 15076 11529 15079
rect 11296 15048 11529 15076
rect 11296 15036 11302 15048
rect 11517 15045 11529 15048
rect 11563 15045 11575 15079
rect 13464 15076 13492 15104
rect 15565 15079 15623 15085
rect 13464 15048 14504 15076
rect 11517 15039 11575 15045
rect 14476 15020 14504 15048
rect 15565 15045 15577 15079
rect 15611 15076 15623 15079
rect 15838 15076 15844 15088
rect 15611 15048 15844 15076
rect 15611 15045 15623 15048
rect 15565 15039 15623 15045
rect 15838 15036 15844 15048
rect 15896 15036 15902 15088
rect 16390 15076 16396 15088
rect 16351 15048 16396 15076
rect 16390 15036 16396 15048
rect 16448 15036 16454 15088
rect 17589 15079 17647 15085
rect 17589 15045 17601 15079
rect 17635 15076 17647 15079
rect 17862 15076 17868 15088
rect 17635 15048 17868 15076
rect 17635 15045 17647 15048
rect 17589 15039 17647 15045
rect 17862 15036 17868 15048
rect 17920 15036 17926 15088
rect 19886 15036 19892 15088
rect 19944 15076 19950 15088
rect 20622 15076 20628 15088
rect 19944 15048 20628 15076
rect 19944 15036 19950 15048
rect 20622 15036 20628 15048
rect 20680 15036 20686 15088
rect 21174 15076 21180 15088
rect 21135 15048 21180 15076
rect 21174 15036 21180 15048
rect 21232 15036 21238 15088
rect 7285 15011 7343 15017
rect 7285 15008 7297 15011
rect 6972 14980 7297 15008
rect 6972 14968 6978 14980
rect 7285 14977 7297 14980
rect 7331 14977 7343 15011
rect 7285 14971 7343 14977
rect 7377 15011 7435 15017
rect 7377 14977 7389 15011
rect 7423 14977 7435 15011
rect 7377 14971 7435 14977
rect 7466 14968 7472 15020
rect 7524 15008 7530 15020
rect 7929 15011 7987 15017
rect 7929 15008 7941 15011
rect 7524 14980 7941 15008
rect 7524 14968 7530 14980
rect 7929 14977 7941 14980
rect 7975 15008 7987 15011
rect 9033 15011 9091 15017
rect 9033 15008 9045 15011
rect 7975 14980 9045 15008
rect 7975 14977 7987 14980
rect 7929 14971 7987 14977
rect 9033 14977 9045 14980
rect 9079 15008 9091 15011
rect 10318 15008 10324 15020
rect 9079 14980 10324 15008
rect 9079 14977 9091 14980
rect 9033 14971 9091 14977
rect 10318 14968 10324 14980
rect 10376 15008 10382 15020
rect 10505 15011 10563 15017
rect 10505 15008 10517 15011
rect 10376 14980 10517 15008
rect 10376 14968 10382 14980
rect 10505 14977 10517 14980
rect 10551 14977 10563 15011
rect 14366 15008 14372 15020
rect 14327 14980 14372 15008
rect 10505 14971 10563 14977
rect 14366 14968 14372 14980
rect 14424 14968 14430 15020
rect 14458 14968 14464 15020
rect 14516 15008 14522 15020
rect 15381 15011 15439 15017
rect 14516 14980 14609 15008
rect 14516 14968 14522 14980
rect 15381 14977 15393 15011
rect 15427 15008 15439 15011
rect 16206 15008 16212 15020
rect 15427 14980 16212 15008
rect 15427 14977 15439 14980
rect 15381 14971 15439 14977
rect 16206 14968 16212 14980
rect 16264 14968 16270 15020
rect 16758 14968 16764 15020
rect 16816 15008 16822 15020
rect 16853 15011 16911 15017
rect 16853 15008 16865 15011
rect 16816 14980 16865 15008
rect 16816 14968 16822 14980
rect 16853 14977 16865 14980
rect 16899 14977 16911 15011
rect 16853 14971 16911 14977
rect 17037 15011 17095 15017
rect 17037 14977 17049 15011
rect 17083 15008 17095 15011
rect 17126 15008 17132 15020
rect 17083 14980 17132 15008
rect 17083 14977 17095 14980
rect 17037 14971 17095 14977
rect 17126 14968 17132 14980
rect 17184 14968 17190 15020
rect 17402 14968 17408 15020
rect 17460 15008 17466 15020
rect 17678 15008 17684 15020
rect 17460 14980 17684 15008
rect 17460 14968 17466 14980
rect 17678 14968 17684 14980
rect 17736 15008 17742 15020
rect 18693 15011 18751 15017
rect 18693 15008 18705 15011
rect 17736 14980 18705 15008
rect 17736 14968 17742 14980
rect 18693 14977 18705 14980
rect 18739 14977 18751 15011
rect 18693 14971 18751 14977
rect 4856 14912 6132 14940
rect 4798 14900 4804 14903
rect 4856 14900 4862 14912
rect 6822 14900 6828 14952
rect 6880 14940 6886 14952
rect 7193 14943 7251 14949
rect 7193 14940 7205 14943
rect 6880 14912 7205 14940
rect 6880 14900 6886 14912
rect 7193 14909 7205 14912
rect 7239 14940 7251 14943
rect 8202 14940 8208 14952
rect 7239 14912 8208 14940
rect 7239 14909 7251 14912
rect 7193 14903 7251 14909
rect 8202 14900 8208 14912
rect 8260 14900 8266 14952
rect 8297 14943 8355 14949
rect 8297 14909 8309 14943
rect 8343 14940 8355 14943
rect 8478 14940 8484 14952
rect 8343 14912 8484 14940
rect 8343 14909 8355 14912
rect 8297 14903 8355 14909
rect 8478 14900 8484 14912
rect 8536 14940 8542 14952
rect 8757 14943 8815 14949
rect 8757 14940 8769 14943
rect 8536 14912 8769 14940
rect 8536 14900 8542 14912
rect 8757 14909 8769 14912
rect 8803 14909 8815 14943
rect 11054 14940 11060 14952
rect 10967 14912 11060 14940
rect 8757 14903 8815 14909
rect 11054 14900 11060 14912
rect 11112 14900 11118 14952
rect 11238 14900 11244 14952
rect 11296 14940 11302 14952
rect 11701 14943 11759 14949
rect 11701 14940 11713 14943
rect 11296 14912 11713 14940
rect 11296 14900 11302 14912
rect 11701 14909 11713 14912
rect 11747 14909 11759 14943
rect 11701 14903 11759 14909
rect 13446 14900 13452 14952
rect 13504 14940 13510 14952
rect 13725 14943 13783 14949
rect 13725 14940 13737 14943
rect 13504 14912 13737 14940
rect 13504 14900 13510 14912
rect 13725 14909 13737 14912
rect 13771 14940 13783 14943
rect 13906 14940 13912 14952
rect 13771 14912 13912 14940
rect 13771 14909 13783 14912
rect 13725 14903 13783 14909
rect 13906 14900 13912 14912
rect 13964 14940 13970 14952
rect 14277 14943 14335 14949
rect 14277 14940 14289 14943
rect 13964 14912 14289 14940
rect 13964 14900 13970 14912
rect 14277 14909 14289 14912
rect 14323 14909 14335 14943
rect 15838 14940 15844 14952
rect 14277 14903 14335 14909
rect 14384 14912 15844 14940
rect 6549 14875 6607 14881
rect 6549 14872 6561 14875
rect 4019 14844 4752 14872
rect 5276 14844 6561 14872
rect 4019 14841 4031 14844
rect 3973 14835 4031 14841
rect 5276 14816 5304 14844
rect 6549 14841 6561 14844
rect 6595 14872 6607 14875
rect 7098 14872 7104 14884
rect 6595 14844 7104 14872
rect 6595 14841 6607 14844
rect 6549 14835 6607 14841
rect 7098 14832 7104 14844
rect 7156 14832 7162 14884
rect 8846 14872 8852 14884
rect 8807 14844 8852 14872
rect 8846 14832 8852 14844
rect 8904 14832 8910 14884
rect 9861 14875 9919 14881
rect 9861 14841 9873 14875
rect 9907 14872 9919 14875
rect 10321 14875 10379 14881
rect 10321 14872 10333 14875
rect 9907 14844 10333 14872
rect 9907 14841 9919 14844
rect 9861 14835 9919 14841
rect 10321 14841 10333 14844
rect 10367 14872 10379 14875
rect 10962 14872 10968 14884
rect 10367 14844 10968 14872
rect 10367 14841 10379 14844
rect 10321 14835 10379 14841
rect 10962 14832 10968 14844
rect 11020 14832 11026 14884
rect 11072 14872 11100 14900
rect 14384 14872 14412 14912
rect 15838 14900 15844 14912
rect 15896 14900 15902 14952
rect 17865 14943 17923 14949
rect 17865 14909 17877 14943
rect 17911 14940 17923 14943
rect 18046 14940 18052 14952
rect 17911 14912 18052 14940
rect 17911 14909 17923 14912
rect 17865 14903 17923 14909
rect 18046 14900 18052 14912
rect 18104 14940 18110 14952
rect 18417 14943 18475 14949
rect 18417 14940 18429 14943
rect 18104 14912 18429 14940
rect 18104 14900 18110 14912
rect 18417 14909 18429 14912
rect 18463 14909 18475 14943
rect 18708 14940 18736 14971
rect 19426 14968 19432 15020
rect 19484 15008 19490 15020
rect 19521 15011 19579 15017
rect 19521 15008 19533 15011
rect 19484 14980 19533 15008
rect 19484 14968 19490 14980
rect 19521 14977 19533 14980
rect 19567 15008 19579 15011
rect 20165 15011 20223 15017
rect 20165 15008 20177 15011
rect 19567 14980 20177 15008
rect 19567 14977 19579 14980
rect 19521 14971 19579 14977
rect 20165 14977 20177 14980
rect 20211 14977 20223 15011
rect 21560 15008 21588 15104
rect 22278 15036 22284 15088
rect 22336 15076 22342 15088
rect 22646 15076 22652 15088
rect 22336 15048 22652 15076
rect 22336 15036 22342 15048
rect 22646 15036 22652 15048
rect 22704 15036 22710 15088
rect 23474 15076 23480 15088
rect 23435 15048 23480 15076
rect 23474 15036 23480 15048
rect 23532 15036 23538 15088
rect 23676 15048 25452 15076
rect 21637 15011 21695 15017
rect 21637 15008 21649 15011
rect 21560 14980 21649 15008
rect 20165 14971 20223 14977
rect 21637 14977 21649 14980
rect 21683 14977 21695 15011
rect 21637 14971 21695 14977
rect 21729 15011 21787 15017
rect 21729 14977 21741 15011
rect 21775 14977 21787 15011
rect 21729 14971 21787 14977
rect 18874 14940 18880 14952
rect 18708 14912 18880 14940
rect 18417 14903 18475 14909
rect 18874 14900 18880 14912
rect 18932 14940 18938 14952
rect 20346 14940 20352 14952
rect 18932 14912 20352 14940
rect 18932 14900 18938 14912
rect 20346 14900 20352 14912
rect 20404 14940 20410 14952
rect 21085 14943 21143 14949
rect 21085 14940 21097 14943
rect 20404 14912 21097 14940
rect 20404 14900 20410 14912
rect 21085 14909 21097 14912
rect 21131 14940 21143 14943
rect 21744 14940 21772 14971
rect 21131 14912 21772 14940
rect 21131 14909 21143 14912
rect 21085 14903 21143 14909
rect 22646 14900 22652 14952
rect 22704 14940 22710 14952
rect 23106 14940 23112 14952
rect 22704 14912 23112 14940
rect 22704 14900 22710 14912
rect 23106 14900 23112 14912
rect 23164 14900 23170 14952
rect 23492 14940 23520 15036
rect 23676 15020 23704 15048
rect 23658 14968 23664 15020
rect 23716 14968 23722 15020
rect 24305 15011 24363 15017
rect 24305 14977 24317 15011
rect 24351 15008 24363 15011
rect 24670 15008 24676 15020
rect 24351 14980 24676 15008
rect 24351 14977 24363 14980
rect 24305 14971 24363 14977
rect 24670 14968 24676 14980
rect 24728 14968 24734 15020
rect 25424 15017 25452 15048
rect 25409 15011 25467 15017
rect 25409 14977 25421 15011
rect 25455 14977 25467 15011
rect 25409 14971 25467 14977
rect 24029 14943 24087 14949
rect 24029 14940 24041 14943
rect 23492 14912 24041 14940
rect 24029 14909 24041 14912
rect 24075 14909 24087 14943
rect 25222 14940 25228 14952
rect 25183 14912 25228 14940
rect 24029 14903 24087 14909
rect 25222 14900 25228 14912
rect 25280 14900 25286 14952
rect 11072 14844 14412 14872
rect 15565 14875 15623 14881
rect 15565 14841 15577 14875
rect 15611 14872 15623 14875
rect 15749 14875 15807 14881
rect 15749 14872 15761 14875
rect 15611 14844 15761 14872
rect 15611 14841 15623 14844
rect 15565 14835 15623 14841
rect 15749 14841 15761 14844
rect 15795 14872 15807 14875
rect 16206 14872 16212 14884
rect 15795 14844 16212 14872
rect 15795 14841 15807 14844
rect 15749 14835 15807 14841
rect 16206 14832 16212 14844
rect 16264 14832 16270 14884
rect 16758 14872 16764 14884
rect 16671 14844 16764 14872
rect 16758 14832 16764 14844
rect 16816 14872 16822 14884
rect 17678 14872 17684 14884
rect 16816 14844 17684 14872
rect 16816 14832 16822 14844
rect 17678 14832 17684 14844
rect 17736 14832 17742 14884
rect 17954 14832 17960 14884
rect 18012 14872 18018 14884
rect 18509 14875 18567 14881
rect 18509 14872 18521 14875
rect 18012 14844 18521 14872
rect 18012 14832 18018 14844
rect 18509 14841 18521 14844
rect 18555 14841 18567 14875
rect 20070 14872 20076 14884
rect 20031 14844 20076 14872
rect 18509 14835 18567 14841
rect 20070 14832 20076 14844
rect 20128 14832 20134 14884
rect 20162 14832 20168 14884
rect 20220 14832 20226 14884
rect 23934 14832 23940 14884
rect 23992 14872 23998 14884
rect 25041 14875 25099 14881
rect 25041 14872 25053 14875
rect 23992 14844 25053 14872
rect 23992 14832 23998 14844
rect 25041 14841 25053 14844
rect 25087 14841 25099 14875
rect 25041 14835 25099 14841
rect 1670 14764 1676 14816
rect 1728 14764 1734 14816
rect 1946 14804 1952 14816
rect 1907 14776 1952 14804
rect 1946 14764 1952 14776
rect 2004 14764 2010 14816
rect 2869 14807 2927 14813
rect 2869 14773 2881 14807
rect 2915 14804 2927 14807
rect 3234 14804 3240 14816
rect 2915 14776 3240 14804
rect 2915 14773 2927 14776
rect 2869 14767 2927 14773
rect 3234 14764 3240 14776
rect 3292 14764 3298 14816
rect 4433 14807 4491 14813
rect 4433 14773 4445 14807
rect 4479 14804 4491 14807
rect 4614 14804 4620 14816
rect 4479 14776 4620 14804
rect 4479 14773 4491 14776
rect 4433 14767 4491 14773
rect 4614 14764 4620 14776
rect 4672 14804 4678 14816
rect 5258 14804 5264 14816
rect 4672 14776 5264 14804
rect 4672 14764 4678 14776
rect 5258 14764 5264 14776
rect 5316 14764 5322 14816
rect 5350 14764 5356 14816
rect 5408 14804 5414 14816
rect 5905 14807 5963 14813
rect 5905 14804 5917 14807
rect 5408 14776 5917 14804
rect 5408 14764 5414 14776
rect 5905 14773 5917 14776
rect 5951 14804 5963 14807
rect 6178 14804 6184 14816
rect 5951 14776 6184 14804
rect 5951 14773 5963 14776
rect 5905 14767 5963 14773
rect 6178 14764 6184 14776
rect 6236 14764 6242 14816
rect 9677 14807 9735 14813
rect 9677 14773 9689 14807
rect 9723 14804 9735 14807
rect 10413 14807 10471 14813
rect 10413 14804 10425 14807
rect 9723 14776 10425 14804
rect 9723 14773 9735 14776
rect 9677 14767 9735 14773
rect 10413 14773 10425 14776
rect 10459 14804 10471 14807
rect 11054 14804 11060 14816
rect 10459 14776 11060 14804
rect 10459 14773 10471 14776
rect 10413 14767 10471 14773
rect 11054 14764 11060 14776
rect 11112 14764 11118 14816
rect 12897 14807 12955 14813
rect 12897 14773 12909 14807
rect 12943 14804 12955 14807
rect 13446 14804 13452 14816
rect 12943 14776 13452 14804
rect 12943 14773 12955 14776
rect 12897 14767 12955 14773
rect 13446 14764 13452 14776
rect 13504 14764 13510 14816
rect 13909 14807 13967 14813
rect 13909 14773 13921 14807
rect 13955 14804 13967 14807
rect 14090 14804 14096 14816
rect 13955 14776 14096 14804
rect 13955 14773 13967 14776
rect 13909 14767 13967 14773
rect 14090 14764 14096 14776
rect 14148 14764 14154 14816
rect 15286 14764 15292 14816
rect 15344 14804 15350 14816
rect 17405 14807 17463 14813
rect 17405 14804 17417 14807
rect 15344 14776 17417 14804
rect 15344 14764 15350 14776
rect 17405 14773 17417 14776
rect 17451 14804 17463 14807
rect 17589 14807 17647 14813
rect 17589 14804 17601 14807
rect 17451 14776 17601 14804
rect 17451 14773 17463 14776
rect 17405 14767 17463 14773
rect 17589 14773 17601 14776
rect 17635 14773 17647 14807
rect 17589 14767 17647 14773
rect 17862 14764 17868 14816
rect 17920 14804 17926 14816
rect 18049 14807 18107 14813
rect 18049 14804 18061 14807
rect 17920 14776 18061 14804
rect 17920 14764 17926 14776
rect 18049 14773 18061 14776
rect 18095 14773 18107 14807
rect 19978 14804 19984 14816
rect 19939 14776 19984 14804
rect 18049 14767 18107 14773
rect 19978 14764 19984 14776
rect 20036 14764 20042 14816
rect 20180 14804 20208 14832
rect 20346 14804 20352 14816
rect 20180 14776 20352 14804
rect 20346 14764 20352 14776
rect 20404 14764 20410 14816
rect 21542 14804 21548 14816
rect 21503 14776 21548 14804
rect 21542 14764 21548 14776
rect 21600 14764 21606 14816
rect 22097 14807 22155 14813
rect 22097 14773 22109 14807
rect 22143 14804 22155 14807
rect 22281 14807 22339 14813
rect 22281 14804 22293 14807
rect 22143 14776 22293 14804
rect 22143 14773 22155 14776
rect 22097 14767 22155 14773
rect 22281 14773 22293 14776
rect 22327 14804 22339 14807
rect 23106 14804 23112 14816
rect 22327 14776 23112 14804
rect 22327 14773 22339 14776
rect 22281 14767 22339 14773
rect 23106 14764 23112 14776
rect 23164 14764 23170 14816
rect 24121 14807 24179 14813
rect 24121 14773 24133 14807
rect 24167 14804 24179 14807
rect 24302 14804 24308 14816
rect 24167 14776 24308 14804
rect 24167 14773 24179 14776
rect 24121 14767 24179 14773
rect 24302 14764 24308 14776
rect 24360 14764 24366 14816
rect 26050 14764 26056 14816
rect 26108 14804 26114 14816
rect 26329 14807 26387 14813
rect 26329 14804 26341 14807
rect 26108 14776 26341 14804
rect 26108 14764 26114 14776
rect 26329 14773 26341 14776
rect 26375 14773 26387 14807
rect 26329 14767 26387 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 2774 14560 2780 14612
rect 2832 14600 2838 14612
rect 2832 14572 2877 14600
rect 2832 14560 2838 14572
rect 3510 14560 3516 14612
rect 3568 14600 3574 14612
rect 5721 14603 5779 14609
rect 5721 14600 5733 14603
rect 3568 14572 5733 14600
rect 3568 14560 3574 14572
rect 5721 14569 5733 14572
rect 5767 14569 5779 14603
rect 5721 14563 5779 14569
rect 6457 14603 6515 14609
rect 6457 14569 6469 14603
rect 6503 14600 6515 14603
rect 6546 14600 6552 14612
rect 6503 14572 6552 14600
rect 6503 14569 6515 14572
rect 6457 14563 6515 14569
rect 6546 14560 6552 14572
rect 6604 14560 6610 14612
rect 8481 14603 8539 14609
rect 8481 14569 8493 14603
rect 8527 14600 8539 14603
rect 8846 14600 8852 14612
rect 8527 14572 8852 14600
rect 8527 14569 8539 14572
rect 8481 14563 8539 14569
rect 8846 14560 8852 14572
rect 8904 14560 8910 14612
rect 9122 14560 9128 14612
rect 9180 14600 9186 14612
rect 10134 14600 10140 14612
rect 9180 14572 9996 14600
rect 10095 14572 10140 14600
rect 9180 14560 9186 14572
rect 1394 14492 1400 14544
rect 1452 14532 1458 14544
rect 1857 14535 1915 14541
rect 1857 14532 1869 14535
rect 1452 14504 1869 14532
rect 1452 14492 1458 14504
rect 1857 14501 1869 14504
rect 1903 14501 1915 14535
rect 1857 14495 1915 14501
rect 2225 14535 2283 14541
rect 2225 14501 2237 14535
rect 2271 14532 2283 14535
rect 3789 14535 3847 14541
rect 3789 14532 3801 14535
rect 2271 14504 3801 14532
rect 2271 14501 2283 14504
rect 2225 14495 2283 14501
rect 3789 14501 3801 14504
rect 3835 14501 3847 14535
rect 4522 14532 4528 14544
rect 3789 14495 3847 14501
rect 4080 14504 4528 14532
rect 1762 14464 1768 14476
rect 1723 14436 1768 14464
rect 1762 14424 1768 14436
rect 1820 14424 1826 14476
rect 1872 14464 1900 14495
rect 4080 14473 4108 14504
rect 4522 14492 4528 14504
rect 4580 14492 4586 14544
rect 4706 14492 4712 14544
rect 4764 14532 4770 14544
rect 6089 14535 6147 14541
rect 6089 14532 6101 14535
rect 4764 14504 6101 14532
rect 4764 14492 4770 14504
rect 6089 14501 6101 14504
rect 6135 14501 6147 14535
rect 6089 14495 6147 14501
rect 6178 14492 6184 14544
rect 6236 14532 6242 14544
rect 6978 14535 7036 14541
rect 6978 14532 6990 14535
rect 6236 14504 6990 14532
rect 6236 14492 6242 14504
rect 6978 14501 6990 14504
rect 7024 14501 7036 14535
rect 9968 14532 9996 14572
rect 10134 14560 10140 14572
rect 10192 14560 10198 14612
rect 11146 14560 11152 14612
rect 11204 14600 11210 14612
rect 12066 14600 12072 14612
rect 11204 14572 12072 14600
rect 11204 14560 11210 14572
rect 12066 14560 12072 14572
rect 12124 14560 12130 14612
rect 12529 14603 12587 14609
rect 12529 14569 12541 14603
rect 12575 14600 12587 14603
rect 12802 14600 12808 14612
rect 12575 14572 12808 14600
rect 12575 14569 12587 14572
rect 12529 14563 12587 14569
rect 12802 14560 12808 14572
rect 12860 14600 12866 14612
rect 12986 14600 12992 14612
rect 12860 14572 12992 14600
rect 12860 14560 12866 14572
rect 12986 14560 12992 14572
rect 13044 14560 13050 14612
rect 14458 14600 14464 14612
rect 14419 14572 14464 14600
rect 14458 14560 14464 14572
rect 14516 14560 14522 14612
rect 15102 14600 15108 14612
rect 15063 14572 15108 14600
rect 15102 14560 15108 14572
rect 15160 14560 15166 14612
rect 15654 14600 15660 14612
rect 15615 14572 15660 14600
rect 15654 14560 15660 14572
rect 15712 14560 15718 14612
rect 16853 14603 16911 14609
rect 16853 14569 16865 14603
rect 16899 14600 16911 14603
rect 17586 14600 17592 14612
rect 16899 14572 17592 14600
rect 16899 14569 16911 14572
rect 16853 14563 16911 14569
rect 17586 14560 17592 14572
rect 17644 14560 17650 14612
rect 18874 14600 18880 14612
rect 18835 14572 18880 14600
rect 18874 14560 18880 14572
rect 18932 14600 18938 14612
rect 19058 14600 19064 14612
rect 18932 14572 19064 14600
rect 18932 14560 18938 14572
rect 19058 14560 19064 14572
rect 19116 14560 19122 14612
rect 20070 14560 20076 14612
rect 20128 14600 20134 14612
rect 20257 14603 20315 14609
rect 20257 14600 20269 14603
rect 20128 14572 20269 14600
rect 20128 14560 20134 14572
rect 20257 14569 20269 14572
rect 20303 14569 20315 14603
rect 20622 14600 20628 14612
rect 20583 14572 20628 14600
rect 20257 14563 20315 14569
rect 20622 14560 20628 14572
rect 20680 14560 20686 14612
rect 23845 14603 23903 14609
rect 23845 14569 23857 14603
rect 23891 14600 23903 14603
rect 23934 14600 23940 14612
rect 23891 14572 23940 14600
rect 23891 14569 23903 14572
rect 23845 14563 23903 14569
rect 23934 14560 23940 14572
rect 23992 14560 23998 14612
rect 24026 14560 24032 14612
rect 24084 14600 24090 14612
rect 24210 14600 24216 14612
rect 24084 14572 24216 14600
rect 24084 14560 24090 14572
rect 24210 14560 24216 14572
rect 24268 14560 24274 14612
rect 24302 14560 24308 14612
rect 24360 14560 24366 14612
rect 25038 14560 25044 14612
rect 25096 14600 25102 14612
rect 25409 14603 25467 14609
rect 25409 14600 25421 14603
rect 25096 14572 25421 14600
rect 25096 14560 25102 14572
rect 25409 14569 25421 14572
rect 25455 14569 25467 14603
rect 25409 14563 25467 14569
rect 10045 14535 10103 14541
rect 10045 14532 10057 14535
rect 9968 14504 10057 14532
rect 6978 14495 7036 14501
rect 10045 14501 10057 14504
rect 10091 14532 10103 14535
rect 10962 14532 10968 14544
rect 10091 14504 10968 14532
rect 10091 14501 10103 14504
rect 10045 14495 10103 14501
rect 10962 14492 10968 14504
rect 11020 14492 11026 14544
rect 11882 14492 11888 14544
rect 11940 14492 11946 14544
rect 12084 14532 12112 14560
rect 13173 14535 13231 14541
rect 13173 14532 13185 14535
rect 12084 14504 13185 14532
rect 13173 14501 13185 14504
rect 13219 14501 13231 14535
rect 13173 14495 13231 14501
rect 13630 14492 13636 14544
rect 13688 14532 13694 14544
rect 13906 14532 13912 14544
rect 13688 14504 13912 14532
rect 13688 14492 13694 14504
rect 13906 14492 13912 14504
rect 13964 14532 13970 14544
rect 15286 14532 15292 14544
rect 13964 14504 15292 14532
rect 13964 14492 13970 14504
rect 15286 14492 15292 14504
rect 15344 14532 15350 14544
rect 15749 14535 15807 14541
rect 15749 14532 15761 14535
rect 15344 14504 15761 14532
rect 15344 14492 15350 14504
rect 15749 14501 15761 14504
rect 15795 14501 15807 14535
rect 15749 14495 15807 14501
rect 16485 14535 16543 14541
rect 16485 14501 16497 14535
rect 16531 14532 16543 14535
rect 17126 14532 17132 14544
rect 16531 14504 17132 14532
rect 16531 14501 16543 14504
rect 16485 14495 16543 14501
rect 17126 14492 17132 14504
rect 17184 14492 17190 14544
rect 17402 14541 17408 14544
rect 17396 14532 17408 14541
rect 17363 14504 17408 14532
rect 17396 14495 17408 14504
rect 17402 14492 17408 14495
rect 17460 14492 17466 14544
rect 23658 14532 23664 14544
rect 20180 14504 23664 14532
rect 4338 14473 4344 14476
rect 3421 14467 3479 14473
rect 3421 14464 3433 14467
rect 1872 14436 3433 14464
rect 3421 14433 3433 14436
rect 3467 14433 3479 14467
rect 3421 14427 3479 14433
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14433 4123 14467
rect 4332 14464 4344 14473
rect 4299 14436 4344 14464
rect 4065 14427 4123 14433
rect 4332 14427 4344 14436
rect 1780 14328 1808 14424
rect 1854 14356 1860 14408
rect 1912 14396 1918 14408
rect 1949 14399 2007 14405
rect 1949 14396 1961 14399
rect 1912 14368 1961 14396
rect 1912 14356 1918 14368
rect 1949 14365 1961 14368
rect 1995 14365 2007 14399
rect 1949 14359 2007 14365
rect 2961 14399 3019 14405
rect 2961 14365 2973 14399
rect 3007 14396 3019 14399
rect 3970 14396 3976 14408
rect 3007 14368 3976 14396
rect 3007 14365 3019 14368
rect 2961 14359 3019 14365
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 2225 14331 2283 14337
rect 2225 14328 2237 14331
rect 1780 14300 2237 14328
rect 2225 14297 2237 14300
rect 2271 14297 2283 14331
rect 2225 14291 2283 14297
rect 2774 14288 2780 14340
rect 2832 14328 2838 14340
rect 4080 14328 4108 14427
rect 4338 14424 4344 14427
rect 4396 14424 4402 14476
rect 6638 14464 6644 14476
rect 6599 14436 6644 14464
rect 6638 14424 6644 14436
rect 6696 14424 6702 14476
rect 9125 14467 9183 14473
rect 9125 14433 9137 14467
rect 9171 14464 9183 14467
rect 9306 14464 9312 14476
rect 9171 14436 9312 14464
rect 9171 14433 9183 14436
rect 9125 14427 9183 14433
rect 9306 14424 9312 14436
rect 9364 14424 9370 14476
rect 11606 14464 11612 14476
rect 11567 14436 11612 14464
rect 11606 14424 11612 14436
rect 11664 14424 11670 14476
rect 11900 14464 11928 14492
rect 13265 14467 13323 14473
rect 11900 14436 12112 14464
rect 6546 14356 6552 14408
rect 6604 14396 6610 14408
rect 6733 14399 6791 14405
rect 6733 14396 6745 14399
rect 6604 14368 6745 14396
rect 6604 14356 6610 14368
rect 6733 14365 6745 14368
rect 6779 14365 6791 14399
rect 6733 14359 6791 14365
rect 8110 14356 8116 14408
rect 8168 14356 8174 14408
rect 10229 14399 10287 14405
rect 10229 14365 10241 14399
rect 10275 14365 10287 14399
rect 10229 14359 10287 14365
rect 2832 14300 4108 14328
rect 2832 14288 2838 14300
rect 7742 14288 7748 14340
rect 7800 14328 7806 14340
rect 8128 14328 8156 14356
rect 8757 14331 8815 14337
rect 8757 14328 8769 14331
rect 7800 14300 8769 14328
rect 7800 14288 7806 14300
rect 8757 14297 8769 14300
rect 8803 14297 8815 14331
rect 8757 14291 8815 14297
rect 9493 14331 9551 14337
rect 9493 14297 9505 14331
rect 9539 14328 9551 14331
rect 9950 14328 9956 14340
rect 9539 14300 9956 14328
rect 9539 14297 9551 14300
rect 9493 14291 9551 14297
rect 9950 14288 9956 14300
rect 10008 14328 10014 14340
rect 10244 14328 10272 14359
rect 11422 14356 11428 14408
rect 11480 14396 11486 14408
rect 11701 14399 11759 14405
rect 11701 14396 11713 14399
rect 11480 14368 11713 14396
rect 11480 14356 11486 14368
rect 11701 14365 11713 14368
rect 11747 14365 11759 14399
rect 11882 14396 11888 14408
rect 11843 14368 11888 14396
rect 11701 14359 11759 14365
rect 11882 14356 11888 14368
rect 11940 14356 11946 14408
rect 12084 14396 12112 14436
rect 13265 14433 13277 14467
rect 13311 14464 13323 14467
rect 13446 14464 13452 14476
rect 13311 14436 13452 14464
rect 13311 14433 13323 14436
rect 13265 14427 13323 14433
rect 13446 14424 13452 14436
rect 13504 14424 13510 14476
rect 16666 14424 16672 14476
rect 16724 14464 16730 14476
rect 16850 14464 16856 14476
rect 16724 14436 16856 14464
rect 16724 14424 16730 14436
rect 16850 14424 16856 14436
rect 16908 14424 16914 14476
rect 17034 14464 17040 14476
rect 16995 14436 17040 14464
rect 17034 14424 17040 14436
rect 17092 14424 17098 14476
rect 18690 14424 18696 14476
rect 18748 14464 18754 14476
rect 19242 14464 19248 14476
rect 18748 14436 19248 14464
rect 18748 14424 18754 14436
rect 19242 14424 19248 14436
rect 19300 14424 19306 14476
rect 19605 14467 19663 14473
rect 19605 14433 19617 14467
rect 19651 14433 19663 14467
rect 19605 14427 19663 14433
rect 13078 14396 13084 14408
rect 12084 14368 13084 14396
rect 13078 14356 13084 14368
rect 13136 14396 13142 14408
rect 13357 14399 13415 14405
rect 13357 14396 13369 14399
rect 13136 14368 13369 14396
rect 13136 14356 13142 14368
rect 13357 14365 13369 14368
rect 13403 14365 13415 14399
rect 13357 14359 13415 14365
rect 14458 14356 14464 14408
rect 14516 14396 14522 14408
rect 15841 14399 15899 14405
rect 15841 14396 15853 14399
rect 14516 14368 15853 14396
rect 14516 14356 14522 14368
rect 15841 14365 15853 14368
rect 15887 14365 15899 14399
rect 15841 14359 15899 14365
rect 17129 14399 17187 14405
rect 17129 14365 17141 14399
rect 17175 14365 17187 14399
rect 19334 14396 19340 14408
rect 19295 14368 19340 14396
rect 17129 14359 17187 14365
rect 15102 14328 15108 14340
rect 10008 14300 10272 14328
rect 14016 14300 15108 14328
rect 10008 14288 10014 14300
rect 1394 14260 1400 14272
rect 1355 14232 1400 14260
rect 1394 14220 1400 14232
rect 1452 14220 1458 14272
rect 1854 14220 1860 14272
rect 1912 14260 1918 14272
rect 2409 14263 2467 14269
rect 2409 14260 2421 14263
rect 1912 14232 2421 14260
rect 1912 14220 1918 14232
rect 2409 14229 2421 14232
rect 2455 14260 2467 14263
rect 2498 14260 2504 14272
rect 2455 14232 2504 14260
rect 2455 14229 2467 14232
rect 2409 14223 2467 14229
rect 2498 14220 2504 14232
rect 2556 14220 2562 14272
rect 5258 14220 5264 14272
rect 5316 14260 5322 14272
rect 5445 14263 5503 14269
rect 5445 14260 5457 14263
rect 5316 14232 5457 14260
rect 5316 14220 5322 14232
rect 5445 14229 5457 14232
rect 5491 14229 5503 14263
rect 5445 14223 5503 14229
rect 8018 14220 8024 14272
rect 8076 14260 8082 14272
rect 8113 14263 8171 14269
rect 8113 14260 8125 14263
rect 8076 14232 8125 14260
rect 8076 14220 8082 14232
rect 8113 14229 8125 14232
rect 8159 14229 8171 14263
rect 8938 14260 8944 14272
rect 8899 14232 8944 14260
rect 8113 14223 8171 14229
rect 8938 14220 8944 14232
rect 8996 14220 9002 14272
rect 9582 14220 9588 14272
rect 9640 14260 9646 14272
rect 9677 14263 9735 14269
rect 9677 14260 9689 14263
rect 9640 14232 9689 14260
rect 9640 14220 9646 14232
rect 9677 14229 9689 14232
rect 9723 14229 9735 14263
rect 10870 14260 10876 14272
rect 10831 14232 10876 14260
rect 9677 14223 9735 14229
rect 10870 14220 10876 14232
rect 10928 14220 10934 14272
rect 11238 14260 11244 14272
rect 11199 14232 11244 14260
rect 11238 14220 11244 14232
rect 11296 14220 11302 14272
rect 12802 14260 12808 14272
rect 12763 14232 12808 14260
rect 12802 14220 12808 14232
rect 12860 14220 12866 14272
rect 13630 14220 13636 14272
rect 13688 14260 13694 14272
rect 14016 14269 14044 14300
rect 15102 14288 15108 14300
rect 15160 14288 15166 14340
rect 15286 14328 15292 14340
rect 15247 14300 15292 14328
rect 15286 14288 15292 14300
rect 15344 14288 15350 14340
rect 14001 14263 14059 14269
rect 14001 14260 14013 14263
rect 13688 14232 14013 14260
rect 13688 14220 13694 14232
rect 14001 14229 14013 14232
rect 14047 14229 14059 14263
rect 17144 14260 17172 14359
rect 19334 14356 19340 14368
rect 19392 14356 19398 14408
rect 19628 14396 19656 14427
rect 19708 14424 19714 14476
rect 19766 14473 19772 14476
rect 19766 14467 19788 14473
rect 19776 14433 19788 14467
rect 19766 14427 19788 14433
rect 19766 14424 19772 14427
rect 20180 14408 20208 14504
rect 23658 14492 23664 14504
rect 23716 14492 23722 14544
rect 23753 14535 23811 14541
rect 23753 14501 23765 14535
rect 23799 14532 23811 14535
rect 24320 14532 24348 14560
rect 23799 14504 24348 14532
rect 24949 14535 25007 14541
rect 23799 14501 23811 14504
rect 23753 14495 23811 14501
rect 24949 14501 24961 14535
rect 24995 14532 25007 14535
rect 25314 14532 25320 14544
rect 24995 14504 25320 14532
rect 24995 14501 25007 14504
rect 24949 14495 25007 14501
rect 25314 14492 25320 14504
rect 25372 14492 25378 14544
rect 21174 14424 21180 14476
rect 21232 14464 21238 14476
rect 21893 14467 21951 14473
rect 21893 14464 21905 14467
rect 21232 14436 21905 14464
rect 21232 14424 21238 14436
rect 21893 14433 21905 14436
rect 21939 14433 21951 14467
rect 24210 14464 24216 14476
rect 24171 14436 24216 14464
rect 21893 14427 21951 14433
rect 24210 14424 24216 14436
rect 24268 14424 24274 14476
rect 24305 14467 24363 14473
rect 24305 14433 24317 14467
rect 24351 14464 24363 14467
rect 24762 14464 24768 14476
rect 24351 14436 24768 14464
rect 24351 14433 24363 14436
rect 24305 14427 24363 14433
rect 24762 14424 24768 14436
rect 24820 14424 24826 14476
rect 25038 14424 25044 14476
rect 25096 14464 25102 14476
rect 25590 14464 25596 14476
rect 25096 14436 25596 14464
rect 25096 14424 25102 14436
rect 25590 14424 25596 14436
rect 25648 14424 25654 14476
rect 19978 14396 19984 14408
rect 19628 14368 19984 14396
rect 19978 14356 19984 14368
rect 20036 14356 20042 14408
rect 20162 14356 20168 14408
rect 20220 14356 20226 14408
rect 20530 14356 20536 14408
rect 20588 14396 20594 14408
rect 21634 14396 21640 14408
rect 20588 14368 21640 14396
rect 20588 14356 20594 14368
rect 21634 14356 21640 14368
rect 21692 14356 21698 14408
rect 23106 14396 23112 14408
rect 23019 14368 23112 14396
rect 19889 14331 19947 14337
rect 19889 14297 19901 14331
rect 19935 14328 19947 14331
rect 20438 14328 20444 14340
rect 19935 14300 20444 14328
rect 19935 14297 19947 14300
rect 19889 14291 19947 14297
rect 20438 14288 20444 14300
rect 20496 14288 20502 14340
rect 18046 14260 18052 14272
rect 17144 14232 18052 14260
rect 14001 14223 14059 14229
rect 18046 14220 18052 14232
rect 18104 14220 18110 14272
rect 18509 14263 18567 14269
rect 18509 14229 18521 14263
rect 18555 14260 18567 14263
rect 18598 14260 18604 14272
rect 18555 14232 18604 14260
rect 18555 14229 18567 14232
rect 18509 14223 18567 14229
rect 18598 14220 18604 14232
rect 18656 14220 18662 14272
rect 19242 14220 19248 14272
rect 19300 14260 19306 14272
rect 19429 14263 19487 14269
rect 19429 14260 19441 14263
rect 19300 14232 19441 14260
rect 19300 14220 19306 14232
rect 19429 14229 19441 14232
rect 19475 14260 19487 14263
rect 20548 14260 20576 14356
rect 23032 14337 23060 14368
rect 23106 14356 23112 14368
rect 23164 14396 23170 14408
rect 23385 14399 23443 14405
rect 23385 14396 23397 14399
rect 23164 14368 23397 14396
rect 23164 14356 23170 14368
rect 23385 14365 23397 14368
rect 23431 14396 23443 14399
rect 24489 14399 24547 14405
rect 24489 14396 24501 14399
rect 23431 14368 24501 14396
rect 23431 14365 23443 14368
rect 23385 14359 23443 14365
rect 24489 14365 24501 14368
rect 24535 14396 24547 14399
rect 24670 14396 24676 14408
rect 24535 14368 24676 14396
rect 24535 14365 24547 14368
rect 24489 14359 24547 14365
rect 24670 14356 24676 14368
rect 24728 14356 24734 14408
rect 23017 14331 23075 14337
rect 23017 14297 23029 14331
rect 23063 14297 23075 14331
rect 23017 14291 23075 14297
rect 21174 14260 21180 14272
rect 19475 14232 20576 14260
rect 21135 14232 21180 14260
rect 19475 14229 19487 14232
rect 19429 14223 19487 14229
rect 21174 14220 21180 14232
rect 21232 14220 21238 14272
rect 21542 14260 21548 14272
rect 21503 14232 21548 14260
rect 21542 14220 21548 14232
rect 21600 14220 21606 14272
rect 22002 14220 22008 14272
rect 22060 14260 22066 14272
rect 23382 14260 23388 14272
rect 22060 14232 23388 14260
rect 22060 14220 22066 14232
rect 23382 14220 23388 14232
rect 23440 14220 23446 14272
rect 23842 14220 23848 14272
rect 23900 14260 23906 14272
rect 24670 14260 24676 14272
rect 23900 14232 24676 14260
rect 23900 14220 23906 14232
rect 24670 14220 24676 14232
rect 24728 14220 24734 14272
rect 25222 14260 25228 14272
rect 25183 14232 25228 14260
rect 25222 14220 25228 14232
rect 25280 14220 25286 14272
rect 25961 14263 26019 14269
rect 25961 14229 25973 14263
rect 26007 14260 26019 14263
rect 26050 14260 26056 14272
rect 26007 14232 26056 14260
rect 26007 14229 26019 14232
rect 25961 14223 26019 14229
rect 26050 14220 26056 14232
rect 26108 14260 26114 14272
rect 26237 14263 26295 14269
rect 26237 14260 26249 14263
rect 26108 14232 26249 14260
rect 26108 14220 26114 14232
rect 26237 14229 26249 14232
rect 26283 14229 26295 14263
rect 26237 14223 26295 14229
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 4798 14056 4804 14068
rect 4759 14028 4804 14056
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 4985 14059 5043 14065
rect 4985 14025 4997 14059
rect 5031 14056 5043 14059
rect 5442 14056 5448 14068
rect 5031 14028 5448 14056
rect 5031 14025 5043 14028
rect 4985 14019 5043 14025
rect 5442 14016 5448 14028
rect 5500 14016 5506 14068
rect 6178 14056 6184 14068
rect 6139 14028 6184 14056
rect 6178 14016 6184 14028
rect 6236 14016 6242 14068
rect 6822 14056 6828 14068
rect 6783 14028 6828 14056
rect 6822 14016 6828 14028
rect 6880 14016 6886 14068
rect 8846 14016 8852 14068
rect 8904 14056 8910 14068
rect 9953 14059 10011 14065
rect 9953 14056 9965 14059
rect 8904 14028 9965 14056
rect 8904 14016 8910 14028
rect 9953 14025 9965 14028
rect 9999 14025 10011 14059
rect 9953 14019 10011 14025
rect 10134 14016 10140 14068
rect 10192 14056 10198 14068
rect 10229 14059 10287 14065
rect 10229 14056 10241 14059
rect 10192 14028 10241 14056
rect 10192 14016 10198 14028
rect 10229 14025 10241 14028
rect 10275 14025 10287 14059
rect 11882 14056 11888 14068
rect 11843 14028 11888 14056
rect 10229 14019 10287 14025
rect 2314 13948 2320 14000
rect 2372 13988 2378 14000
rect 2774 13988 2780 14000
rect 2372 13960 2780 13988
rect 2372 13948 2378 13960
rect 2774 13948 2780 13960
rect 2832 13948 2838 14000
rect 4157 13991 4215 13997
rect 4157 13957 4169 13991
rect 4203 13957 4215 13991
rect 4157 13951 4215 13957
rect 1670 13920 1676 13932
rect 1631 13892 1676 13920
rect 1670 13880 1676 13892
rect 1728 13880 1734 13932
rect 1489 13855 1547 13861
rect 1489 13821 1501 13855
rect 1535 13852 1547 13855
rect 1762 13852 1768 13864
rect 1535 13824 1768 13852
rect 1535 13821 1547 13824
rect 1489 13815 1547 13821
rect 1762 13812 1768 13824
rect 1820 13812 1826 13864
rect 2774 13812 2780 13864
rect 2832 13852 2838 13864
rect 4172 13852 4200 13951
rect 4816 13920 4844 14016
rect 5537 13923 5595 13929
rect 5537 13920 5549 13923
rect 4816 13892 5549 13920
rect 5537 13889 5549 13892
rect 5583 13889 5595 13923
rect 5537 13883 5595 13889
rect 7098 13880 7104 13932
rect 7156 13920 7162 13932
rect 7377 13923 7435 13929
rect 7377 13920 7389 13923
rect 7156 13892 7389 13920
rect 7156 13880 7162 13892
rect 7377 13889 7389 13892
rect 7423 13920 7435 13923
rect 7837 13923 7895 13929
rect 7837 13920 7849 13923
rect 7423 13892 7849 13920
rect 7423 13889 7435 13892
rect 7377 13883 7435 13889
rect 7837 13889 7849 13892
rect 7883 13889 7895 13923
rect 7837 13883 7895 13889
rect 8018 13880 8024 13932
rect 8076 13920 8082 13932
rect 8481 13923 8539 13929
rect 8481 13920 8493 13923
rect 8076 13892 8493 13920
rect 8076 13880 8082 13892
rect 8481 13889 8493 13892
rect 8527 13920 8539 13923
rect 8527 13892 8708 13920
rect 8527 13889 8539 13892
rect 8481 13883 8539 13889
rect 4338 13852 4344 13864
rect 2832 13824 2877 13852
rect 4172 13824 4344 13852
rect 2832 13812 2838 13824
rect 4338 13812 4344 13824
rect 4396 13852 4402 13864
rect 4525 13855 4583 13861
rect 4525 13852 4537 13855
rect 4396 13824 4537 13852
rect 4396 13812 4402 13824
rect 4525 13821 4537 13824
rect 4571 13852 4583 13855
rect 6641 13855 6699 13861
rect 4571 13824 5488 13852
rect 4571 13821 4583 13824
rect 4525 13815 4583 13821
rect 2130 13744 2136 13796
rect 2188 13784 2194 13796
rect 2593 13787 2651 13793
rect 2593 13784 2605 13787
rect 2188 13756 2605 13784
rect 2188 13744 2194 13756
rect 2593 13753 2605 13756
rect 2639 13753 2651 13787
rect 2593 13747 2651 13753
rect 2866 13744 2872 13796
rect 2924 13784 2930 13796
rect 3022 13787 3080 13793
rect 3022 13784 3034 13787
rect 2924 13756 3034 13784
rect 2924 13744 2930 13756
rect 3022 13753 3034 13756
rect 3068 13753 3080 13787
rect 5460 13784 5488 13824
rect 6641 13821 6653 13855
rect 6687 13852 6699 13855
rect 6687 13824 6776 13852
rect 6687 13821 6699 13824
rect 6641 13815 6699 13821
rect 5994 13784 6000 13796
rect 5460 13756 6000 13784
rect 3022 13747 3080 13753
rect 5994 13744 6000 13756
rect 6052 13744 6058 13796
rect 6748 13784 6776 13824
rect 6822 13812 6828 13864
rect 6880 13852 6886 13864
rect 7285 13855 7343 13861
rect 7285 13852 7297 13855
rect 6880 13824 7297 13852
rect 6880 13812 6886 13824
rect 7285 13821 7297 13824
rect 7331 13821 7343 13855
rect 8570 13852 8576 13864
rect 8531 13824 8576 13852
rect 7285 13815 7343 13821
rect 8570 13812 8576 13824
rect 8628 13812 8634 13864
rect 8680 13852 8708 13892
rect 8840 13855 8898 13861
rect 8840 13852 8852 13855
rect 8680 13824 8852 13852
rect 8840 13821 8852 13824
rect 8886 13852 8898 13855
rect 9950 13852 9956 13864
rect 8886 13824 9956 13852
rect 8886 13821 8898 13824
rect 8840 13815 8898 13821
rect 9950 13812 9956 13824
rect 10008 13812 10014 13864
rect 10244 13852 10272 14019
rect 11882 14016 11888 14028
rect 11940 14016 11946 14068
rect 12066 14016 12072 14068
rect 12124 14056 12130 14068
rect 12161 14059 12219 14065
rect 12161 14056 12173 14059
rect 12124 14028 12173 14056
rect 12124 14016 12130 14028
rect 12161 14025 12173 14028
rect 12207 14056 12219 14059
rect 12342 14056 12348 14068
rect 12207 14028 12348 14056
rect 12207 14025 12219 14028
rect 12161 14019 12219 14025
rect 12342 14016 12348 14028
rect 12400 14016 12406 14068
rect 12437 14059 12495 14065
rect 12437 14025 12449 14059
rect 12483 14056 12495 14059
rect 12618 14056 12624 14068
rect 12483 14028 12624 14056
rect 12483 14025 12495 14028
rect 12437 14019 12495 14025
rect 12618 14016 12624 14028
rect 12676 14016 12682 14068
rect 13630 14056 13636 14068
rect 13591 14028 13636 14056
rect 13630 14016 13636 14028
rect 13688 14016 13694 14068
rect 14001 14059 14059 14065
rect 14001 14025 14013 14059
rect 14047 14056 14059 14059
rect 14642 14056 14648 14068
rect 14047 14028 14648 14056
rect 14047 14025 14059 14028
rect 14001 14019 14059 14025
rect 14642 14016 14648 14028
rect 14700 14016 14706 14068
rect 15654 14056 15660 14068
rect 15615 14028 15660 14056
rect 15654 14016 15660 14028
rect 15712 14016 15718 14068
rect 16390 14056 16396 14068
rect 16351 14028 16396 14056
rect 16390 14016 16396 14028
rect 16448 14016 16454 14068
rect 17402 14056 17408 14068
rect 17363 14028 17408 14056
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 19426 14056 19432 14068
rect 19387 14028 19432 14056
rect 19426 14016 19432 14028
rect 19484 14016 19490 14068
rect 19702 14056 19708 14068
rect 19663 14028 19708 14056
rect 19702 14016 19708 14028
rect 19760 14016 19766 14068
rect 20346 14016 20352 14068
rect 20404 14056 20410 14068
rect 20714 14056 20720 14068
rect 20404 14028 20720 14056
rect 20404 14016 20410 14028
rect 20714 14016 20720 14028
rect 20772 14016 20778 14068
rect 20898 14056 20904 14068
rect 20859 14028 20904 14056
rect 20898 14016 20904 14028
rect 20956 14016 20962 14068
rect 22649 14059 22707 14065
rect 22649 14025 22661 14059
rect 22695 14056 22707 14059
rect 22738 14056 22744 14068
rect 22695 14028 22744 14056
rect 22695 14025 22707 14028
rect 22649 14019 22707 14025
rect 22738 14016 22744 14028
rect 22796 14016 22802 14068
rect 23014 14056 23020 14068
rect 22975 14028 23020 14056
rect 23014 14016 23020 14028
rect 23072 14016 23078 14068
rect 23658 14056 23664 14068
rect 23619 14028 23664 14056
rect 23658 14016 23664 14028
rect 23716 14016 23722 14068
rect 24210 14016 24216 14068
rect 24268 14056 24274 14068
rect 24673 14059 24731 14065
rect 24673 14056 24685 14059
rect 24268 14028 24685 14056
rect 24268 14016 24274 14028
rect 24673 14025 24685 14028
rect 24719 14025 24731 14059
rect 24673 14019 24731 14025
rect 10781 13991 10839 13997
rect 10781 13957 10793 13991
rect 10827 13988 10839 13991
rect 10962 13988 10968 14000
rect 10827 13960 10968 13988
rect 10827 13957 10839 13960
rect 10781 13951 10839 13957
rect 10962 13948 10968 13960
rect 11020 13948 11026 14000
rect 11146 13948 11152 14000
rect 11204 13988 11210 14000
rect 13446 13988 13452 14000
rect 11204 13960 12195 13988
rect 13407 13960 13452 13988
rect 11204 13948 11210 13960
rect 10870 13880 10876 13932
rect 10928 13920 10934 13932
rect 11425 13923 11483 13929
rect 11425 13920 11437 13923
rect 10928 13892 11437 13920
rect 10928 13880 10934 13892
rect 11425 13889 11437 13892
rect 11471 13920 11483 13923
rect 12066 13920 12072 13932
rect 11471 13892 12072 13920
rect 11471 13889 11483 13892
rect 11425 13883 11483 13889
rect 12066 13880 12072 13892
rect 12124 13880 12130 13932
rect 10689 13855 10747 13861
rect 10244 13824 10640 13852
rect 7193 13787 7251 13793
rect 7193 13784 7205 13787
rect 6748 13756 7205 13784
rect 7193 13753 7205 13756
rect 7239 13784 7251 13787
rect 8754 13784 8760 13796
rect 7239 13756 8760 13784
rect 7239 13753 7251 13756
rect 7193 13747 7251 13753
rect 8754 13744 8760 13756
rect 8812 13744 8818 13796
rect 9398 13744 9404 13796
rect 9456 13784 9462 13796
rect 9674 13784 9680 13796
rect 9456 13756 9680 13784
rect 9456 13744 9462 13756
rect 9674 13744 9680 13756
rect 9732 13744 9738 13796
rect 10612 13784 10640 13824
rect 10689 13821 10701 13855
rect 10735 13852 10747 13855
rect 10778 13852 10784 13864
rect 10735 13824 10784 13852
rect 10735 13821 10747 13824
rect 10689 13815 10747 13821
rect 10778 13812 10784 13824
rect 10836 13852 10842 13864
rect 11241 13855 11299 13861
rect 11241 13852 11253 13855
rect 10836 13824 11253 13852
rect 10836 13812 10842 13824
rect 11241 13821 11253 13824
rect 11287 13821 11299 13855
rect 12167 13852 12195 13960
rect 13446 13948 13452 13960
rect 13504 13948 13510 14000
rect 13906 13948 13912 14000
rect 13964 13988 13970 14000
rect 15289 13991 15347 13997
rect 15289 13988 15301 13991
rect 13964 13960 15301 13988
rect 13964 13948 13970 13960
rect 15289 13957 15301 13960
rect 15335 13957 15347 13991
rect 15289 13951 15347 13957
rect 21174 13948 21180 14000
rect 21232 13988 21238 14000
rect 21821 13991 21879 13997
rect 21821 13988 21833 13991
rect 21232 13960 21833 13988
rect 21232 13948 21238 13960
rect 12894 13920 12900 13932
rect 12855 13892 12900 13920
rect 12894 13880 12900 13892
rect 12952 13880 12958 13932
rect 12986 13880 12992 13932
rect 13044 13920 13050 13932
rect 14642 13920 14648 13932
rect 13044 13892 13089 13920
rect 14603 13892 14648 13920
rect 13044 13880 13050 13892
rect 14642 13880 14648 13892
rect 14700 13880 14706 13932
rect 16301 13923 16359 13929
rect 16301 13889 16313 13923
rect 16347 13920 16359 13923
rect 17037 13923 17095 13929
rect 17037 13920 17049 13923
rect 16347 13892 17049 13920
rect 16347 13889 16359 13892
rect 16301 13883 16359 13889
rect 17037 13889 17049 13892
rect 17083 13920 17095 13923
rect 17126 13920 17132 13932
rect 17083 13892 17132 13920
rect 17083 13889 17095 13892
rect 17037 13883 17095 13889
rect 17126 13880 17132 13892
rect 17184 13920 17190 13932
rect 21468 13929 21496 13960
rect 21821 13957 21833 13960
rect 21867 13988 21879 13991
rect 21913 13991 21971 13997
rect 21913 13988 21925 13991
rect 21867 13960 21925 13988
rect 21867 13957 21879 13960
rect 21821 13951 21879 13957
rect 21913 13957 21925 13960
rect 21959 13957 21971 13991
rect 21913 13951 21971 13957
rect 22373 13991 22431 13997
rect 22373 13957 22385 13991
rect 22419 13988 22431 13991
rect 22922 13988 22928 14000
rect 22419 13960 22928 13988
rect 22419 13957 22431 13960
rect 22373 13951 22431 13957
rect 22922 13948 22928 13960
rect 22980 13948 22986 14000
rect 17773 13923 17831 13929
rect 17773 13920 17785 13923
rect 17184 13892 17785 13920
rect 17184 13880 17190 13892
rect 17773 13889 17785 13892
rect 17819 13920 17831 13923
rect 21453 13923 21511 13929
rect 17819 13892 18184 13920
rect 17819 13889 17831 13892
rect 17773 13883 17831 13889
rect 13909 13855 13967 13861
rect 12167 13824 12480 13852
rect 11241 13815 11299 13821
rect 10870 13784 10876 13796
rect 10612 13756 10876 13784
rect 10870 13744 10876 13756
rect 10928 13744 10934 13796
rect 11149 13787 11207 13793
rect 11149 13753 11161 13787
rect 11195 13784 11207 13787
rect 11330 13784 11336 13796
rect 11195 13756 11336 13784
rect 11195 13753 11207 13756
rect 11149 13747 11207 13753
rect 11330 13744 11336 13756
rect 11388 13744 11394 13796
rect 12452 13784 12480 13824
rect 13909 13821 13921 13855
rect 13955 13852 13967 13855
rect 14458 13852 14464 13864
rect 13955 13824 14464 13852
rect 13955 13821 13967 13824
rect 13909 13815 13967 13821
rect 14458 13812 14464 13824
rect 14516 13812 14522 13864
rect 16850 13852 16856 13864
rect 16763 13824 16856 13852
rect 16850 13812 16856 13824
rect 16908 13852 16914 13864
rect 17862 13852 17868 13864
rect 16908 13824 17868 13852
rect 16908 13812 16914 13824
rect 17862 13812 17868 13824
rect 17920 13812 17926 13864
rect 18046 13852 18052 13864
rect 18007 13824 18052 13852
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 18156 13852 18184 13892
rect 21453 13889 21465 13923
rect 21499 13889 21511 13923
rect 24213 13923 24271 13929
rect 24213 13920 24225 13923
rect 21453 13883 21511 13889
rect 23400 13892 24225 13920
rect 18316 13855 18374 13861
rect 18316 13852 18328 13855
rect 18156 13824 18328 13852
rect 18316 13821 18328 13824
rect 18362 13852 18374 13855
rect 18598 13852 18604 13864
rect 18362 13824 18604 13852
rect 18362 13821 18374 13824
rect 18316 13815 18374 13821
rect 18598 13812 18604 13824
rect 18656 13812 18662 13864
rect 20714 13852 20720 13864
rect 20675 13824 20720 13852
rect 20714 13812 20720 13824
rect 20772 13852 20778 13864
rect 21361 13855 21419 13861
rect 21361 13852 21373 13855
rect 20772 13824 21373 13852
rect 20772 13812 20778 13824
rect 21361 13821 21373 13824
rect 21407 13821 21419 13855
rect 21361 13815 21419 13821
rect 21818 13812 21824 13864
rect 21876 13812 21882 13864
rect 22465 13855 22523 13861
rect 22465 13821 22477 13855
rect 22511 13852 22523 13855
rect 23014 13852 23020 13864
rect 22511 13824 23020 13852
rect 22511 13821 22523 13824
rect 22465 13815 22523 13821
rect 23014 13812 23020 13824
rect 23072 13812 23078 13864
rect 12452 13756 15240 13784
rect 1854 13676 1860 13728
rect 1912 13716 1918 13728
rect 2225 13719 2283 13725
rect 2225 13716 2237 13719
rect 1912 13688 2237 13716
rect 1912 13676 1918 13688
rect 2225 13685 2237 13688
rect 2271 13685 2283 13719
rect 5350 13716 5356 13728
rect 5311 13688 5356 13716
rect 2225 13679 2283 13685
rect 5350 13676 5356 13688
rect 5408 13676 5414 13728
rect 5445 13719 5503 13725
rect 5445 13685 5457 13719
rect 5491 13716 5503 13719
rect 5534 13716 5540 13728
rect 5491 13688 5540 13716
rect 5491 13685 5503 13688
rect 5445 13679 5503 13685
rect 5534 13676 5540 13688
rect 5592 13676 5598 13728
rect 8570 13676 8576 13728
rect 8628 13716 8634 13728
rect 11238 13716 11244 13728
rect 8628 13688 11244 13716
rect 8628 13676 8634 13688
rect 11238 13676 11244 13688
rect 11296 13676 11302 13728
rect 12802 13716 12808 13728
rect 12763 13688 12808 13716
rect 12802 13676 12808 13688
rect 12860 13676 12866 13728
rect 12894 13676 12900 13728
rect 12952 13716 12958 13728
rect 13633 13719 13691 13725
rect 13633 13716 13645 13719
rect 12952 13688 13645 13716
rect 12952 13676 12958 13688
rect 13633 13685 13645 13688
rect 13679 13716 13691 13719
rect 14369 13719 14427 13725
rect 14369 13716 14381 13719
rect 13679 13688 14381 13716
rect 13679 13685 13691 13688
rect 13633 13679 13691 13685
rect 14369 13685 14381 13688
rect 14415 13685 14427 13719
rect 15212 13716 15240 13756
rect 16390 13744 16396 13796
rect 16448 13784 16454 13796
rect 16666 13784 16672 13796
rect 16448 13756 16672 13784
rect 16448 13744 16454 13756
rect 16666 13744 16672 13756
rect 16724 13744 16730 13796
rect 16761 13787 16819 13793
rect 16761 13753 16773 13787
rect 16807 13784 16819 13787
rect 16942 13784 16948 13796
rect 16807 13756 16948 13784
rect 16807 13753 16819 13756
rect 16761 13747 16819 13753
rect 16942 13744 16948 13756
rect 17000 13744 17006 13796
rect 17126 13744 17132 13796
rect 17184 13784 17190 13796
rect 20441 13787 20499 13793
rect 20441 13784 20453 13787
rect 17184 13756 20453 13784
rect 17184 13744 17190 13756
rect 20441 13753 20453 13756
rect 20487 13784 20499 13787
rect 21269 13787 21327 13793
rect 21269 13784 21281 13787
rect 20487 13756 21281 13784
rect 20487 13753 20499 13756
rect 20441 13747 20499 13753
rect 21269 13753 21281 13756
rect 21315 13784 21327 13787
rect 21836 13784 21864 13812
rect 21315 13756 21864 13784
rect 21315 13753 21327 13756
rect 21269 13747 21327 13753
rect 23290 13744 23296 13796
rect 23348 13784 23354 13796
rect 23400 13784 23428 13892
rect 24213 13889 24225 13892
rect 24259 13889 24271 13923
rect 24213 13883 24271 13889
rect 25130 13880 25136 13932
rect 25188 13920 25194 13932
rect 25409 13923 25467 13929
rect 25409 13920 25421 13923
rect 25188 13892 25421 13920
rect 25188 13880 25194 13892
rect 25409 13889 25421 13892
rect 25455 13889 25467 13923
rect 25409 13883 25467 13889
rect 25222 13852 25228 13864
rect 25183 13824 25228 13852
rect 25222 13812 25228 13824
rect 25280 13852 25286 13864
rect 25961 13855 26019 13861
rect 25961 13852 25973 13855
rect 25280 13824 25973 13852
rect 25280 13812 25286 13824
rect 25961 13821 25973 13824
rect 26007 13821 26019 13855
rect 25961 13815 26019 13821
rect 24121 13787 24179 13793
rect 24121 13784 24133 13787
rect 23348 13756 23428 13784
rect 23492 13756 24133 13784
rect 23348 13744 23354 13756
rect 18690 13716 18696 13728
rect 15212 13688 18696 13716
rect 14369 13679 14427 13685
rect 18690 13676 18696 13688
rect 18748 13676 18754 13728
rect 21821 13719 21879 13725
rect 21821 13685 21833 13719
rect 21867 13716 21879 13719
rect 22186 13716 22192 13728
rect 21867 13688 22192 13716
rect 21867 13685 21879 13688
rect 21821 13679 21879 13685
rect 22186 13676 22192 13688
rect 22244 13676 22250 13728
rect 22738 13676 22744 13728
rect 22796 13716 22802 13728
rect 23385 13719 23443 13725
rect 23385 13716 23397 13719
rect 22796 13688 23397 13716
rect 22796 13676 22802 13688
rect 23385 13685 23397 13688
rect 23431 13716 23443 13719
rect 23492 13716 23520 13756
rect 24121 13753 24133 13756
rect 24167 13753 24179 13787
rect 24121 13747 24179 13753
rect 23431 13688 23520 13716
rect 23431 13685 23443 13688
rect 23385 13679 23443 13685
rect 23934 13676 23940 13728
rect 23992 13716 23998 13728
rect 24029 13719 24087 13725
rect 24029 13716 24041 13719
rect 23992 13688 24041 13716
rect 23992 13676 23998 13688
rect 24029 13685 24041 13688
rect 24075 13716 24087 13719
rect 25041 13719 25099 13725
rect 25041 13716 25053 13719
rect 24075 13688 25053 13716
rect 24075 13685 24087 13688
rect 24029 13679 24087 13685
rect 25041 13685 25053 13688
rect 25087 13685 25099 13719
rect 25041 13679 25099 13685
rect 26050 13676 26056 13728
rect 26108 13716 26114 13728
rect 26329 13719 26387 13725
rect 26329 13716 26341 13719
rect 26108 13688 26341 13716
rect 26108 13676 26114 13688
rect 26329 13685 26341 13688
rect 26375 13685 26387 13719
rect 26329 13679 26387 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 2409 13515 2467 13521
rect 2409 13481 2421 13515
rect 2455 13512 2467 13515
rect 3142 13512 3148 13524
rect 2455 13484 3148 13512
rect 2455 13481 2467 13484
rect 2409 13475 2467 13481
rect 3142 13472 3148 13484
rect 3200 13472 3206 13524
rect 4154 13472 4160 13524
rect 4212 13512 4218 13524
rect 4433 13515 4491 13521
rect 4433 13512 4445 13515
rect 4212 13484 4445 13512
rect 4212 13472 4218 13484
rect 4433 13481 4445 13484
rect 4479 13481 4491 13515
rect 4433 13475 4491 13481
rect 5537 13515 5595 13521
rect 5537 13481 5549 13515
rect 5583 13512 5595 13515
rect 5626 13512 5632 13524
rect 5583 13484 5632 13512
rect 5583 13481 5595 13484
rect 5537 13475 5595 13481
rect 5626 13472 5632 13484
rect 5684 13472 5690 13524
rect 6365 13515 6423 13521
rect 6365 13481 6377 13515
rect 6411 13512 6423 13515
rect 6457 13515 6515 13521
rect 6457 13512 6469 13515
rect 6411 13484 6469 13512
rect 6411 13481 6423 13484
rect 6365 13475 6423 13481
rect 6457 13481 6469 13484
rect 6503 13512 6515 13515
rect 6822 13512 6828 13524
rect 6503 13484 6828 13512
rect 6503 13481 6515 13484
rect 6457 13475 6515 13481
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 6917 13515 6975 13521
rect 6917 13481 6929 13515
rect 6963 13512 6975 13515
rect 7006 13512 7012 13524
rect 6963 13484 7012 13512
rect 6963 13481 6975 13484
rect 6917 13475 6975 13481
rect 2590 13404 2596 13456
rect 2648 13444 2654 13456
rect 2774 13444 2780 13456
rect 2648 13416 2780 13444
rect 2648 13404 2654 13416
rect 2774 13404 2780 13416
rect 2832 13444 2838 13456
rect 6932 13444 6960 13475
rect 7006 13472 7012 13484
rect 7064 13472 7070 13524
rect 8018 13512 8024 13524
rect 7979 13484 8024 13512
rect 8018 13472 8024 13484
rect 8076 13472 8082 13524
rect 8389 13515 8447 13521
rect 8389 13481 8401 13515
rect 8435 13512 8447 13515
rect 8662 13512 8668 13524
rect 8435 13484 8668 13512
rect 8435 13481 8447 13484
rect 8389 13475 8447 13481
rect 8662 13472 8668 13484
rect 8720 13512 8726 13524
rect 9677 13515 9735 13521
rect 9677 13512 9689 13515
rect 8720 13484 9689 13512
rect 8720 13472 8726 13484
rect 9677 13481 9689 13484
rect 9723 13481 9735 13515
rect 9677 13475 9735 13481
rect 9766 13472 9772 13524
rect 9824 13512 9830 13524
rect 10137 13515 10195 13521
rect 10137 13512 10149 13515
rect 9824 13484 10149 13512
rect 9824 13472 9830 13484
rect 10137 13481 10149 13484
rect 10183 13512 10195 13515
rect 10778 13512 10784 13524
rect 10183 13484 10784 13512
rect 10183 13481 10195 13484
rect 10137 13475 10195 13481
rect 10778 13472 10784 13484
rect 10836 13472 10842 13524
rect 10873 13515 10931 13521
rect 10873 13481 10885 13515
rect 10919 13512 10931 13515
rect 11330 13512 11336 13524
rect 10919 13484 11336 13512
rect 10919 13481 10931 13484
rect 10873 13475 10931 13481
rect 11330 13472 11336 13484
rect 11388 13472 11394 13524
rect 12250 13472 12256 13524
rect 12308 13512 12314 13524
rect 12434 13512 12440 13524
rect 12308 13484 12440 13512
rect 12308 13472 12314 13484
rect 12434 13472 12440 13484
rect 12492 13472 12498 13524
rect 12802 13472 12808 13524
rect 12860 13512 12866 13524
rect 14645 13515 14703 13521
rect 14645 13512 14657 13515
rect 12860 13484 14657 13512
rect 12860 13472 12866 13484
rect 14645 13481 14657 13484
rect 14691 13481 14703 13515
rect 15930 13512 15936 13524
rect 14645 13475 14703 13481
rect 14752 13484 15936 13512
rect 2832 13416 2925 13444
rect 6656 13416 6960 13444
rect 2832 13404 2838 13416
rect 2869 13379 2927 13385
rect 2869 13345 2881 13379
rect 2915 13376 2927 13379
rect 3142 13376 3148 13388
rect 2915 13348 3148 13376
rect 2915 13345 2927 13348
rect 2869 13339 2927 13345
rect 3142 13336 3148 13348
rect 3200 13376 3206 13388
rect 3878 13376 3884 13388
rect 3200 13348 3884 13376
rect 3200 13336 3206 13348
rect 3878 13336 3884 13348
rect 3936 13336 3942 13388
rect 3970 13336 3976 13388
rect 4028 13376 4034 13388
rect 5077 13379 5135 13385
rect 5077 13376 5089 13379
rect 4028 13348 5089 13376
rect 4028 13336 4034 13348
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13277 3111 13311
rect 3510 13308 3516 13320
rect 3471 13280 3516 13308
rect 3053 13271 3111 13277
rect 1673 13175 1731 13181
rect 1673 13141 1685 13175
rect 1719 13172 1731 13175
rect 1762 13172 1768 13184
rect 1719 13144 1768 13172
rect 1719 13141 1731 13144
rect 1673 13135 1731 13141
rect 1762 13132 1768 13144
rect 1820 13132 1826 13184
rect 2038 13132 2044 13184
rect 2096 13172 2102 13184
rect 2317 13175 2375 13181
rect 2317 13172 2329 13175
rect 2096 13144 2329 13172
rect 2096 13132 2102 13144
rect 2317 13141 2329 13144
rect 2363 13172 2375 13175
rect 3068 13172 3096 13271
rect 3510 13268 3516 13280
rect 3568 13268 3574 13320
rect 4522 13308 4528 13320
rect 4483 13280 4528 13308
rect 4522 13268 4528 13280
rect 4580 13268 4586 13320
rect 4632 13317 4660 13348
rect 5077 13345 5089 13348
rect 5123 13376 5135 13379
rect 5258 13376 5264 13388
rect 5123 13348 5264 13376
rect 5123 13345 5135 13348
rect 5077 13339 5135 13345
rect 5258 13336 5264 13348
rect 5316 13336 5322 13388
rect 4617 13311 4675 13317
rect 4617 13277 4629 13311
rect 4663 13277 4675 13311
rect 4617 13271 4675 13277
rect 6454 13268 6460 13320
rect 6512 13308 6518 13320
rect 6656 13308 6684 13416
rect 8294 13404 8300 13456
rect 8352 13444 8358 13456
rect 8481 13447 8539 13453
rect 8481 13444 8493 13447
rect 8352 13416 8493 13444
rect 8352 13404 8358 13416
rect 8481 13413 8493 13416
rect 8527 13444 8539 13447
rect 9582 13444 9588 13456
rect 8527 13416 9588 13444
rect 8527 13413 8539 13416
rect 8481 13407 8539 13413
rect 9582 13404 9588 13416
rect 9640 13404 9646 13456
rect 11514 13404 11520 13456
rect 11572 13444 11578 13456
rect 11698 13453 11704 13456
rect 11670 13447 11704 13453
rect 11670 13444 11682 13447
rect 11572 13416 11682 13444
rect 11572 13404 11578 13416
rect 11670 13413 11682 13416
rect 11756 13444 11762 13456
rect 13078 13444 13084 13456
rect 11756 13416 11818 13444
rect 13039 13416 13084 13444
rect 11670 13407 11704 13413
rect 11698 13404 11704 13407
rect 11756 13404 11762 13416
rect 13078 13404 13084 13416
rect 13136 13404 13142 13456
rect 13446 13444 13452 13456
rect 13407 13416 13452 13444
rect 13446 13404 13452 13416
rect 13504 13404 13510 13456
rect 14001 13447 14059 13453
rect 14001 13413 14013 13447
rect 14047 13444 14059 13447
rect 14090 13444 14096 13456
rect 14047 13416 14096 13444
rect 14047 13413 14059 13416
rect 14001 13407 14059 13413
rect 14090 13404 14096 13416
rect 14148 13404 14154 13456
rect 14274 13404 14280 13456
rect 14332 13444 14338 13456
rect 14752 13444 14780 13484
rect 15930 13472 15936 13484
rect 15988 13472 15994 13524
rect 16850 13472 16856 13524
rect 16908 13512 16914 13524
rect 16945 13515 17003 13521
rect 16945 13512 16957 13515
rect 16908 13484 16957 13512
rect 16908 13472 16914 13484
rect 16945 13481 16957 13484
rect 16991 13481 17003 13515
rect 16945 13475 17003 13481
rect 17034 13472 17040 13524
rect 17092 13512 17098 13524
rect 17313 13515 17371 13521
rect 17313 13512 17325 13515
rect 17092 13484 17325 13512
rect 17092 13472 17098 13484
rect 17313 13481 17325 13484
rect 17359 13512 17371 13515
rect 17402 13512 17408 13524
rect 17359 13484 17408 13512
rect 17359 13481 17371 13484
rect 17313 13475 17371 13481
rect 17402 13472 17408 13484
rect 17460 13472 17466 13524
rect 17586 13472 17592 13524
rect 17644 13512 17650 13524
rect 18141 13515 18199 13521
rect 18141 13512 18153 13515
rect 17644 13484 18153 13512
rect 17644 13472 17650 13484
rect 18141 13481 18153 13484
rect 18187 13512 18199 13515
rect 19978 13512 19984 13524
rect 18187 13484 19984 13512
rect 18187 13481 18199 13484
rect 18141 13475 18199 13481
rect 19978 13472 19984 13484
rect 20036 13512 20042 13524
rect 20257 13515 20315 13521
rect 20257 13512 20269 13515
rect 20036 13484 20269 13512
rect 20036 13472 20042 13484
rect 20257 13481 20269 13484
rect 20303 13481 20315 13515
rect 22002 13512 22008 13524
rect 20257 13475 20315 13481
rect 20640 13484 22008 13512
rect 17954 13444 17960 13456
rect 14332 13416 14780 13444
rect 15304 13416 17960 13444
rect 14332 13404 14338 13416
rect 6730 13336 6736 13388
rect 6788 13376 6794 13388
rect 6825 13379 6883 13385
rect 6825 13376 6837 13379
rect 6788 13348 6837 13376
rect 6788 13336 6794 13348
rect 6825 13345 6837 13348
rect 6871 13345 6883 13379
rect 6825 13339 6883 13345
rect 9122 13336 9128 13388
rect 9180 13376 9186 13388
rect 9401 13379 9459 13385
rect 9401 13376 9413 13379
rect 9180 13348 9413 13376
rect 9180 13336 9186 13348
rect 9401 13345 9413 13348
rect 9447 13345 9459 13379
rect 9401 13339 9459 13345
rect 9490 13336 9496 13388
rect 9548 13336 9554 13388
rect 9674 13336 9680 13388
rect 9732 13376 9738 13388
rect 10045 13379 10103 13385
rect 10045 13376 10057 13379
rect 9732 13348 10057 13376
rect 9732 13336 9738 13348
rect 10045 13345 10057 13348
rect 10091 13376 10103 13379
rect 10318 13376 10324 13388
rect 10091 13348 10324 13376
rect 10091 13345 10103 13348
rect 10045 13339 10103 13345
rect 10318 13336 10324 13348
rect 10376 13336 10382 13388
rect 11238 13336 11244 13388
rect 11296 13376 11302 13388
rect 11425 13379 11483 13385
rect 11425 13376 11437 13379
rect 11296 13348 11437 13376
rect 11296 13336 11302 13348
rect 11425 13345 11437 13348
rect 11471 13376 11483 13379
rect 12434 13376 12440 13388
rect 11471 13348 12440 13376
rect 11471 13345 11483 13348
rect 11425 13339 11483 13345
rect 12434 13336 12440 13348
rect 12492 13336 12498 13388
rect 13906 13336 13912 13388
rect 13964 13376 13970 13388
rect 15304 13376 15332 13416
rect 17954 13404 17960 13416
rect 18012 13404 18018 13456
rect 18868 13447 18926 13453
rect 18868 13413 18880 13447
rect 18914 13444 18926 13447
rect 19426 13444 19432 13456
rect 18914 13416 19432 13444
rect 18914 13413 18926 13416
rect 18868 13407 18926 13413
rect 19426 13404 19432 13416
rect 19484 13404 19490 13456
rect 13964 13348 15332 13376
rect 15556 13379 15614 13385
rect 13964 13336 13970 13348
rect 15556 13345 15568 13379
rect 15602 13376 15614 13379
rect 16390 13376 16396 13388
rect 15602 13348 16396 13376
rect 15602 13345 15614 13348
rect 15556 13339 15614 13345
rect 16390 13336 16396 13348
rect 16448 13336 16454 13388
rect 17126 13336 17132 13388
rect 17184 13376 17190 13388
rect 17497 13379 17555 13385
rect 17497 13376 17509 13379
rect 17184 13348 17509 13376
rect 17184 13336 17190 13348
rect 17497 13345 17509 13348
rect 17543 13345 17555 13379
rect 17497 13339 17555 13345
rect 18046 13336 18052 13388
rect 18104 13376 18110 13388
rect 18601 13379 18659 13385
rect 18601 13376 18613 13379
rect 18104 13348 18613 13376
rect 18104 13336 18110 13348
rect 18601 13345 18613 13348
rect 18647 13376 18659 13379
rect 19242 13376 19248 13388
rect 18647 13348 19248 13376
rect 18647 13345 18659 13348
rect 18601 13339 18659 13345
rect 19242 13336 19248 13348
rect 19300 13336 19306 13388
rect 19334 13336 19340 13388
rect 19392 13376 19398 13388
rect 20640 13376 20668 13484
rect 22002 13472 22008 13484
rect 22060 13512 22066 13524
rect 22097 13515 22155 13521
rect 22097 13512 22109 13515
rect 22060 13484 22109 13512
rect 22060 13472 22066 13484
rect 22097 13481 22109 13484
rect 22143 13481 22155 13515
rect 22097 13475 22155 13481
rect 22741 13515 22799 13521
rect 22741 13481 22753 13515
rect 22787 13512 22799 13515
rect 22922 13512 22928 13524
rect 22787 13484 22928 13512
rect 22787 13481 22799 13484
rect 22741 13475 22799 13481
rect 22922 13472 22928 13484
rect 22980 13472 22986 13524
rect 25409 13515 25467 13521
rect 25409 13481 25421 13515
rect 25455 13512 25467 13515
rect 25958 13512 25964 13524
rect 25455 13484 25964 13512
rect 25455 13481 25467 13484
rect 25409 13475 25467 13481
rect 25958 13472 25964 13484
rect 26016 13472 26022 13524
rect 20990 13404 20996 13456
rect 21048 13444 21054 13456
rect 21177 13447 21235 13453
rect 21177 13444 21189 13447
rect 21048 13416 21189 13444
rect 21048 13404 21054 13416
rect 21177 13413 21189 13416
rect 21223 13444 21235 13447
rect 21634 13444 21640 13456
rect 21223 13416 21640 13444
rect 21223 13413 21235 13416
rect 21177 13407 21235 13413
rect 21634 13404 21640 13416
rect 21692 13404 21698 13456
rect 22462 13404 22468 13456
rect 22520 13444 22526 13456
rect 23017 13447 23075 13453
rect 23017 13444 23029 13447
rect 22520 13416 23029 13444
rect 22520 13404 22526 13416
rect 23017 13413 23029 13416
rect 23063 13444 23075 13447
rect 23290 13444 23296 13456
rect 23063 13416 23296 13444
rect 23063 13413 23075 13416
rect 23017 13407 23075 13413
rect 23290 13404 23296 13416
rect 23348 13404 23354 13456
rect 25225 13447 25283 13453
rect 25225 13444 25237 13447
rect 23400 13416 25237 13444
rect 19392 13348 20668 13376
rect 19392 13336 19398 13348
rect 21542 13336 21548 13388
rect 21600 13376 21606 13388
rect 22005 13379 22063 13385
rect 22005 13376 22017 13379
rect 21600 13348 22017 13376
rect 21600 13336 21606 13348
rect 22005 13345 22017 13348
rect 22051 13345 22063 13379
rect 22005 13339 22063 13345
rect 23106 13336 23112 13388
rect 23164 13376 23170 13388
rect 23201 13379 23259 13385
rect 23201 13376 23213 13379
rect 23164 13348 23213 13376
rect 23164 13336 23170 13348
rect 23201 13345 23213 13348
rect 23247 13376 23259 13379
rect 23400 13376 23428 13416
rect 25225 13413 25237 13416
rect 25271 13444 25283 13447
rect 25869 13447 25927 13453
rect 25869 13444 25881 13447
rect 25271 13416 25881 13444
rect 25271 13413 25283 13416
rect 25225 13407 25283 13413
rect 25869 13413 25881 13416
rect 25915 13444 25927 13447
rect 26050 13444 26056 13456
rect 25915 13416 26056 13444
rect 25915 13413 25927 13416
rect 25869 13407 25927 13413
rect 26050 13404 26056 13416
rect 26108 13444 26114 13456
rect 26237 13447 26295 13453
rect 26237 13444 26249 13447
rect 26108 13416 26249 13444
rect 26108 13404 26114 13416
rect 26237 13413 26249 13416
rect 26283 13413 26295 13447
rect 26237 13407 26295 13413
rect 23474 13385 23480 13388
rect 23247 13348 23428 13376
rect 23247 13345 23259 13348
rect 23201 13339 23259 13345
rect 23468 13339 23480 13385
rect 23532 13376 23538 13388
rect 24026 13376 24032 13388
rect 23532 13348 24032 13376
rect 23474 13336 23480 13339
rect 23532 13336 23538 13348
rect 24026 13336 24032 13348
rect 24084 13336 24090 13388
rect 6512 13280 6684 13308
rect 7101 13311 7159 13317
rect 6512 13268 6518 13280
rect 7101 13277 7113 13311
rect 7147 13308 7159 13311
rect 7466 13308 7472 13320
rect 7147 13280 7472 13308
rect 7147 13277 7159 13280
rect 7101 13271 7159 13277
rect 4065 13243 4123 13249
rect 4065 13209 4077 13243
rect 4111 13240 4123 13243
rect 5350 13240 5356 13252
rect 4111 13212 5356 13240
rect 4111 13209 4123 13212
rect 4065 13203 4123 13209
rect 5350 13200 5356 13212
rect 5408 13200 5414 13252
rect 5994 13200 6000 13252
rect 6052 13240 6058 13252
rect 7116 13240 7144 13271
rect 7466 13268 7472 13280
rect 7524 13268 7530 13320
rect 8665 13311 8723 13317
rect 8665 13277 8677 13311
rect 8711 13277 8723 13311
rect 8665 13271 8723 13277
rect 6052 13212 7144 13240
rect 6052 13200 6058 13212
rect 3234 13172 3240 13184
rect 2363 13144 3240 13172
rect 2363 13141 2375 13144
rect 2317 13135 2375 13141
rect 3234 13132 3240 13144
rect 3292 13132 3298 13184
rect 3510 13132 3516 13184
rect 3568 13172 3574 13184
rect 3789 13175 3847 13181
rect 3789 13172 3801 13175
rect 3568 13144 3801 13172
rect 3568 13132 3574 13144
rect 3789 13141 3801 13144
rect 3835 13141 3847 13175
rect 3789 13135 3847 13141
rect 5534 13132 5540 13184
rect 5592 13172 5598 13184
rect 5813 13175 5871 13181
rect 5813 13172 5825 13175
rect 5592 13144 5825 13172
rect 5592 13132 5598 13144
rect 5813 13141 5825 13144
rect 5859 13141 5871 13175
rect 7466 13172 7472 13184
rect 7427 13144 7472 13172
rect 5813 13135 5871 13141
rect 7466 13132 7472 13144
rect 7524 13132 7530 13184
rect 7926 13172 7932 13184
rect 7887 13144 7932 13172
rect 7926 13132 7932 13144
rect 7984 13132 7990 13184
rect 8680 13172 8708 13271
rect 9508 13184 9536 13336
rect 10229 13311 10287 13317
rect 10229 13277 10241 13311
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 9950 13200 9956 13252
rect 10008 13240 10014 13252
rect 10244 13240 10272 13271
rect 13814 13268 13820 13320
rect 13872 13308 13878 13320
rect 14093 13311 14151 13317
rect 14093 13308 14105 13311
rect 13872 13280 14105 13308
rect 13872 13268 13878 13280
rect 14093 13277 14105 13280
rect 14139 13277 14151 13311
rect 14093 13271 14151 13277
rect 14277 13311 14335 13317
rect 14277 13277 14289 13311
rect 14323 13308 14335 13311
rect 14550 13308 14556 13320
rect 14323 13280 14556 13308
rect 14323 13277 14335 13280
rect 14277 13271 14335 13277
rect 14550 13268 14556 13280
rect 14608 13268 14614 13320
rect 14642 13268 14648 13320
rect 14700 13308 14706 13320
rect 15013 13311 15071 13317
rect 15013 13308 15025 13311
rect 14700 13280 15025 13308
rect 14700 13268 14706 13280
rect 15013 13277 15025 13280
rect 15059 13277 15071 13311
rect 15286 13308 15292 13320
rect 15247 13280 15292 13308
rect 15013 13271 15071 13277
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 18230 13308 18236 13320
rect 16408 13280 18236 13308
rect 10008 13212 10272 13240
rect 10008 13200 10014 13212
rect 10870 13200 10876 13252
rect 10928 13240 10934 13252
rect 12802 13240 12808 13252
rect 10928 13212 11376 13240
rect 12763 13212 12808 13240
rect 10928 13200 10934 13212
rect 8846 13172 8852 13184
rect 8680 13144 8852 13172
rect 8846 13132 8852 13144
rect 8904 13172 8910 13184
rect 9122 13172 9128 13184
rect 8904 13144 9128 13172
rect 8904 13132 8910 13144
rect 9122 13132 9128 13144
rect 9180 13132 9186 13184
rect 9490 13132 9496 13184
rect 9548 13132 9554 13184
rect 11238 13172 11244 13184
rect 11199 13144 11244 13172
rect 11238 13132 11244 13144
rect 11296 13132 11302 13184
rect 11348 13172 11376 13212
rect 12802 13200 12808 13212
rect 12860 13200 12866 13252
rect 13633 13243 13691 13249
rect 13633 13209 13645 13243
rect 13679 13240 13691 13243
rect 13722 13240 13728 13252
rect 13679 13212 13728 13240
rect 13679 13209 13691 13212
rect 13633 13203 13691 13209
rect 13722 13200 13728 13212
rect 13780 13200 13786 13252
rect 16408 13172 16436 13280
rect 18230 13268 18236 13280
rect 18288 13268 18294 13320
rect 22186 13268 22192 13320
rect 22244 13308 22250 13320
rect 22281 13311 22339 13317
rect 22281 13308 22293 13311
rect 22244 13280 22293 13308
rect 22244 13268 22250 13280
rect 22281 13277 22293 13280
rect 22327 13277 22339 13311
rect 22281 13271 22339 13277
rect 16669 13243 16727 13249
rect 16669 13209 16681 13243
rect 16715 13240 16727 13243
rect 16850 13240 16856 13252
rect 16715 13212 16856 13240
rect 16715 13209 16727 13212
rect 16669 13203 16727 13209
rect 16850 13200 16856 13212
rect 16908 13240 16914 13252
rect 17586 13240 17592 13252
rect 16908 13212 17592 13240
rect 16908 13200 16914 13212
rect 17586 13200 17592 13212
rect 17644 13200 17650 13252
rect 21358 13200 21364 13252
rect 21416 13240 21422 13252
rect 21637 13243 21695 13249
rect 21637 13240 21649 13243
rect 21416 13212 21649 13240
rect 21416 13200 21422 13212
rect 21637 13209 21649 13212
rect 21683 13209 21695 13243
rect 21637 13203 21695 13209
rect 11348 13144 16436 13172
rect 17218 13132 17224 13184
rect 17276 13172 17282 13184
rect 17681 13175 17739 13181
rect 17681 13172 17693 13175
rect 17276 13144 17693 13172
rect 17276 13132 17282 13144
rect 17681 13141 17693 13144
rect 17727 13141 17739 13175
rect 17681 13135 17739 13141
rect 18509 13175 18567 13181
rect 18509 13141 18521 13175
rect 18555 13172 18567 13175
rect 18874 13172 18880 13184
rect 18555 13144 18880 13172
rect 18555 13141 18567 13144
rect 18509 13135 18567 13141
rect 18874 13132 18880 13144
rect 18932 13132 18938 13184
rect 19981 13175 20039 13181
rect 19981 13141 19993 13175
rect 20027 13172 20039 13175
rect 20438 13172 20444 13184
rect 20027 13144 20444 13172
rect 20027 13141 20039 13144
rect 19981 13135 20039 13141
rect 20438 13132 20444 13144
rect 20496 13132 20502 13184
rect 20714 13172 20720 13184
rect 20675 13144 20720 13172
rect 20714 13132 20720 13144
rect 20772 13132 20778 13184
rect 22296 13172 22324 13271
rect 24762 13268 24768 13320
rect 24820 13308 24826 13320
rect 24857 13311 24915 13317
rect 24857 13308 24869 13311
rect 24820 13280 24869 13308
rect 24820 13268 24826 13280
rect 24857 13277 24869 13280
rect 24903 13277 24915 13311
rect 24857 13271 24915 13277
rect 22922 13172 22928 13184
rect 22296 13144 22928 13172
rect 22922 13132 22928 13144
rect 22980 13172 22986 13184
rect 24581 13175 24639 13181
rect 24581 13172 24593 13175
rect 22980 13144 24593 13172
rect 22980 13132 22986 13144
rect 24581 13141 24593 13144
rect 24627 13141 24639 13175
rect 24581 13135 24639 13141
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12968 1639 12971
rect 2958 12968 2964 12980
rect 1627 12940 2964 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 2958 12928 2964 12940
rect 3016 12928 3022 12980
rect 4709 12971 4767 12977
rect 4709 12937 4721 12971
rect 4755 12968 4767 12971
rect 5534 12968 5540 12980
rect 4755 12940 5540 12968
rect 4755 12937 4767 12940
rect 4709 12931 4767 12937
rect 5534 12928 5540 12940
rect 5592 12928 5598 12980
rect 5813 12971 5871 12977
rect 5813 12937 5825 12971
rect 5859 12968 5871 12971
rect 5994 12968 6000 12980
rect 5859 12940 6000 12968
rect 5859 12937 5871 12940
rect 5813 12931 5871 12937
rect 5994 12928 6000 12940
rect 6052 12928 6058 12980
rect 6181 12971 6239 12977
rect 6181 12937 6193 12971
rect 6227 12968 6239 12971
rect 6730 12968 6736 12980
rect 6227 12940 6736 12968
rect 6227 12937 6239 12940
rect 6181 12931 6239 12937
rect 6730 12928 6736 12940
rect 6788 12928 6794 12980
rect 9030 12968 9036 12980
rect 8991 12940 9036 12968
rect 9030 12928 9036 12940
rect 9088 12928 9094 12980
rect 9766 12928 9772 12980
rect 9824 12968 9830 12980
rect 10134 12968 10140 12980
rect 9824 12940 10140 12968
rect 9824 12928 9830 12940
rect 10134 12928 10140 12940
rect 10192 12928 10198 12980
rect 13354 12928 13360 12980
rect 13412 12968 13418 12980
rect 13630 12968 13636 12980
rect 13412 12940 13636 12968
rect 13412 12928 13418 12940
rect 13630 12928 13636 12940
rect 13688 12928 13694 12980
rect 14185 12971 14243 12977
rect 14185 12937 14197 12971
rect 14231 12968 14243 12971
rect 14550 12968 14556 12980
rect 14231 12940 14556 12968
rect 14231 12937 14243 12940
rect 14185 12931 14243 12937
rect 14550 12928 14556 12940
rect 14608 12928 14614 12980
rect 15746 12928 15752 12980
rect 15804 12968 15810 12980
rect 16025 12971 16083 12977
rect 16025 12968 16037 12971
rect 15804 12940 16037 12968
rect 15804 12928 15810 12940
rect 16025 12937 16037 12940
rect 16071 12937 16083 12971
rect 16025 12931 16083 12937
rect 16761 12971 16819 12977
rect 16761 12937 16773 12971
rect 16807 12968 16819 12971
rect 16942 12968 16948 12980
rect 16807 12940 16948 12968
rect 16807 12937 16819 12940
rect 16761 12931 16819 12937
rect 16942 12928 16948 12940
rect 17000 12928 17006 12980
rect 17126 12928 17132 12980
rect 17184 12968 17190 12980
rect 17497 12971 17555 12977
rect 17497 12968 17509 12971
rect 17184 12940 17509 12968
rect 17184 12928 17190 12940
rect 17497 12937 17509 12940
rect 17543 12937 17555 12971
rect 17497 12931 17555 12937
rect 17678 12928 17684 12980
rect 17736 12968 17742 12980
rect 18417 12971 18475 12977
rect 18417 12968 18429 12971
rect 17736 12940 18429 12968
rect 17736 12928 17742 12940
rect 18417 12937 18429 12940
rect 18463 12937 18475 12971
rect 19426 12968 19432 12980
rect 19387 12940 19432 12968
rect 18417 12931 18475 12937
rect 19426 12928 19432 12940
rect 19484 12928 19490 12980
rect 20254 12968 20260 12980
rect 20215 12940 20260 12968
rect 20254 12928 20260 12940
rect 20312 12928 20318 12980
rect 21174 12968 21180 12980
rect 21135 12940 21180 12968
rect 21174 12928 21180 12940
rect 21232 12928 21238 12980
rect 21910 12928 21916 12980
rect 21968 12968 21974 12980
rect 22189 12971 22247 12977
rect 22189 12968 22201 12971
rect 21968 12940 22201 12968
rect 21968 12928 21974 12940
rect 22189 12937 22201 12940
rect 22235 12937 22247 12971
rect 22189 12931 22247 12937
rect 22649 12971 22707 12977
rect 22649 12937 22661 12971
rect 22695 12968 22707 12971
rect 22922 12968 22928 12980
rect 22695 12940 22928 12968
rect 22695 12937 22707 12940
rect 22649 12931 22707 12937
rect 1118 12860 1124 12912
rect 1176 12900 1182 12912
rect 2685 12903 2743 12909
rect 1176 12872 1900 12900
rect 1176 12860 1182 12872
rect 1872 12832 1900 12872
rect 2685 12869 2697 12903
rect 2731 12900 2743 12903
rect 2774 12900 2780 12912
rect 2731 12872 2780 12900
rect 2731 12869 2743 12872
rect 2685 12863 2743 12869
rect 2774 12860 2780 12872
rect 2832 12860 2838 12912
rect 3145 12903 3203 12909
rect 3145 12869 3157 12903
rect 3191 12900 3203 12903
rect 4062 12900 4068 12912
rect 3191 12872 4068 12900
rect 3191 12869 3203 12872
rect 3145 12863 3203 12869
rect 4062 12860 4068 12872
rect 4120 12860 4126 12912
rect 6454 12900 6460 12912
rect 6415 12872 6460 12900
rect 6454 12860 6460 12872
rect 6512 12860 6518 12912
rect 8389 12903 8447 12909
rect 8389 12869 8401 12903
rect 8435 12900 8447 12903
rect 8573 12903 8631 12909
rect 8573 12900 8585 12903
rect 8435 12872 8585 12900
rect 8435 12869 8447 12872
rect 8389 12863 8447 12869
rect 8573 12869 8585 12872
rect 8619 12900 8631 12903
rect 9122 12900 9128 12912
rect 8619 12872 9128 12900
rect 8619 12869 8631 12872
rect 8573 12863 8631 12869
rect 9122 12860 9128 12872
rect 9180 12900 9186 12912
rect 9180 12872 9628 12900
rect 9180 12860 9186 12872
rect 2130 12832 2136 12844
rect 1872 12804 2136 12832
rect 2130 12792 2136 12804
rect 2188 12792 2194 12844
rect 3418 12792 3424 12844
rect 3476 12832 3482 12844
rect 3605 12835 3663 12841
rect 3605 12832 3617 12835
rect 3476 12804 3617 12832
rect 3476 12792 3482 12804
rect 3605 12801 3617 12804
rect 3651 12801 3663 12835
rect 3786 12832 3792 12844
rect 3699 12804 3792 12832
rect 3605 12795 3663 12801
rect 3786 12792 3792 12804
rect 3844 12832 3850 12844
rect 4617 12835 4675 12841
rect 3844 12804 4108 12832
rect 3844 12792 3850 12804
rect 1210 12724 1216 12776
rect 1268 12764 1274 12776
rect 1268 12736 2084 12764
rect 1268 12724 1274 12736
rect 2056 12705 2084 12736
rect 2590 12724 2596 12776
rect 2648 12764 2654 12776
rect 3510 12764 3516 12776
rect 2648 12736 3516 12764
rect 2648 12724 2654 12736
rect 3510 12724 3516 12736
rect 3568 12724 3574 12776
rect 2041 12699 2099 12705
rect 2041 12665 2053 12699
rect 2087 12696 2099 12699
rect 2087 12668 2636 12696
rect 2087 12665 2099 12668
rect 2041 12659 2099 12665
rect 1394 12588 1400 12640
rect 1452 12628 1458 12640
rect 1949 12631 2007 12637
rect 1949 12628 1961 12631
rect 1452 12600 1961 12628
rect 1452 12588 1458 12600
rect 1949 12597 1961 12600
rect 1995 12628 2007 12631
rect 2498 12628 2504 12640
rect 1995 12600 2504 12628
rect 1995 12597 2007 12600
rect 1949 12591 2007 12597
rect 2498 12588 2504 12600
rect 2556 12588 2562 12640
rect 2608 12628 2636 12668
rect 2774 12628 2780 12640
rect 2608 12600 2780 12628
rect 2774 12588 2780 12600
rect 2832 12588 2838 12640
rect 3053 12631 3111 12637
rect 3053 12597 3065 12631
rect 3099 12628 3111 12631
rect 3142 12628 3148 12640
rect 3099 12600 3148 12628
rect 3099 12597 3111 12600
rect 3053 12591 3111 12597
rect 3142 12588 3148 12600
rect 3200 12588 3206 12640
rect 4080 12628 4108 12804
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 5166 12832 5172 12844
rect 4663 12804 5172 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 5166 12792 5172 12804
rect 5224 12792 5230 12844
rect 5258 12792 5264 12844
rect 5316 12832 5322 12844
rect 5316 12804 5361 12832
rect 5316 12792 5322 12804
rect 6546 12792 6552 12844
rect 6604 12832 6610 12844
rect 6825 12835 6883 12841
rect 6825 12832 6837 12835
rect 6604 12804 6837 12832
rect 6604 12792 6610 12804
rect 6825 12801 6837 12804
rect 6871 12801 6883 12835
rect 6825 12795 6883 12801
rect 7926 12792 7932 12844
rect 7984 12832 7990 12844
rect 9600 12841 9628 12872
rect 10042 12860 10048 12912
rect 10100 12900 10106 12912
rect 10597 12903 10655 12909
rect 10597 12900 10609 12903
rect 10100 12872 10609 12900
rect 10100 12860 10106 12872
rect 10597 12869 10609 12872
rect 10643 12869 10655 12903
rect 10597 12863 10655 12869
rect 16206 12860 16212 12912
rect 16264 12900 16270 12912
rect 18233 12903 18291 12909
rect 18233 12900 18245 12903
rect 16264 12872 18245 12900
rect 16264 12860 16270 12872
rect 18233 12869 18245 12872
rect 18279 12869 18291 12903
rect 18233 12863 18291 12869
rect 19981 12903 20039 12909
rect 19981 12869 19993 12903
rect 20027 12900 20039 12903
rect 20162 12900 20168 12912
rect 20027 12872 20168 12900
rect 20027 12869 20039 12872
rect 19981 12863 20039 12869
rect 9493 12835 9551 12841
rect 9493 12832 9505 12835
rect 7984 12804 9505 12832
rect 7984 12792 7990 12804
rect 9493 12801 9505 12804
rect 9539 12801 9551 12835
rect 9493 12795 9551 12801
rect 9585 12835 9643 12841
rect 9585 12801 9597 12835
rect 9631 12832 9643 12835
rect 10137 12835 10195 12841
rect 9631 12804 9904 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 4706 12724 4712 12776
rect 4764 12764 4770 12776
rect 5074 12764 5080 12776
rect 4764 12736 5080 12764
rect 4764 12724 4770 12736
rect 5074 12724 5080 12736
rect 5132 12724 5138 12776
rect 8849 12767 8907 12773
rect 8849 12733 8861 12767
rect 8895 12764 8907 12767
rect 9122 12764 9128 12776
rect 8895 12736 9128 12764
rect 8895 12733 8907 12736
rect 8849 12727 8907 12733
rect 9122 12724 9128 12736
rect 9180 12764 9186 12776
rect 9398 12764 9404 12776
rect 9180 12736 9404 12764
rect 9180 12724 9186 12736
rect 9398 12724 9404 12736
rect 9456 12724 9462 12776
rect 9508 12764 9536 12795
rect 9674 12764 9680 12776
rect 9508 12736 9680 12764
rect 9674 12724 9680 12736
rect 9732 12724 9738 12776
rect 9876 12764 9904 12804
rect 10137 12801 10149 12835
rect 10183 12832 10195 12835
rect 10318 12832 10324 12844
rect 10183 12804 10324 12832
rect 10183 12801 10195 12804
rect 10137 12795 10195 12801
rect 10318 12792 10324 12804
rect 10376 12792 10382 12844
rect 10686 12792 10692 12844
rect 10744 12832 10750 12844
rect 11057 12835 11115 12841
rect 11057 12832 11069 12835
rect 10744 12804 11069 12832
rect 10744 12792 10750 12804
rect 11057 12801 11069 12804
rect 11103 12801 11115 12835
rect 11238 12832 11244 12844
rect 11151 12804 11244 12832
rect 11057 12795 11115 12801
rect 11238 12792 11244 12804
rect 11296 12832 11302 12844
rect 11698 12832 11704 12844
rect 11296 12804 11704 12832
rect 11296 12792 11302 12804
rect 11698 12792 11704 12804
rect 11756 12792 11762 12844
rect 12434 12832 12440 12844
rect 12395 12804 12440 12832
rect 12434 12792 12440 12804
rect 12492 12792 12498 12844
rect 16574 12792 16580 12844
rect 16632 12832 16638 12844
rect 16945 12835 17003 12841
rect 16945 12832 16957 12835
rect 16632 12804 16957 12832
rect 16632 12792 16638 12804
rect 16945 12801 16957 12804
rect 16991 12801 17003 12835
rect 16945 12795 17003 12801
rect 9876 12736 11275 12764
rect 4249 12699 4307 12705
rect 4249 12665 4261 12699
rect 4295 12696 4307 12699
rect 4522 12696 4528 12708
rect 4295 12668 4528 12696
rect 4295 12665 4307 12668
rect 4249 12659 4307 12665
rect 4522 12656 4528 12668
rect 4580 12696 4586 12708
rect 5258 12696 5264 12708
rect 4580 12668 5264 12696
rect 4580 12656 4586 12668
rect 5258 12656 5264 12668
rect 5316 12656 5322 12708
rect 5350 12656 5356 12708
rect 5408 12696 5414 12708
rect 7070 12699 7128 12705
rect 7070 12696 7082 12699
rect 5408 12668 7082 12696
rect 5408 12656 5414 12668
rect 7070 12665 7082 12668
rect 7116 12696 7128 12699
rect 7466 12696 7472 12708
rect 7116 12668 7472 12696
rect 7116 12665 7128 12668
rect 7070 12659 7128 12665
rect 7466 12656 7472 12668
rect 7524 12696 7530 12708
rect 8389 12699 8447 12705
rect 8389 12696 8401 12699
rect 7524 12668 8401 12696
rect 7524 12656 7530 12668
rect 8389 12665 8401 12668
rect 8435 12665 8447 12699
rect 9858 12696 9864 12708
rect 8389 12659 8447 12665
rect 8864 12668 9864 12696
rect 8864 12640 8892 12668
rect 9858 12656 9864 12668
rect 9916 12656 9922 12708
rect 10226 12656 10232 12708
rect 10284 12696 10290 12708
rect 11146 12696 11152 12708
rect 10284 12668 11152 12696
rect 10284 12656 10290 12668
rect 11146 12656 11152 12668
rect 11204 12656 11210 12708
rect 11247 12696 11275 12736
rect 11606 12724 11612 12776
rect 11664 12764 11670 12776
rect 11974 12764 11980 12776
rect 11664 12736 11980 12764
rect 11664 12724 11670 12736
rect 11974 12724 11980 12736
rect 12032 12724 12038 12776
rect 13814 12764 13820 12776
rect 12084 12736 13820 12764
rect 12084 12696 12112 12736
rect 13814 12724 13820 12736
rect 13872 12724 13878 12776
rect 14645 12767 14703 12773
rect 14645 12733 14657 12767
rect 14691 12764 14703 12767
rect 15286 12764 15292 12776
rect 14691 12736 15292 12764
rect 14691 12733 14703 12736
rect 14645 12727 14703 12733
rect 15286 12724 15292 12736
rect 15344 12724 15350 12776
rect 16390 12724 16396 12776
rect 16448 12724 16454 12776
rect 18248 12764 18276 12863
rect 18874 12832 18880 12844
rect 18835 12804 18880 12832
rect 18874 12792 18880 12804
rect 18932 12792 18938 12844
rect 19058 12832 19064 12844
rect 19019 12804 19064 12832
rect 19058 12792 19064 12804
rect 19116 12792 19122 12844
rect 20088 12773 20116 12872
rect 20162 12860 20168 12872
rect 20220 12860 20226 12912
rect 20717 12835 20775 12841
rect 20717 12801 20729 12835
rect 20763 12832 20775 12835
rect 21729 12835 21787 12841
rect 21729 12832 21741 12835
rect 20763 12804 21741 12832
rect 20763 12801 20775 12804
rect 20717 12795 20775 12801
rect 21729 12801 21741 12804
rect 21775 12832 21787 12835
rect 22664 12832 22692 12931
rect 22922 12928 22928 12940
rect 22980 12928 22986 12980
rect 23293 12971 23351 12977
rect 23293 12937 23305 12971
rect 23339 12968 23351 12971
rect 23474 12968 23480 12980
rect 23339 12940 23480 12968
rect 23339 12937 23351 12940
rect 23293 12931 23351 12937
rect 23474 12928 23480 12940
rect 23532 12968 23538 12980
rect 25041 12971 25099 12977
rect 25041 12968 25053 12971
rect 23532 12940 25053 12968
rect 23532 12928 23538 12940
rect 25041 12937 25053 12940
rect 25087 12937 25099 12971
rect 25314 12968 25320 12980
rect 25275 12940 25320 12968
rect 25041 12931 25099 12937
rect 25314 12928 25320 12940
rect 25372 12968 25378 12980
rect 25685 12971 25743 12977
rect 25685 12968 25697 12971
rect 25372 12940 25697 12968
rect 25372 12928 25378 12940
rect 25685 12937 25697 12940
rect 25731 12937 25743 12971
rect 26050 12968 26056 12980
rect 26011 12940 26056 12968
rect 25685 12931 25743 12937
rect 26050 12928 26056 12940
rect 26108 12968 26114 12980
rect 26421 12971 26479 12977
rect 26421 12968 26433 12971
rect 26108 12940 26433 12968
rect 26108 12928 26114 12940
rect 26421 12937 26433 12940
rect 26467 12937 26479 12971
rect 26421 12931 26479 12937
rect 21775 12804 22692 12832
rect 21775 12801 21787 12804
rect 21729 12795 21787 12801
rect 23014 12792 23020 12844
rect 23072 12832 23078 12844
rect 23661 12835 23719 12841
rect 23661 12832 23673 12835
rect 23072 12804 23673 12832
rect 23072 12792 23078 12804
rect 23661 12801 23673 12804
rect 23707 12801 23719 12835
rect 23661 12795 23719 12801
rect 18785 12767 18843 12773
rect 18785 12764 18797 12767
rect 18248 12736 18797 12764
rect 18785 12733 18797 12736
rect 18831 12733 18843 12767
rect 18785 12727 18843 12733
rect 20073 12767 20131 12773
rect 20073 12733 20085 12767
rect 20119 12733 20131 12767
rect 21634 12764 21640 12776
rect 21595 12736 21640 12764
rect 20073 12727 20131 12733
rect 21634 12724 21640 12736
rect 21692 12764 21698 12776
rect 23106 12764 23112 12776
rect 21692 12736 23112 12764
rect 21692 12724 21698 12736
rect 23106 12724 23112 12736
rect 23164 12724 23170 12776
rect 11247 12668 12112 12696
rect 12253 12699 12311 12705
rect 12253 12665 12265 12699
rect 12299 12696 12311 12699
rect 12704 12699 12762 12705
rect 12704 12696 12716 12699
rect 12299 12668 12716 12696
rect 12299 12665 12311 12668
rect 12253 12659 12311 12665
rect 12704 12665 12716 12668
rect 12750 12696 12762 12699
rect 12802 12696 12808 12708
rect 12750 12668 12808 12696
rect 12750 12665 12762 12668
rect 12704 12659 12762 12665
rect 12802 12656 12808 12668
rect 12860 12656 12866 12708
rect 14918 12705 14924 12708
rect 14553 12699 14611 12705
rect 14553 12696 14565 12699
rect 13832 12668 14565 12696
rect 6546 12628 6552 12640
rect 4080 12600 6552 12628
rect 6546 12588 6552 12600
rect 6604 12628 6610 12640
rect 8018 12628 8024 12640
rect 6604 12600 8024 12628
rect 6604 12588 6610 12600
rect 8018 12588 8024 12600
rect 8076 12628 8082 12640
rect 8205 12631 8263 12637
rect 8205 12628 8217 12631
rect 8076 12600 8217 12628
rect 8076 12588 8082 12600
rect 8205 12597 8217 12600
rect 8251 12597 8263 12631
rect 8205 12591 8263 12597
rect 8846 12588 8852 12640
rect 8904 12588 8910 12640
rect 10505 12631 10563 12637
rect 10505 12597 10517 12631
rect 10551 12628 10563 12631
rect 10870 12628 10876 12640
rect 10551 12600 10876 12628
rect 10551 12597 10563 12600
rect 10505 12591 10563 12597
rect 10870 12588 10876 12600
rect 10928 12628 10934 12640
rect 10965 12631 11023 12637
rect 10965 12628 10977 12631
rect 10928 12600 10977 12628
rect 10928 12588 10934 12600
rect 10965 12597 10977 12600
rect 11011 12597 11023 12631
rect 10965 12591 11023 12597
rect 11514 12588 11520 12640
rect 11572 12628 11578 12640
rect 11701 12631 11759 12637
rect 11701 12628 11713 12631
rect 11572 12600 11713 12628
rect 11572 12588 11578 12600
rect 11701 12597 11713 12600
rect 11747 12628 11759 12631
rect 11974 12628 11980 12640
rect 11747 12600 11980 12628
rect 11747 12597 11759 12600
rect 11701 12591 11759 12597
rect 11974 12588 11980 12600
rect 12032 12588 12038 12640
rect 13832 12637 13860 12668
rect 14553 12665 14565 12668
rect 14599 12696 14611 12699
rect 14912 12696 14924 12705
rect 14599 12668 14924 12696
rect 14599 12665 14611 12668
rect 14553 12659 14611 12665
rect 14912 12659 14924 12668
rect 14918 12656 14924 12659
rect 14976 12656 14982 12708
rect 16301 12699 16359 12705
rect 16301 12665 16313 12699
rect 16347 12696 16359 12699
rect 16408 12696 16436 12724
rect 16574 12696 16580 12708
rect 16347 12668 16580 12696
rect 16347 12665 16359 12668
rect 16301 12659 16359 12665
rect 16574 12656 16580 12668
rect 16632 12656 16638 12708
rect 16666 12656 16672 12708
rect 16724 12696 16730 12708
rect 16942 12696 16948 12708
rect 16724 12668 16948 12696
rect 16724 12656 16730 12668
rect 16942 12656 16948 12668
rect 17000 12656 17006 12708
rect 17678 12656 17684 12708
rect 17736 12696 17742 12708
rect 18414 12696 18420 12708
rect 17736 12668 18420 12696
rect 17736 12656 17742 12668
rect 18414 12656 18420 12668
rect 18472 12656 18478 12708
rect 20990 12696 20996 12708
rect 20951 12668 20996 12696
rect 20990 12656 20996 12668
rect 21048 12696 21054 12708
rect 21545 12699 21603 12705
rect 21545 12696 21557 12699
rect 21048 12668 21557 12696
rect 21048 12656 21054 12668
rect 21545 12665 21557 12668
rect 21591 12665 21603 12699
rect 21545 12659 21603 12665
rect 22646 12656 22652 12708
rect 22704 12696 22710 12708
rect 23014 12696 23020 12708
rect 22704 12668 23020 12696
rect 22704 12656 22710 12668
rect 23014 12656 23020 12668
rect 23072 12656 23078 12708
rect 23290 12656 23296 12708
rect 23348 12696 23354 12708
rect 23566 12696 23572 12708
rect 23348 12668 23572 12696
rect 23348 12656 23354 12668
rect 23566 12656 23572 12668
rect 23624 12656 23630 12708
rect 23842 12656 23848 12708
rect 23900 12705 23906 12708
rect 23900 12699 23964 12705
rect 23900 12665 23918 12699
rect 23952 12696 23964 12699
rect 23952 12668 24532 12696
rect 23952 12665 23964 12668
rect 23900 12659 23964 12665
rect 23900 12656 23906 12659
rect 13817 12631 13875 12637
rect 13817 12597 13829 12631
rect 13863 12597 13875 12631
rect 13817 12591 13875 12597
rect 14458 12588 14464 12640
rect 14516 12628 14522 12640
rect 16206 12628 16212 12640
rect 14516 12600 16212 12628
rect 14516 12588 14522 12600
rect 16206 12588 16212 12600
rect 16264 12588 16270 12640
rect 16390 12588 16396 12640
rect 16448 12628 16454 12640
rect 17310 12628 17316 12640
rect 16448 12600 17316 12628
rect 16448 12588 16454 12600
rect 17310 12588 17316 12600
rect 17368 12588 17374 12640
rect 22462 12588 22468 12640
rect 22520 12628 22526 12640
rect 22830 12628 22836 12640
rect 22520 12600 22836 12628
rect 22520 12588 22526 12600
rect 22830 12588 22836 12600
rect 22888 12588 22894 12640
rect 24504 12628 24532 12668
rect 24762 12628 24768 12640
rect 24504 12600 24768 12628
rect 24762 12588 24768 12600
rect 24820 12588 24826 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1118 12384 1124 12436
rect 1176 12424 1182 12436
rect 1673 12427 1731 12433
rect 1673 12424 1685 12427
rect 1176 12396 1685 12424
rect 1176 12384 1182 12396
rect 1673 12393 1685 12396
rect 1719 12424 1731 12427
rect 3145 12427 3203 12433
rect 3145 12424 3157 12427
rect 1719 12396 3157 12424
rect 1719 12393 1731 12396
rect 1673 12387 1731 12393
rect 3145 12393 3157 12396
rect 3191 12393 3203 12427
rect 3145 12387 3203 12393
rect 3513 12427 3571 12433
rect 3513 12393 3525 12427
rect 3559 12424 3571 12427
rect 3786 12424 3792 12436
rect 3559 12396 3792 12424
rect 3559 12393 3571 12396
rect 3513 12387 3571 12393
rect 3786 12384 3792 12396
rect 3844 12384 3850 12436
rect 3881 12427 3939 12433
rect 3881 12393 3893 12427
rect 3927 12424 3939 12427
rect 3970 12424 3976 12436
rect 3927 12396 3976 12424
rect 3927 12393 3939 12396
rect 3881 12387 3939 12393
rect 3970 12384 3976 12396
rect 4028 12384 4034 12436
rect 4154 12384 4160 12436
rect 4212 12424 4218 12436
rect 4249 12427 4307 12433
rect 4249 12424 4261 12427
rect 4212 12396 4261 12424
rect 4212 12384 4218 12396
rect 4249 12393 4261 12396
rect 4295 12393 4307 12427
rect 4249 12387 4307 12393
rect 4338 12384 4344 12436
rect 4396 12424 4402 12436
rect 4985 12427 5043 12433
rect 4985 12424 4997 12427
rect 4396 12396 4997 12424
rect 4396 12384 4402 12396
rect 4985 12393 4997 12396
rect 5031 12393 5043 12427
rect 4985 12387 5043 12393
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 6365 12427 6423 12433
rect 6365 12424 6377 12427
rect 5592 12396 6377 12424
rect 5592 12384 5598 12396
rect 6365 12393 6377 12396
rect 6411 12393 6423 12427
rect 8294 12424 8300 12436
rect 8255 12396 8300 12424
rect 6365 12387 6423 12393
rect 8294 12384 8300 12396
rect 8352 12384 8358 12436
rect 8662 12424 8668 12436
rect 8623 12396 8668 12424
rect 8662 12384 8668 12396
rect 8720 12384 8726 12436
rect 9674 12424 9680 12436
rect 9635 12396 9680 12424
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 9858 12384 9864 12436
rect 9916 12424 9922 12436
rect 10137 12427 10195 12433
rect 10137 12424 10149 12427
rect 9916 12396 10149 12424
rect 9916 12384 9922 12396
rect 10137 12393 10149 12396
rect 10183 12393 10195 12427
rect 10137 12387 10195 12393
rect 10778 12384 10784 12436
rect 10836 12424 10842 12436
rect 12250 12424 12256 12436
rect 10836 12396 12256 12424
rect 10836 12384 10842 12396
rect 12250 12384 12256 12396
rect 12308 12424 12314 12436
rect 14090 12424 14096 12436
rect 12308 12396 14096 12424
rect 12308 12384 12314 12396
rect 14090 12384 14096 12396
rect 14148 12384 14154 12436
rect 15838 12384 15844 12436
rect 15896 12424 15902 12436
rect 16206 12424 16212 12436
rect 15896 12396 16212 12424
rect 15896 12384 15902 12396
rect 16206 12384 16212 12396
rect 16264 12384 16270 12436
rect 16574 12384 16580 12436
rect 16632 12424 16638 12436
rect 16669 12427 16727 12433
rect 16669 12424 16681 12427
rect 16632 12396 16681 12424
rect 16632 12384 16638 12396
rect 16669 12393 16681 12396
rect 16715 12393 16727 12427
rect 16942 12424 16948 12436
rect 16903 12396 16948 12424
rect 16669 12387 16727 12393
rect 16942 12384 16948 12396
rect 17000 12384 17006 12436
rect 17310 12424 17316 12436
rect 17271 12396 17316 12424
rect 17310 12384 17316 12396
rect 17368 12384 17374 12436
rect 18509 12427 18567 12433
rect 18509 12393 18521 12427
rect 18555 12424 18567 12427
rect 19058 12424 19064 12436
rect 18555 12396 19064 12424
rect 18555 12393 18567 12396
rect 18509 12387 18567 12393
rect 19058 12384 19064 12396
rect 19116 12384 19122 12436
rect 19150 12384 19156 12436
rect 19208 12424 19214 12436
rect 20990 12424 20996 12436
rect 19208 12396 20996 12424
rect 19208 12384 19214 12396
rect 20990 12384 20996 12396
rect 21048 12384 21054 12436
rect 22278 12384 22284 12436
rect 22336 12424 22342 12436
rect 22462 12424 22468 12436
rect 22336 12396 22468 12424
rect 22336 12384 22342 12396
rect 22462 12384 22468 12396
rect 22520 12384 22526 12436
rect 23385 12427 23443 12433
rect 23385 12393 23397 12427
rect 23431 12424 23443 12427
rect 23753 12427 23811 12433
rect 23753 12424 23765 12427
rect 23431 12396 23765 12424
rect 23431 12393 23443 12396
rect 23385 12387 23443 12393
rect 23753 12393 23765 12396
rect 23799 12424 23811 12427
rect 23842 12424 23848 12436
rect 23799 12396 23848 12424
rect 23799 12393 23811 12396
rect 23753 12387 23811 12393
rect 23842 12384 23848 12396
rect 23900 12384 23906 12436
rect 24118 12424 24124 12436
rect 24079 12396 24124 12424
rect 24118 12384 24124 12396
rect 24176 12384 24182 12436
rect 25317 12427 25375 12433
rect 25317 12393 25329 12427
rect 25363 12424 25375 12427
rect 25406 12424 25412 12436
rect 25363 12396 25412 12424
rect 25363 12393 25375 12396
rect 25317 12387 25375 12393
rect 25406 12384 25412 12396
rect 25464 12384 25470 12436
rect 26050 12424 26056 12436
rect 26011 12396 26056 12424
rect 26050 12384 26056 12396
rect 26108 12384 26114 12436
rect 845 12359 903 12365
rect 845 12325 857 12359
rect 891 12356 903 12359
rect 1394 12356 1400 12368
rect 891 12328 1400 12356
rect 891 12325 903 12328
rect 845 12319 903 12325
rect 1394 12316 1400 12328
rect 1452 12316 1458 12368
rect 2314 12356 2320 12368
rect 1780 12328 2320 12356
rect 1780 12297 1808 12328
rect 2314 12316 2320 12328
rect 2372 12316 2378 12368
rect 4706 12356 4712 12368
rect 4667 12328 4712 12356
rect 4706 12316 4712 12328
rect 4764 12316 4770 12368
rect 6546 12316 6552 12368
rect 6604 12356 6610 12368
rect 6794 12359 6852 12365
rect 6794 12356 6806 12359
rect 6604 12328 6806 12356
rect 6604 12316 6610 12328
rect 6794 12325 6806 12328
rect 6840 12325 6852 12359
rect 6794 12319 6852 12325
rect 9493 12359 9551 12365
rect 9493 12325 9505 12359
rect 9539 12356 9551 12359
rect 9582 12356 9588 12368
rect 9539 12328 9588 12356
rect 9539 12325 9551 12328
rect 9493 12319 9551 12325
rect 9582 12316 9588 12328
rect 9640 12316 9646 12368
rect 12621 12359 12679 12365
rect 12621 12325 12633 12359
rect 12667 12356 12679 12359
rect 12713 12359 12771 12365
rect 12713 12356 12725 12359
rect 12667 12328 12725 12356
rect 12667 12325 12679 12328
rect 12621 12319 12679 12325
rect 12713 12325 12725 12328
rect 12759 12325 12771 12359
rect 12713 12319 12771 12325
rect 13998 12316 14004 12368
rect 14056 12356 14062 12368
rect 15556 12359 15614 12365
rect 14056 12328 15516 12356
rect 14056 12316 14062 12328
rect 1765 12291 1823 12297
rect 1765 12257 1777 12291
rect 1811 12257 1823 12291
rect 1765 12251 1823 12257
rect 1854 12248 1860 12300
rect 1912 12288 1918 12300
rect 2021 12291 2079 12297
rect 2021 12288 2033 12291
rect 1912 12260 2033 12288
rect 1912 12248 1918 12260
rect 2021 12257 2033 12260
rect 2067 12257 2079 12291
rect 2021 12251 2079 12257
rect 4154 12248 4160 12300
rect 4212 12288 4218 12300
rect 5353 12291 5411 12297
rect 5353 12288 5365 12291
rect 4212 12260 5365 12288
rect 4212 12248 4218 12260
rect 5353 12257 5365 12260
rect 5399 12288 5411 12291
rect 6178 12288 6184 12300
rect 5399 12260 6184 12288
rect 5399 12257 5411 12260
rect 5353 12251 5411 12257
rect 6178 12248 6184 12260
rect 6236 12248 6242 12300
rect 10045 12291 10103 12297
rect 10045 12257 10057 12291
rect 10091 12288 10103 12291
rect 10318 12288 10324 12300
rect 10091 12260 10324 12288
rect 10091 12257 10103 12260
rect 10045 12251 10103 12257
rect 10318 12248 10324 12260
rect 10376 12248 10382 12300
rect 11514 12288 11520 12300
rect 11475 12260 11520 12288
rect 11514 12248 11520 12260
rect 11572 12248 11578 12300
rect 15286 12288 15292 12300
rect 15247 12260 15292 12288
rect 15286 12248 15292 12260
rect 15344 12248 15350 12300
rect 15488 12288 15516 12328
rect 15556 12325 15568 12359
rect 15602 12356 15614 12359
rect 15746 12356 15752 12368
rect 15602 12328 15752 12356
rect 15602 12325 15614 12328
rect 15556 12319 15614 12325
rect 15746 12316 15752 12328
rect 15804 12316 15810 12368
rect 17034 12316 17040 12368
rect 17092 12356 17098 12368
rect 20806 12356 20812 12368
rect 17092 12328 20812 12356
rect 17092 12316 17098 12328
rect 20806 12316 20812 12328
rect 20864 12316 20870 12368
rect 21910 12316 21916 12368
rect 21968 12356 21974 12368
rect 22646 12356 22652 12368
rect 21968 12328 22652 12356
rect 21968 12316 21974 12328
rect 22646 12316 22652 12328
rect 22704 12316 22710 12368
rect 24673 12359 24731 12365
rect 24673 12325 24685 12359
rect 24719 12356 24731 12359
rect 24946 12356 24952 12368
rect 24719 12328 24952 12356
rect 24719 12325 24731 12328
rect 24673 12319 24731 12325
rect 24946 12316 24952 12328
rect 25004 12316 25010 12368
rect 17494 12288 17500 12300
rect 15488 12260 17500 12288
rect 17494 12248 17500 12260
rect 17552 12248 17558 12300
rect 18969 12291 19027 12297
rect 18969 12257 18981 12291
rect 19015 12288 19027 12291
rect 19429 12291 19487 12297
rect 19429 12288 19441 12291
rect 19015 12260 19441 12288
rect 19015 12257 19027 12260
rect 18969 12251 19027 12257
rect 19429 12257 19441 12260
rect 19475 12257 19487 12291
rect 19429 12251 19487 12257
rect 20717 12291 20775 12297
rect 20717 12257 20729 12291
rect 20763 12288 20775 12291
rect 20898 12288 20904 12300
rect 20763 12260 20904 12288
rect 20763 12257 20775 12260
rect 20717 12251 20775 12257
rect 20898 12248 20904 12260
rect 20956 12248 20962 12300
rect 22272 12291 22330 12297
rect 22272 12257 22284 12291
rect 22318 12288 22330 12291
rect 23014 12288 23020 12300
rect 22318 12260 23020 12288
rect 22318 12257 22330 12260
rect 22272 12251 22330 12257
rect 23014 12248 23020 12260
rect 23072 12248 23078 12300
rect 23382 12248 23388 12300
rect 23440 12288 23446 12300
rect 23842 12288 23848 12300
rect 23440 12260 23848 12288
rect 23440 12248 23446 12260
rect 23842 12248 23848 12260
rect 23900 12248 23906 12300
rect 24581 12291 24639 12297
rect 24581 12257 24593 12291
rect 24627 12288 24639 12291
rect 25222 12288 25228 12300
rect 24627 12260 25228 12288
rect 24627 12257 24639 12260
rect 24581 12251 24639 12257
rect 25222 12248 25228 12260
rect 25280 12248 25286 12300
rect 5442 12220 5448 12232
rect 5403 12192 5448 12220
rect 5442 12180 5448 12192
rect 5500 12180 5506 12232
rect 5537 12223 5595 12229
rect 5537 12189 5549 12223
rect 5583 12189 5595 12223
rect 5537 12183 5595 12189
rect 5074 12112 5080 12164
rect 5132 12152 5138 12164
rect 5552 12152 5580 12183
rect 6454 12180 6460 12232
rect 6512 12220 6518 12232
rect 6549 12223 6607 12229
rect 6549 12220 6561 12223
rect 6512 12192 6561 12220
rect 6512 12180 6518 12192
rect 6549 12189 6561 12192
rect 6595 12189 6607 12223
rect 6549 12183 6607 12189
rect 9950 12180 9956 12232
rect 10008 12220 10014 12232
rect 10229 12223 10287 12229
rect 10229 12220 10241 12223
rect 10008 12192 10241 12220
rect 10008 12180 10014 12192
rect 10229 12189 10241 12192
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 10502 12180 10508 12232
rect 10560 12220 10566 12232
rect 10778 12220 10784 12232
rect 10560 12192 10784 12220
rect 10560 12180 10566 12192
rect 10778 12180 10784 12192
rect 10836 12180 10842 12232
rect 10962 12180 10968 12232
rect 11020 12220 11026 12232
rect 11330 12220 11336 12232
rect 11020 12192 11336 12220
rect 11020 12180 11026 12192
rect 11330 12180 11336 12192
rect 11388 12220 11394 12232
rect 11609 12223 11667 12229
rect 11609 12220 11621 12223
rect 11388 12192 11621 12220
rect 11388 12180 11394 12192
rect 11609 12189 11621 12192
rect 11655 12189 11667 12223
rect 11609 12183 11667 12189
rect 11698 12180 11704 12232
rect 11756 12220 11762 12232
rect 14458 12220 14464 12232
rect 11756 12192 11849 12220
rect 14419 12192 14464 12220
rect 11756 12180 11762 12192
rect 14458 12180 14464 12192
rect 14516 12180 14522 12232
rect 16574 12180 16580 12232
rect 16632 12220 16638 12232
rect 17586 12220 17592 12232
rect 16632 12192 17592 12220
rect 16632 12180 16638 12192
rect 17586 12180 17592 12192
rect 17644 12180 17650 12232
rect 17770 12180 17776 12232
rect 17828 12220 17834 12232
rect 19061 12223 19119 12229
rect 19061 12220 19073 12223
rect 17828 12192 19073 12220
rect 17828 12180 17834 12192
rect 19061 12189 19073 12192
rect 19107 12189 19119 12223
rect 19061 12183 19119 12189
rect 19245 12223 19303 12229
rect 19245 12189 19257 12223
rect 19291 12220 19303 12223
rect 19334 12220 19340 12232
rect 19291 12192 19340 12220
rect 19291 12189 19303 12192
rect 19245 12183 19303 12189
rect 19334 12180 19340 12192
rect 19392 12180 19398 12232
rect 21910 12180 21916 12232
rect 21968 12220 21974 12232
rect 22005 12223 22063 12229
rect 22005 12220 22017 12223
rect 21968 12192 22017 12220
rect 21968 12180 21974 12192
rect 22005 12189 22017 12192
rect 22051 12189 22063 12223
rect 22005 12183 22063 12189
rect 24765 12223 24823 12229
rect 24765 12189 24777 12223
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 5132 12124 5580 12152
rect 5132 12112 5138 12124
rect 9674 12112 9680 12164
rect 9732 12152 9738 12164
rect 10134 12152 10140 12164
rect 9732 12124 10140 12152
rect 9732 12112 9738 12124
rect 10134 12112 10140 12124
rect 10192 12112 10198 12164
rect 11716 12152 11744 12180
rect 10704 12124 11744 12152
rect 10704 12096 10732 12124
rect 12250 12112 12256 12164
rect 12308 12152 12314 12164
rect 12621 12155 12679 12161
rect 12621 12152 12633 12155
rect 12308 12124 12633 12152
rect 12308 12112 12314 12124
rect 12621 12121 12633 12124
rect 12667 12121 12679 12155
rect 12621 12115 12679 12121
rect 18601 12155 18659 12161
rect 18601 12121 18613 12155
rect 18647 12152 18659 12155
rect 20254 12152 20260 12164
rect 18647 12124 20260 12152
rect 18647 12121 18659 12124
rect 18601 12115 18659 12121
rect 20254 12112 20260 12124
rect 20312 12112 20318 12164
rect 21082 12152 21088 12164
rect 21043 12124 21088 12152
rect 21082 12112 21088 12124
rect 21140 12112 21146 12164
rect 24780 12152 24808 12183
rect 23860 12124 24808 12152
rect 6086 12084 6092 12096
rect 6047 12056 6092 12084
rect 6086 12044 6092 12056
rect 6144 12044 6150 12096
rect 7926 12084 7932 12096
rect 7887 12056 7932 12084
rect 7926 12044 7932 12056
rect 7984 12044 7990 12096
rect 9125 12087 9183 12093
rect 9125 12053 9137 12087
rect 9171 12084 9183 12087
rect 9398 12084 9404 12096
rect 9171 12056 9404 12084
rect 9171 12053 9183 12056
rect 9125 12047 9183 12053
rect 9398 12044 9404 12056
rect 9456 12084 9462 12096
rect 9950 12084 9956 12096
rect 9456 12056 9956 12084
rect 9456 12044 9462 12056
rect 9950 12044 9956 12056
rect 10008 12044 10014 12096
rect 10686 12084 10692 12096
rect 10647 12056 10692 12084
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 10778 12044 10784 12096
rect 10836 12084 10842 12096
rect 11149 12087 11207 12093
rect 11149 12084 11161 12087
rect 10836 12056 11161 12084
rect 10836 12044 10842 12056
rect 11149 12053 11161 12056
rect 11195 12053 11207 12087
rect 12526 12084 12532 12096
rect 12487 12056 12532 12084
rect 11149 12047 11207 12053
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 14921 12087 14979 12093
rect 14921 12053 14933 12087
rect 14967 12084 14979 12087
rect 15286 12084 15292 12096
rect 14967 12056 15292 12084
rect 14967 12053 14979 12056
rect 14921 12047 14979 12053
rect 15286 12044 15292 12056
rect 15344 12084 15350 12096
rect 16390 12084 16396 12096
rect 15344 12056 16396 12084
rect 15344 12044 15350 12056
rect 16390 12044 16396 12056
rect 16448 12044 16454 12096
rect 17586 12044 17592 12096
rect 17644 12084 17650 12096
rect 17681 12087 17739 12093
rect 17681 12084 17693 12087
rect 17644 12056 17693 12084
rect 17644 12044 17650 12056
rect 17681 12053 17693 12056
rect 17727 12053 17739 12087
rect 17681 12047 17739 12053
rect 17954 12044 17960 12096
rect 18012 12084 18018 12096
rect 18049 12087 18107 12093
rect 18049 12084 18061 12087
rect 18012 12056 18061 12084
rect 18012 12044 18018 12056
rect 18049 12053 18061 12056
rect 18095 12053 18107 12087
rect 18049 12047 18107 12053
rect 19429 12087 19487 12093
rect 19429 12053 19441 12087
rect 19475 12084 19487 12087
rect 19705 12087 19763 12093
rect 19705 12084 19717 12087
rect 19475 12056 19717 12084
rect 19475 12053 19487 12056
rect 19429 12047 19487 12053
rect 19705 12053 19717 12056
rect 19751 12084 19763 12087
rect 19978 12084 19984 12096
rect 19751 12056 19984 12084
rect 19751 12053 19763 12056
rect 19705 12047 19763 12053
rect 19978 12044 19984 12056
rect 20036 12044 20042 12096
rect 21634 12084 21640 12096
rect 21595 12056 21640 12084
rect 21634 12044 21640 12056
rect 21692 12044 21698 12096
rect 22002 12044 22008 12096
rect 22060 12084 22066 12096
rect 23860 12084 23888 12124
rect 24688 12096 24716 12124
rect 22060 12056 23888 12084
rect 22060 12044 22066 12056
rect 23934 12044 23940 12096
rect 23992 12084 23998 12096
rect 24213 12087 24271 12093
rect 24213 12084 24225 12087
rect 23992 12056 24225 12084
rect 23992 12044 23998 12056
rect 24213 12053 24225 12056
rect 24259 12053 24271 12087
rect 24213 12047 24271 12053
rect 24670 12044 24676 12096
rect 24728 12044 24734 12096
rect 25590 12084 25596 12096
rect 25551 12056 25596 12084
rect 25590 12044 25596 12056
rect 25648 12044 25654 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2314 11880 2320 11892
rect 2148 11852 2320 11880
rect 2148 11753 2176 11852
rect 2314 11840 2320 11852
rect 2372 11840 2378 11892
rect 2498 11840 2504 11892
rect 2556 11880 2562 11892
rect 3789 11883 3847 11889
rect 3789 11880 3801 11883
rect 2556 11852 3801 11880
rect 2556 11840 2562 11852
rect 3789 11849 3801 11852
rect 3835 11849 3847 11883
rect 3789 11843 3847 11849
rect 4341 11883 4399 11889
rect 4341 11849 4353 11883
rect 4387 11880 4399 11883
rect 5442 11880 5448 11892
rect 4387 11852 5448 11880
rect 4387 11849 4399 11852
rect 4341 11843 4399 11849
rect 5442 11840 5448 11852
rect 5500 11840 5506 11892
rect 6178 11880 6184 11892
rect 6139 11852 6184 11880
rect 6178 11840 6184 11852
rect 6236 11840 6242 11892
rect 6546 11880 6552 11892
rect 6507 11852 6552 11880
rect 6546 11840 6552 11852
rect 6604 11840 6610 11892
rect 7558 11880 7564 11892
rect 7519 11852 7564 11880
rect 7558 11840 7564 11852
rect 7616 11840 7622 11892
rect 9769 11883 9827 11889
rect 9769 11849 9781 11883
rect 9815 11880 9827 11883
rect 9858 11880 9864 11892
rect 9815 11852 9864 11880
rect 9815 11849 9827 11852
rect 9769 11843 9827 11849
rect 9858 11840 9864 11852
rect 9916 11840 9922 11892
rect 10226 11880 10232 11892
rect 10187 11852 10232 11880
rect 10226 11840 10232 11852
rect 10284 11840 10290 11892
rect 10594 11840 10600 11892
rect 10652 11880 10658 11892
rect 11238 11880 11244 11892
rect 10652 11852 11244 11880
rect 10652 11840 10658 11852
rect 11238 11840 11244 11852
rect 11296 11840 11302 11892
rect 13078 11840 13084 11892
rect 13136 11880 13142 11892
rect 13538 11880 13544 11892
rect 13136 11852 13544 11880
rect 13136 11840 13142 11852
rect 13538 11840 13544 11852
rect 13596 11840 13602 11892
rect 13722 11840 13728 11892
rect 13780 11880 13786 11892
rect 14645 11883 14703 11889
rect 14645 11880 14657 11883
rect 13780 11852 14657 11880
rect 13780 11840 13786 11852
rect 14645 11849 14657 11852
rect 14691 11849 14703 11883
rect 16390 11880 16396 11892
rect 16351 11852 16396 11880
rect 14645 11843 14703 11849
rect 16390 11840 16396 11852
rect 16448 11840 16454 11892
rect 17494 11880 17500 11892
rect 17455 11852 17500 11880
rect 17494 11840 17500 11852
rect 17552 11840 17558 11892
rect 20257 11883 20315 11889
rect 20257 11849 20269 11883
rect 20303 11880 20315 11883
rect 20622 11880 20628 11892
rect 20303 11852 20628 11880
rect 20303 11849 20315 11852
rect 20257 11843 20315 11849
rect 20622 11840 20628 11852
rect 20680 11840 20686 11892
rect 21818 11880 21824 11892
rect 21779 11852 21824 11880
rect 21818 11840 21824 11852
rect 21876 11840 21882 11892
rect 23198 11840 23204 11892
rect 23256 11880 23262 11892
rect 23477 11883 23535 11889
rect 23477 11880 23489 11883
rect 23256 11852 23489 11880
rect 23256 11840 23262 11852
rect 23477 11849 23489 11852
rect 23523 11880 23535 11883
rect 23566 11880 23572 11892
rect 23523 11852 23572 11880
rect 23523 11849 23535 11852
rect 23477 11843 23535 11849
rect 23566 11840 23572 11852
rect 23624 11880 23630 11892
rect 24489 11883 24547 11889
rect 24489 11880 24501 11883
rect 23624 11852 24501 11880
rect 23624 11840 23630 11852
rect 24489 11849 24501 11852
rect 24535 11849 24547 11883
rect 24670 11880 24676 11892
rect 24631 11852 24676 11880
rect 24489 11843 24547 11849
rect 24670 11840 24676 11852
rect 24728 11840 24734 11892
rect 25409 11883 25467 11889
rect 25409 11849 25421 11883
rect 25455 11880 25467 11883
rect 26418 11880 26424 11892
rect 25455 11852 26424 11880
rect 25455 11849 25467 11852
rect 25409 11843 25467 11849
rect 26418 11840 26424 11852
rect 26476 11840 26482 11892
rect 5074 11812 5080 11824
rect 5035 11784 5080 11812
rect 5074 11772 5080 11784
rect 5132 11812 5138 11824
rect 7837 11815 7895 11821
rect 7837 11812 7849 11815
rect 5132 11784 7849 11812
rect 5132 11772 5138 11784
rect 7837 11781 7849 11784
rect 7883 11812 7895 11815
rect 7926 11812 7932 11824
rect 7883 11784 7932 11812
rect 7883 11781 7895 11784
rect 7837 11775 7895 11781
rect 7926 11772 7932 11784
rect 7984 11772 7990 11824
rect 9122 11772 9128 11824
rect 9180 11812 9186 11824
rect 9950 11812 9956 11824
rect 9180 11784 9956 11812
rect 9180 11772 9186 11784
rect 9950 11772 9956 11784
rect 10008 11772 10014 11824
rect 10686 11772 10692 11824
rect 10744 11812 10750 11824
rect 14550 11812 14556 11824
rect 10744 11784 10824 11812
rect 14511 11784 14556 11812
rect 10744 11772 10750 11784
rect 2133 11747 2191 11753
rect 2133 11713 2145 11747
rect 2179 11713 2191 11747
rect 2133 11707 2191 11713
rect 4709 11747 4767 11753
rect 4709 11713 4721 11747
rect 4755 11744 4767 11747
rect 5721 11747 5779 11753
rect 5721 11744 5733 11747
rect 4755 11716 5733 11744
rect 4755 11713 4767 11716
rect 4709 11707 4767 11713
rect 5721 11713 5733 11716
rect 5767 11744 5779 11747
rect 6178 11744 6184 11756
rect 5767 11716 6184 11744
rect 5767 11713 5779 11716
rect 5721 11707 5779 11713
rect 6178 11704 6184 11716
rect 6236 11704 6242 11756
rect 6454 11704 6460 11756
rect 6512 11744 6518 11756
rect 8021 11747 8079 11753
rect 8021 11744 8033 11747
rect 6512 11716 8033 11744
rect 6512 11704 6518 11716
rect 8021 11713 8033 11716
rect 8067 11713 8079 11747
rect 8021 11707 8079 11713
rect 9858 11704 9864 11756
rect 9916 11744 9922 11756
rect 10502 11744 10508 11756
rect 9916 11716 10508 11744
rect 9916 11704 9922 11716
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 10796 11753 10824 11784
rect 14550 11772 14556 11784
rect 14608 11772 14614 11824
rect 23661 11815 23719 11821
rect 23661 11781 23673 11815
rect 23707 11812 23719 11815
rect 25222 11812 25228 11824
rect 23707 11784 25228 11812
rect 23707 11781 23719 11784
rect 23661 11775 23719 11781
rect 25222 11772 25228 11784
rect 25280 11772 25286 11824
rect 10781 11747 10839 11753
rect 10781 11713 10793 11747
rect 10827 11744 10839 11747
rect 10962 11744 10968 11756
rect 10827 11716 10968 11744
rect 10827 11713 10839 11716
rect 10781 11707 10839 11713
rect 10962 11704 10968 11716
rect 11020 11744 11026 11756
rect 11609 11747 11667 11753
rect 11609 11744 11621 11747
rect 11020 11716 11621 11744
rect 11020 11704 11026 11716
rect 11609 11713 11621 11716
rect 11655 11713 11667 11747
rect 12434 11744 12440 11756
rect 12395 11716 12440 11744
rect 11609 11707 11667 11713
rect 12434 11704 12440 11716
rect 12492 11704 12498 11756
rect 13814 11704 13820 11756
rect 13872 11744 13878 11756
rect 14185 11747 14243 11753
rect 14185 11744 14197 11747
rect 13872 11716 14197 11744
rect 13872 11704 13878 11716
rect 14185 11713 14197 11716
rect 14231 11744 14243 11747
rect 15197 11747 15255 11753
rect 15197 11744 15209 11747
rect 14231 11716 15209 11744
rect 14231 11713 14243 11716
rect 14185 11707 14243 11713
rect 15197 11713 15209 11716
rect 15243 11713 15255 11747
rect 16942 11744 16948 11756
rect 16903 11716 16948 11744
rect 15197 11707 15255 11713
rect 16942 11704 16948 11716
rect 17000 11744 17006 11756
rect 17954 11744 17960 11756
rect 17000 11716 17960 11744
rect 17000 11704 17006 11716
rect 17954 11704 17960 11716
rect 18012 11744 18018 11756
rect 18012 11716 18184 11744
rect 18012 11704 18018 11716
rect 5629 11679 5687 11685
rect 5629 11645 5641 11679
rect 5675 11676 5687 11679
rect 6086 11676 6092 11688
rect 5675 11648 6092 11676
rect 5675 11645 5687 11648
rect 5629 11639 5687 11645
rect 6086 11636 6092 11648
rect 6144 11636 6150 11688
rect 7926 11636 7932 11688
rect 7984 11676 7990 11688
rect 8277 11679 8335 11685
rect 8277 11676 8289 11679
rect 7984 11648 8289 11676
rect 7984 11636 7990 11648
rect 8277 11645 8289 11648
rect 8323 11645 8335 11679
rect 8277 11639 8335 11645
rect 10137 11679 10195 11685
rect 10137 11645 10149 11679
rect 10183 11676 10195 11679
rect 10689 11679 10747 11685
rect 10689 11676 10701 11679
rect 10183 11648 10701 11676
rect 10183 11645 10195 11648
rect 10137 11639 10195 11645
rect 10689 11645 10701 11648
rect 10735 11676 10747 11679
rect 11698 11676 11704 11688
rect 10735 11648 11704 11676
rect 10735 11645 10747 11648
rect 10689 11639 10747 11645
rect 11698 11636 11704 11648
rect 11756 11636 11762 11688
rect 13262 11636 13268 11688
rect 13320 11676 13326 11688
rect 13906 11676 13912 11688
rect 13320 11648 13912 11676
rect 13320 11636 13326 11648
rect 13906 11636 13912 11648
rect 13964 11636 13970 11688
rect 14550 11636 14556 11688
rect 14608 11676 14614 11688
rect 15105 11679 15163 11685
rect 15105 11676 15117 11679
rect 14608 11648 15117 11676
rect 14608 11636 14614 11648
rect 15105 11645 15117 11648
rect 15151 11645 15163 11679
rect 18049 11679 18107 11685
rect 18049 11676 18061 11679
rect 15105 11639 15163 11645
rect 15212 11648 18061 11676
rect 15212 11620 15240 11648
rect 18049 11645 18061 11648
rect 18095 11645 18107 11679
rect 18156 11676 18184 11716
rect 20254 11704 20260 11756
rect 20312 11744 20318 11756
rect 20717 11747 20775 11753
rect 20717 11744 20729 11747
rect 20312 11716 20729 11744
rect 20312 11704 20318 11716
rect 20717 11713 20729 11716
rect 20763 11713 20775 11747
rect 20717 11707 20775 11713
rect 20809 11747 20867 11753
rect 20809 11713 20821 11747
rect 20855 11713 20867 11747
rect 20809 11707 20867 11713
rect 18305 11679 18363 11685
rect 18305 11676 18317 11679
rect 18156 11648 18317 11676
rect 18049 11639 18107 11645
rect 18305 11645 18317 11648
rect 18351 11676 18363 11679
rect 19518 11676 19524 11688
rect 18351 11648 19524 11676
rect 18351 11645 18363 11648
rect 18305 11639 18363 11645
rect 2041 11611 2099 11617
rect 2041 11577 2053 11611
rect 2087 11608 2099 11611
rect 2130 11608 2136 11620
rect 2087 11580 2136 11608
rect 2087 11577 2099 11580
rect 2041 11571 2099 11577
rect 2130 11568 2136 11580
rect 2188 11608 2194 11620
rect 2400 11611 2458 11617
rect 2400 11608 2412 11611
rect 2188 11580 2412 11608
rect 2188 11568 2194 11580
rect 2400 11577 2412 11580
rect 2446 11608 2458 11611
rect 2682 11608 2688 11620
rect 2446 11580 2688 11608
rect 2446 11577 2458 11580
rect 2400 11571 2458 11577
rect 2682 11568 2688 11580
rect 2740 11568 2746 11620
rect 5534 11608 5540 11620
rect 5495 11580 5540 11608
rect 5534 11568 5540 11580
rect 5592 11568 5598 11620
rect 10318 11568 10324 11620
rect 10376 11608 10382 11620
rect 10376 11580 10916 11608
rect 10376 11568 10382 11580
rect 10888 11552 10916 11580
rect 12526 11568 12532 11620
rect 12584 11608 12590 11620
rect 12704 11611 12762 11617
rect 12704 11608 12716 11611
rect 12584 11580 12716 11608
rect 12584 11568 12590 11580
rect 12704 11577 12716 11580
rect 12750 11608 12762 11611
rect 13538 11608 13544 11620
rect 12750 11580 13544 11608
rect 12750 11577 12762 11580
rect 12704 11571 12762 11577
rect 13538 11568 13544 11580
rect 13596 11568 13602 11620
rect 15194 11568 15200 11620
rect 15252 11568 15258 11620
rect 16853 11611 16911 11617
rect 16853 11608 16865 11611
rect 15948 11580 16865 11608
rect 15948 11552 15976 11580
rect 16853 11577 16865 11580
rect 16899 11577 16911 11611
rect 16853 11571 16911 11577
rect 17954 11568 17960 11620
rect 18012 11608 18018 11620
rect 18064 11608 18092 11639
rect 19518 11636 19524 11648
rect 19576 11636 19582 11688
rect 20165 11679 20223 11685
rect 20165 11645 20177 11679
rect 20211 11676 20223 11679
rect 20622 11676 20628 11688
rect 20211 11648 20628 11676
rect 20211 11645 20223 11648
rect 20165 11639 20223 11645
rect 20622 11636 20628 11648
rect 20680 11676 20686 11688
rect 20824 11676 20852 11707
rect 22002 11704 22008 11756
rect 22060 11744 22066 11756
rect 22465 11747 22523 11753
rect 22465 11744 22477 11747
rect 22060 11716 22477 11744
rect 22060 11704 22066 11716
rect 22465 11713 22477 11716
rect 22511 11744 22523 11747
rect 22830 11744 22836 11756
rect 22511 11716 22836 11744
rect 22511 11713 22523 11716
rect 22465 11707 22523 11713
rect 22830 11704 22836 11716
rect 22888 11704 22894 11756
rect 23014 11704 23020 11756
rect 23072 11704 23078 11756
rect 24118 11744 24124 11756
rect 24079 11716 24124 11744
rect 24118 11704 24124 11716
rect 24176 11704 24182 11756
rect 24305 11747 24363 11753
rect 24305 11713 24317 11747
rect 24351 11744 24363 11747
rect 24489 11747 24547 11753
rect 24489 11744 24501 11747
rect 24351 11716 24501 11744
rect 24351 11713 24363 11716
rect 24305 11707 24363 11713
rect 24489 11713 24501 11716
rect 24535 11713 24547 11747
rect 24489 11707 24547 11713
rect 25133 11747 25191 11753
rect 25133 11713 25145 11747
rect 25179 11744 25191 11747
rect 25866 11744 25872 11756
rect 25179 11716 25872 11744
rect 25179 11713 25191 11716
rect 25133 11707 25191 11713
rect 20680 11648 20852 11676
rect 22925 11679 22983 11685
rect 20680 11636 20686 11648
rect 22925 11645 22937 11679
rect 22971 11676 22983 11679
rect 23032 11676 23060 11704
rect 23198 11676 23204 11688
rect 22971 11648 23204 11676
rect 22971 11645 22983 11648
rect 22925 11639 22983 11645
rect 23198 11636 23204 11648
rect 23256 11636 23262 11688
rect 24029 11679 24087 11685
rect 24029 11645 24041 11679
rect 24075 11676 24087 11679
rect 25148 11676 25176 11707
rect 25866 11704 25872 11716
rect 25924 11704 25930 11756
rect 24075 11648 25176 11676
rect 25225 11679 25283 11685
rect 24075 11645 24087 11648
rect 24029 11639 24087 11645
rect 25225 11645 25237 11679
rect 25271 11676 25283 11679
rect 25406 11676 25412 11688
rect 25271 11648 25412 11676
rect 25271 11645 25283 11648
rect 25225 11639 25283 11645
rect 25406 11636 25412 11648
rect 25464 11636 25470 11688
rect 18012 11580 18092 11608
rect 18012 11568 18018 11580
rect 19334 11568 19340 11620
rect 19392 11608 19398 11620
rect 19705 11611 19763 11617
rect 19705 11608 19717 11611
rect 19392 11580 19717 11608
rect 19392 11568 19398 11580
rect 19705 11577 19717 11580
rect 19751 11577 19763 11611
rect 19705 11571 19763 11577
rect 21361 11611 21419 11617
rect 21361 11577 21373 11611
rect 21407 11608 21419 11611
rect 21726 11608 21732 11620
rect 21407 11580 21732 11608
rect 21407 11577 21419 11580
rect 21361 11571 21419 11577
rect 21726 11568 21732 11580
rect 21784 11608 21790 11620
rect 22281 11611 22339 11617
rect 22281 11608 22293 11611
rect 21784 11580 22293 11608
rect 21784 11568 21790 11580
rect 22281 11577 22293 11580
rect 22327 11608 22339 11611
rect 22830 11608 22836 11620
rect 22327 11580 22836 11608
rect 22327 11577 22339 11580
rect 22281 11571 22339 11577
rect 22830 11568 22836 11580
rect 22888 11568 22894 11620
rect 24210 11568 24216 11620
rect 24268 11608 24274 11620
rect 24854 11608 24860 11620
rect 24268 11580 24860 11608
rect 24268 11568 24274 11580
rect 24854 11568 24860 11580
rect 24912 11608 24918 11620
rect 25777 11611 25835 11617
rect 25777 11608 25789 11611
rect 24912 11580 25789 11608
rect 24912 11568 24918 11580
rect 25777 11577 25789 11580
rect 25823 11577 25835 11611
rect 25777 11571 25835 11577
rect 1673 11543 1731 11549
rect 1673 11509 1685 11543
rect 1719 11540 1731 11543
rect 1854 11540 1860 11552
rect 1719 11512 1860 11540
rect 1719 11509 1731 11512
rect 1673 11503 1731 11509
rect 1854 11500 1860 11512
rect 1912 11540 1918 11552
rect 2958 11540 2964 11552
rect 1912 11512 2964 11540
rect 1912 11500 1918 11512
rect 2958 11500 2964 11512
rect 3016 11500 3022 11552
rect 3510 11540 3516 11552
rect 3471 11512 3516 11540
rect 3510 11500 3516 11512
rect 3568 11500 3574 11552
rect 5166 11540 5172 11552
rect 5127 11512 5172 11540
rect 5166 11500 5172 11512
rect 5224 11500 5230 11552
rect 6822 11540 6828 11552
rect 6783 11512 6828 11540
rect 6822 11500 6828 11512
rect 6880 11500 6886 11552
rect 9401 11543 9459 11549
rect 9401 11509 9413 11543
rect 9447 11540 9459 11543
rect 9490 11540 9496 11552
rect 9447 11512 9496 11540
rect 9447 11509 9459 11512
rect 9401 11503 9459 11509
rect 9490 11500 9496 11512
rect 9548 11500 9554 11552
rect 10134 11500 10140 11552
rect 10192 11540 10198 11552
rect 10597 11543 10655 11549
rect 10597 11540 10609 11543
rect 10192 11512 10609 11540
rect 10192 11500 10198 11512
rect 10597 11509 10609 11512
rect 10643 11509 10655 11543
rect 10597 11503 10655 11509
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 11238 11540 11244 11552
rect 10928 11512 11244 11540
rect 10928 11500 10934 11512
rect 11238 11500 11244 11512
rect 11296 11500 11302 11552
rect 11330 11500 11336 11552
rect 11388 11540 11394 11552
rect 12161 11543 12219 11549
rect 12161 11540 12173 11543
rect 11388 11512 12173 11540
rect 11388 11500 11394 11512
rect 12161 11509 12173 11512
rect 12207 11540 12219 11543
rect 12250 11540 12256 11552
rect 12207 11512 12256 11540
rect 12207 11509 12219 11512
rect 12161 11503 12219 11509
rect 12250 11500 12256 11512
rect 12308 11500 12314 11552
rect 13814 11540 13820 11552
rect 13775 11512 13820 11540
rect 13814 11500 13820 11512
rect 13872 11500 13878 11552
rect 14642 11500 14648 11552
rect 14700 11540 14706 11552
rect 15013 11543 15071 11549
rect 15013 11540 15025 11543
rect 14700 11512 15025 11540
rect 14700 11500 14706 11512
rect 15013 11509 15025 11512
rect 15059 11509 15071 11543
rect 15930 11540 15936 11552
rect 15891 11512 15936 11540
rect 15013 11503 15071 11509
rect 15930 11500 15936 11512
rect 15988 11500 15994 11552
rect 16301 11543 16359 11549
rect 16301 11509 16313 11543
rect 16347 11540 16359 11543
rect 16761 11543 16819 11549
rect 16761 11540 16773 11543
rect 16347 11512 16773 11540
rect 16347 11509 16359 11512
rect 16301 11503 16359 11509
rect 16761 11509 16773 11512
rect 16807 11540 16819 11543
rect 17310 11540 17316 11552
rect 16807 11512 17316 11540
rect 16807 11509 16819 11512
rect 16761 11503 16819 11509
rect 17310 11500 17316 11512
rect 17368 11500 17374 11552
rect 19429 11543 19487 11549
rect 19429 11509 19441 11543
rect 19475 11540 19487 11543
rect 19518 11540 19524 11552
rect 19475 11512 19524 11540
rect 19475 11509 19487 11512
rect 19429 11503 19487 11509
rect 19518 11500 19524 11512
rect 19576 11500 19582 11552
rect 20254 11500 20260 11552
rect 20312 11540 20318 11552
rect 20625 11543 20683 11549
rect 20625 11540 20637 11543
rect 20312 11512 20637 11540
rect 20312 11500 20318 11512
rect 20625 11509 20637 11512
rect 20671 11509 20683 11543
rect 20625 11503 20683 11509
rect 21637 11543 21695 11549
rect 21637 11509 21649 11543
rect 21683 11540 21695 11543
rect 21818 11540 21824 11552
rect 21683 11512 21824 11540
rect 21683 11509 21695 11512
rect 21637 11503 21695 11509
rect 21818 11500 21824 11512
rect 21876 11540 21882 11552
rect 22189 11543 22247 11549
rect 22189 11540 22201 11543
rect 21876 11512 22201 11540
rect 21876 11500 21882 11512
rect 22189 11509 22201 11512
rect 22235 11509 22247 11543
rect 26234 11540 26240 11552
rect 26195 11512 26240 11540
rect 22189 11503 22247 11509
rect 26234 11500 26240 11512
rect 26292 11500 26298 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1762 11296 1768 11348
rect 1820 11336 1826 11348
rect 2130 11336 2136 11348
rect 1820 11308 2136 11336
rect 1820 11296 1826 11308
rect 2130 11296 2136 11308
rect 2188 11296 2194 11348
rect 2958 11336 2964 11348
rect 2919 11308 2964 11336
rect 2958 11296 2964 11308
rect 3016 11296 3022 11348
rect 4617 11339 4675 11345
rect 4617 11305 4629 11339
rect 4663 11336 4675 11339
rect 5534 11336 5540 11348
rect 4663 11308 5540 11336
rect 4663 11305 4675 11308
rect 4617 11299 4675 11305
rect 5534 11296 5540 11308
rect 5592 11296 5598 11348
rect 6822 11296 6828 11348
rect 6880 11336 6886 11348
rect 7285 11339 7343 11345
rect 7285 11336 7297 11339
rect 6880 11308 7297 11336
rect 6880 11296 6886 11308
rect 7285 11305 7297 11308
rect 7331 11336 7343 11339
rect 7374 11336 7380 11348
rect 7331 11308 7380 11336
rect 7331 11305 7343 11308
rect 7285 11299 7343 11305
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 8110 11336 8116 11348
rect 8071 11308 8116 11336
rect 8110 11296 8116 11308
rect 8168 11296 8174 11348
rect 8478 11336 8484 11348
rect 8439 11308 8484 11336
rect 8478 11296 8484 11308
rect 8536 11296 8542 11348
rect 8573 11339 8631 11345
rect 8573 11305 8585 11339
rect 8619 11336 8631 11339
rect 9214 11336 9220 11348
rect 8619 11308 9220 11336
rect 8619 11305 8631 11308
rect 8573 11299 8631 11305
rect 9214 11296 9220 11308
rect 9272 11296 9278 11348
rect 9398 11336 9404 11348
rect 9359 11308 9404 11336
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 9674 11336 9680 11348
rect 9635 11308 9680 11336
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 10134 11296 10140 11348
rect 10192 11336 10198 11348
rect 10689 11339 10747 11345
rect 10689 11336 10701 11339
rect 10192 11308 10701 11336
rect 10192 11296 10198 11308
rect 10689 11305 10701 11308
rect 10735 11305 10747 11339
rect 10689 11299 10747 11305
rect 11514 11296 11520 11348
rect 11572 11336 11578 11348
rect 12805 11339 12863 11345
rect 12805 11336 12817 11339
rect 11572 11308 12817 11336
rect 11572 11296 11578 11308
rect 12805 11305 12817 11308
rect 12851 11305 12863 11339
rect 13630 11336 13636 11348
rect 13591 11308 13636 11336
rect 12805 11299 12863 11305
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 13906 11296 13912 11348
rect 13964 11336 13970 11348
rect 14093 11339 14151 11345
rect 14093 11336 14105 11339
rect 13964 11308 14105 11336
rect 13964 11296 13970 11308
rect 14093 11305 14105 11308
rect 14139 11305 14151 11339
rect 14642 11336 14648 11348
rect 14603 11308 14648 11336
rect 14093 11299 14151 11305
rect 14642 11296 14648 11308
rect 14700 11296 14706 11348
rect 15105 11339 15163 11345
rect 15105 11305 15117 11339
rect 15151 11336 15163 11339
rect 15746 11336 15752 11348
rect 15151 11308 15752 11336
rect 15151 11305 15163 11308
rect 15105 11299 15163 11305
rect 15746 11296 15752 11308
rect 15804 11296 15810 11348
rect 16669 11339 16727 11345
rect 16669 11305 16681 11339
rect 16715 11336 16727 11339
rect 17034 11336 17040 11348
rect 16715 11308 17040 11336
rect 16715 11305 16727 11308
rect 16669 11299 16727 11305
rect 17034 11296 17040 11308
rect 17092 11336 17098 11348
rect 17310 11336 17316 11348
rect 17092 11308 17316 11336
rect 17092 11296 17098 11308
rect 17310 11296 17316 11308
rect 17368 11296 17374 11348
rect 19978 11296 19984 11348
rect 20036 11336 20042 11348
rect 20901 11339 20959 11345
rect 20901 11336 20913 11339
rect 20036 11308 20913 11336
rect 20036 11296 20042 11308
rect 20901 11305 20913 11308
rect 20947 11305 20959 11339
rect 22002 11336 22008 11348
rect 21963 11308 22008 11336
rect 20901 11299 20959 11305
rect 22002 11296 22008 11308
rect 22060 11296 22066 11348
rect 22738 11296 22744 11348
rect 22796 11336 22802 11348
rect 23014 11336 23020 11348
rect 22796 11308 22876 11336
rect 22975 11308 23020 11336
rect 22796 11296 22802 11308
rect 4976 11271 5034 11277
rect 1596 11240 3832 11268
rect 1596 11209 1624 11240
rect 1854 11209 1860 11212
rect 1581 11203 1639 11209
rect 1581 11169 1593 11203
rect 1627 11169 1639 11203
rect 1848 11200 1860 11209
rect 1815 11172 1860 11200
rect 1581 11163 1639 11169
rect 1848 11163 1860 11172
rect 1912 11200 1918 11212
rect 2130 11200 2136 11212
rect 1912 11172 2136 11200
rect 1854 11160 1860 11163
rect 1912 11160 1918 11172
rect 2130 11160 2136 11172
rect 2188 11200 2194 11212
rect 3510 11200 3516 11212
rect 2188 11172 3516 11200
rect 2188 11160 2194 11172
rect 3510 11160 3516 11172
rect 3568 11160 3574 11212
rect 2774 11092 2780 11144
rect 2832 11132 2838 11144
rect 3237 11135 3295 11141
rect 3237 11132 3249 11135
rect 2832 11104 3249 11132
rect 2832 11092 2838 11104
rect 3237 11101 3249 11104
rect 3283 11101 3295 11135
rect 3237 11095 3295 11101
rect 3804 11132 3832 11240
rect 4976 11237 4988 11271
rect 5022 11268 5034 11271
rect 5074 11268 5080 11280
rect 5022 11240 5080 11268
rect 5022 11237 5034 11240
rect 4976 11231 5034 11237
rect 5074 11228 5080 11240
rect 5132 11228 5138 11280
rect 6086 11160 6092 11212
rect 6144 11200 6150 11212
rect 6365 11203 6423 11209
rect 6365 11200 6377 11203
rect 6144 11172 6377 11200
rect 6144 11160 6150 11172
rect 6365 11169 6377 11172
rect 6411 11200 6423 11203
rect 6733 11203 6791 11209
rect 6733 11200 6745 11203
rect 6411 11172 6745 11200
rect 6411 11169 6423 11172
rect 6365 11163 6423 11169
rect 6733 11169 6745 11172
rect 6779 11169 6791 11203
rect 7374 11200 7380 11212
rect 7335 11172 7380 11200
rect 6733 11163 6791 11169
rect 4709 11135 4767 11141
rect 4709 11132 4721 11135
rect 3804 11104 4721 11132
rect 3804 11008 3832 11104
rect 4709 11101 4721 11104
rect 4755 11101 4767 11135
rect 6748 11132 6776 11163
rect 7374 11160 7380 11172
rect 7432 11200 7438 11212
rect 7834 11200 7840 11212
rect 7432 11172 7840 11200
rect 7432 11160 7438 11172
rect 7834 11160 7840 11172
rect 7892 11160 7898 11212
rect 8128 11200 8156 11296
rect 11790 11228 11796 11280
rect 11848 11268 11854 11280
rect 12069 11271 12127 11277
rect 12069 11268 12081 11271
rect 11848 11240 12081 11268
rect 11848 11228 11854 11240
rect 12069 11237 12081 11240
rect 12115 11237 12127 11271
rect 12069 11231 12127 11237
rect 13265 11271 13323 11277
rect 13265 11237 13277 11271
rect 13311 11268 13323 11271
rect 14274 11268 14280 11280
rect 13311 11240 14280 11268
rect 13311 11237 13323 11240
rect 13265 11231 13323 11237
rect 13648 11212 13676 11240
rect 14274 11228 14280 11240
rect 14332 11268 14338 11280
rect 15556 11271 15614 11277
rect 14332 11240 15516 11268
rect 14332 11228 14338 11240
rect 8478 11200 8484 11212
rect 8128 11172 8484 11200
rect 8478 11160 8484 11172
rect 8536 11160 8542 11212
rect 9674 11160 9680 11212
rect 9732 11200 9738 11212
rect 10045 11203 10103 11209
rect 10045 11200 10057 11203
rect 9732 11172 10057 11200
rect 9732 11160 9738 11172
rect 10045 11169 10057 11172
rect 10091 11169 10103 11203
rect 10045 11163 10103 11169
rect 10137 11203 10195 11209
rect 10137 11169 10149 11203
rect 10183 11200 10195 11203
rect 10594 11200 10600 11212
rect 10183 11172 10600 11200
rect 10183 11169 10195 11172
rect 10137 11163 10195 11169
rect 10594 11160 10600 11172
rect 10652 11160 10658 11212
rect 11698 11160 11704 11212
rect 11756 11200 11762 11212
rect 12161 11203 12219 11209
rect 12161 11200 12173 11203
rect 11756 11172 12173 11200
rect 11756 11160 11762 11172
rect 12161 11169 12173 11172
rect 12207 11200 12219 11203
rect 12342 11200 12348 11212
rect 12207 11172 12348 11200
rect 12207 11169 12219 11172
rect 12161 11163 12219 11169
rect 12342 11160 12348 11172
rect 12400 11160 12406 11212
rect 13170 11200 13176 11212
rect 13131 11172 13176 11200
rect 13170 11160 13176 11172
rect 13228 11160 13234 11212
rect 13630 11160 13636 11212
rect 13688 11160 13694 11212
rect 14001 11203 14059 11209
rect 14001 11169 14013 11203
rect 14047 11200 14059 11203
rect 14366 11200 14372 11212
rect 14047 11172 14372 11200
rect 14047 11169 14059 11172
rect 14001 11163 14059 11169
rect 14366 11160 14372 11172
rect 14424 11160 14430 11212
rect 15488 11200 15516 11240
rect 15556 11237 15568 11271
rect 15602 11268 15614 11271
rect 15654 11268 15660 11280
rect 15602 11240 15660 11268
rect 15602 11237 15614 11240
rect 15556 11231 15614 11237
rect 15654 11228 15660 11240
rect 15712 11268 15718 11280
rect 16850 11268 16856 11280
rect 15712 11240 16856 11268
rect 15712 11228 15718 11240
rect 16850 11228 16856 11240
rect 16908 11228 16914 11280
rect 18046 11200 18052 11212
rect 15488 11172 18052 11200
rect 18046 11160 18052 11172
rect 18104 11160 18110 11212
rect 18230 11209 18236 11212
rect 18224 11200 18236 11209
rect 18143 11172 18236 11200
rect 18224 11163 18236 11172
rect 18288 11200 18294 11212
rect 19981 11203 20039 11209
rect 18288 11172 19564 11200
rect 18230 11160 18236 11163
rect 18288 11160 18294 11172
rect 19536 11144 19564 11172
rect 19981 11169 19993 11203
rect 20027 11200 20039 11203
rect 20070 11200 20076 11212
rect 20027 11172 20076 11200
rect 20027 11169 20039 11172
rect 19981 11163 20039 11169
rect 20070 11160 20076 11172
rect 20128 11200 20134 11212
rect 21269 11203 21327 11209
rect 21269 11200 21281 11203
rect 20128 11172 21281 11200
rect 20128 11160 20134 11172
rect 21269 11169 21281 11172
rect 21315 11169 21327 11203
rect 22281 11203 22339 11209
rect 22281 11200 22293 11203
rect 21269 11163 21327 11169
rect 21376 11172 22293 11200
rect 21376 11144 21404 11172
rect 22281 11169 22293 11172
rect 22327 11169 22339 11203
rect 22281 11163 22339 11169
rect 22465 11203 22523 11209
rect 22465 11169 22477 11203
rect 22511 11200 22523 11203
rect 22738 11200 22744 11212
rect 22511 11172 22744 11200
rect 22511 11169 22523 11172
rect 22465 11163 22523 11169
rect 22738 11160 22744 11172
rect 22796 11160 22802 11212
rect 22848 11200 22876 11308
rect 23014 11296 23020 11308
rect 23072 11296 23078 11348
rect 23198 11296 23204 11348
rect 23256 11336 23262 11348
rect 24026 11336 24032 11348
rect 23256 11308 24032 11336
rect 23256 11296 23262 11308
rect 24026 11296 24032 11308
rect 24084 11296 24090 11348
rect 24946 11336 24952 11348
rect 24907 11308 24952 11336
rect 24946 11296 24952 11308
rect 25004 11296 25010 11348
rect 25222 11336 25228 11348
rect 25183 11308 25228 11336
rect 25222 11296 25228 11308
rect 25280 11296 25286 11348
rect 25314 11296 25320 11348
rect 25372 11336 25378 11348
rect 25961 11339 26019 11345
rect 25961 11336 25973 11339
rect 25372 11308 25973 11336
rect 25372 11296 25378 11308
rect 25961 11305 25973 11308
rect 26007 11305 26019 11339
rect 25961 11299 26019 11305
rect 23382 11228 23388 11280
rect 23440 11268 23446 11280
rect 23814 11271 23872 11277
rect 23814 11268 23826 11271
rect 23440 11240 23826 11268
rect 23440 11228 23446 11240
rect 23814 11237 23826 11240
rect 23860 11268 23872 11271
rect 24670 11268 24676 11280
rect 23860 11240 24676 11268
rect 23860 11237 23872 11240
rect 23814 11231 23872 11237
rect 24670 11228 24676 11240
rect 24728 11228 24734 11280
rect 23014 11200 23020 11212
rect 22848 11172 23020 11200
rect 23014 11160 23020 11172
rect 23072 11160 23078 11212
rect 7469 11135 7527 11141
rect 7469 11132 7481 11135
rect 6748 11104 7481 11132
rect 4709 11095 4767 11101
rect 7469 11101 7481 11104
rect 7515 11132 7527 11135
rect 7558 11132 7564 11144
rect 7515 11104 7564 11132
rect 7515 11101 7527 11104
rect 7469 11095 7527 11101
rect 7558 11092 7564 11104
rect 7616 11092 7622 11144
rect 10229 11135 10287 11141
rect 10229 11101 10241 11135
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 11241 11135 11299 11141
rect 11241 11101 11253 11135
rect 11287 11132 11299 11135
rect 12066 11132 12072 11144
rect 11287 11104 12072 11132
rect 11287 11101 11299 11104
rect 11241 11095 11299 11101
rect 6914 11064 6920 11076
rect 6875 11036 6920 11064
rect 6914 11024 6920 11036
rect 6972 11024 6978 11076
rect 8110 11024 8116 11076
rect 8168 11064 8174 11076
rect 9033 11067 9091 11073
rect 9033 11064 9045 11067
rect 8168 11036 9045 11064
rect 8168 11024 8174 11036
rect 9033 11033 9045 11036
rect 9079 11064 9091 11067
rect 10244 11064 10272 11095
rect 12066 11092 12072 11104
rect 12124 11092 12130 11144
rect 12253 11135 12311 11141
rect 12253 11101 12265 11135
rect 12299 11101 12311 11135
rect 12253 11095 12311 11101
rect 13357 11135 13415 11141
rect 13357 11101 13369 11135
rect 13403 11132 13415 11135
rect 13906 11132 13912 11144
rect 13403 11104 13912 11132
rect 13403 11101 13415 11104
rect 13357 11095 13415 11101
rect 10318 11064 10324 11076
rect 9079 11036 10324 11064
rect 9079 11033 9091 11036
rect 9033 11027 9091 11033
rect 10318 11024 10324 11036
rect 10376 11064 10382 11076
rect 10962 11064 10968 11076
rect 10376 11036 10968 11064
rect 10376 11024 10382 11036
rect 10962 11024 10968 11036
rect 11020 11024 11026 11076
rect 11054 11024 11060 11076
rect 11112 11064 11118 11076
rect 11701 11067 11759 11073
rect 11701 11064 11713 11067
rect 11112 11036 11713 11064
rect 11112 11024 11118 11036
rect 11701 11033 11713 11036
rect 11747 11033 11759 11067
rect 12268 11064 12296 11095
rect 11701 11027 11759 11033
rect 12176 11036 12296 11064
rect 3697 10999 3755 11005
rect 3697 10965 3709 10999
rect 3743 10996 3755 10999
rect 3786 10996 3792 11008
rect 3743 10968 3792 10996
rect 3743 10965 3755 10968
rect 3697 10959 3755 10965
rect 3786 10956 3792 10968
rect 3844 10956 3850 11008
rect 3970 10956 3976 11008
rect 4028 10996 4034 11008
rect 6089 10999 6147 11005
rect 6089 10996 6101 10999
rect 4028 10968 6101 10996
rect 4028 10956 4034 10968
rect 6089 10965 6101 10968
rect 6135 10996 6147 10999
rect 6454 10996 6460 11008
rect 6135 10968 6460 10996
rect 6135 10965 6147 10968
rect 6089 10959 6147 10965
rect 6454 10956 6460 10968
rect 6512 10956 6518 11008
rect 11422 10956 11428 11008
rect 11480 10996 11486 11008
rect 11517 10999 11575 11005
rect 11517 10996 11529 10999
rect 11480 10968 11529 10996
rect 11480 10956 11486 10968
rect 11517 10965 11529 10968
rect 11563 10996 11575 10999
rect 12176 10996 12204 11036
rect 12342 11024 12348 11076
rect 12400 11064 12406 11076
rect 13372 11064 13400 11095
rect 13906 11092 13912 11104
rect 13964 11132 13970 11144
rect 14185 11135 14243 11141
rect 14185 11132 14197 11135
rect 13964 11104 14197 11132
rect 13964 11092 13970 11104
rect 14185 11101 14197 11104
rect 14231 11101 14243 11135
rect 14185 11095 14243 11101
rect 15194 11092 15200 11144
rect 15252 11132 15258 11144
rect 15289 11135 15347 11141
rect 15289 11132 15301 11135
rect 15252 11104 15301 11132
rect 15252 11092 15258 11104
rect 15289 11101 15301 11104
rect 15335 11101 15347 11135
rect 17954 11132 17960 11144
rect 17915 11104 17960 11132
rect 15289 11095 15347 11101
rect 17954 11092 17960 11104
rect 18012 11092 18018 11144
rect 19518 11092 19524 11144
rect 19576 11132 19582 11144
rect 21358 11132 21364 11144
rect 19576 11104 20760 11132
rect 21319 11104 21364 11132
rect 19576 11092 19582 11104
rect 12400 11036 13400 11064
rect 12400 11024 12406 11036
rect 14274 11024 14280 11076
rect 14332 11064 14338 11076
rect 14332 11036 14955 11064
rect 14332 11024 14338 11036
rect 11563 10968 12204 10996
rect 11563 10965 11575 10968
rect 11517 10959 11575 10965
rect 13998 10956 14004 11008
rect 14056 10996 14062 11008
rect 14826 10996 14832 11008
rect 14056 10968 14832 10996
rect 14056 10956 14062 10968
rect 14826 10956 14832 10968
rect 14884 10956 14890 11008
rect 14927 10996 14955 11036
rect 16850 11024 16856 11076
rect 16908 11064 16914 11076
rect 16945 11067 17003 11073
rect 16945 11064 16957 11067
rect 16908 11036 16957 11064
rect 16908 11024 16914 11036
rect 16945 11033 16957 11036
rect 16991 11033 17003 11067
rect 17402 11064 17408 11076
rect 17363 11036 17408 11064
rect 16945 11027 17003 11033
rect 17402 11024 17408 11036
rect 17460 11024 17466 11076
rect 17770 11064 17776 11076
rect 17731 11036 17776 11064
rect 17770 11024 17776 11036
rect 17828 11024 17834 11076
rect 19426 11024 19432 11076
rect 19484 11064 19490 11076
rect 20254 11064 20260 11076
rect 19484 11036 20260 11064
rect 19484 11024 19490 11036
rect 20254 11024 20260 11036
rect 20312 11024 20318 11076
rect 20732 11073 20760 11104
rect 21358 11092 21364 11104
rect 21416 11092 21422 11144
rect 21453 11135 21511 11141
rect 21453 11101 21465 11135
rect 21499 11101 21511 11135
rect 21453 11095 21511 11101
rect 20717 11067 20775 11073
rect 20717 11033 20729 11067
rect 20763 11064 20775 11067
rect 21468 11064 21496 11095
rect 23474 11092 23480 11144
rect 23532 11132 23538 11144
rect 23569 11135 23627 11141
rect 23569 11132 23581 11135
rect 23532 11104 23581 11132
rect 23532 11092 23538 11104
rect 23569 11101 23581 11104
rect 23615 11101 23627 11135
rect 23569 11095 23627 11101
rect 20763 11036 21496 11064
rect 22649 11067 22707 11073
rect 20763 11033 20775 11036
rect 20717 11027 20775 11033
rect 22649 11033 22661 11067
rect 22695 11064 22707 11067
rect 23290 11064 23296 11076
rect 22695 11036 23296 11064
rect 22695 11033 22707 11036
rect 22649 11027 22707 11033
rect 23290 11024 23296 11036
rect 23348 11024 23354 11076
rect 18138 10996 18144 11008
rect 14927 10968 18144 10996
rect 18138 10956 18144 10968
rect 18196 10956 18202 11008
rect 19334 10996 19340 11008
rect 19295 10968 19340 10996
rect 19334 10956 19340 10968
rect 19392 10956 19398 11008
rect 23474 10996 23480 11008
rect 23435 10968 23480 10996
rect 23474 10956 23480 10968
rect 23532 10956 23538 11008
rect 25590 10996 25596 11008
rect 25551 10968 25596 10996
rect 25590 10956 25596 10968
rect 25648 10956 25654 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 2225 10795 2283 10801
rect 2225 10761 2237 10795
rect 2271 10792 2283 10795
rect 2590 10792 2596 10804
rect 2271 10764 2596 10792
rect 2271 10761 2283 10764
rect 2225 10755 2283 10761
rect 2590 10752 2596 10764
rect 2648 10752 2654 10804
rect 5350 10792 5356 10804
rect 2792 10764 5356 10792
rect 1026 10616 1032 10668
rect 1084 10656 1090 10668
rect 1578 10656 1584 10668
rect 1084 10628 1584 10656
rect 1084 10616 1090 10628
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 2792 10665 2820 10764
rect 5350 10752 5356 10764
rect 5408 10752 5414 10804
rect 5905 10795 5963 10801
rect 5905 10761 5917 10795
rect 5951 10792 5963 10795
rect 6638 10792 6644 10804
rect 5951 10764 6644 10792
rect 5951 10761 5963 10764
rect 5905 10755 5963 10761
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 8294 10792 8300 10804
rect 8255 10764 8300 10792
rect 8294 10752 8300 10764
rect 8352 10752 8358 10804
rect 10318 10792 10324 10804
rect 10279 10764 10324 10792
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 13722 10792 13728 10804
rect 13683 10764 13728 10792
rect 13722 10752 13728 10764
rect 13780 10752 13786 10804
rect 14093 10795 14151 10801
rect 14093 10761 14105 10795
rect 14139 10792 14151 10795
rect 16022 10792 16028 10804
rect 14139 10764 16028 10792
rect 14139 10761 14151 10764
rect 14093 10755 14151 10761
rect 5074 10684 5080 10736
rect 5132 10724 5138 10736
rect 5169 10727 5227 10733
rect 5169 10724 5181 10727
rect 5132 10696 5181 10724
rect 5132 10684 5138 10696
rect 5169 10693 5181 10696
rect 5215 10724 5227 10727
rect 5537 10727 5595 10733
rect 5537 10724 5549 10727
rect 5215 10696 5549 10724
rect 5215 10693 5227 10696
rect 5169 10687 5227 10693
rect 5537 10693 5549 10696
rect 5583 10724 5595 10727
rect 6270 10724 6276 10736
rect 5583 10696 6276 10724
rect 5583 10693 5595 10696
rect 5537 10687 5595 10693
rect 6270 10684 6276 10696
rect 6328 10684 6334 10736
rect 7374 10684 7380 10736
rect 7432 10724 7438 10736
rect 7742 10724 7748 10736
rect 7432 10696 7748 10724
rect 7432 10684 7438 10696
rect 7742 10684 7748 10696
rect 7800 10684 7806 10736
rect 11790 10724 11796 10736
rect 11751 10696 11796 10724
rect 11790 10684 11796 10696
rect 11848 10684 11854 10736
rect 13170 10684 13176 10736
rect 13228 10724 13234 10736
rect 14108 10724 14136 10755
rect 16022 10752 16028 10764
rect 16080 10752 16086 10804
rect 16298 10792 16304 10804
rect 16259 10764 16304 10792
rect 16298 10752 16304 10764
rect 16356 10792 16362 10804
rect 17497 10795 17555 10801
rect 16356 10764 16896 10792
rect 16356 10752 16362 10764
rect 14826 10724 14832 10736
rect 13228 10696 14136 10724
rect 14787 10696 14832 10724
rect 13228 10684 13234 10696
rect 14826 10684 14832 10696
rect 14884 10684 14890 10736
rect 15194 10684 15200 10736
rect 15252 10724 15258 10736
rect 15746 10724 15752 10736
rect 15252 10696 15752 10724
rect 15252 10684 15258 10696
rect 15746 10684 15752 10696
rect 15804 10684 15810 10736
rect 1765 10659 1823 10665
rect 1765 10625 1777 10659
rect 1811 10656 1823 10659
rect 2777 10659 2835 10665
rect 2777 10656 2789 10659
rect 1811 10628 2789 10656
rect 1811 10625 1823 10628
rect 1765 10619 1823 10625
rect 2777 10625 2789 10628
rect 2823 10625 2835 10659
rect 2777 10619 2835 10625
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10656 6699 10659
rect 7469 10659 7527 10665
rect 6687 10628 7236 10656
rect 6687 10625 6699 10628
rect 6641 10619 6699 10625
rect 7208 10600 7236 10628
rect 7469 10625 7481 10659
rect 7515 10656 7527 10659
rect 7558 10656 7564 10668
rect 7515 10628 7564 10656
rect 7515 10625 7527 10628
rect 7469 10619 7527 10625
rect 7558 10616 7564 10628
rect 7616 10616 7622 10668
rect 8846 10616 8852 10668
rect 8904 10656 8910 10668
rect 8941 10659 8999 10665
rect 8941 10656 8953 10659
rect 8904 10628 8953 10656
rect 8904 10616 8910 10628
rect 8941 10625 8953 10628
rect 8987 10625 8999 10659
rect 10594 10656 10600 10668
rect 10555 10628 10600 10656
rect 8941 10619 8999 10625
rect 10594 10616 10600 10628
rect 10652 10616 10658 10668
rect 11422 10616 11428 10668
rect 11480 10656 11486 10668
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 11480 10628 13001 10656
rect 11480 10616 11486 10628
rect 12989 10625 13001 10628
rect 13035 10625 13047 10659
rect 15286 10656 15292 10668
rect 15247 10628 15292 10656
rect 12989 10619 13047 10625
rect 15286 10616 15292 10628
rect 15344 10616 15350 10668
rect 16868 10665 16896 10764
rect 17497 10761 17509 10795
rect 17543 10792 17555 10795
rect 18230 10792 18236 10804
rect 17543 10764 18236 10792
rect 17543 10761 17555 10764
rect 17497 10755 17555 10761
rect 15473 10659 15531 10665
rect 15473 10625 15485 10659
rect 15519 10625 15531 10659
rect 15473 10619 15531 10625
rect 16853 10659 16911 10665
rect 16853 10625 16865 10659
rect 16899 10625 16911 10659
rect 17034 10656 17040 10668
rect 16947 10628 17040 10656
rect 16853 10619 16911 10625
rect 2593 10591 2651 10597
rect 2593 10557 2605 10591
rect 2639 10588 2651 10591
rect 2682 10588 2688 10600
rect 2639 10560 2688 10588
rect 2639 10557 2651 10560
rect 2593 10551 2651 10557
rect 2682 10548 2688 10560
rect 2740 10548 2746 10600
rect 3786 10588 3792 10600
rect 3747 10560 3792 10588
rect 3786 10548 3792 10560
rect 3844 10548 3850 10600
rect 6273 10591 6331 10597
rect 6273 10557 6285 10591
rect 6319 10588 6331 10591
rect 6822 10588 6828 10600
rect 6319 10560 6828 10588
rect 6319 10557 6331 10560
rect 6273 10551 6331 10557
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 7190 10588 7196 10600
rect 7151 10560 7196 10588
rect 7190 10548 7196 10560
rect 7248 10548 7254 10600
rect 8294 10548 8300 10600
rect 8352 10588 8358 10600
rect 8478 10588 8484 10600
rect 8352 10560 8484 10588
rect 8352 10548 8358 10560
rect 8478 10548 8484 10560
rect 8536 10588 8542 10600
rect 8573 10591 8631 10597
rect 8573 10588 8585 10591
rect 8536 10560 8585 10588
rect 8536 10548 8542 10560
rect 8573 10557 8585 10560
rect 8619 10557 8631 10591
rect 8573 10551 8631 10557
rect 9208 10591 9266 10597
rect 9208 10557 9220 10591
rect 9254 10588 9266 10591
rect 9490 10588 9496 10600
rect 9254 10560 9496 10588
rect 9254 10557 9266 10560
rect 9208 10551 9266 10557
rect 9490 10548 9496 10560
rect 9548 10548 9554 10600
rect 11146 10548 11152 10600
rect 11204 10588 11210 10600
rect 12253 10591 12311 10597
rect 12253 10588 12265 10591
rect 11204 10560 12265 10588
rect 11204 10548 11210 10560
rect 12253 10557 12265 10560
rect 12299 10588 12311 10591
rect 12897 10591 12955 10597
rect 12897 10588 12909 10591
rect 12299 10560 12909 10588
rect 12299 10557 12311 10560
rect 12253 10551 12311 10557
rect 12897 10557 12909 10560
rect 12943 10588 12955 10591
rect 14274 10588 14280 10600
rect 12943 10560 14280 10588
rect 12943 10557 12955 10560
rect 12897 10551 12955 10557
rect 14274 10548 14280 10560
rect 14332 10548 14338 10600
rect 15488 10588 15516 10619
rect 17034 10616 17040 10628
rect 17092 10656 17098 10668
rect 17512 10656 17540 10755
rect 18230 10752 18236 10764
rect 18288 10752 18294 10804
rect 18690 10752 18696 10804
rect 18748 10792 18754 10804
rect 18969 10795 19027 10801
rect 18969 10792 18981 10795
rect 18748 10764 18981 10792
rect 18748 10752 18754 10764
rect 18969 10761 18981 10764
rect 19015 10761 19027 10795
rect 18969 10755 19027 10761
rect 20714 10752 20720 10804
rect 20772 10792 20778 10804
rect 20901 10795 20959 10801
rect 20901 10792 20913 10795
rect 20772 10764 20913 10792
rect 20772 10752 20778 10764
rect 20901 10761 20913 10764
rect 20947 10761 20959 10795
rect 20901 10755 20959 10761
rect 21082 10752 21088 10804
rect 21140 10792 21146 10804
rect 21177 10795 21235 10801
rect 21177 10792 21189 10795
rect 21140 10764 21189 10792
rect 21140 10752 21146 10764
rect 21177 10761 21189 10764
rect 21223 10792 21235 10795
rect 23477 10795 23535 10801
rect 21223 10764 21680 10792
rect 21223 10761 21235 10764
rect 21177 10755 21235 10761
rect 17092 10628 17540 10656
rect 20732 10656 20760 10752
rect 20806 10684 20812 10736
rect 20864 10724 20870 10736
rect 21545 10727 21603 10733
rect 21545 10724 21557 10727
rect 20864 10696 21557 10724
rect 20864 10684 20870 10696
rect 21545 10693 21557 10696
rect 21591 10693 21603 10727
rect 21545 10687 21603 10693
rect 21082 10656 21088 10668
rect 20732 10628 21088 10656
rect 17092 10616 17098 10628
rect 21082 10616 21088 10628
rect 21140 10616 21146 10668
rect 17052 10588 17080 10616
rect 15488 10560 17080 10588
rect 17494 10548 17500 10600
rect 17552 10588 17558 10600
rect 17773 10591 17831 10597
rect 17773 10588 17785 10591
rect 17552 10560 17785 10588
rect 17552 10548 17558 10560
rect 17773 10557 17785 10560
rect 17819 10557 17831 10591
rect 17773 10551 17831 10557
rect 18417 10591 18475 10597
rect 18417 10557 18429 10591
rect 18463 10588 18475 10591
rect 18690 10588 18696 10600
rect 18463 10560 18696 10588
rect 18463 10557 18475 10560
rect 18417 10551 18475 10557
rect 18690 10548 18696 10560
rect 18748 10548 18754 10600
rect 19521 10591 19579 10597
rect 19521 10557 19533 10591
rect 19567 10588 19579 10591
rect 20254 10588 20260 10600
rect 19567 10560 20260 10588
rect 19567 10557 19579 10560
rect 19521 10551 19579 10557
rect 20254 10548 20260 10560
rect 20312 10548 20318 10600
rect 20806 10548 20812 10600
rect 20864 10588 20870 10600
rect 21450 10588 21456 10600
rect 20864 10560 21456 10588
rect 20864 10548 20870 10560
rect 21450 10548 21456 10560
rect 21508 10548 21514 10600
rect 21560 10588 21588 10687
rect 21652 10656 21680 10764
rect 23477 10761 23489 10795
rect 23523 10792 23535 10795
rect 23566 10792 23572 10804
rect 23523 10764 23572 10792
rect 23523 10761 23535 10764
rect 23477 10755 23535 10761
rect 23566 10752 23572 10764
rect 23624 10752 23630 10804
rect 23661 10795 23719 10801
rect 23661 10761 23673 10795
rect 23707 10792 23719 10795
rect 24210 10792 24216 10804
rect 23707 10764 24216 10792
rect 23707 10761 23719 10764
rect 23661 10755 23719 10761
rect 24210 10752 24216 10764
rect 24268 10752 24274 10804
rect 24670 10792 24676 10804
rect 24631 10764 24676 10792
rect 24670 10752 24676 10764
rect 24728 10792 24734 10804
rect 24854 10792 24860 10804
rect 24728 10764 24860 10792
rect 24728 10752 24734 10764
rect 24854 10752 24860 10764
rect 24912 10752 24918 10804
rect 25774 10752 25780 10804
rect 25832 10792 25838 10804
rect 25961 10795 26019 10801
rect 25961 10792 25973 10795
rect 25832 10764 25973 10792
rect 25832 10752 25838 10764
rect 25961 10761 25973 10764
rect 26007 10761 26019 10795
rect 25961 10755 26019 10761
rect 21729 10727 21787 10733
rect 21729 10693 21741 10727
rect 21775 10724 21787 10727
rect 22002 10724 22008 10736
rect 21775 10696 22008 10724
rect 21775 10693 21787 10696
rect 21729 10687 21787 10693
rect 22002 10684 22008 10696
rect 22060 10684 22066 10736
rect 22738 10724 22744 10736
rect 22699 10696 22744 10724
rect 22738 10684 22744 10696
rect 22796 10684 22802 10736
rect 22373 10659 22431 10665
rect 22373 10656 22385 10659
rect 21652 10628 22385 10656
rect 22373 10625 22385 10628
rect 22419 10656 22431 10659
rect 23290 10656 23296 10668
rect 22419 10628 23296 10656
rect 22419 10625 22431 10628
rect 22373 10619 22431 10625
rect 23290 10616 23296 10628
rect 23348 10616 23354 10668
rect 23584 10656 23612 10752
rect 24213 10659 24271 10665
rect 24213 10656 24225 10659
rect 23584 10628 24225 10656
rect 24213 10625 24225 10628
rect 24259 10625 24271 10659
rect 25406 10656 25412 10668
rect 25367 10628 25412 10656
rect 24213 10619 24271 10625
rect 25406 10616 25412 10628
rect 25464 10616 25470 10668
rect 22097 10591 22155 10597
rect 22097 10588 22109 10591
rect 21560 10560 22109 10588
rect 22097 10557 22109 10560
rect 22143 10557 22155 10591
rect 22097 10551 22155 10557
rect 23474 10548 23480 10600
rect 23532 10588 23538 10600
rect 24029 10591 24087 10597
rect 24029 10588 24041 10591
rect 23532 10560 24041 10588
rect 23532 10548 23538 10560
rect 24029 10557 24041 10560
rect 24075 10557 24087 10591
rect 24029 10551 24087 10557
rect 25225 10591 25283 10597
rect 25225 10557 25237 10591
rect 25271 10588 25283 10591
rect 25774 10588 25780 10600
rect 25271 10560 25780 10588
rect 25271 10557 25283 10560
rect 25225 10551 25283 10557
rect 25774 10548 25780 10560
rect 25832 10548 25838 10600
rect 4062 10529 4068 10532
rect 3697 10523 3755 10529
rect 3697 10489 3709 10523
rect 3743 10520 3755 10523
rect 4056 10520 4068 10529
rect 3743 10492 4068 10520
rect 3743 10489 3755 10492
rect 3697 10483 3755 10489
rect 4056 10483 4068 10492
rect 4062 10480 4068 10483
rect 4120 10480 4126 10532
rect 7285 10523 7343 10529
rect 7285 10489 7297 10523
rect 7331 10520 7343 10523
rect 7926 10520 7932 10532
rect 7331 10492 7932 10520
rect 7331 10489 7343 10492
rect 7285 10483 7343 10489
rect 7926 10480 7932 10492
rect 7984 10480 7990 10532
rect 12805 10523 12863 10529
rect 12805 10520 12817 10523
rect 11164 10492 12817 10520
rect 11164 10464 11192 10492
rect 12805 10489 12817 10492
rect 12851 10489 12863 10523
rect 12805 10483 12863 10489
rect 15562 10480 15568 10532
rect 15620 10520 15626 10532
rect 15746 10520 15752 10532
rect 15620 10492 15752 10520
rect 15620 10480 15626 10492
rect 15746 10480 15752 10492
rect 15804 10480 15810 10532
rect 16761 10523 16819 10529
rect 16761 10520 16773 10523
rect 15856 10492 16773 10520
rect 15856 10464 15884 10492
rect 16761 10489 16773 10492
rect 16807 10489 16819 10523
rect 19766 10523 19824 10529
rect 19766 10520 19778 10523
rect 16761 10483 16819 10489
rect 19352 10492 19778 10520
rect 19352 10464 19380 10492
rect 19766 10489 19778 10492
rect 19812 10489 19824 10523
rect 25041 10523 25099 10529
rect 25041 10520 25053 10523
rect 19766 10483 19824 10489
rect 24136 10492 25053 10520
rect 2133 10455 2191 10461
rect 2133 10421 2145 10455
rect 2179 10452 2191 10455
rect 2590 10452 2596 10464
rect 2179 10424 2596 10452
rect 2179 10421 2191 10424
rect 2133 10415 2191 10421
rect 2590 10412 2596 10424
rect 2648 10452 2654 10464
rect 2685 10455 2743 10461
rect 2685 10452 2697 10455
rect 2648 10424 2697 10452
rect 2648 10412 2654 10424
rect 2685 10421 2697 10424
rect 2731 10421 2743 10455
rect 3234 10452 3240 10464
rect 3195 10424 3240 10452
rect 2685 10415 2743 10421
rect 3234 10412 3240 10424
rect 3292 10412 3298 10464
rect 6822 10452 6828 10464
rect 6783 10424 6828 10452
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 8389 10455 8447 10461
rect 8389 10421 8401 10455
rect 8435 10452 8447 10455
rect 8478 10452 8484 10464
rect 8435 10424 8484 10452
rect 8435 10421 8447 10424
rect 8389 10415 8447 10421
rect 8478 10412 8484 10424
rect 8536 10412 8542 10464
rect 11146 10452 11152 10464
rect 11107 10424 11152 10452
rect 11146 10412 11152 10424
rect 11204 10412 11210 10464
rect 11330 10452 11336 10464
rect 11291 10424 11336 10452
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 12342 10412 12348 10464
rect 12400 10452 12406 10464
rect 12437 10455 12495 10461
rect 12437 10452 12449 10455
rect 12400 10424 12449 10452
rect 12400 10412 12406 10424
rect 12437 10421 12449 10424
rect 12483 10421 12495 10455
rect 14366 10452 14372 10464
rect 14327 10424 14372 10452
rect 12437 10415 12495 10421
rect 14366 10412 14372 10424
rect 14424 10412 14430 10464
rect 15194 10452 15200 10464
rect 15155 10424 15200 10452
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 15838 10452 15844 10464
rect 15799 10424 15844 10452
rect 15838 10412 15844 10424
rect 15896 10412 15902 10464
rect 16390 10452 16396 10464
rect 16351 10424 16396 10452
rect 16390 10412 16396 10424
rect 16448 10412 16454 10464
rect 16666 10412 16672 10464
rect 16724 10452 16730 10464
rect 16942 10452 16948 10464
rect 16724 10424 16948 10452
rect 16724 10412 16730 10424
rect 16942 10412 16948 10424
rect 17000 10412 17006 10464
rect 18601 10455 18659 10461
rect 18601 10421 18613 10455
rect 18647 10452 18659 10455
rect 18690 10452 18696 10464
rect 18647 10424 18696 10452
rect 18647 10421 18659 10424
rect 18601 10415 18659 10421
rect 18690 10412 18696 10424
rect 18748 10412 18754 10464
rect 19334 10452 19340 10464
rect 19295 10424 19340 10452
rect 19334 10412 19340 10424
rect 19392 10412 19398 10464
rect 22186 10452 22192 10464
rect 22147 10424 22192 10452
rect 22186 10412 22192 10424
rect 22244 10412 22250 10464
rect 24026 10412 24032 10464
rect 24084 10452 24090 10464
rect 24136 10461 24164 10492
rect 25041 10489 25053 10492
rect 25087 10489 25099 10523
rect 25041 10483 25099 10489
rect 24121 10455 24179 10461
rect 24121 10452 24133 10455
rect 24084 10424 24133 10452
rect 24084 10412 24090 10424
rect 24121 10421 24133 10424
rect 24167 10421 24179 10455
rect 24121 10415 24179 10421
rect 25590 10412 25596 10464
rect 25648 10452 25654 10464
rect 26329 10455 26387 10461
rect 26329 10452 26341 10455
rect 25648 10424 26341 10452
rect 25648 10412 25654 10424
rect 26329 10421 26341 10424
rect 26375 10421 26387 10455
rect 26329 10415 26387 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1673 10251 1731 10257
rect 1673 10217 1685 10251
rect 1719 10248 1731 10251
rect 1854 10248 1860 10260
rect 1719 10220 1860 10248
rect 1719 10217 1731 10220
rect 1673 10211 1731 10217
rect 1854 10208 1860 10220
rect 1912 10208 1918 10260
rect 2317 10251 2375 10257
rect 2317 10217 2329 10251
rect 2363 10248 2375 10251
rect 2682 10248 2688 10260
rect 2363 10220 2688 10248
rect 2363 10217 2375 10220
rect 2317 10211 2375 10217
rect 2682 10208 2688 10220
rect 2740 10208 2746 10260
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 3234 10248 3240 10260
rect 2832 10220 3240 10248
rect 2832 10208 2838 10220
rect 3234 10208 3240 10220
rect 3292 10208 3298 10260
rect 4617 10251 4675 10257
rect 4617 10217 4629 10251
rect 4663 10248 4675 10251
rect 4798 10248 4804 10260
rect 4663 10220 4804 10248
rect 4663 10217 4675 10220
rect 4617 10211 4675 10217
rect 4798 10208 4804 10220
rect 4856 10208 4862 10260
rect 4985 10251 5043 10257
rect 4985 10217 4997 10251
rect 5031 10248 5043 10251
rect 5166 10248 5172 10260
rect 5031 10220 5172 10248
rect 5031 10217 5043 10220
rect 4985 10211 5043 10217
rect 4525 10183 4583 10189
rect 4525 10149 4537 10183
rect 4571 10180 4583 10183
rect 5000 10180 5028 10211
rect 5166 10208 5172 10220
rect 5224 10208 5230 10260
rect 8294 10248 8300 10260
rect 8255 10220 8300 10248
rect 8294 10208 8300 10220
rect 8352 10208 8358 10260
rect 8389 10251 8447 10257
rect 8389 10217 8401 10251
rect 8435 10248 8447 10251
rect 9493 10251 9551 10257
rect 9493 10248 9505 10251
rect 8435 10220 9505 10248
rect 8435 10217 8447 10220
rect 8389 10211 8447 10217
rect 9493 10217 9505 10220
rect 9539 10248 9551 10251
rect 9674 10248 9680 10260
rect 9539 10220 9680 10248
rect 9539 10217 9551 10220
rect 9493 10211 9551 10217
rect 9674 10208 9680 10220
rect 9732 10208 9738 10260
rect 10042 10248 10048 10260
rect 10003 10220 10048 10248
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 10134 10208 10140 10260
rect 10192 10248 10198 10260
rect 10778 10248 10784 10260
rect 10192 10220 10784 10248
rect 10192 10208 10198 10220
rect 10778 10208 10784 10220
rect 10836 10208 10842 10260
rect 10873 10251 10931 10257
rect 10873 10217 10885 10251
rect 10919 10248 10931 10251
rect 10962 10248 10968 10260
rect 10919 10220 10968 10248
rect 10919 10217 10931 10220
rect 10873 10211 10931 10217
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 13630 10248 13636 10260
rect 13591 10220 13636 10248
rect 13630 10208 13636 10220
rect 13688 10208 13694 10260
rect 13906 10248 13912 10260
rect 13867 10220 13912 10248
rect 13906 10208 13912 10220
rect 13964 10208 13970 10260
rect 15194 10208 15200 10260
rect 15252 10248 15258 10260
rect 17221 10251 17279 10257
rect 17221 10248 17233 10251
rect 15252 10220 17233 10248
rect 15252 10208 15258 10220
rect 17221 10217 17233 10220
rect 17267 10248 17279 10251
rect 17773 10251 17831 10257
rect 17773 10248 17785 10251
rect 17267 10220 17785 10248
rect 17267 10217 17279 10220
rect 17221 10211 17279 10217
rect 17773 10217 17785 10220
rect 17819 10217 17831 10251
rect 17773 10211 17831 10217
rect 18046 10208 18052 10260
rect 18104 10248 18110 10260
rect 18233 10251 18291 10257
rect 18233 10248 18245 10251
rect 18104 10220 18245 10248
rect 18104 10208 18110 10220
rect 18233 10217 18245 10220
rect 18279 10217 18291 10251
rect 19150 10248 19156 10260
rect 19111 10220 19156 10248
rect 18233 10211 18291 10217
rect 19150 10208 19156 10220
rect 19208 10208 19214 10260
rect 20901 10251 20959 10257
rect 20901 10217 20913 10251
rect 20947 10248 20959 10251
rect 21358 10248 21364 10260
rect 20947 10220 21364 10248
rect 20947 10217 20959 10220
rect 20901 10211 20959 10217
rect 21358 10208 21364 10220
rect 21416 10208 21422 10260
rect 22465 10251 22523 10257
rect 22465 10217 22477 10251
rect 22511 10248 22523 10251
rect 22738 10248 22744 10260
rect 22511 10220 22744 10248
rect 22511 10217 22523 10220
rect 22465 10211 22523 10217
rect 22738 10208 22744 10220
rect 22796 10208 22802 10260
rect 22833 10251 22891 10257
rect 22833 10217 22845 10251
rect 22879 10248 22891 10251
rect 23014 10248 23020 10260
rect 22879 10220 23020 10248
rect 22879 10217 22891 10220
rect 22833 10211 22891 10217
rect 23014 10208 23020 10220
rect 23072 10248 23078 10260
rect 24854 10248 24860 10260
rect 23072 10220 24348 10248
rect 24815 10220 24860 10248
rect 23072 10208 23078 10220
rect 4571 10152 5028 10180
rect 4571 10149 4583 10152
rect 4525 10143 4583 10149
rect 6178 10140 6184 10192
rect 6236 10180 6242 10192
rect 6426 10183 6484 10189
rect 6426 10180 6438 10183
rect 6236 10152 6438 10180
rect 6236 10140 6242 10152
rect 6426 10149 6438 10152
rect 6472 10149 6484 10183
rect 11698 10180 11704 10192
rect 11659 10152 11704 10180
rect 6426 10143 6484 10149
rect 11698 10140 11704 10152
rect 11756 10140 11762 10192
rect 15565 10183 15623 10189
rect 15565 10149 15577 10183
rect 15611 10180 15623 10183
rect 15654 10180 15660 10192
rect 15611 10152 15660 10180
rect 15611 10149 15623 10152
rect 15565 10143 15623 10149
rect 15654 10140 15660 10152
rect 15712 10140 15718 10192
rect 16574 10180 16580 10192
rect 16487 10152 16580 10180
rect 16574 10140 16580 10152
rect 16632 10180 16638 10192
rect 16758 10180 16764 10192
rect 16632 10152 16764 10180
rect 16632 10140 16638 10152
rect 16758 10140 16764 10152
rect 16816 10140 16822 10192
rect 18141 10183 18199 10189
rect 18141 10149 18153 10183
rect 18187 10180 18199 10183
rect 18322 10180 18328 10192
rect 18187 10152 18328 10180
rect 18187 10149 18199 10152
rect 18141 10143 18199 10149
rect 18322 10140 18328 10152
rect 18380 10140 18386 10192
rect 20717 10183 20775 10189
rect 20717 10149 20729 10183
rect 20763 10180 20775 10183
rect 21269 10183 21327 10189
rect 21269 10180 21281 10183
rect 20763 10152 21281 10180
rect 20763 10149 20775 10152
rect 20717 10143 20775 10149
rect 21269 10149 21281 10152
rect 21315 10180 21327 10183
rect 23744 10183 23802 10189
rect 21315 10152 22508 10180
rect 21315 10149 21327 10152
rect 21269 10143 21327 10149
rect 22480 10124 22508 10152
rect 23744 10149 23756 10183
rect 23790 10180 23802 10183
rect 24210 10180 24216 10192
rect 23790 10152 24216 10180
rect 23790 10149 23802 10152
rect 23744 10143 23802 10149
rect 24210 10140 24216 10152
rect 24268 10140 24274 10192
rect 24320 10180 24348 10220
rect 24854 10208 24860 10220
rect 24912 10208 24918 10260
rect 26050 10180 26056 10192
rect 24320 10152 26056 10180
rect 26050 10140 26056 10152
rect 26108 10140 26114 10192
rect 2498 10072 2504 10124
rect 2556 10112 2562 10124
rect 2682 10112 2688 10124
rect 2556 10084 2688 10112
rect 2556 10072 2562 10084
rect 2682 10072 2688 10084
rect 2740 10072 2746 10124
rect 2869 10115 2927 10121
rect 2869 10112 2881 10115
rect 2792 10084 2881 10112
rect 2792 10044 2820 10084
rect 2869 10081 2881 10084
rect 2915 10112 2927 10115
rect 3421 10115 3479 10121
rect 3421 10112 3433 10115
rect 2915 10084 3433 10112
rect 2915 10081 2927 10084
rect 2869 10075 2927 10081
rect 3421 10081 3433 10084
rect 3467 10081 3479 10115
rect 3421 10075 3479 10081
rect 5077 10115 5135 10121
rect 5077 10081 5089 10115
rect 5123 10112 5135 10115
rect 5442 10112 5448 10124
rect 5123 10084 5448 10112
rect 5123 10081 5135 10084
rect 5077 10075 5135 10081
rect 5442 10072 5448 10084
rect 5500 10072 5506 10124
rect 5721 10115 5779 10121
rect 5721 10081 5733 10115
rect 5767 10112 5779 10115
rect 6086 10112 6092 10124
rect 5767 10084 6092 10112
rect 5767 10081 5779 10084
rect 5721 10075 5779 10081
rect 6086 10072 6092 10084
rect 6144 10112 6150 10124
rect 6270 10112 6276 10124
rect 6144 10084 6276 10112
rect 6144 10072 6150 10084
rect 6270 10072 6276 10084
rect 6328 10072 6334 10124
rect 9033 10115 9091 10121
rect 9033 10081 9045 10115
rect 9079 10112 9091 10115
rect 9490 10112 9496 10124
rect 9079 10084 9496 10112
rect 9079 10081 9091 10084
rect 9033 10075 9091 10081
rect 9490 10072 9496 10084
rect 9548 10072 9554 10124
rect 12158 10121 12164 10124
rect 12152 10112 12164 10121
rect 12119 10084 12164 10112
rect 12152 10075 12164 10084
rect 12158 10072 12164 10075
rect 12216 10072 12222 10124
rect 14093 10115 14151 10121
rect 14093 10081 14105 10115
rect 14139 10112 14151 10115
rect 14274 10112 14280 10124
rect 14139 10084 14280 10112
rect 14139 10081 14151 10084
rect 14093 10075 14151 10081
rect 14274 10072 14280 10084
rect 14332 10112 14338 10124
rect 14642 10112 14648 10124
rect 14332 10084 14648 10112
rect 14332 10072 14338 10084
rect 14642 10072 14648 10084
rect 14700 10072 14706 10124
rect 16669 10115 16727 10121
rect 16669 10081 16681 10115
rect 16715 10112 16727 10115
rect 17129 10115 17187 10121
rect 17129 10112 17141 10115
rect 16715 10084 17141 10112
rect 16715 10081 16727 10084
rect 16669 10075 16727 10081
rect 17129 10081 17141 10084
rect 17175 10112 17187 10115
rect 17589 10115 17647 10121
rect 17589 10112 17601 10115
rect 17175 10084 17601 10112
rect 17175 10081 17187 10084
rect 17129 10075 17187 10081
rect 17589 10081 17601 10084
rect 17635 10081 17647 10115
rect 17589 10075 17647 10081
rect 17770 10072 17776 10124
rect 17828 10112 17834 10124
rect 19518 10112 19524 10124
rect 17828 10084 18460 10112
rect 19479 10084 19524 10112
rect 17828 10072 17834 10084
rect 2958 10044 2964 10056
rect 2700 10016 2820 10044
rect 2919 10016 2964 10044
rect 2406 9976 2412 9988
rect 2367 9948 2412 9976
rect 2406 9936 2412 9948
rect 2464 9936 2470 9988
rect 2700 9920 2728 10016
rect 2958 10004 2964 10016
rect 3016 10004 3022 10056
rect 5261 10047 5319 10053
rect 5261 10013 5273 10047
rect 5307 10013 5319 10047
rect 5261 10007 5319 10013
rect 5537 10047 5595 10053
rect 5537 10013 5549 10047
rect 5583 10044 5595 10047
rect 5994 10044 6000 10056
rect 5583 10016 6000 10044
rect 5583 10013 5595 10016
rect 5537 10007 5595 10013
rect 4798 9936 4804 9988
rect 4856 9976 4862 9988
rect 5276 9976 5304 10007
rect 5994 10004 6000 10016
rect 6052 10044 6058 10056
rect 6181 10047 6239 10053
rect 6181 10044 6193 10047
rect 6052 10016 6193 10044
rect 6052 10004 6058 10016
rect 6181 10013 6193 10016
rect 6227 10013 6239 10047
rect 10226 10044 10232 10056
rect 10187 10016 10232 10044
rect 6181 10007 6239 10013
rect 10226 10004 10232 10016
rect 10284 10004 10290 10056
rect 11882 10044 11888 10056
rect 11843 10016 11888 10044
rect 11882 10004 11888 10016
rect 11940 10004 11946 10056
rect 14921 10047 14979 10053
rect 14921 10013 14933 10047
rect 14967 10044 14979 10047
rect 16117 10047 16175 10053
rect 16117 10044 16129 10047
rect 14967 10016 16129 10044
rect 14967 10013 14979 10016
rect 14921 10007 14979 10013
rect 16117 10013 16129 10016
rect 16163 10044 16175 10047
rect 16853 10047 16911 10053
rect 16853 10044 16865 10047
rect 16163 10016 16865 10044
rect 16163 10013 16175 10016
rect 16117 10007 16175 10013
rect 16853 10013 16865 10016
rect 16899 10044 16911 10047
rect 17034 10044 17040 10056
rect 16899 10016 17040 10044
rect 16899 10013 16911 10016
rect 16853 10007 16911 10013
rect 17034 10004 17040 10016
rect 17092 10004 17098 10056
rect 18432 10053 18460 10084
rect 19518 10072 19524 10084
rect 19576 10072 19582 10124
rect 19610 10072 19616 10124
rect 19668 10112 19674 10124
rect 19705 10115 19763 10121
rect 19705 10112 19717 10115
rect 19668 10084 19717 10112
rect 19668 10072 19674 10084
rect 19705 10081 19717 10084
rect 19751 10081 19763 10115
rect 19705 10075 19763 10081
rect 20349 10115 20407 10121
rect 20349 10081 20361 10115
rect 20395 10112 20407 10115
rect 20622 10112 20628 10124
rect 20395 10084 20628 10112
rect 20395 10081 20407 10084
rect 20349 10075 20407 10081
rect 18417 10047 18475 10053
rect 18417 10013 18429 10047
rect 18463 10044 18475 10047
rect 20364 10044 20392 10075
rect 20622 10072 20628 10084
rect 20680 10112 20686 10124
rect 20680 10084 21588 10112
rect 20680 10072 20686 10084
rect 21560 10053 21588 10084
rect 22462 10072 22468 10124
rect 22520 10072 22526 10124
rect 22738 10072 22744 10124
rect 22796 10112 22802 10124
rect 23198 10112 23204 10124
rect 22796 10084 23204 10112
rect 22796 10072 22802 10084
rect 23198 10072 23204 10084
rect 23256 10072 23262 10124
rect 23566 10072 23572 10124
rect 23624 10072 23630 10124
rect 18463 10016 20392 10044
rect 21361 10047 21419 10053
rect 18463 10013 18475 10016
rect 18417 10007 18475 10013
rect 21361 10013 21373 10047
rect 21407 10013 21419 10047
rect 21361 10007 21419 10013
rect 21545 10047 21603 10053
rect 21545 10013 21557 10047
rect 21591 10044 21603 10047
rect 21913 10047 21971 10053
rect 21913 10044 21925 10047
rect 21591 10016 21925 10044
rect 21591 10013 21603 10016
rect 21545 10007 21603 10013
rect 21913 10013 21925 10016
rect 21959 10013 21971 10047
rect 22756 10044 22784 10072
rect 21913 10007 21971 10013
rect 22020 10016 22784 10044
rect 13265 9979 13323 9985
rect 4856 9948 6132 9976
rect 4856 9936 4862 9948
rect 6104 9920 6132 9948
rect 13265 9945 13277 9979
rect 13311 9976 13323 9979
rect 13538 9976 13544 9988
rect 13311 9948 13544 9976
rect 13311 9945 13323 9948
rect 13265 9939 13323 9945
rect 13538 9936 13544 9948
rect 13596 9936 13602 9988
rect 16209 9979 16267 9985
rect 16209 9945 16221 9979
rect 16255 9976 16267 9979
rect 18785 9979 18843 9985
rect 18785 9976 18797 9979
rect 16255 9948 18797 9976
rect 16255 9945 16267 9948
rect 16209 9939 16267 9945
rect 18785 9945 18797 9948
rect 18831 9976 18843 9979
rect 18966 9976 18972 9988
rect 18831 9948 18972 9976
rect 18831 9945 18843 9948
rect 18785 9939 18843 9945
rect 18966 9936 18972 9948
rect 19024 9936 19030 9988
rect 19889 9979 19947 9985
rect 19889 9945 19901 9979
rect 19935 9976 19947 9979
rect 20438 9976 20444 9988
rect 19935 9948 20444 9976
rect 19935 9945 19947 9948
rect 19889 9939 19947 9945
rect 20438 9936 20444 9948
rect 20496 9936 20502 9988
rect 21376 9976 21404 10007
rect 22020 9976 22048 10016
rect 23014 10004 23020 10056
rect 23072 10044 23078 10056
rect 23293 10047 23351 10053
rect 23293 10044 23305 10047
rect 23072 10016 23305 10044
rect 23072 10004 23078 10016
rect 23293 10013 23305 10016
rect 23339 10013 23351 10047
rect 23293 10007 23351 10013
rect 23477 10047 23535 10053
rect 23477 10013 23489 10047
rect 23523 10044 23535 10047
rect 23584 10044 23612 10072
rect 23523 10016 23612 10044
rect 23523 10013 23535 10016
rect 23477 10007 23535 10013
rect 21376 9948 22048 9976
rect 22186 9936 22192 9988
rect 22244 9976 22250 9988
rect 22373 9979 22431 9985
rect 22373 9976 22385 9979
rect 22244 9948 22385 9976
rect 22244 9936 22250 9948
rect 22373 9945 22385 9948
rect 22419 9976 22431 9979
rect 23382 9976 23388 9988
rect 22419 9948 23388 9976
rect 22419 9945 22431 9948
rect 22373 9939 22431 9945
rect 23382 9936 23388 9948
rect 23440 9936 23446 9988
rect 25130 9976 25136 9988
rect 25091 9948 25136 9976
rect 25130 9936 25136 9948
rect 25188 9976 25194 9988
rect 25501 9979 25559 9985
rect 25501 9976 25513 9979
rect 25188 9948 25513 9976
rect 25188 9936 25194 9948
rect 25501 9945 25513 9948
rect 25547 9976 25559 9979
rect 26234 9976 26240 9988
rect 25547 9948 26240 9976
rect 25547 9945 25559 9948
rect 25501 9939 25559 9945
rect 26234 9936 26240 9948
rect 26292 9936 26298 9988
rect 2682 9868 2688 9920
rect 2740 9868 2746 9920
rect 3786 9868 3792 9920
rect 3844 9908 3850 9920
rect 3881 9911 3939 9917
rect 3881 9908 3893 9911
rect 3844 9880 3893 9908
rect 3844 9868 3850 9880
rect 3881 9877 3893 9880
rect 3927 9908 3939 9911
rect 5537 9911 5595 9917
rect 5537 9908 5549 9911
rect 3927 9880 5549 9908
rect 3927 9877 3939 9880
rect 3881 9871 3939 9877
rect 5537 9877 5549 9880
rect 5583 9877 5595 9911
rect 5994 9908 6000 9920
rect 5955 9880 6000 9908
rect 5537 9871 5595 9877
rect 5994 9868 6000 9880
rect 6052 9868 6058 9920
rect 6086 9868 6092 9920
rect 6144 9908 6150 9920
rect 7561 9911 7619 9917
rect 7561 9908 7573 9911
rect 6144 9880 7573 9908
rect 6144 9868 6150 9880
rect 7561 9877 7573 9880
rect 7607 9877 7619 9911
rect 7561 9871 7619 9877
rect 7929 9911 7987 9917
rect 7929 9877 7941 9911
rect 7975 9908 7987 9911
rect 8018 9908 8024 9920
rect 7975 9880 8024 9908
rect 7975 9877 7987 9880
rect 7929 9871 7987 9877
rect 8018 9868 8024 9880
rect 8076 9868 8082 9920
rect 9674 9908 9680 9920
rect 9635 9880 9680 9908
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 11422 9908 11428 9920
rect 11383 9880 11428 9908
rect 11422 9868 11428 9880
rect 11480 9868 11486 9920
rect 14277 9911 14335 9917
rect 14277 9877 14289 9911
rect 14323 9908 14335 9911
rect 14458 9908 14464 9920
rect 14323 9880 14464 9908
rect 14323 9877 14335 9880
rect 14277 9871 14335 9877
rect 14458 9868 14464 9880
rect 14516 9868 14522 9920
rect 16666 9868 16672 9920
rect 16724 9908 16730 9920
rect 17129 9911 17187 9917
rect 17129 9908 17141 9911
rect 16724 9880 17141 9908
rect 16724 9868 16730 9880
rect 17129 9877 17141 9880
rect 17175 9877 17187 9911
rect 17129 9871 17187 9877
rect 19337 9911 19395 9917
rect 19337 9877 19349 9911
rect 19383 9908 19395 9911
rect 19978 9908 19984 9920
rect 19383 9880 19984 9908
rect 19383 9877 19395 9880
rect 19337 9871 19395 9877
rect 19978 9868 19984 9880
rect 20036 9868 20042 9920
rect 20898 9868 20904 9920
rect 20956 9908 20962 9920
rect 22833 9911 22891 9917
rect 22833 9908 22845 9911
rect 20956 9880 22845 9908
rect 20956 9868 20962 9880
rect 22833 9877 22845 9880
rect 22879 9877 22891 9911
rect 23014 9908 23020 9920
rect 22975 9880 23020 9908
rect 22833 9871 22891 9877
rect 23014 9868 23020 9880
rect 23072 9868 23078 9920
rect 25590 9868 25596 9920
rect 25648 9908 25654 9920
rect 25869 9911 25927 9917
rect 25869 9908 25881 9911
rect 25648 9880 25881 9908
rect 25648 9868 25654 9880
rect 25869 9877 25881 9880
rect 25915 9877 25927 9911
rect 25869 9871 25927 9877
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 937 9707 995 9713
rect 937 9673 949 9707
rect 983 9704 995 9707
rect 4709 9707 4767 9713
rect 983 9676 2084 9704
rect 983 9673 995 9676
rect 937 9667 995 9673
rect 1578 9636 1584 9648
rect 1539 9608 1584 9636
rect 1578 9596 1584 9608
rect 1636 9596 1642 9648
rect 1854 9596 1860 9648
rect 1912 9636 1918 9648
rect 2056 9636 2084 9676
rect 4709 9673 4721 9707
rect 4755 9704 4767 9707
rect 4798 9704 4804 9716
rect 4755 9676 4804 9704
rect 4755 9673 4767 9676
rect 4709 9667 4767 9673
rect 4798 9664 4804 9676
rect 4856 9664 4862 9716
rect 6178 9704 6184 9716
rect 6139 9676 6184 9704
rect 6178 9664 6184 9676
rect 6236 9704 6242 9716
rect 10042 9704 10048 9716
rect 6236 9676 8432 9704
rect 6236 9664 6242 9676
rect 4982 9636 4988 9648
rect 1912 9608 2084 9636
rect 4943 9608 4988 9636
rect 1912 9596 1918 9608
rect 4982 9596 4988 9608
rect 5040 9636 5046 9648
rect 8404 9636 8432 9676
rect 9600 9676 10048 9704
rect 8849 9639 8907 9645
rect 8849 9636 8861 9639
rect 5040 9608 5672 9636
rect 8404 9608 8861 9636
rect 5040 9596 5046 9608
rect 5644 9577 5672 9608
rect 8849 9605 8861 9608
rect 8895 9605 8907 9639
rect 8849 9599 8907 9605
rect 9309 9639 9367 9645
rect 9309 9605 9321 9639
rect 9355 9636 9367 9639
rect 9600 9636 9628 9676
rect 10042 9664 10048 9676
rect 10100 9664 10106 9716
rect 11146 9704 11152 9716
rect 10612 9676 11152 9704
rect 9355 9608 9628 9636
rect 9677 9639 9735 9645
rect 9355 9605 9367 9608
rect 9309 9599 9367 9605
rect 9677 9605 9689 9639
rect 9723 9636 9735 9639
rect 10134 9636 10140 9648
rect 9723 9608 10140 9636
rect 9723 9605 9735 9608
rect 9677 9599 9735 9605
rect 5629 9571 5687 9577
rect 5629 9537 5641 9571
rect 5675 9537 5687 9571
rect 5629 9531 5687 9537
rect 5813 9571 5871 9577
rect 5813 9537 5825 9571
rect 5859 9568 5871 9571
rect 6270 9568 6276 9580
rect 5859 9540 6276 9568
rect 5859 9537 5871 9540
rect 5813 9531 5871 9537
rect 6270 9528 6276 9540
rect 6328 9528 6334 9580
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 1670 9500 1676 9512
rect 1443 9472 1676 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1670 9460 1676 9472
rect 1728 9460 1734 9512
rect 2406 9460 2412 9512
rect 2464 9500 2470 9512
rect 2685 9503 2743 9509
rect 2685 9500 2697 9503
rect 2464 9472 2697 9500
rect 2464 9460 2470 9472
rect 2685 9469 2697 9472
rect 2731 9500 2743 9503
rect 3786 9500 3792 9512
rect 2731 9472 3792 9500
rect 2731 9469 2743 9472
rect 2685 9463 2743 9469
rect 3786 9460 3792 9472
rect 3844 9460 3850 9512
rect 5994 9460 6000 9512
rect 6052 9500 6058 9512
rect 6641 9503 6699 9509
rect 6641 9500 6653 9503
rect 6052 9472 6653 9500
rect 6052 9460 6058 9472
rect 6641 9469 6653 9472
rect 6687 9500 6699 9503
rect 7469 9503 7527 9509
rect 7469 9500 7481 9503
rect 6687 9472 7481 9500
rect 6687 9469 6699 9472
rect 6641 9463 6699 9469
rect 7469 9469 7481 9472
rect 7515 9500 7527 9503
rect 8018 9500 8024 9512
rect 7515 9472 8024 9500
rect 7515 9469 7527 9472
rect 7469 9463 7527 9469
rect 8018 9460 8024 9472
rect 8076 9460 8082 9512
rect 8864 9500 8892 9599
rect 10134 9596 10140 9608
rect 10192 9596 10198 9648
rect 9769 9571 9827 9577
rect 9769 9537 9781 9571
rect 9815 9568 9827 9571
rect 10612 9568 10640 9676
rect 11146 9664 11152 9676
rect 11204 9664 11210 9716
rect 12434 9664 12440 9716
rect 12492 9664 12498 9716
rect 14093 9707 14151 9713
rect 14093 9673 14105 9707
rect 14139 9704 14151 9707
rect 14274 9704 14280 9716
rect 14139 9676 14280 9704
rect 14139 9673 14151 9676
rect 14093 9667 14151 9673
rect 14274 9664 14280 9676
rect 14332 9664 14338 9716
rect 16666 9704 16672 9716
rect 16592 9676 16672 9704
rect 10689 9639 10747 9645
rect 10689 9605 10701 9639
rect 10735 9636 10747 9639
rect 10735 9608 11468 9636
rect 10735 9605 10747 9608
rect 10689 9599 10747 9605
rect 9815 9540 10640 9568
rect 9815 9537 9827 9540
rect 9769 9531 9827 9537
rect 11054 9528 11060 9580
rect 11112 9568 11118 9580
rect 11440 9577 11468 9608
rect 11241 9571 11299 9577
rect 11241 9568 11253 9571
rect 11112 9540 11253 9568
rect 11112 9528 11118 9540
rect 11241 9537 11253 9540
rect 11287 9537 11299 9571
rect 11241 9531 11299 9537
rect 11425 9571 11483 9577
rect 11425 9537 11437 9571
rect 11471 9568 11483 9571
rect 11790 9568 11796 9580
rect 11471 9540 11796 9568
rect 11471 9537 11483 9540
rect 11425 9531 11483 9537
rect 11790 9528 11796 9540
rect 11848 9528 11854 9580
rect 12452 9577 12480 9664
rect 14182 9596 14188 9648
rect 14240 9636 14246 9648
rect 14461 9639 14519 9645
rect 14461 9636 14473 9639
rect 14240 9608 14473 9636
rect 14240 9596 14246 9608
rect 14461 9605 14473 9608
rect 14507 9605 14519 9639
rect 14461 9599 14519 9605
rect 14645 9639 14703 9645
rect 14645 9605 14657 9639
rect 14691 9636 14703 9639
rect 14734 9636 14740 9648
rect 14691 9608 14740 9636
rect 14691 9605 14703 9608
rect 14645 9599 14703 9605
rect 12437 9571 12495 9577
rect 12437 9537 12449 9571
rect 12483 9537 12495 9571
rect 12437 9531 12495 9537
rect 10226 9500 10232 9512
rect 8864 9472 10232 9500
rect 10226 9460 10232 9472
rect 10284 9460 10290 9512
rect 2958 9441 2964 9444
rect 2952 9432 2964 9441
rect 2871 9404 2964 9432
rect 2952 9395 2964 9404
rect 2958 9392 2964 9395
rect 3016 9392 3022 9444
rect 4522 9392 4528 9444
rect 4580 9432 4586 9444
rect 6546 9432 6552 9444
rect 4580 9404 6552 9432
rect 4580 9392 4586 9404
rect 6546 9392 6552 9404
rect 6604 9392 6610 9444
rect 7377 9435 7435 9441
rect 7377 9401 7389 9435
rect 7423 9432 7435 9435
rect 7714 9435 7772 9441
rect 7714 9432 7726 9435
rect 7423 9404 7726 9432
rect 7423 9401 7435 9404
rect 7377 9395 7435 9401
rect 7714 9401 7726 9404
rect 7760 9432 7772 9435
rect 8110 9432 8116 9444
rect 7760 9404 8116 9432
rect 7760 9401 7772 9404
rect 7714 9395 7772 9401
rect 8110 9392 8116 9404
rect 8168 9392 8174 9444
rect 11146 9432 11152 9444
rect 11059 9404 11152 9432
rect 11146 9392 11152 9404
rect 11204 9432 11210 9444
rect 12342 9432 12348 9444
rect 11204 9404 12348 9432
rect 11204 9392 11210 9404
rect 12342 9392 12348 9404
rect 12400 9392 12406 9444
rect 12710 9441 12716 9444
rect 12704 9432 12716 9441
rect 12671 9404 12716 9432
rect 12704 9395 12716 9404
rect 12710 9392 12716 9395
rect 12768 9392 12774 9444
rect 14476 9432 14504 9599
rect 14734 9596 14740 9608
rect 14792 9596 14798 9648
rect 16393 9639 16451 9645
rect 16393 9605 16405 9639
rect 16439 9636 16451 9639
rect 16592 9636 16620 9676
rect 16666 9664 16672 9676
rect 16724 9664 16730 9716
rect 18046 9704 18052 9716
rect 17880 9676 18052 9704
rect 17497 9639 17555 9645
rect 17497 9636 17509 9639
rect 16439 9608 16620 9636
rect 17052 9608 17509 9636
rect 16439 9605 16451 9608
rect 16393 9599 16451 9605
rect 15197 9571 15255 9577
rect 15197 9568 15209 9571
rect 14660 9540 15209 9568
rect 14660 9512 14688 9540
rect 15197 9537 15209 9540
rect 15243 9537 15255 9571
rect 15197 9531 15255 9537
rect 16301 9571 16359 9577
rect 16301 9537 16313 9571
rect 16347 9568 16359 9571
rect 16482 9568 16488 9580
rect 16347 9540 16488 9568
rect 16347 9537 16359 9540
rect 16301 9531 16359 9537
rect 16482 9528 16488 9540
rect 16540 9528 16546 9580
rect 16850 9528 16856 9580
rect 16908 9568 16914 9580
rect 17052 9577 17080 9608
rect 17497 9605 17509 9608
rect 17543 9636 17555 9639
rect 17770 9636 17776 9648
rect 17543 9608 17776 9636
rect 17543 9605 17555 9608
rect 17497 9599 17555 9605
rect 17770 9596 17776 9608
rect 17828 9596 17834 9648
rect 17880 9645 17908 9676
rect 18046 9664 18052 9676
rect 18104 9664 18110 9716
rect 18322 9704 18328 9716
rect 18283 9676 18328 9704
rect 18322 9664 18328 9676
rect 18380 9664 18386 9716
rect 21174 9664 21180 9716
rect 21232 9704 21238 9716
rect 21637 9707 21695 9713
rect 21637 9704 21649 9707
rect 21232 9676 21649 9704
rect 21232 9664 21238 9676
rect 21637 9673 21649 9676
rect 21683 9673 21695 9707
rect 22738 9704 22744 9716
rect 22699 9676 22744 9704
rect 21637 9667 21695 9673
rect 22738 9664 22744 9676
rect 22796 9664 22802 9716
rect 23477 9707 23535 9713
rect 23477 9673 23489 9707
rect 23523 9704 23535 9707
rect 24946 9704 24952 9716
rect 23523 9676 24952 9704
rect 23523 9673 23535 9676
rect 23477 9667 23535 9673
rect 24946 9664 24952 9676
rect 25004 9704 25010 9716
rect 25041 9707 25099 9713
rect 25041 9704 25053 9707
rect 25004 9676 25053 9704
rect 25004 9664 25010 9676
rect 25041 9673 25053 9676
rect 25087 9673 25099 9707
rect 25041 9667 25099 9673
rect 17865 9639 17923 9645
rect 17865 9605 17877 9639
rect 17911 9605 17923 9639
rect 17865 9599 17923 9605
rect 18509 9639 18567 9645
rect 18509 9605 18521 9639
rect 18555 9636 18567 9639
rect 19426 9636 19432 9648
rect 18555 9608 19432 9636
rect 18555 9605 18567 9608
rect 18509 9599 18567 9605
rect 19426 9596 19432 9608
rect 19484 9596 19490 9648
rect 20070 9636 20076 9648
rect 20031 9608 20076 9636
rect 20070 9596 20076 9608
rect 20128 9596 20134 9648
rect 21818 9596 21824 9648
rect 21876 9636 21882 9648
rect 21910 9636 21916 9648
rect 21876 9608 21916 9636
rect 21876 9596 21882 9608
rect 21910 9596 21916 9608
rect 21968 9596 21974 9648
rect 22278 9636 22284 9648
rect 22195 9608 22284 9636
rect 17037 9571 17095 9577
rect 17037 9568 17049 9571
rect 16908 9540 17049 9568
rect 16908 9528 16914 9540
rect 17037 9537 17049 9540
rect 17083 9537 17095 9571
rect 18966 9568 18972 9580
rect 18927 9540 18972 9568
rect 17037 9531 17095 9537
rect 18966 9528 18972 9540
rect 19024 9528 19030 9580
rect 19061 9571 19119 9577
rect 19061 9537 19073 9571
rect 19107 9568 19119 9571
rect 19242 9568 19248 9580
rect 19107 9540 19248 9568
rect 19107 9537 19119 9540
rect 19061 9531 19119 9537
rect 14642 9460 14648 9512
rect 14700 9460 14706 9512
rect 15102 9500 15108 9512
rect 15063 9472 15108 9500
rect 15102 9460 15108 9472
rect 15160 9460 15166 9512
rect 16206 9460 16212 9512
rect 16264 9500 16270 9512
rect 18322 9500 18328 9512
rect 16264 9472 18328 9500
rect 16264 9460 16270 9472
rect 18322 9460 18328 9472
rect 18380 9460 18386 9512
rect 18598 9460 18604 9512
rect 18656 9500 18662 9512
rect 19076 9500 19104 9531
rect 19242 9528 19248 9540
rect 19300 9528 19306 9580
rect 20622 9568 20628 9580
rect 20583 9540 20628 9568
rect 20622 9528 20628 9540
rect 20680 9528 20686 9580
rect 21266 9568 21272 9580
rect 21227 9540 21272 9568
rect 21266 9528 21272 9540
rect 21324 9528 21330 9580
rect 22195 9577 22223 9608
rect 22278 9596 22284 9608
rect 22336 9596 22342 9648
rect 22189 9571 22247 9577
rect 22189 9537 22201 9571
rect 22235 9537 22247 9571
rect 22189 9531 22247 9537
rect 23109 9571 23167 9577
rect 23109 9537 23121 9571
rect 23155 9568 23167 9571
rect 23155 9540 23796 9568
rect 23155 9537 23167 9540
rect 23109 9531 23167 9537
rect 19886 9500 19892 9512
rect 18656 9472 19104 9500
rect 19847 9472 19892 9500
rect 18656 9460 18662 9472
rect 19886 9460 19892 9472
rect 19944 9500 19950 9512
rect 20441 9503 20499 9509
rect 20441 9500 20453 9503
rect 19944 9472 20453 9500
rect 19944 9460 19950 9472
rect 20441 9469 20453 9472
rect 20487 9469 20499 9503
rect 20441 9463 20499 9469
rect 22738 9460 22744 9512
rect 22796 9500 22802 9512
rect 23382 9500 23388 9512
rect 22796 9472 23388 9500
rect 22796 9460 22802 9472
rect 23382 9460 23388 9472
rect 23440 9460 23446 9512
rect 23566 9460 23572 9512
rect 23624 9500 23630 9512
rect 23661 9503 23719 9509
rect 23661 9500 23673 9503
rect 23624 9472 23673 9500
rect 23624 9460 23630 9472
rect 23661 9469 23673 9472
rect 23707 9469 23719 9503
rect 23768 9500 23796 9540
rect 23934 9509 23940 9512
rect 23928 9500 23940 9509
rect 23768 9472 23940 9500
rect 23661 9463 23719 9469
rect 23928 9463 23940 9472
rect 15010 9432 15016 9444
rect 14476 9404 15016 9432
rect 15010 9392 15016 9404
rect 15068 9392 15074 9444
rect 16482 9392 16488 9444
rect 16540 9432 16546 9444
rect 16853 9435 16911 9441
rect 16853 9432 16865 9435
rect 16540 9404 16865 9432
rect 16540 9392 16546 9404
rect 16853 9401 16865 9404
rect 16899 9432 16911 9435
rect 18138 9432 18144 9444
rect 16899 9404 18144 9432
rect 16899 9401 16911 9404
rect 16853 9395 16911 9401
rect 18138 9392 18144 9404
rect 18196 9392 18202 9444
rect 18877 9435 18935 9441
rect 18877 9401 18889 9435
rect 18923 9432 18935 9435
rect 19150 9432 19156 9444
rect 18923 9404 19156 9432
rect 18923 9401 18935 9404
rect 18877 9395 18935 9401
rect 19150 9392 19156 9404
rect 19208 9392 19214 9444
rect 20898 9392 20904 9444
rect 20956 9432 20962 9444
rect 21453 9435 21511 9441
rect 21453 9432 21465 9435
rect 20956 9404 21465 9432
rect 20956 9392 20962 9404
rect 21453 9401 21465 9404
rect 21499 9401 21511 9435
rect 23676 9432 23704 9463
rect 23934 9460 23940 9463
rect 23992 9460 23998 9512
rect 25317 9435 25375 9441
rect 25317 9432 25329 9435
rect 23676 9404 25329 9432
rect 21453 9395 21511 9401
rect 25317 9401 25329 9404
rect 25363 9432 25375 9435
rect 25590 9432 25596 9444
rect 25363 9404 25596 9432
rect 25363 9401 25375 9404
rect 25317 9395 25375 9401
rect 2133 9367 2191 9373
rect 2133 9333 2145 9367
rect 2179 9364 2191 9367
rect 2409 9367 2467 9373
rect 2409 9364 2421 9367
rect 2179 9336 2421 9364
rect 2179 9333 2191 9336
rect 2133 9327 2191 9333
rect 2409 9333 2421 9336
rect 2455 9364 2467 9367
rect 2976 9364 3004 9392
rect 3510 9364 3516 9376
rect 2455 9336 3516 9364
rect 2455 9333 2467 9336
rect 2409 9327 2467 9333
rect 3510 9324 3516 9336
rect 3568 9324 3574 9376
rect 4062 9364 4068 9376
rect 4023 9336 4068 9364
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 5166 9364 5172 9376
rect 5127 9336 5172 9364
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 5537 9367 5595 9373
rect 5537 9333 5549 9367
rect 5583 9364 5595 9367
rect 5994 9364 6000 9376
rect 5583 9336 6000 9364
rect 5583 9333 5595 9336
rect 5537 9327 5595 9333
rect 5994 9324 6000 9336
rect 6052 9324 6058 9376
rect 10778 9364 10784 9376
rect 10739 9336 10784 9364
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 11977 9367 12035 9373
rect 11977 9333 11989 9367
rect 12023 9364 12035 9367
rect 12158 9364 12164 9376
rect 12023 9336 12164 9364
rect 12023 9333 12035 9336
rect 11977 9327 12035 9333
rect 12158 9324 12164 9336
rect 12216 9364 12222 9376
rect 13538 9364 13544 9376
rect 12216 9336 13544 9364
rect 12216 9324 12222 9336
rect 13538 9324 13544 9336
rect 13596 9364 13602 9376
rect 13817 9367 13875 9373
rect 13817 9364 13829 9367
rect 13596 9336 13829 9364
rect 13596 9324 13602 9336
rect 13817 9333 13829 9336
rect 13863 9333 13875 9367
rect 13817 9327 13875 9333
rect 15933 9367 15991 9373
rect 15933 9333 15945 9367
rect 15979 9364 15991 9367
rect 16574 9364 16580 9376
rect 15979 9336 16580 9364
rect 15979 9333 15991 9336
rect 15933 9327 15991 9333
rect 16574 9324 16580 9336
rect 16632 9364 16638 9376
rect 16761 9367 16819 9373
rect 16761 9364 16773 9367
rect 16632 9336 16773 9364
rect 16632 9324 16638 9336
rect 16761 9333 16773 9336
rect 16807 9333 16819 9367
rect 16761 9327 16819 9333
rect 19426 9324 19432 9376
rect 19484 9364 19490 9376
rect 19521 9367 19579 9373
rect 19521 9364 19533 9367
rect 19484 9336 19533 9364
rect 19484 9324 19490 9336
rect 19521 9333 19533 9336
rect 19567 9333 19579 9367
rect 19521 9327 19579 9333
rect 20530 9324 20536 9376
rect 20588 9364 20594 9376
rect 20588 9336 20633 9364
rect 20588 9324 20594 9336
rect 20990 9324 20996 9376
rect 21048 9364 21054 9376
rect 21174 9364 21180 9376
rect 21048 9336 21180 9364
rect 21048 9324 21054 9336
rect 21174 9324 21180 9336
rect 21232 9324 21238 9376
rect 21269 9367 21327 9373
rect 21269 9333 21281 9367
rect 21315 9364 21327 9367
rect 21358 9364 21364 9376
rect 21315 9336 21364 9364
rect 21315 9333 21327 9336
rect 21269 9327 21327 9333
rect 21358 9324 21364 9336
rect 21416 9324 21422 9376
rect 21468 9364 21496 9395
rect 25590 9392 25596 9404
rect 25648 9432 25654 9444
rect 25685 9435 25743 9441
rect 25685 9432 25697 9435
rect 25648 9404 25697 9432
rect 25648 9392 25654 9404
rect 25685 9401 25697 9404
rect 25731 9432 25743 9435
rect 26053 9435 26111 9441
rect 26053 9432 26065 9435
rect 25731 9404 26065 9432
rect 25731 9401 25743 9404
rect 25685 9395 25743 9401
rect 26053 9401 26065 9404
rect 26099 9401 26111 9435
rect 26053 9395 26111 9401
rect 22005 9367 22063 9373
rect 22005 9364 22017 9367
rect 21468 9336 22017 9364
rect 22005 9333 22017 9336
rect 22051 9333 22063 9367
rect 22005 9327 22063 9333
rect 22097 9367 22155 9373
rect 22097 9333 22109 9367
rect 22143 9364 22155 9367
rect 22186 9364 22192 9376
rect 22143 9336 22192 9364
rect 22143 9333 22155 9336
rect 22097 9327 22155 9333
rect 22186 9324 22192 9336
rect 22244 9364 22250 9376
rect 24946 9364 24952 9376
rect 22244 9336 24952 9364
rect 22244 9324 22250 9336
rect 24946 9324 24952 9336
rect 25004 9324 25010 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1670 9120 1676 9172
rect 1728 9160 1734 9172
rect 1857 9163 1915 9169
rect 1857 9160 1869 9163
rect 1728 9132 1869 9160
rect 1728 9120 1734 9132
rect 1857 9129 1869 9132
rect 1903 9129 1915 9163
rect 1857 9123 1915 9129
rect 2409 9163 2467 9169
rect 2409 9129 2421 9163
rect 2455 9160 2467 9163
rect 2682 9160 2688 9172
rect 2455 9132 2688 9160
rect 2455 9129 2467 9132
rect 2409 9123 2467 9129
rect 2682 9120 2688 9132
rect 2740 9120 2746 9172
rect 4709 9163 4767 9169
rect 4709 9129 4721 9163
rect 4755 9160 4767 9163
rect 5442 9160 5448 9172
rect 4755 9132 5448 9160
rect 4755 9129 4767 9132
rect 4709 9123 4767 9129
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 6549 9163 6607 9169
rect 6549 9129 6561 9163
rect 6595 9160 6607 9163
rect 6822 9160 6828 9172
rect 6595 9132 6828 9160
rect 6595 9129 6607 9132
rect 6549 9123 6607 9129
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 9766 9160 9772 9172
rect 9727 9132 9772 9160
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 10321 9163 10379 9169
rect 10321 9129 10333 9163
rect 10367 9160 10379 9163
rect 11146 9160 11152 9172
rect 10367 9132 11152 9160
rect 10367 9129 10379 9132
rect 10321 9123 10379 9129
rect 11146 9120 11152 9132
rect 11204 9120 11210 9172
rect 11790 9120 11796 9172
rect 11848 9160 11854 9172
rect 12161 9163 12219 9169
rect 12161 9160 12173 9163
rect 11848 9132 12173 9160
rect 11848 9120 11854 9132
rect 12161 9129 12173 9132
rect 12207 9160 12219 9163
rect 12710 9160 12716 9172
rect 12207 9132 12716 9160
rect 12207 9129 12219 9132
rect 12161 9123 12219 9129
rect 12710 9120 12716 9132
rect 12768 9160 12774 9172
rect 12805 9163 12863 9169
rect 12805 9160 12817 9163
rect 12768 9132 12817 9160
rect 12768 9120 12774 9132
rect 12805 9129 12817 9132
rect 12851 9129 12863 9163
rect 12805 9123 12863 9129
rect 13262 9120 13268 9172
rect 13320 9160 13326 9172
rect 13446 9160 13452 9172
rect 13320 9132 13452 9160
rect 13320 9120 13326 9132
rect 13446 9120 13452 9132
rect 13504 9120 13510 9172
rect 14642 9160 14648 9172
rect 14603 9132 14648 9160
rect 14642 9120 14648 9132
rect 14700 9120 14706 9172
rect 15102 9160 15108 9172
rect 15063 9132 15108 9160
rect 15102 9120 15108 9132
rect 15160 9120 15166 9172
rect 15289 9163 15347 9169
rect 15289 9129 15301 9163
rect 15335 9160 15347 9163
rect 15378 9160 15384 9172
rect 15335 9132 15384 9160
rect 15335 9129 15347 9132
rect 15289 9123 15347 9129
rect 15378 9120 15384 9132
rect 15436 9120 15442 9172
rect 15654 9160 15660 9172
rect 15615 9132 15660 9160
rect 15654 9120 15660 9132
rect 15712 9160 15718 9172
rect 16206 9160 16212 9172
rect 15712 9132 16212 9160
rect 15712 9120 15718 9132
rect 16206 9120 16212 9132
rect 16264 9120 16270 9172
rect 16482 9160 16488 9172
rect 16443 9132 16488 9160
rect 16482 9120 16488 9132
rect 16540 9120 16546 9172
rect 16850 9160 16856 9172
rect 16811 9132 16856 9160
rect 16850 9120 16856 9132
rect 16908 9120 16914 9172
rect 17494 9160 17500 9172
rect 17455 9132 17500 9160
rect 17494 9120 17500 9132
rect 17552 9120 17558 9172
rect 18598 9160 18604 9172
rect 18559 9132 18604 9160
rect 18598 9120 18604 9132
rect 18656 9120 18662 9172
rect 18693 9163 18751 9169
rect 18693 9129 18705 9163
rect 18739 9160 18751 9163
rect 18782 9160 18788 9172
rect 18739 9132 18788 9160
rect 18739 9129 18751 9132
rect 18693 9123 18751 9129
rect 18782 9120 18788 9132
rect 18840 9120 18846 9172
rect 20165 9163 20223 9169
rect 20165 9129 20177 9163
rect 20211 9160 20223 9163
rect 20530 9160 20536 9172
rect 20211 9132 20536 9160
rect 20211 9129 20223 9132
rect 20165 9123 20223 9129
rect 20530 9120 20536 9132
rect 20588 9120 20594 9172
rect 21174 9120 21180 9172
rect 21232 9160 21238 9172
rect 22186 9160 22192 9172
rect 21232 9132 22192 9160
rect 21232 9120 21238 9132
rect 22186 9120 22192 9132
rect 22244 9120 22250 9172
rect 23934 9120 23940 9172
rect 23992 9160 23998 9172
rect 24121 9163 24179 9169
rect 24121 9160 24133 9163
rect 23992 9132 24133 9160
rect 23992 9120 23998 9132
rect 24121 9129 24133 9132
rect 24167 9129 24179 9163
rect 24121 9123 24179 9129
rect 24857 9163 24915 9169
rect 24857 9129 24869 9163
rect 24903 9160 24915 9163
rect 25130 9160 25136 9172
rect 24903 9132 25136 9160
rect 24903 9129 24915 9132
rect 24857 9123 24915 9129
rect 25130 9120 25136 9132
rect 25188 9120 25194 9172
rect 25590 9160 25596 9172
rect 25551 9132 25596 9160
rect 25590 9120 25596 9132
rect 25648 9160 25654 9172
rect 25869 9163 25927 9169
rect 25869 9160 25881 9163
rect 25648 9132 25881 9160
rect 25648 9120 25654 9132
rect 25869 9129 25881 9132
rect 25915 9160 25927 9163
rect 26142 9160 26148 9172
rect 25915 9132 26148 9160
rect 25915 9129 25927 9132
rect 25869 9123 25927 9129
rect 26142 9120 26148 9132
rect 26200 9160 26206 9172
rect 26237 9163 26295 9169
rect 26237 9160 26249 9163
rect 26200 9132 26249 9160
rect 26200 9120 26206 9132
rect 26237 9129 26249 9132
rect 26283 9129 26295 9163
rect 26237 9123 26295 9129
rect 2869 9095 2927 9101
rect 2869 9092 2881 9095
rect 2240 9064 2881 9092
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8956 1455 8959
rect 1578 8956 1584 8968
rect 1443 8928 1584 8956
rect 1443 8925 1455 8928
rect 1397 8919 1455 8925
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 2240 8897 2268 9064
rect 2869 9061 2881 9064
rect 2915 9061 2927 9095
rect 2869 9055 2927 9061
rect 5261 9095 5319 9101
rect 5261 9061 5273 9095
rect 5307 9092 5319 9095
rect 5994 9092 6000 9104
rect 5307 9064 6000 9092
rect 5307 9061 5319 9064
rect 5261 9055 5319 9061
rect 5994 9052 6000 9064
rect 6052 9052 6058 9104
rect 7377 9095 7435 9101
rect 7377 9061 7389 9095
rect 7423 9092 7435 9095
rect 7926 9092 7932 9104
rect 7423 9064 7932 9092
rect 7423 9061 7435 9064
rect 7377 9055 7435 9061
rect 7926 9052 7932 9064
rect 7984 9052 7990 9104
rect 8846 9052 8852 9104
rect 8904 9092 8910 9104
rect 9398 9092 9404 9104
rect 8904 9064 9404 9092
rect 8904 9052 8910 9064
rect 9398 9052 9404 9064
rect 9456 9052 9462 9104
rect 10689 9095 10747 9101
rect 10689 9061 10701 9095
rect 10735 9092 10747 9095
rect 11026 9095 11084 9101
rect 11026 9092 11038 9095
rect 10735 9064 11038 9092
rect 10735 9061 10747 9064
rect 10689 9055 10747 9061
rect 11026 9061 11038 9064
rect 11072 9092 11084 9095
rect 11422 9092 11428 9104
rect 11072 9064 11428 9092
rect 11072 9061 11084 9064
rect 11026 9055 11084 9061
rect 11422 9052 11428 9064
rect 11480 9092 11486 9104
rect 11480 9064 12572 9092
rect 11480 9052 11486 9064
rect 2682 8984 2688 9036
rect 2740 9024 2746 9036
rect 2777 9027 2835 9033
rect 2777 9024 2789 9027
rect 2740 8996 2789 9024
rect 2740 8984 2746 8996
rect 2777 8993 2789 8996
rect 2823 8993 2835 9027
rect 2777 8987 2835 8993
rect 5534 8984 5540 9036
rect 5592 9024 5598 9036
rect 5813 9027 5871 9033
rect 5813 9024 5825 9027
rect 5592 8996 5825 9024
rect 5592 8984 5598 8996
rect 5813 8993 5825 8996
rect 5859 9024 5871 9027
rect 7469 9027 7527 9033
rect 5859 8996 6132 9024
rect 5859 8993 5871 8996
rect 5813 8987 5871 8993
rect 2958 8916 2964 8968
rect 3016 8956 3022 8968
rect 3421 8959 3479 8965
rect 3421 8956 3433 8959
rect 3016 8928 3433 8956
rect 3016 8916 3022 8928
rect 3421 8925 3433 8928
rect 3467 8925 3479 8959
rect 3421 8919 3479 8925
rect 5166 8916 5172 8968
rect 5224 8956 5230 8968
rect 5905 8959 5963 8965
rect 5905 8956 5917 8959
rect 5224 8928 5917 8956
rect 5224 8916 5230 8928
rect 5905 8925 5917 8928
rect 5951 8925 5963 8959
rect 5905 8919 5963 8925
rect 5997 8959 6055 8965
rect 5997 8925 6009 8959
rect 6043 8925 6055 8959
rect 5997 8919 6055 8925
rect 2225 8891 2283 8897
rect 2225 8888 2237 8891
rect 2056 8860 2237 8888
rect 2056 8832 2084 8860
rect 2225 8857 2237 8860
rect 2271 8857 2283 8891
rect 2225 8851 2283 8857
rect 3881 8891 3939 8897
rect 3881 8857 3893 8891
rect 3927 8888 3939 8891
rect 5442 8888 5448 8900
rect 3927 8860 5448 8888
rect 3927 8857 3939 8860
rect 3881 8851 3939 8857
rect 5442 8848 5448 8860
rect 5500 8848 5506 8900
rect 2038 8780 2044 8832
rect 2096 8780 2102 8832
rect 4338 8820 4344 8832
rect 4299 8792 4344 8820
rect 4338 8780 4344 8792
rect 4396 8780 4402 8832
rect 4890 8780 4896 8832
rect 4948 8820 4954 8832
rect 6012 8820 6040 8919
rect 6104 8888 6132 8996
rect 7469 8993 7481 9027
rect 7515 9024 7527 9027
rect 7650 9024 7656 9036
rect 7515 8996 7656 9024
rect 7515 8993 7527 8996
rect 7469 8987 7527 8993
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 6270 8916 6276 8968
rect 6328 8956 6334 8968
rect 6454 8956 6460 8968
rect 6328 8928 6460 8956
rect 6328 8916 6334 8928
rect 6454 8916 6460 8928
rect 6512 8956 6518 8968
rect 7561 8959 7619 8965
rect 7561 8956 7573 8959
rect 6512 8928 7573 8956
rect 6512 8916 6518 8928
rect 7561 8925 7573 8928
rect 7607 8925 7619 8959
rect 8570 8956 8576 8968
rect 8531 8928 8576 8956
rect 7561 8919 7619 8925
rect 8570 8916 8576 8928
rect 8628 8916 8634 8968
rect 9398 8916 9404 8968
rect 9456 8956 9462 8968
rect 12544 8965 12572 9064
rect 13170 9052 13176 9104
rect 13228 9092 13234 9104
rect 13357 9095 13415 9101
rect 13357 9092 13369 9095
rect 13228 9064 13369 9092
rect 13228 9052 13234 9064
rect 13357 9061 13369 9064
rect 13403 9092 13415 9095
rect 13906 9092 13912 9104
rect 13403 9064 13912 9092
rect 13403 9061 13415 9064
rect 13357 9055 13415 9061
rect 13906 9052 13912 9064
rect 13964 9052 13970 9104
rect 22922 9052 22928 9104
rect 22980 9101 22986 9104
rect 22980 9095 23044 9101
rect 22980 9061 22998 9095
rect 23032 9061 23044 9095
rect 22980 9055 23044 9061
rect 22980 9052 22986 9055
rect 13446 8984 13452 9036
rect 13504 9024 13510 9036
rect 14001 9027 14059 9033
rect 14001 9024 14013 9027
rect 13504 8996 14013 9024
rect 13504 8984 13510 8996
rect 14001 8993 14013 8996
rect 14047 8993 14059 9027
rect 14001 8987 14059 8993
rect 16942 8984 16948 9036
rect 17000 9024 17006 9036
rect 17000 8996 17632 9024
rect 17000 8984 17006 8996
rect 10781 8959 10839 8965
rect 10781 8956 10793 8959
rect 9456 8928 10793 8956
rect 9456 8916 9462 8928
rect 10781 8925 10793 8928
rect 10827 8925 10839 8959
rect 10781 8919 10839 8925
rect 12529 8959 12587 8965
rect 12529 8925 12541 8959
rect 12575 8956 12587 8959
rect 12986 8956 12992 8968
rect 12575 8928 12992 8956
rect 12575 8925 12587 8928
rect 12529 8919 12587 8925
rect 7009 8891 7067 8897
rect 7009 8888 7021 8891
rect 6104 8860 7021 8888
rect 7009 8857 7021 8860
rect 7055 8857 7067 8891
rect 7009 8851 7067 8857
rect 8018 8848 8024 8900
rect 8076 8888 8082 8900
rect 8113 8891 8171 8897
rect 8113 8888 8125 8891
rect 8076 8860 8125 8888
rect 8076 8848 8082 8860
rect 8113 8857 8125 8860
rect 8159 8888 8171 8891
rect 8159 8860 9168 8888
rect 8159 8857 8171 8860
rect 8113 8851 8171 8857
rect 9140 8832 9168 8860
rect 6270 8820 6276 8832
rect 4948 8792 6276 8820
rect 4948 8780 4954 8792
rect 6270 8780 6276 8792
rect 6328 8820 6334 8832
rect 6825 8823 6883 8829
rect 6825 8820 6837 8823
rect 6328 8792 6837 8820
rect 6328 8780 6334 8792
rect 6825 8789 6837 8792
rect 6871 8789 6883 8823
rect 6825 8783 6883 8789
rect 7834 8780 7840 8832
rect 7892 8820 7898 8832
rect 8481 8823 8539 8829
rect 8481 8820 8493 8823
rect 7892 8792 8493 8820
rect 7892 8780 7898 8792
rect 8481 8789 8493 8792
rect 8527 8820 8539 8823
rect 8662 8820 8668 8832
rect 8527 8792 8668 8820
rect 8527 8789 8539 8792
rect 8481 8783 8539 8789
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 9122 8820 9128 8832
rect 9083 8792 9128 8820
rect 9122 8780 9128 8792
rect 9180 8780 9186 8832
rect 10796 8820 10824 8919
rect 12986 8916 12992 8928
rect 13044 8916 13050 8968
rect 13538 8956 13544 8968
rect 13499 8928 13544 8956
rect 13538 8916 13544 8928
rect 13596 8916 13602 8968
rect 15746 8956 15752 8968
rect 15707 8928 15752 8956
rect 15746 8916 15752 8928
rect 15804 8916 15810 8968
rect 15841 8959 15899 8965
rect 15841 8925 15853 8959
rect 15887 8925 15899 8959
rect 15841 8919 15899 8925
rect 11882 8848 11888 8900
rect 11940 8888 11946 8900
rect 11940 8860 13768 8888
rect 11940 8848 11946 8860
rect 10962 8820 10968 8832
rect 10796 8792 10968 8820
rect 10962 8780 10968 8792
rect 11020 8780 11026 8832
rect 12989 8823 13047 8829
rect 12989 8789 13001 8823
rect 13035 8820 13047 8823
rect 13630 8820 13636 8832
rect 13035 8792 13636 8820
rect 13035 8789 13047 8792
rect 12989 8783 13047 8789
rect 13630 8780 13636 8792
rect 13688 8780 13694 8832
rect 13740 8820 13768 8860
rect 14366 8848 14372 8900
rect 14424 8888 14430 8900
rect 15856 8888 15884 8919
rect 17218 8916 17224 8968
rect 17276 8916 17282 8968
rect 17604 8965 17632 8996
rect 17954 8984 17960 9036
rect 18012 9024 18018 9036
rect 19061 9027 19119 9033
rect 19061 9024 19073 9027
rect 18012 8996 19073 9024
rect 18012 8984 18018 8996
rect 19061 8993 19073 8996
rect 19107 9024 19119 9027
rect 19705 9027 19763 9033
rect 19705 9024 19717 9027
rect 19107 8996 19717 9024
rect 19107 8993 19119 8996
rect 19061 8987 19119 8993
rect 19705 8993 19717 8996
rect 19751 8993 19763 9027
rect 19705 8987 19763 8993
rect 19978 8984 19984 9036
rect 20036 9024 20042 9036
rect 20441 9027 20499 9033
rect 20441 9024 20453 9027
rect 20036 8996 20453 9024
rect 20036 8984 20042 8996
rect 20441 8993 20453 8996
rect 20487 9024 20499 9027
rect 20530 9024 20536 9036
rect 20487 8996 20536 9024
rect 20487 8993 20499 8996
rect 20441 8987 20499 8993
rect 20530 8984 20536 8996
rect 20588 8984 20594 9036
rect 20898 8984 20904 9036
rect 20956 9024 20962 9036
rect 21269 9027 21327 9033
rect 21269 9024 21281 9027
rect 20956 8996 21281 9024
rect 20956 8984 20962 8996
rect 21269 8993 21281 8996
rect 21315 8993 21327 9027
rect 23566 9024 23572 9036
rect 21269 8987 21327 8993
rect 22756 8996 23572 9024
rect 17589 8959 17647 8965
rect 17589 8925 17601 8959
rect 17635 8956 17647 8959
rect 17678 8956 17684 8968
rect 17635 8928 17684 8956
rect 17635 8925 17647 8928
rect 17589 8919 17647 8925
rect 17678 8916 17684 8928
rect 17736 8916 17742 8968
rect 17773 8959 17831 8965
rect 17773 8925 17785 8959
rect 17819 8956 17831 8959
rect 18046 8956 18052 8968
rect 17819 8928 18052 8956
rect 17819 8925 17831 8928
rect 17773 8919 17831 8925
rect 18046 8916 18052 8928
rect 18104 8916 18110 8968
rect 18233 8959 18291 8965
rect 18233 8925 18245 8959
rect 18279 8956 18291 8959
rect 19150 8956 19156 8968
rect 18279 8928 19156 8956
rect 18279 8925 18291 8928
rect 18233 8919 18291 8925
rect 19150 8916 19156 8928
rect 19208 8916 19214 8968
rect 19337 8959 19395 8965
rect 19337 8925 19349 8959
rect 19383 8956 19395 8959
rect 19518 8956 19524 8968
rect 19383 8928 19524 8956
rect 19383 8925 19395 8928
rect 19337 8919 19395 8925
rect 19518 8916 19524 8928
rect 19576 8916 19582 8968
rect 21174 8916 21180 8968
rect 21232 8956 21238 8968
rect 21361 8959 21419 8965
rect 21361 8956 21373 8959
rect 21232 8928 21373 8956
rect 21232 8916 21238 8928
rect 21361 8925 21373 8928
rect 21407 8925 21419 8959
rect 21361 8919 21419 8925
rect 21453 8959 21511 8965
rect 21453 8925 21465 8959
rect 21499 8925 21511 8959
rect 21453 8919 21511 8925
rect 14424 8860 15884 8888
rect 17236 8888 17264 8916
rect 17236 8860 18000 8888
rect 14424 8848 14430 8860
rect 17972 8832 18000 8860
rect 20622 8848 20628 8900
rect 20680 8888 20686 8900
rect 21468 8888 21496 8919
rect 21818 8916 21824 8968
rect 21876 8956 21882 8968
rect 22756 8965 22784 8996
rect 23566 8984 23572 8996
rect 23624 8984 23630 9036
rect 24946 9024 24952 9036
rect 24907 8996 24952 9024
rect 24946 8984 24952 8996
rect 25004 8984 25010 9036
rect 22741 8959 22799 8965
rect 22741 8956 22753 8959
rect 21876 8928 22753 8956
rect 21876 8916 21882 8928
rect 22741 8925 22753 8928
rect 22787 8925 22799 8959
rect 22741 8919 22799 8925
rect 21542 8888 21548 8900
rect 20680 8860 21548 8888
rect 20680 8848 20686 8860
rect 21542 8848 21548 8860
rect 21600 8848 21606 8900
rect 25590 8888 25596 8900
rect 24412 8860 25596 8888
rect 16390 8820 16396 8832
rect 13740 8792 16396 8820
rect 16390 8780 16396 8792
rect 16448 8780 16454 8832
rect 17129 8823 17187 8829
rect 17129 8789 17141 8823
rect 17175 8820 17187 8823
rect 17218 8820 17224 8832
rect 17175 8792 17224 8820
rect 17175 8789 17187 8792
rect 17129 8783 17187 8789
rect 17218 8780 17224 8792
rect 17276 8780 17282 8832
rect 17954 8780 17960 8832
rect 18012 8780 18018 8832
rect 20254 8820 20260 8832
rect 20215 8792 20260 8820
rect 20254 8780 20260 8792
rect 20312 8780 20318 8832
rect 20806 8780 20812 8832
rect 20864 8820 20870 8832
rect 20901 8823 20959 8829
rect 20901 8820 20913 8823
rect 20864 8792 20913 8820
rect 20864 8780 20870 8792
rect 20901 8789 20913 8792
rect 20947 8789 20959 8823
rect 20901 8783 20959 8789
rect 21450 8780 21456 8832
rect 21508 8820 21514 8832
rect 22002 8820 22008 8832
rect 21508 8792 22008 8820
rect 21508 8780 21514 8792
rect 22002 8780 22008 8792
rect 22060 8780 22066 8832
rect 22186 8780 22192 8832
rect 22244 8820 22250 8832
rect 22281 8823 22339 8829
rect 22281 8820 22293 8823
rect 22244 8792 22293 8820
rect 22244 8780 22250 8792
rect 22281 8789 22293 8792
rect 22327 8820 22339 8823
rect 23014 8820 23020 8832
rect 22327 8792 23020 8820
rect 22327 8789 22339 8792
rect 22281 8783 22339 8789
rect 23014 8780 23020 8792
rect 23072 8820 23078 8832
rect 24412 8829 24440 8860
rect 25590 8848 25596 8860
rect 25648 8848 25654 8900
rect 24397 8823 24455 8829
rect 24397 8820 24409 8823
rect 23072 8792 24409 8820
rect 23072 8780 23078 8792
rect 24397 8789 24409 8792
rect 24443 8789 24455 8823
rect 25130 8820 25136 8832
rect 25091 8792 25136 8820
rect 24397 8783 24455 8789
rect 25130 8780 25136 8792
rect 25188 8780 25194 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 5074 8616 5080 8628
rect 5035 8588 5080 8616
rect 5074 8576 5080 8588
rect 5132 8576 5138 8628
rect 6273 8619 6331 8625
rect 6273 8585 6285 8619
rect 6319 8616 6331 8619
rect 6454 8616 6460 8628
rect 6319 8588 6460 8616
rect 6319 8585 6331 8588
rect 6273 8579 6331 8585
rect 6454 8576 6460 8588
rect 6512 8576 6518 8628
rect 6641 8619 6699 8625
rect 6641 8585 6653 8619
rect 6687 8616 6699 8619
rect 7650 8616 7656 8628
rect 6687 8588 7656 8616
rect 6687 8585 6699 8588
rect 6641 8579 6699 8585
rect 7650 8576 7656 8588
rect 7708 8576 7714 8628
rect 7926 8616 7932 8628
rect 7887 8588 7932 8616
rect 7926 8576 7932 8588
rect 7984 8576 7990 8628
rect 8297 8619 8355 8625
rect 8297 8585 8309 8619
rect 8343 8616 8355 8619
rect 8386 8616 8392 8628
rect 8343 8588 8392 8616
rect 8343 8585 8355 8588
rect 8297 8579 8355 8585
rect 8386 8576 8392 8588
rect 8444 8576 8450 8628
rect 9398 8576 9404 8628
rect 9456 8616 9462 8628
rect 9953 8619 10011 8625
rect 9953 8616 9965 8619
rect 9456 8588 9965 8616
rect 9456 8576 9462 8588
rect 9953 8585 9965 8588
rect 9999 8616 10011 8619
rect 10134 8616 10140 8628
rect 9999 8588 10140 8616
rect 9999 8585 10011 8588
rect 9953 8579 10011 8585
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 13538 8616 13544 8628
rect 13499 8588 13544 8616
rect 13538 8576 13544 8588
rect 13596 8576 13602 8628
rect 14734 8576 14740 8628
rect 14792 8616 14798 8628
rect 15838 8616 15844 8628
rect 14792 8588 15844 8616
rect 14792 8576 14798 8588
rect 15838 8576 15844 8588
rect 15896 8616 15902 8628
rect 16301 8619 16359 8625
rect 16301 8616 16313 8619
rect 15896 8588 16313 8616
rect 15896 8576 15902 8588
rect 16301 8585 16313 8588
rect 16347 8585 16359 8619
rect 16301 8579 16359 8585
rect 17129 8619 17187 8625
rect 17129 8585 17141 8619
rect 17175 8616 17187 8619
rect 17494 8616 17500 8628
rect 17175 8588 17500 8616
rect 17175 8585 17187 8588
rect 17129 8579 17187 8585
rect 17494 8576 17500 8588
rect 17552 8576 17558 8628
rect 17678 8576 17684 8628
rect 17736 8616 17742 8628
rect 17773 8619 17831 8625
rect 17773 8616 17785 8619
rect 17736 8588 17785 8616
rect 17736 8576 17742 8588
rect 17773 8585 17785 8588
rect 17819 8616 17831 8619
rect 18414 8616 18420 8628
rect 17819 8588 18420 8616
rect 17819 8585 17831 8588
rect 17773 8579 17831 8585
rect 18414 8576 18420 8588
rect 18472 8576 18478 8628
rect 19426 8616 19432 8628
rect 19387 8588 19432 8616
rect 19426 8576 19432 8588
rect 19484 8576 19490 8628
rect 21174 8616 21180 8628
rect 20364 8588 21180 8616
rect 6825 8551 6883 8557
rect 6825 8548 6837 8551
rect 5552 8520 6837 8548
rect 1210 8440 1216 8492
rect 1268 8480 1274 8492
rect 1762 8480 1768 8492
rect 1268 8452 1768 8480
rect 1268 8440 1274 8452
rect 1762 8440 1768 8452
rect 1820 8440 1826 8492
rect 4338 8440 4344 8492
rect 4396 8480 4402 8492
rect 5552 8489 5580 8520
rect 6825 8517 6837 8520
rect 6871 8517 6883 8551
rect 6825 8511 6883 8517
rect 10781 8551 10839 8557
rect 10781 8517 10793 8551
rect 10827 8548 10839 8551
rect 14366 8548 14372 8560
rect 10827 8520 12940 8548
rect 14327 8520 14372 8548
rect 10827 8517 10839 8520
rect 10781 8511 10839 8517
rect 5537 8483 5595 8489
rect 5537 8480 5549 8483
rect 4396 8452 5549 8480
rect 4396 8440 4402 8452
rect 5537 8449 5549 8452
rect 5583 8449 5595 8483
rect 5537 8443 5595 8449
rect 5629 8483 5687 8489
rect 5629 8449 5641 8483
rect 5675 8449 5687 8483
rect 5629 8443 5687 8449
rect 1670 8372 1676 8424
rect 1728 8412 1734 8424
rect 2406 8412 2412 8424
rect 1728 8384 2412 8412
rect 1728 8372 1734 8384
rect 2406 8372 2412 8384
rect 2464 8412 2470 8424
rect 2869 8415 2927 8421
rect 2869 8412 2881 8415
rect 2464 8384 2881 8412
rect 2464 8372 2470 8384
rect 2869 8381 2881 8384
rect 2915 8381 2927 8415
rect 4890 8412 4896 8424
rect 2869 8375 2927 8381
rect 3436 8384 4896 8412
rect 1762 8344 1768 8356
rect 1723 8316 1768 8344
rect 1762 8304 1768 8316
rect 1820 8304 1826 8356
rect 1857 8347 1915 8353
rect 1857 8313 1869 8347
rect 1903 8344 1915 8347
rect 1903 8316 2820 8344
rect 1903 8313 1915 8316
rect 1857 8307 1915 8313
rect 2792 8288 2820 8316
rect 2958 8304 2964 8356
rect 3016 8344 3022 8356
rect 3114 8347 3172 8353
rect 3114 8344 3126 8347
rect 3016 8316 3126 8344
rect 3016 8304 3022 8316
rect 3114 8313 3126 8316
rect 3160 8344 3172 8347
rect 3436 8344 3464 8384
rect 4890 8372 4896 8384
rect 4948 8372 4954 8424
rect 5442 8412 5448 8424
rect 5403 8384 5448 8412
rect 5442 8372 5448 8384
rect 5500 8372 5506 8424
rect 3160 8316 3464 8344
rect 3160 8313 3172 8316
rect 3114 8307 3172 8313
rect 3510 8304 3516 8356
rect 3568 8344 3574 8356
rect 4617 8347 4675 8353
rect 4617 8344 4629 8347
rect 3568 8316 4629 8344
rect 3568 8304 3574 8316
rect 1302 8236 1308 8288
rect 1360 8276 1366 8288
rect 2409 8279 2467 8285
rect 2409 8276 2421 8279
rect 1360 8248 2421 8276
rect 1360 8236 1366 8248
rect 2409 8245 2421 8248
rect 2455 8276 2467 8279
rect 2682 8276 2688 8288
rect 2455 8248 2688 8276
rect 2455 8245 2467 8248
rect 2409 8239 2467 8245
rect 2682 8236 2688 8248
rect 2740 8236 2746 8288
rect 2774 8236 2780 8288
rect 2832 8236 2838 8288
rect 4264 8285 4292 8316
rect 4617 8313 4629 8316
rect 4663 8344 4675 8347
rect 5644 8344 5672 8443
rect 6270 8440 6276 8492
rect 6328 8480 6334 8492
rect 7377 8483 7435 8489
rect 7377 8480 7389 8483
rect 6328 8452 7389 8480
rect 6328 8440 6334 8452
rect 7377 8449 7389 8452
rect 7423 8449 7435 8483
rect 7377 8443 7435 8449
rect 9033 8483 9091 8489
rect 9033 8449 9045 8483
rect 9079 8480 9091 8483
rect 11238 8480 11244 8492
rect 9079 8452 9113 8480
rect 11199 8452 11244 8480
rect 9079 8449 9091 8452
rect 9033 8443 9091 8449
rect 6822 8372 6828 8424
rect 6880 8412 6886 8424
rect 7193 8415 7251 8421
rect 7193 8412 7205 8415
rect 6880 8384 7205 8412
rect 6880 8372 6886 8384
rect 7193 8381 7205 8384
rect 7239 8381 7251 8415
rect 7193 8375 7251 8381
rect 8386 8372 8392 8424
rect 8444 8412 8450 8424
rect 8757 8415 8815 8421
rect 8757 8412 8769 8415
rect 8444 8384 8769 8412
rect 8444 8372 8450 8384
rect 8757 8381 8769 8384
rect 8803 8381 8815 8415
rect 8757 8375 8815 8381
rect 8846 8372 8852 8424
rect 8904 8412 8910 8424
rect 9048 8412 9076 8443
rect 11238 8440 11244 8452
rect 11296 8440 11302 8492
rect 11422 8480 11428 8492
rect 11335 8452 11428 8480
rect 11422 8440 11428 8452
rect 11480 8480 11486 8492
rect 11793 8483 11851 8489
rect 11793 8480 11805 8483
rect 11480 8452 11805 8480
rect 11480 8440 11486 8452
rect 11793 8449 11805 8452
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 9401 8415 9459 8421
rect 9401 8412 9413 8415
rect 8904 8384 9413 8412
rect 8904 8372 8910 8384
rect 9401 8381 9413 8384
rect 9447 8381 9459 8415
rect 10137 8415 10195 8421
rect 10137 8412 10149 8415
rect 9401 8375 9459 8381
rect 9784 8384 10149 8412
rect 9784 8356 9812 8384
rect 10137 8381 10149 8384
rect 10183 8381 10195 8415
rect 10137 8375 10195 8381
rect 10689 8415 10747 8421
rect 10689 8381 10701 8415
rect 10735 8412 10747 8415
rect 11146 8412 11152 8424
rect 10735 8384 11152 8412
rect 10735 8381 10747 8384
rect 10689 8375 10747 8381
rect 11146 8372 11152 8384
rect 11204 8372 11210 8424
rect 4663 8316 5672 8344
rect 4663 8313 4675 8316
rect 4617 8307 4675 8313
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 7285 8347 7343 8353
rect 7285 8344 7297 8347
rect 6972 8316 7297 8344
rect 6972 8304 6978 8316
rect 7285 8313 7297 8316
rect 7331 8344 7343 8347
rect 7558 8344 7564 8356
rect 7331 8316 7564 8344
rect 7331 8313 7343 8316
rect 7285 8307 7343 8313
rect 7558 8304 7564 8316
rect 7616 8304 7622 8356
rect 8662 8304 8668 8356
rect 8720 8344 8726 8356
rect 9214 8344 9220 8356
rect 8720 8316 9220 8344
rect 8720 8304 8726 8316
rect 4249 8279 4307 8285
rect 4249 8245 4261 8279
rect 4295 8245 4307 8279
rect 8386 8276 8392 8288
rect 8347 8248 8392 8276
rect 4249 8239 4307 8245
rect 8386 8236 8392 8248
rect 8444 8236 8450 8288
rect 8864 8285 8892 8316
rect 9214 8304 9220 8316
rect 9272 8304 9278 8356
rect 9766 8344 9772 8356
rect 9727 8316 9772 8344
rect 9766 8304 9772 8316
rect 9824 8304 9830 8356
rect 11256 8344 11284 8440
rect 12253 8415 12311 8421
rect 12253 8381 12265 8415
rect 12299 8412 12311 8415
rect 12434 8412 12440 8424
rect 12299 8384 12440 8412
rect 12299 8381 12311 8384
rect 12253 8375 12311 8381
rect 12434 8372 12440 8384
rect 12492 8412 12498 8424
rect 12805 8415 12863 8421
rect 12805 8412 12817 8415
rect 12492 8384 12817 8412
rect 12492 8372 12498 8384
rect 12805 8381 12817 8384
rect 12851 8381 12863 8415
rect 12805 8375 12863 8381
rect 12912 8353 12940 8520
rect 14366 8508 14372 8520
rect 14424 8508 14430 8560
rect 17221 8551 17279 8557
rect 17221 8517 17233 8551
rect 17267 8548 17279 8551
rect 17267 8520 18092 8548
rect 17267 8517 17279 8520
rect 17221 8511 17279 8517
rect 12986 8440 12992 8492
rect 13044 8480 13050 8492
rect 13044 8452 13089 8480
rect 13044 8440 13050 8452
rect 14918 8412 14924 8424
rect 14879 8384 14924 8412
rect 14918 8372 14924 8384
rect 14976 8372 14982 8424
rect 15188 8415 15246 8421
rect 15188 8381 15200 8415
rect 15234 8412 15246 8415
rect 16022 8412 16028 8424
rect 15234 8384 16028 8412
rect 15234 8381 15246 8384
rect 15188 8375 15246 8381
rect 10980 8316 11284 8344
rect 12897 8347 12955 8353
rect 8849 8279 8907 8285
rect 8849 8245 8861 8279
rect 8895 8245 8907 8279
rect 8849 8239 8907 8245
rect 10778 8236 10784 8288
rect 10836 8276 10842 8288
rect 10980 8276 11008 8316
rect 12897 8313 12909 8347
rect 12943 8344 12955 8347
rect 13817 8347 13875 8353
rect 13817 8344 13829 8347
rect 12943 8316 13829 8344
rect 12943 8313 12955 8316
rect 12897 8307 12955 8313
rect 13817 8313 13829 8316
rect 13863 8313 13875 8347
rect 13817 8307 13875 8313
rect 14829 8347 14887 8353
rect 14829 8313 14841 8347
rect 14875 8344 14887 8347
rect 15203 8344 15231 8375
rect 16022 8372 16028 8384
rect 16080 8372 16086 8424
rect 17402 8412 17408 8424
rect 17363 8384 17408 8412
rect 17402 8372 17408 8384
rect 17460 8372 17466 8424
rect 18064 8421 18092 8520
rect 19334 8508 19340 8560
rect 19392 8548 19398 8560
rect 20364 8557 20392 8588
rect 21174 8576 21180 8588
rect 21232 8576 21238 8628
rect 22186 8616 22192 8628
rect 22147 8588 22192 8616
rect 22186 8576 22192 8588
rect 22244 8576 22250 8628
rect 22741 8619 22799 8625
rect 22741 8585 22753 8619
rect 22787 8616 22799 8619
rect 22922 8616 22928 8628
rect 22787 8588 22928 8616
rect 22787 8585 22799 8588
rect 22741 8579 22799 8585
rect 22922 8576 22928 8588
rect 22980 8576 22986 8628
rect 23658 8616 23664 8628
rect 23619 8588 23664 8616
rect 23658 8576 23664 8588
rect 23716 8576 23722 8628
rect 24946 8616 24952 8628
rect 24907 8588 24952 8616
rect 24946 8576 24952 8588
rect 25004 8576 25010 8628
rect 26142 8616 26148 8628
rect 26103 8588 26148 8616
rect 26142 8576 26148 8588
rect 26200 8576 26206 8628
rect 20349 8551 20407 8557
rect 20349 8548 20361 8551
rect 19392 8520 20361 8548
rect 19392 8508 19398 8520
rect 20349 8517 20361 8520
rect 20395 8517 20407 8551
rect 20349 8511 20407 8517
rect 22002 8440 22008 8492
rect 22060 8480 22066 8492
rect 22278 8480 22284 8492
rect 22060 8452 22284 8480
rect 22060 8440 22066 8452
rect 22278 8440 22284 8452
rect 22336 8480 22342 8492
rect 23109 8483 23167 8489
rect 23109 8480 23121 8483
rect 22336 8452 23121 8480
rect 22336 8440 22342 8452
rect 23109 8449 23121 8452
rect 23155 8480 23167 8483
rect 24213 8483 24271 8489
rect 24213 8480 24225 8483
rect 23155 8452 24225 8480
rect 23155 8449 23167 8452
rect 23109 8443 23167 8449
rect 24213 8449 24225 8452
rect 24259 8449 24271 8483
rect 24213 8443 24271 8449
rect 18049 8415 18107 8421
rect 18049 8381 18061 8415
rect 18095 8412 18107 8415
rect 18095 8384 18552 8412
rect 18095 8381 18107 8384
rect 18049 8375 18107 8381
rect 18524 8356 18552 8384
rect 20254 8372 20260 8424
rect 20312 8412 20318 8424
rect 20533 8415 20591 8421
rect 20533 8412 20545 8415
rect 20312 8384 20545 8412
rect 20312 8372 20318 8384
rect 20533 8381 20545 8384
rect 20579 8381 20591 8415
rect 20800 8415 20858 8421
rect 20800 8412 20812 8415
rect 20533 8375 20591 8381
rect 20732 8384 20812 8412
rect 14875 8316 15231 8344
rect 16761 8347 16819 8353
rect 14875 8313 14887 8316
rect 14829 8307 14887 8313
rect 16761 8313 16773 8347
rect 16807 8344 16819 8347
rect 16807 8316 17908 8344
rect 16807 8313 16819 8316
rect 16761 8307 16819 8313
rect 11146 8276 11152 8288
rect 10836 8248 11008 8276
rect 11107 8248 11152 8276
rect 10836 8236 10842 8248
rect 11146 8236 11152 8248
rect 11204 8236 11210 8288
rect 12434 8236 12440 8288
rect 12492 8276 12498 8288
rect 12492 8248 12537 8276
rect 12492 8236 12498 8248
rect 13906 8236 13912 8288
rect 13964 8276 13970 8288
rect 14090 8276 14096 8288
rect 13964 8248 14096 8276
rect 13964 8236 13970 8248
rect 14090 8236 14096 8248
rect 14148 8236 14154 8288
rect 14550 8236 14556 8288
rect 14608 8276 14614 8288
rect 15378 8276 15384 8288
rect 14608 8248 15384 8276
rect 14608 8236 14614 8248
rect 15378 8236 15384 8248
rect 15436 8236 15442 8288
rect 15746 8236 15752 8288
rect 15804 8276 15810 8288
rect 17310 8276 17316 8288
rect 15804 8248 17316 8276
rect 15804 8236 15810 8248
rect 17310 8236 17316 8248
rect 17368 8236 17374 8288
rect 17880 8276 17908 8316
rect 18138 8304 18144 8356
rect 18196 8344 18202 8356
rect 18294 8347 18352 8353
rect 18294 8344 18306 8347
rect 18196 8316 18306 8344
rect 18196 8304 18202 8316
rect 18294 8313 18306 8316
rect 18340 8313 18352 8347
rect 18294 8307 18352 8313
rect 18506 8304 18512 8356
rect 18564 8304 18570 8356
rect 18046 8276 18052 8288
rect 17880 8248 18052 8276
rect 18046 8236 18052 8248
rect 18104 8236 18110 8288
rect 19518 8236 19524 8288
rect 19576 8276 19582 8288
rect 19705 8279 19763 8285
rect 19705 8276 19717 8279
rect 19576 8248 19717 8276
rect 19576 8236 19582 8248
rect 19705 8245 19717 8248
rect 19751 8245 19763 8279
rect 20548 8276 20576 8375
rect 20732 8356 20760 8384
rect 20800 8381 20812 8384
rect 20846 8412 20858 8415
rect 21082 8412 21088 8424
rect 20846 8384 21088 8412
rect 20846 8381 20858 8384
rect 20800 8375 20858 8381
rect 21082 8372 21088 8384
rect 21140 8372 21146 8424
rect 24029 8415 24087 8421
rect 24029 8381 24041 8415
rect 24075 8412 24087 8415
rect 24118 8412 24124 8424
rect 24075 8384 24124 8412
rect 24075 8381 24087 8384
rect 24029 8375 24087 8381
rect 24118 8372 24124 8384
rect 24176 8372 24182 8424
rect 25130 8372 25136 8424
rect 25188 8412 25194 8424
rect 25225 8415 25283 8421
rect 25225 8412 25237 8415
rect 25188 8384 25237 8412
rect 25188 8372 25194 8384
rect 25225 8381 25237 8384
rect 25271 8412 25283 8415
rect 25777 8415 25835 8421
rect 25777 8412 25789 8415
rect 25271 8384 25789 8412
rect 25271 8381 25283 8384
rect 25225 8375 25283 8381
rect 25777 8381 25789 8384
rect 25823 8381 25835 8415
rect 25777 8375 25835 8381
rect 20714 8304 20720 8356
rect 20772 8304 20778 8356
rect 23477 8347 23535 8353
rect 23477 8313 23489 8347
rect 23523 8344 23535 8347
rect 23566 8344 23572 8356
rect 23523 8316 23572 8344
rect 23523 8313 23535 8316
rect 23477 8307 23535 8313
rect 23566 8304 23572 8316
rect 23624 8344 23630 8356
rect 24762 8344 24768 8356
rect 23624 8316 24768 8344
rect 23624 8304 23630 8316
rect 21726 8276 21732 8288
rect 20548 8248 21732 8276
rect 19705 8239 19763 8245
rect 21726 8236 21732 8248
rect 21784 8236 21790 8288
rect 21910 8276 21916 8288
rect 21871 8248 21916 8276
rect 21910 8236 21916 8248
rect 21968 8236 21974 8288
rect 24136 8285 24164 8316
rect 24762 8304 24768 8316
rect 24820 8304 24826 8356
rect 24121 8279 24179 8285
rect 24121 8245 24133 8279
rect 24167 8245 24179 8279
rect 24121 8239 24179 8245
rect 25409 8279 25467 8285
rect 25409 8245 25421 8279
rect 25455 8276 25467 8279
rect 25866 8276 25872 8288
rect 25455 8248 25872 8276
rect 25455 8245 25467 8248
rect 25409 8239 25467 8245
rect 25866 8236 25872 8248
rect 25924 8236 25930 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 2409 8075 2467 8081
rect 2409 8041 2421 8075
rect 2455 8072 2467 8075
rect 2498 8072 2504 8084
rect 2455 8044 2504 8072
rect 2455 8041 2467 8044
rect 2409 8035 2467 8041
rect 2498 8032 2504 8044
rect 2556 8032 2562 8084
rect 4801 8075 4859 8081
rect 4801 8041 4813 8075
rect 4847 8072 4859 8075
rect 5166 8072 5172 8084
rect 4847 8044 5172 8072
rect 4847 8041 4859 8044
rect 4801 8035 4859 8041
rect 5166 8032 5172 8044
rect 5224 8032 5230 8084
rect 6270 8072 6276 8084
rect 6231 8044 6276 8072
rect 6270 8032 6276 8044
rect 6328 8032 6334 8084
rect 7558 8072 7564 8084
rect 7519 8044 7564 8072
rect 7558 8032 7564 8044
rect 7616 8032 7622 8084
rect 7650 8032 7656 8084
rect 7708 8072 7714 8084
rect 8481 8075 8539 8081
rect 8481 8072 8493 8075
rect 7708 8044 8493 8072
rect 7708 8032 7714 8044
rect 8481 8041 8493 8044
rect 8527 8041 8539 8075
rect 8481 8035 8539 8041
rect 9122 8032 9128 8084
rect 9180 8072 9186 8084
rect 9401 8075 9459 8081
rect 9401 8072 9413 8075
rect 9180 8044 9413 8072
rect 9180 8032 9186 8044
rect 9401 8041 9413 8044
rect 9447 8041 9459 8075
rect 9401 8035 9459 8041
rect 10134 8032 10140 8084
rect 10192 8072 10198 8084
rect 10413 8075 10471 8081
rect 10413 8072 10425 8075
rect 10192 8044 10425 8072
rect 10192 8032 10198 8044
rect 10413 8041 10425 8044
rect 10459 8041 10471 8075
rect 10778 8072 10784 8084
rect 10739 8044 10784 8072
rect 10413 8035 10471 8041
rect 2774 7964 2780 8016
rect 2832 8004 2838 8016
rect 4433 8007 4491 8013
rect 2832 7976 2877 8004
rect 2832 7964 2838 7976
rect 4433 7973 4445 8007
rect 4479 8004 4491 8007
rect 5442 8004 5448 8016
rect 4479 7976 5448 8004
rect 4479 7973 4491 7976
rect 4433 7967 4491 7973
rect 5442 7964 5448 7976
rect 5500 7964 5506 8016
rect 8294 7964 8300 8016
rect 8352 8004 8358 8016
rect 8389 8007 8447 8013
rect 8389 8004 8401 8007
rect 8352 7976 8401 8004
rect 8352 7964 8358 7976
rect 8389 7973 8401 7976
rect 8435 8004 8447 8007
rect 9582 8004 9588 8016
rect 8435 7976 9588 8004
rect 8435 7973 8447 7976
rect 8389 7967 8447 7973
rect 9582 7964 9588 7976
rect 9640 7964 9646 8016
rect 2869 7939 2927 7945
rect 2869 7905 2881 7939
rect 2915 7936 2927 7939
rect 2915 7908 3188 7936
rect 2915 7905 2927 7908
rect 2869 7899 2927 7905
rect 3160 7880 3188 7908
rect 4982 7896 4988 7948
rect 5040 7936 5046 7948
rect 5160 7939 5218 7945
rect 5160 7936 5172 7939
rect 5040 7908 5172 7936
rect 5040 7896 5046 7908
rect 5160 7905 5172 7908
rect 5206 7936 5218 7939
rect 6454 7936 6460 7948
rect 5206 7908 6460 7936
rect 5206 7905 5218 7908
rect 5160 7899 5218 7905
rect 6454 7896 6460 7908
rect 6512 7896 6518 7948
rect 6914 7936 6920 7948
rect 6875 7908 6920 7936
rect 6914 7896 6920 7908
rect 6972 7896 6978 7948
rect 7098 7896 7104 7948
rect 7156 7936 7162 7948
rect 7285 7939 7343 7945
rect 7285 7936 7297 7939
rect 7156 7908 7297 7936
rect 7156 7896 7162 7908
rect 7285 7905 7297 7908
rect 7331 7905 7343 7939
rect 7285 7899 7343 7905
rect 8754 7896 8760 7948
rect 8812 7936 8818 7948
rect 9490 7936 9496 7948
rect 8812 7908 9496 7936
rect 8812 7896 8818 7908
rect 9490 7896 9496 7908
rect 9548 7896 9554 7948
rect 9858 7936 9864 7948
rect 9819 7908 9864 7936
rect 9858 7896 9864 7908
rect 9916 7896 9922 7948
rect 10428 7936 10456 8035
rect 10778 8032 10784 8044
rect 10836 8032 10842 8084
rect 12250 8032 12256 8084
rect 12308 8072 12314 8084
rect 12986 8072 12992 8084
rect 12308 8044 12992 8072
rect 12308 8032 12314 8044
rect 12986 8032 12992 8044
rect 13044 8032 13050 8084
rect 13173 8075 13231 8081
rect 13173 8041 13185 8075
rect 13219 8072 13231 8075
rect 13446 8072 13452 8084
rect 13219 8044 13452 8072
rect 13219 8041 13231 8044
rect 13173 8035 13231 8041
rect 13446 8032 13452 8044
rect 13504 8032 13510 8084
rect 14090 8032 14096 8084
rect 14148 8072 14154 8084
rect 14553 8075 14611 8081
rect 14553 8072 14565 8075
rect 14148 8044 14565 8072
rect 14148 8032 14154 8044
rect 14553 8041 14565 8044
rect 14599 8041 14611 8075
rect 14553 8035 14611 8041
rect 14826 8032 14832 8084
rect 14884 8072 14890 8084
rect 15013 8075 15071 8081
rect 15013 8072 15025 8075
rect 14884 8044 15025 8072
rect 14884 8032 14890 8044
rect 15013 8041 15025 8044
rect 15059 8041 15071 8075
rect 15013 8035 15071 8041
rect 15286 8032 15292 8084
rect 15344 8072 15350 8084
rect 15654 8072 15660 8084
rect 15344 8044 15660 8072
rect 15344 8032 15350 8044
rect 15654 8032 15660 8044
rect 15712 8032 15718 8084
rect 16117 8075 16175 8081
rect 16117 8041 16129 8075
rect 16163 8072 16175 8075
rect 16206 8072 16212 8084
rect 16163 8044 16212 8072
rect 16163 8041 16175 8044
rect 16117 8035 16175 8041
rect 16206 8032 16212 8044
rect 16264 8032 16270 8084
rect 16761 8075 16819 8081
rect 16761 8041 16773 8075
rect 16807 8072 16819 8075
rect 17862 8072 17868 8084
rect 16807 8044 17868 8072
rect 16807 8041 16819 8044
rect 16761 8035 16819 8041
rect 17862 8032 17868 8044
rect 17920 8032 17926 8084
rect 18138 8072 18144 8084
rect 18099 8044 18144 8072
rect 18138 8032 18144 8044
rect 18196 8072 18202 8084
rect 19518 8072 19524 8084
rect 18196 8044 19524 8072
rect 18196 8032 18202 8044
rect 19518 8032 19524 8044
rect 19576 8072 19582 8084
rect 19705 8075 19763 8081
rect 19705 8072 19717 8075
rect 19576 8044 19717 8072
rect 19576 8032 19582 8044
rect 19705 8041 19717 8044
rect 19751 8041 19763 8075
rect 20622 8072 20628 8084
rect 20583 8044 20628 8072
rect 19705 8035 19763 8041
rect 20622 8032 20628 8044
rect 20680 8032 20686 8084
rect 21542 8072 21548 8084
rect 21503 8044 21548 8072
rect 21542 8032 21548 8044
rect 21600 8032 21606 8084
rect 22922 8032 22928 8084
rect 22980 8072 22986 8084
rect 23201 8075 23259 8081
rect 23201 8072 23213 8075
rect 22980 8044 23213 8072
rect 22980 8032 22986 8044
rect 23201 8041 23213 8044
rect 23247 8041 23259 8075
rect 24026 8072 24032 8084
rect 23987 8044 24032 8072
rect 23201 8035 23259 8041
rect 24026 8032 24032 8044
rect 24084 8032 24090 8084
rect 25222 8032 25228 8084
rect 25280 8072 25286 8084
rect 25409 8075 25467 8081
rect 25409 8072 25421 8075
rect 25280 8044 25421 8072
rect 25280 8032 25286 8044
rect 25409 8041 25421 8044
rect 25455 8072 25467 8075
rect 25777 8075 25835 8081
rect 25777 8072 25789 8075
rect 25455 8044 25789 8072
rect 25455 8041 25467 8044
rect 25409 8035 25467 8041
rect 25777 8041 25789 8044
rect 25823 8072 25835 8075
rect 26142 8072 26148 8084
rect 25823 8044 26148 8072
rect 25823 8041 25835 8044
rect 25777 8035 25835 8041
rect 26142 8032 26148 8044
rect 26200 8032 26206 8084
rect 11232 8007 11290 8013
rect 11232 7973 11244 8007
rect 11278 8004 11290 8007
rect 11422 8004 11428 8016
rect 11278 7976 11428 8004
rect 11278 7973 11290 7976
rect 11232 7967 11290 7973
rect 11422 7964 11428 7976
rect 11480 7964 11486 8016
rect 12434 7964 12440 8016
rect 12492 8004 12498 8016
rect 13541 8007 13599 8013
rect 13541 8004 13553 8007
rect 12492 7976 13553 8004
rect 12492 7964 12498 7976
rect 13541 7973 13553 7976
rect 13587 8004 13599 8007
rect 13814 8004 13820 8016
rect 13587 7976 13820 8004
rect 13587 7973 13599 7976
rect 13541 7967 13599 7973
rect 13814 7964 13820 7976
rect 13872 7964 13878 8016
rect 16669 8007 16727 8013
rect 16669 7973 16681 8007
rect 16715 8004 16727 8007
rect 17126 8004 17132 8016
rect 16715 7976 17132 8004
rect 16715 7973 16727 7976
rect 16669 7967 16727 7973
rect 17126 7964 17132 7976
rect 17184 7964 17190 8016
rect 22094 8013 22100 8016
rect 22088 8004 22100 8013
rect 22055 7976 22100 8004
rect 22088 7967 22100 7976
rect 22094 7964 22100 7967
rect 22152 7964 22158 8016
rect 23750 7964 23756 8016
rect 23808 8004 23814 8016
rect 24489 8007 24547 8013
rect 24489 8004 24501 8007
rect 23808 7976 24501 8004
rect 23808 7964 23814 7976
rect 24489 7973 24501 7976
rect 24535 8004 24547 8007
rect 25041 8007 25099 8013
rect 25041 8004 25053 8007
rect 24535 7976 25053 8004
rect 24535 7973 24547 7976
rect 24489 7967 24547 7973
rect 25041 7973 25053 7976
rect 25087 7973 25099 8007
rect 25041 7967 25099 7973
rect 10778 7936 10784 7948
rect 10428 7908 10784 7936
rect 10778 7896 10784 7908
rect 10836 7936 10842 7948
rect 10965 7939 11023 7945
rect 10965 7936 10977 7939
rect 10836 7908 10977 7936
rect 10836 7896 10842 7908
rect 10965 7905 10977 7908
rect 11011 7905 11023 7939
rect 12342 7936 12348 7948
rect 10965 7899 11023 7905
rect 11072 7908 12348 7936
rect 2130 7828 2136 7880
rect 2188 7868 2194 7880
rect 2498 7868 2504 7880
rect 2188 7840 2504 7868
rect 2188 7828 2194 7840
rect 2498 7828 2504 7840
rect 2556 7828 2562 7880
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7837 3111 7871
rect 3053 7831 3111 7837
rect 2958 7760 2964 7812
rect 3016 7800 3022 7812
rect 3068 7800 3096 7831
rect 3142 7828 3148 7880
rect 3200 7828 3206 7880
rect 4890 7868 4896 7880
rect 4851 7840 4896 7868
rect 4890 7828 4896 7840
rect 4948 7828 4954 7880
rect 8665 7871 8723 7877
rect 8665 7837 8677 7871
rect 8711 7868 8723 7871
rect 8846 7868 8852 7880
rect 8711 7840 8852 7868
rect 8711 7837 8723 7840
rect 8665 7831 8723 7837
rect 8846 7828 8852 7840
rect 8904 7828 8910 7880
rect 11072 7868 11100 7908
rect 12342 7896 12348 7908
rect 12400 7896 12406 7948
rect 12710 7896 12716 7948
rect 12768 7936 12774 7948
rect 13446 7936 13452 7948
rect 12768 7908 13452 7936
rect 12768 7896 12774 7908
rect 13446 7896 13452 7908
rect 13504 7936 13510 7948
rect 15289 7939 15347 7945
rect 13504 7908 13768 7936
rect 13504 7896 13510 7908
rect 13630 7868 13636 7880
rect 10060 7840 11100 7868
rect 13591 7840 13636 7868
rect 3016 7772 3096 7800
rect 3016 7760 3022 7772
rect 7006 7760 7012 7812
rect 7064 7800 7070 7812
rect 7101 7803 7159 7809
rect 7101 7800 7113 7803
rect 7064 7772 7113 7800
rect 7064 7760 7070 7772
rect 7101 7769 7113 7772
rect 7147 7800 7159 7803
rect 9122 7800 9128 7812
rect 7147 7772 9128 7800
rect 7147 7769 7159 7772
rect 7101 7763 7159 7769
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 10060 7809 10088 7840
rect 13630 7828 13636 7840
rect 13688 7828 13694 7880
rect 13740 7877 13768 7908
rect 15289 7905 15301 7939
rect 15335 7936 15347 7939
rect 16022 7936 16028 7948
rect 15335 7908 16028 7936
rect 15335 7905 15347 7908
rect 15289 7899 15347 7905
rect 16022 7896 16028 7908
rect 16080 7896 16086 7948
rect 17221 7939 17279 7945
rect 17221 7905 17233 7939
rect 17267 7936 17279 7939
rect 17402 7936 17408 7948
rect 17267 7908 17408 7936
rect 17267 7905 17279 7908
rect 17221 7899 17279 7905
rect 17402 7896 17408 7908
rect 17460 7896 17466 7948
rect 18581 7939 18639 7945
rect 18581 7936 18593 7939
rect 18248 7908 18593 7936
rect 13725 7871 13783 7877
rect 13725 7837 13737 7871
rect 13771 7837 13783 7871
rect 15470 7868 15476 7880
rect 15431 7840 15476 7868
rect 13725 7831 13783 7837
rect 15470 7828 15476 7840
rect 15528 7828 15534 7880
rect 17310 7868 17316 7880
rect 17271 7840 17316 7868
rect 17310 7828 17316 7840
rect 17368 7868 17374 7880
rect 18248 7868 18276 7908
rect 18581 7905 18593 7908
rect 18627 7905 18639 7939
rect 18581 7899 18639 7905
rect 23290 7896 23296 7948
rect 23348 7936 23354 7948
rect 24397 7939 24455 7945
rect 23348 7908 24256 7936
rect 23348 7896 23354 7908
rect 17368 7840 18276 7868
rect 18325 7871 18383 7877
rect 17368 7828 17374 7840
rect 18325 7837 18337 7871
rect 18371 7837 18383 7871
rect 18325 7831 18383 7837
rect 10045 7803 10103 7809
rect 10045 7769 10057 7803
rect 10091 7769 10103 7803
rect 13648 7800 13676 7828
rect 14185 7803 14243 7809
rect 14185 7800 14197 7803
rect 13648 7772 14197 7800
rect 10045 7763 10103 7769
rect 14185 7769 14197 7772
rect 14231 7769 14243 7803
rect 14185 7763 14243 7769
rect 14274 7760 14280 7812
rect 14332 7800 14338 7812
rect 15286 7800 15292 7812
rect 14332 7772 15292 7800
rect 14332 7760 14338 7772
rect 15286 7760 15292 7772
rect 15344 7760 15350 7812
rect 1670 7732 1676 7744
rect 1631 7704 1676 7732
rect 1670 7692 1676 7704
rect 1728 7692 1734 7744
rect 2130 7732 2136 7744
rect 2091 7704 2136 7732
rect 2130 7692 2136 7704
rect 2188 7692 2194 7744
rect 3694 7732 3700 7744
rect 3655 7704 3700 7732
rect 3694 7692 3700 7704
rect 3752 7692 3758 7744
rect 7742 7692 7748 7744
rect 7800 7732 7806 7744
rect 8021 7735 8079 7741
rect 8021 7732 8033 7735
rect 7800 7704 8033 7732
rect 7800 7692 7806 7704
rect 8021 7701 8033 7704
rect 8067 7701 8079 7735
rect 8021 7695 8079 7701
rect 8846 7692 8852 7744
rect 8904 7732 8910 7744
rect 9033 7735 9091 7741
rect 9033 7732 9045 7735
rect 8904 7704 9045 7732
rect 8904 7692 8910 7704
rect 9033 7701 9045 7704
rect 9079 7701 9091 7735
rect 9033 7695 9091 7701
rect 12250 7692 12256 7744
rect 12308 7732 12314 7744
rect 12345 7735 12403 7741
rect 12345 7732 12357 7735
rect 12308 7704 12357 7732
rect 12308 7692 12314 7704
rect 12345 7701 12357 7704
rect 12391 7701 12403 7735
rect 12618 7732 12624 7744
rect 12579 7704 12624 7732
rect 12345 7695 12403 7701
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 12802 7692 12808 7744
rect 12860 7732 12866 7744
rect 12989 7735 13047 7741
rect 12989 7732 13001 7735
rect 12860 7704 13001 7732
rect 12860 7692 12866 7704
rect 12989 7701 13001 7704
rect 13035 7701 13047 7735
rect 18340 7732 18368 7831
rect 21726 7828 21732 7880
rect 21784 7868 21790 7880
rect 21821 7871 21879 7877
rect 21821 7868 21833 7871
rect 21784 7840 21833 7868
rect 21784 7828 21790 7840
rect 21821 7837 21833 7840
rect 21867 7837 21879 7871
rect 21821 7831 21879 7837
rect 23753 7871 23811 7877
rect 23753 7837 23765 7871
rect 23799 7868 23811 7871
rect 24118 7868 24124 7880
rect 23799 7840 24124 7868
rect 23799 7837 23811 7840
rect 23753 7831 23811 7837
rect 24118 7828 24124 7840
rect 24176 7828 24182 7880
rect 24228 7868 24256 7908
rect 24397 7905 24409 7939
rect 24443 7936 24455 7939
rect 24670 7936 24676 7948
rect 24443 7908 24676 7936
rect 24443 7905 24455 7908
rect 24397 7899 24455 7905
rect 24670 7896 24676 7908
rect 24728 7896 24734 7948
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 24228 7840 24593 7868
rect 24581 7837 24593 7840
rect 24627 7868 24639 7871
rect 24762 7868 24768 7880
rect 24627 7840 24768 7868
rect 24627 7837 24639 7840
rect 24581 7831 24639 7837
rect 24762 7828 24768 7840
rect 24820 7828 24826 7880
rect 18506 7732 18512 7744
rect 18340 7704 18512 7732
rect 12989 7695 13047 7701
rect 18506 7692 18512 7704
rect 18564 7692 18570 7744
rect 19426 7692 19432 7744
rect 19484 7732 19490 7744
rect 19981 7735 20039 7741
rect 19981 7732 19993 7735
rect 19484 7704 19993 7732
rect 19484 7692 19490 7704
rect 19981 7701 19993 7704
rect 20027 7701 20039 7735
rect 19981 7695 20039 7701
rect 20898 7692 20904 7744
rect 20956 7732 20962 7744
rect 21085 7735 21143 7741
rect 21085 7732 21097 7735
rect 20956 7704 21097 7732
rect 20956 7692 20962 7704
rect 21085 7701 21097 7704
rect 21131 7701 21143 7735
rect 21085 7695 21143 7701
rect 23934 7692 23940 7744
rect 23992 7732 23998 7744
rect 26234 7732 26240 7744
rect 23992 7704 26240 7732
rect 23992 7692 23998 7704
rect 26234 7692 26240 7704
rect 26292 7692 26298 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 2038 7528 2044 7540
rect 1999 7500 2044 7528
rect 2038 7488 2044 7500
rect 2096 7488 2102 7540
rect 7650 7488 7656 7540
rect 7708 7528 7714 7540
rect 7929 7531 7987 7537
rect 7929 7528 7941 7531
rect 7708 7500 7941 7528
rect 7708 7488 7714 7500
rect 7929 7497 7941 7500
rect 7975 7497 7987 7531
rect 9582 7528 9588 7540
rect 9543 7500 9588 7528
rect 7929 7491 7987 7497
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 9858 7528 9864 7540
rect 9819 7500 9864 7528
rect 9858 7488 9864 7500
rect 9916 7488 9922 7540
rect 10778 7528 10784 7540
rect 10739 7500 10784 7528
rect 10778 7488 10784 7500
rect 10836 7488 10842 7540
rect 11422 7488 11428 7540
rect 11480 7528 11486 7540
rect 11793 7531 11851 7537
rect 11793 7528 11805 7531
rect 11480 7500 11805 7528
rect 11480 7488 11486 7500
rect 11793 7497 11805 7500
rect 11839 7528 11851 7531
rect 11882 7528 11888 7540
rect 11839 7500 11888 7528
rect 11839 7497 11851 7500
rect 11793 7491 11851 7497
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 12250 7528 12256 7540
rect 12211 7500 12256 7528
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 12437 7531 12495 7537
rect 12437 7497 12449 7531
rect 12483 7528 12495 7531
rect 13630 7528 13636 7540
rect 12483 7500 13636 7528
rect 12483 7497 12495 7500
rect 12437 7491 12495 7497
rect 13630 7488 13636 7500
rect 13688 7488 13694 7540
rect 16022 7528 16028 7540
rect 15983 7500 16028 7528
rect 16022 7488 16028 7500
rect 16080 7488 16086 7540
rect 16393 7531 16451 7537
rect 16393 7497 16405 7531
rect 16439 7528 16451 7531
rect 17034 7528 17040 7540
rect 16439 7500 17040 7528
rect 16439 7497 16451 7500
rect 16393 7491 16451 7497
rect 658 7420 664 7472
rect 716 7460 722 7472
rect 1946 7460 1952 7472
rect 716 7432 1952 7460
rect 716 7420 722 7432
rect 1946 7420 1952 7432
rect 2004 7420 2010 7472
rect 2130 7420 2136 7472
rect 2188 7460 2194 7472
rect 4982 7460 4988 7472
rect 2188 7432 4988 7460
rect 2188 7420 2194 7432
rect 2700 7401 2728 7432
rect 4982 7420 4988 7432
rect 5040 7420 5046 7472
rect 6273 7463 6331 7469
rect 6273 7460 6285 7463
rect 5828 7432 6285 7460
rect 2685 7395 2743 7401
rect 2685 7361 2697 7395
rect 2731 7361 2743 7395
rect 2685 7355 2743 7361
rect 3694 7352 3700 7404
rect 3752 7392 3758 7404
rect 4249 7395 4307 7401
rect 4249 7392 4261 7395
rect 3752 7364 4261 7392
rect 3752 7352 3758 7364
rect 4249 7361 4261 7364
rect 4295 7392 4307 7395
rect 4890 7392 4896 7404
rect 4295 7364 4896 7392
rect 4295 7361 4307 7364
rect 4249 7355 4307 7361
rect 4890 7352 4896 7364
rect 4948 7392 4954 7404
rect 5828 7401 5856 7432
rect 6273 7429 6285 7432
rect 6319 7460 6331 7463
rect 6319 7432 7420 7460
rect 6319 7429 6331 7432
rect 6273 7423 6331 7429
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 4948 7364 5825 7392
rect 4948 7352 4954 7364
rect 5813 7361 5825 7364
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 6914 7352 6920 7404
rect 6972 7392 6978 7404
rect 7392 7401 7420 7432
rect 8294 7420 8300 7472
rect 8352 7460 8358 7472
rect 8846 7460 8852 7472
rect 8352 7432 8852 7460
rect 8352 7420 8358 7432
rect 8846 7420 8852 7432
rect 8904 7460 8910 7472
rect 8904 7432 9076 7460
rect 8904 7420 8910 7432
rect 7285 7395 7343 7401
rect 7285 7392 7297 7395
rect 6972 7364 7297 7392
rect 6972 7352 6978 7364
rect 7285 7361 7297 7364
rect 7331 7361 7343 7395
rect 7285 7355 7343 7361
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7392 7435 7395
rect 7558 7392 7564 7404
rect 7423 7364 7564 7392
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 7558 7352 7564 7364
rect 7616 7352 7622 7404
rect 8389 7395 8447 7401
rect 8389 7361 8401 7395
rect 8435 7392 8447 7395
rect 8938 7392 8944 7404
rect 8435 7364 8944 7392
rect 8435 7361 8447 7364
rect 8389 7355 8447 7361
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 9048 7401 9076 7432
rect 10042 7420 10048 7472
rect 10100 7460 10106 7472
rect 11054 7460 11060 7472
rect 10100 7432 11060 7460
rect 10100 7420 10106 7432
rect 11054 7420 11060 7432
rect 11112 7420 11118 7472
rect 11440 7401 11468 7488
rect 13446 7460 13452 7472
rect 13407 7432 13452 7460
rect 13446 7420 13452 7432
rect 13504 7420 13510 7472
rect 9033 7395 9091 7401
rect 9033 7361 9045 7395
rect 9079 7361 9091 7395
rect 9033 7355 9091 7361
rect 10321 7395 10379 7401
rect 10321 7361 10333 7395
rect 10367 7392 10379 7395
rect 11425 7395 11483 7401
rect 11425 7392 11437 7395
rect 10367 7364 11437 7392
rect 10367 7361 10379 7364
rect 10321 7355 10379 7361
rect 11425 7361 11437 7364
rect 11471 7361 11483 7395
rect 11425 7355 11483 7361
rect 12618 7352 12624 7404
rect 12676 7392 12682 7404
rect 12897 7395 12955 7401
rect 12897 7392 12909 7395
rect 12676 7364 12909 7392
rect 12676 7352 12682 7364
rect 12897 7361 12909 7364
rect 12943 7361 12955 7395
rect 12897 7355 12955 7361
rect 12986 7352 12992 7404
rect 13044 7392 13050 7404
rect 13044 7364 13089 7392
rect 13044 7352 13050 7364
rect 1949 7327 2007 7333
rect 1949 7293 1961 7327
rect 1995 7324 2007 7327
rect 2498 7324 2504 7336
rect 1995 7296 2504 7324
rect 1995 7293 2007 7296
rect 1949 7287 2007 7293
rect 2498 7284 2504 7296
rect 2556 7284 2562 7336
rect 3513 7327 3571 7333
rect 3513 7293 3525 7327
rect 3559 7324 3571 7327
rect 4062 7324 4068 7336
rect 3559 7296 4068 7324
rect 3559 7293 3571 7296
rect 3513 7287 3571 7293
rect 4062 7284 4068 7296
rect 4120 7284 4126 7336
rect 5077 7327 5135 7333
rect 5077 7293 5089 7327
rect 5123 7324 5135 7327
rect 5629 7327 5687 7333
rect 5629 7324 5641 7327
rect 5123 7296 5641 7324
rect 5123 7293 5135 7296
rect 5077 7287 5135 7293
rect 5629 7293 5641 7296
rect 5675 7324 5687 7327
rect 6362 7324 6368 7336
rect 5675 7296 6368 7324
rect 5675 7293 5687 7296
rect 5629 7287 5687 7293
rect 6362 7284 6368 7296
rect 6420 7284 6426 7336
rect 8570 7284 8576 7336
rect 8628 7324 8634 7336
rect 8849 7327 8907 7333
rect 8849 7324 8861 7327
rect 8628 7296 8861 7324
rect 8628 7284 8634 7296
rect 8849 7293 8861 7296
rect 8895 7293 8907 7327
rect 8849 7287 8907 7293
rect 10686 7284 10692 7336
rect 10744 7324 10750 7336
rect 11241 7327 11299 7333
rect 11241 7324 11253 7327
rect 10744 7296 11253 7324
rect 10744 7284 10750 7296
rect 11241 7293 11253 7296
rect 11287 7293 11299 7327
rect 11241 7287 11299 7293
rect 11330 7284 11336 7336
rect 11388 7324 11394 7336
rect 12802 7324 12808 7336
rect 11388 7296 12808 7324
rect 11388 7284 11394 7296
rect 12802 7284 12808 7296
rect 12860 7284 12866 7336
rect 14277 7327 14335 7333
rect 14277 7293 14289 7327
rect 14323 7324 14335 7327
rect 14826 7324 14832 7336
rect 14323 7296 14832 7324
rect 14323 7293 14335 7296
rect 14277 7287 14335 7293
rect 14826 7284 14832 7296
rect 14884 7284 14890 7336
rect 15010 7284 15016 7336
rect 15068 7324 15074 7336
rect 16390 7324 16396 7336
rect 15068 7296 16396 7324
rect 15068 7284 15074 7296
rect 16390 7284 16396 7296
rect 16448 7284 16454 7336
rect 16500 7333 16528 7500
rect 17034 7488 17040 7500
rect 17092 7488 17098 7540
rect 20806 7528 20812 7540
rect 20767 7500 20812 7528
rect 20806 7488 20812 7500
rect 20864 7488 20870 7540
rect 22094 7488 22100 7540
rect 22152 7528 22158 7540
rect 22189 7531 22247 7537
rect 22189 7528 22201 7531
rect 22152 7500 22201 7528
rect 22152 7488 22158 7500
rect 22189 7497 22201 7500
rect 22235 7497 22247 7531
rect 22189 7491 22247 7497
rect 23474 7488 23480 7540
rect 23532 7528 23538 7540
rect 23661 7531 23719 7537
rect 23661 7528 23673 7531
rect 23532 7500 23673 7528
rect 23532 7488 23538 7500
rect 23661 7497 23673 7500
rect 23707 7497 23719 7531
rect 23661 7491 23719 7497
rect 24762 7488 24768 7540
rect 24820 7528 24826 7540
rect 25041 7531 25099 7537
rect 25041 7528 25053 7531
rect 24820 7500 25053 7528
rect 24820 7488 24826 7500
rect 25041 7497 25053 7500
rect 25087 7497 25099 7531
rect 26142 7528 26148 7540
rect 26103 7500 26148 7528
rect 25041 7491 25099 7497
rect 26142 7488 26148 7500
rect 26200 7488 26206 7540
rect 20714 7460 20720 7472
rect 20675 7432 20720 7460
rect 20714 7420 20720 7432
rect 20772 7460 20778 7472
rect 20772 7432 21312 7460
rect 20772 7420 20778 7432
rect 18046 7352 18052 7404
rect 18104 7392 18110 7404
rect 21284 7401 21312 7432
rect 22462 7420 22468 7472
rect 22520 7460 22526 7472
rect 26602 7460 26608 7472
rect 22520 7432 26608 7460
rect 22520 7420 22526 7432
rect 26602 7420 26608 7432
rect 26660 7420 26666 7472
rect 18509 7395 18567 7401
rect 18509 7392 18521 7395
rect 18104 7364 18521 7392
rect 18104 7352 18110 7364
rect 18509 7361 18521 7364
rect 18555 7392 18567 7395
rect 21269 7395 21327 7401
rect 18555 7364 18736 7392
rect 18555 7361 18567 7364
rect 18509 7355 18567 7361
rect 16485 7327 16543 7333
rect 16485 7293 16497 7327
rect 16531 7293 16543 7327
rect 18598 7324 18604 7336
rect 18559 7296 18604 7324
rect 16485 7287 16543 7293
rect 18598 7284 18604 7296
rect 18656 7284 18662 7336
rect 18708 7324 18736 7364
rect 21269 7361 21281 7395
rect 21315 7361 21327 7395
rect 21269 7355 21327 7361
rect 21453 7395 21511 7401
rect 21453 7361 21465 7395
rect 21499 7392 21511 7395
rect 21542 7392 21548 7404
rect 21499 7364 21548 7392
rect 21499 7361 21511 7364
rect 21453 7355 21511 7361
rect 18868 7327 18926 7333
rect 18868 7324 18880 7327
rect 18708 7296 18880 7324
rect 18868 7293 18880 7296
rect 18914 7324 18926 7327
rect 21468 7324 21496 7355
rect 21542 7352 21548 7364
rect 21600 7392 21606 7404
rect 21821 7395 21879 7401
rect 21821 7392 21833 7395
rect 21600 7364 21833 7392
rect 21600 7352 21606 7364
rect 21821 7361 21833 7364
rect 21867 7392 21879 7395
rect 22094 7392 22100 7404
rect 21867 7364 22100 7392
rect 21867 7361 21879 7364
rect 21821 7355 21879 7361
rect 22094 7352 22100 7364
rect 22152 7352 22158 7404
rect 22554 7352 22560 7404
rect 22612 7392 22618 7404
rect 23290 7392 23296 7404
rect 22612 7364 23296 7392
rect 22612 7352 22618 7364
rect 23290 7352 23296 7364
rect 23348 7352 23354 7404
rect 23842 7352 23848 7404
rect 23900 7392 23906 7404
rect 24121 7395 24179 7401
rect 24121 7392 24133 7395
rect 23900 7364 24133 7392
rect 23900 7352 23906 7364
rect 24121 7361 24133 7364
rect 24167 7361 24179 7395
rect 24305 7395 24363 7401
rect 24305 7392 24317 7395
rect 24121 7355 24179 7361
rect 24228 7364 24317 7392
rect 18914 7296 21496 7324
rect 18914 7293 18926 7296
rect 18868 7287 18926 7293
rect 22002 7284 22008 7336
rect 22060 7324 22066 7336
rect 22465 7327 22523 7333
rect 22465 7324 22477 7327
rect 22060 7296 22477 7324
rect 22060 7284 22066 7296
rect 22465 7293 22477 7296
rect 22511 7324 22523 7327
rect 23017 7327 23075 7333
rect 23017 7324 23029 7327
rect 22511 7296 23029 7324
rect 22511 7293 22523 7296
rect 22465 7287 22523 7293
rect 23017 7293 23029 7296
rect 23063 7293 23075 7327
rect 23017 7287 23075 7293
rect 23750 7284 23756 7336
rect 23808 7324 23814 7336
rect 24228 7324 24256 7364
rect 24305 7361 24317 7364
rect 24351 7392 24363 7395
rect 24762 7392 24768 7404
rect 24351 7364 24768 7392
rect 24351 7361 24363 7364
rect 24305 7355 24363 7361
rect 24762 7352 24768 7364
rect 24820 7352 24826 7404
rect 23808 7296 24256 7324
rect 25225 7327 25283 7333
rect 23808 7284 23814 7296
rect 25225 7293 25237 7327
rect 25271 7324 25283 7327
rect 25777 7327 25835 7333
rect 25777 7324 25789 7327
rect 25271 7296 25789 7324
rect 25271 7293 25283 7296
rect 25225 7287 25283 7293
rect 25777 7293 25789 7296
rect 25823 7293 25835 7327
rect 25777 7287 25835 7293
rect 4154 7256 4160 7268
rect 3620 7228 4160 7256
rect 1946 7148 1952 7200
rect 2004 7188 2010 7200
rect 2409 7191 2467 7197
rect 2409 7188 2421 7191
rect 2004 7160 2421 7188
rect 2004 7148 2010 7160
rect 2409 7157 2421 7160
rect 2455 7157 2467 7191
rect 3142 7188 3148 7200
rect 3103 7160 3148 7188
rect 2409 7151 2467 7157
rect 3142 7148 3148 7160
rect 3200 7148 3206 7200
rect 3620 7197 3648 7228
rect 4154 7216 4160 7228
rect 4212 7216 4218 7268
rect 4709 7259 4767 7265
rect 4709 7225 4721 7259
rect 4755 7256 4767 7259
rect 5537 7259 5595 7265
rect 5537 7256 5549 7259
rect 4755 7228 5549 7256
rect 4755 7225 4767 7228
rect 4709 7219 4767 7225
rect 5537 7225 5549 7228
rect 5583 7256 5595 7259
rect 5994 7256 6000 7268
rect 5583 7228 6000 7256
rect 5583 7225 5595 7228
rect 5537 7219 5595 7225
rect 5994 7216 6000 7228
rect 6052 7216 6058 7268
rect 6549 7259 6607 7265
rect 6549 7225 6561 7259
rect 6595 7256 6607 7259
rect 7193 7259 7251 7265
rect 7193 7256 7205 7259
rect 6595 7228 7205 7256
rect 6595 7225 6607 7228
rect 6549 7219 6607 7225
rect 7193 7225 7205 7228
rect 7239 7256 7251 7259
rect 7374 7256 7380 7268
rect 7239 7228 7380 7256
rect 7239 7225 7251 7228
rect 7193 7219 7251 7225
rect 7374 7216 7380 7228
rect 7432 7216 7438 7268
rect 10597 7259 10655 7265
rect 10597 7225 10609 7259
rect 10643 7256 10655 7259
rect 11149 7259 11207 7265
rect 11149 7256 11161 7259
rect 10643 7228 11161 7256
rect 10643 7225 10655 7228
rect 10597 7219 10655 7225
rect 11149 7225 11161 7228
rect 11195 7256 11207 7259
rect 12066 7256 12072 7268
rect 11195 7228 12072 7256
rect 11195 7225 11207 7228
rect 11149 7219 11207 7225
rect 12066 7216 12072 7228
rect 12124 7216 12130 7268
rect 14185 7259 14243 7265
rect 14185 7225 14197 7259
rect 14231 7256 14243 7259
rect 14544 7259 14602 7265
rect 14544 7256 14556 7259
rect 14231 7228 14556 7256
rect 14231 7225 14243 7228
rect 14185 7219 14243 7225
rect 14544 7225 14556 7228
rect 14590 7256 14602 7259
rect 14734 7256 14740 7268
rect 14590 7228 14740 7256
rect 14590 7225 14602 7228
rect 14544 7219 14602 7225
rect 14734 7216 14740 7228
rect 14792 7216 14798 7268
rect 16758 7256 16764 7268
rect 16719 7228 16764 7256
rect 16758 7216 16764 7228
rect 16816 7216 16822 7268
rect 17310 7256 17316 7268
rect 17223 7228 17316 7256
rect 17310 7216 17316 7228
rect 17368 7256 17374 7268
rect 17865 7259 17923 7265
rect 17865 7256 17877 7259
rect 17368 7228 17877 7256
rect 17368 7216 17374 7228
rect 17865 7225 17877 7228
rect 17911 7256 17923 7259
rect 24029 7259 24087 7265
rect 24029 7256 24041 7259
rect 17911 7228 18644 7256
rect 17911 7225 17923 7228
rect 17865 7219 17923 7225
rect 3605 7191 3663 7197
rect 3605 7157 3617 7191
rect 3651 7157 3663 7191
rect 3970 7188 3976 7200
rect 3931 7160 3976 7188
rect 3605 7151 3663 7157
rect 3970 7148 3976 7160
rect 4028 7148 4034 7200
rect 5166 7188 5172 7200
rect 5127 7160 5172 7188
rect 5166 7148 5172 7160
rect 5224 7148 5230 7200
rect 6638 7148 6644 7200
rect 6696 7188 6702 7200
rect 6825 7191 6883 7197
rect 6825 7188 6837 7191
rect 6696 7160 6837 7188
rect 6696 7148 6702 7160
rect 6825 7157 6837 7160
rect 6871 7157 6883 7191
rect 8478 7188 8484 7200
rect 8439 7160 8484 7188
rect 6825 7151 6883 7157
rect 8478 7148 8484 7160
rect 8536 7148 8542 7200
rect 15194 7148 15200 7200
rect 15252 7188 15258 7200
rect 15654 7188 15660 7200
rect 15252 7160 15660 7188
rect 15252 7148 15258 7160
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 18616 7188 18644 7228
rect 23492 7228 24041 7256
rect 23492 7200 23520 7228
rect 24029 7225 24041 7228
rect 24075 7225 24087 7259
rect 24029 7219 24087 7225
rect 24118 7216 24124 7268
rect 24176 7256 24182 7268
rect 25240 7256 25268 7287
rect 24176 7228 25268 7256
rect 24176 7216 24182 7228
rect 19981 7191 20039 7197
rect 19981 7188 19993 7191
rect 18616 7160 19993 7188
rect 19981 7157 19993 7160
rect 20027 7188 20039 7191
rect 20070 7188 20076 7200
rect 20027 7160 20076 7188
rect 20027 7157 20039 7160
rect 19981 7151 20039 7157
rect 20070 7148 20076 7160
rect 20128 7148 20134 7200
rect 20346 7188 20352 7200
rect 20259 7160 20352 7188
rect 20346 7148 20352 7160
rect 20404 7188 20410 7200
rect 21177 7191 21235 7197
rect 21177 7188 21189 7191
rect 20404 7160 21189 7188
rect 20404 7148 20410 7160
rect 21177 7157 21189 7160
rect 21223 7157 21235 7191
rect 22646 7188 22652 7200
rect 22607 7160 22652 7188
rect 21177 7151 21235 7157
rect 22646 7148 22652 7160
rect 22704 7148 22710 7200
rect 23474 7188 23480 7200
rect 23435 7160 23480 7188
rect 23474 7148 23480 7160
rect 23532 7148 23538 7200
rect 25222 7148 25228 7200
rect 25280 7188 25286 7200
rect 25409 7191 25467 7197
rect 25409 7188 25421 7191
rect 25280 7160 25421 7188
rect 25280 7148 25286 7160
rect 25409 7157 25421 7160
rect 25455 7157 25467 7191
rect 25409 7151 25467 7157
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1762 6984 1768 6996
rect 1723 6956 1768 6984
rect 1762 6944 1768 6956
rect 1820 6944 1826 6996
rect 2774 6944 2780 6996
rect 2832 6984 2838 6996
rect 3237 6987 3295 6993
rect 3237 6984 3249 6987
rect 2832 6956 3249 6984
rect 2832 6944 2838 6956
rect 3237 6953 3249 6956
rect 3283 6953 3295 6987
rect 3237 6947 3295 6953
rect 3697 6987 3755 6993
rect 3697 6953 3709 6987
rect 3743 6984 3755 6987
rect 3970 6984 3976 6996
rect 3743 6956 3976 6984
rect 3743 6953 3755 6956
rect 3697 6947 3755 6953
rect 3970 6944 3976 6956
rect 4028 6944 4034 6996
rect 4982 6984 4988 6996
rect 4943 6956 4988 6984
rect 4982 6944 4988 6956
rect 5040 6944 5046 6996
rect 8570 6944 8576 6996
rect 8628 6984 8634 6996
rect 9033 6987 9091 6993
rect 9033 6984 9045 6987
rect 8628 6956 9045 6984
rect 8628 6944 8634 6956
rect 9033 6953 9045 6956
rect 9079 6953 9091 6987
rect 9033 6947 9091 6953
rect 9674 6944 9680 6996
rect 9732 6984 9738 6996
rect 10042 6984 10048 6996
rect 9732 6956 10048 6984
rect 9732 6944 9738 6956
rect 10042 6944 10048 6956
rect 10100 6944 10106 6996
rect 10870 6944 10876 6996
rect 10928 6984 10934 6996
rect 11149 6987 11207 6993
rect 11149 6984 11161 6987
rect 10928 6956 11161 6984
rect 10928 6944 10934 6956
rect 11149 6953 11161 6956
rect 11195 6953 11207 6987
rect 11330 6984 11336 6996
rect 11291 6956 11336 6984
rect 11149 6947 11207 6953
rect 11330 6944 11336 6956
rect 11388 6944 11394 6996
rect 11698 6984 11704 6996
rect 11659 6956 11704 6984
rect 11698 6944 11704 6956
rect 11756 6944 11762 6996
rect 11790 6944 11796 6996
rect 11848 6984 11854 6996
rect 12250 6984 12256 6996
rect 11848 6956 12256 6984
rect 11848 6944 11854 6956
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 14737 6987 14795 6993
rect 12912 6956 13860 6984
rect 6638 6916 6644 6928
rect 5552 6888 6644 6916
rect 2590 6848 2596 6860
rect 2551 6820 2596 6848
rect 2590 6808 2596 6820
rect 2648 6808 2654 6860
rect 4617 6851 4675 6857
rect 4617 6817 4629 6851
rect 4663 6848 4675 6851
rect 5350 6848 5356 6860
rect 4663 6820 5356 6848
rect 4663 6817 4675 6820
rect 4617 6811 4675 6817
rect 5350 6808 5356 6820
rect 5408 6848 5414 6860
rect 5552 6848 5580 6888
rect 6638 6876 6644 6888
rect 6696 6876 6702 6928
rect 8389 6919 8447 6925
rect 8389 6916 8401 6919
rect 6840 6888 8401 6916
rect 5408 6820 5580 6848
rect 5408 6808 5414 6820
rect 5626 6808 5632 6860
rect 5684 6848 5690 6860
rect 6840 6857 6868 6888
rect 8389 6885 8401 6888
rect 8435 6916 8447 6919
rect 8478 6916 8484 6928
rect 8435 6888 8484 6916
rect 8435 6885 8447 6888
rect 8389 6879 8447 6885
rect 8478 6876 8484 6888
rect 8536 6876 8542 6928
rect 12912 6860 12940 6956
rect 13265 6919 13323 6925
rect 13265 6885 13277 6919
rect 13311 6916 13323 6919
rect 13722 6916 13728 6928
rect 13311 6888 13728 6916
rect 13311 6885 13323 6888
rect 13265 6879 13323 6885
rect 13722 6876 13728 6888
rect 13780 6876 13786 6928
rect 13832 6916 13860 6956
rect 14737 6953 14749 6987
rect 14783 6984 14795 6987
rect 15010 6984 15016 6996
rect 14783 6956 15016 6984
rect 14783 6953 14795 6956
rect 14737 6947 14795 6953
rect 15010 6944 15016 6956
rect 15068 6944 15074 6996
rect 15105 6987 15163 6993
rect 15105 6953 15117 6987
rect 15151 6984 15163 6987
rect 15657 6987 15715 6993
rect 15657 6984 15669 6987
rect 15151 6956 15669 6984
rect 15151 6953 15163 6956
rect 15105 6947 15163 6953
rect 15657 6953 15669 6956
rect 15703 6984 15715 6987
rect 16206 6984 16212 6996
rect 15703 6956 16212 6984
rect 15703 6953 15715 6956
rect 15657 6947 15715 6953
rect 16206 6944 16212 6956
rect 16264 6944 16270 6996
rect 16853 6987 16911 6993
rect 16853 6953 16865 6987
rect 16899 6984 16911 6987
rect 17402 6984 17408 6996
rect 16899 6956 17408 6984
rect 16899 6953 16911 6956
rect 16853 6947 16911 6953
rect 17402 6944 17408 6956
rect 17460 6944 17466 6996
rect 17770 6984 17776 6996
rect 17731 6956 17776 6984
rect 17770 6944 17776 6956
rect 17828 6944 17834 6996
rect 20714 6984 20720 6996
rect 17972 6956 20720 6984
rect 14921 6919 14979 6925
rect 14921 6916 14933 6919
rect 13832 6888 14933 6916
rect 14921 6885 14933 6888
rect 14967 6885 14979 6919
rect 17972 6916 18000 6956
rect 20714 6944 20720 6956
rect 20772 6944 20778 6996
rect 23753 6987 23811 6993
rect 23753 6953 23765 6987
rect 23799 6984 23811 6987
rect 23842 6984 23848 6996
rect 23799 6956 23848 6984
rect 23799 6953 23811 6956
rect 23753 6947 23811 6953
rect 23842 6944 23848 6956
rect 23900 6944 23906 6996
rect 25869 6987 25927 6993
rect 25869 6953 25881 6987
rect 25915 6984 25927 6987
rect 26142 6984 26148 6996
rect 25915 6956 26148 6984
rect 25915 6953 25927 6956
rect 25869 6947 25927 6953
rect 26142 6944 26148 6956
rect 26200 6944 26206 6996
rect 19426 6916 19432 6928
rect 14921 6879 14979 6885
rect 15120 6888 18000 6916
rect 19387 6888 19432 6916
rect 6825 6851 6883 6857
rect 5684 6820 5729 6848
rect 5684 6808 5690 6820
rect 6825 6817 6837 6851
rect 6871 6817 6883 6851
rect 6825 6811 6883 6817
rect 6917 6851 6975 6857
rect 6917 6817 6929 6851
rect 6963 6848 6975 6851
rect 7006 6848 7012 6860
rect 6963 6820 7012 6848
rect 6963 6817 6975 6820
rect 6917 6811 6975 6817
rect 7006 6808 7012 6820
rect 7064 6808 7070 6860
rect 10686 6808 10692 6860
rect 10744 6848 10750 6860
rect 10781 6851 10839 6857
rect 10781 6848 10793 6851
rect 10744 6820 10793 6848
rect 10744 6808 10750 6820
rect 10781 6817 10793 6820
rect 10827 6817 10839 6851
rect 10781 6811 10839 6817
rect 11514 6808 11520 6860
rect 11572 6848 11578 6860
rect 11793 6851 11851 6857
rect 11793 6848 11805 6851
rect 11572 6820 11805 6848
rect 11572 6808 11578 6820
rect 11793 6817 11805 6820
rect 11839 6817 11851 6851
rect 11793 6811 11851 6817
rect 12618 6808 12624 6860
rect 12676 6848 12682 6860
rect 12894 6848 12900 6860
rect 12676 6820 12900 6848
rect 12676 6808 12682 6820
rect 12894 6808 12900 6820
rect 12952 6808 12958 6860
rect 13354 6808 13360 6860
rect 13412 6848 13418 6860
rect 13412 6820 13457 6848
rect 13412 6808 13418 6820
rect 13814 6808 13820 6860
rect 13872 6848 13878 6860
rect 14277 6851 14335 6857
rect 14277 6848 14289 6851
rect 13872 6820 14289 6848
rect 13872 6808 13878 6820
rect 14277 6817 14289 6820
rect 14323 6817 14335 6851
rect 14277 6811 14335 6817
rect 14829 6851 14887 6857
rect 14829 6817 14841 6851
rect 14875 6848 14887 6851
rect 15120 6848 15148 6888
rect 19426 6876 19432 6888
rect 19484 6876 19490 6928
rect 21358 6876 21364 6928
rect 21416 6916 21422 6928
rect 21416 6888 22324 6916
rect 21416 6876 21422 6888
rect 22296 6860 22324 6888
rect 22646 6876 22652 6928
rect 22704 6916 22710 6928
rect 24946 6916 24952 6928
rect 22704 6888 24952 6916
rect 22704 6876 22710 6888
rect 24946 6876 24952 6888
rect 25004 6876 25010 6928
rect 14875 6820 15148 6848
rect 15749 6851 15807 6857
rect 14875 6817 14887 6820
rect 14829 6811 14887 6817
rect 15749 6817 15761 6851
rect 15795 6848 15807 6851
rect 15930 6848 15936 6860
rect 15795 6820 15936 6848
rect 15795 6817 15807 6820
rect 15749 6811 15807 6817
rect 15930 6808 15936 6820
rect 15988 6848 15994 6860
rect 16482 6848 16488 6860
rect 15988 6820 16488 6848
rect 15988 6808 15994 6820
rect 16482 6808 16488 6820
rect 16540 6808 16546 6860
rect 17218 6848 17224 6860
rect 17179 6820 17224 6848
rect 17218 6808 17224 6820
rect 17276 6808 17282 6860
rect 17862 6848 17868 6860
rect 17823 6820 17868 6848
rect 17862 6808 17868 6820
rect 17920 6808 17926 6860
rect 21269 6851 21327 6857
rect 21269 6817 21281 6851
rect 21315 6848 21327 6851
rect 21818 6848 21824 6860
rect 21315 6820 21824 6848
rect 21315 6817 21327 6820
rect 21269 6811 21327 6817
rect 21818 6808 21824 6820
rect 21876 6808 21882 6860
rect 22278 6808 22284 6860
rect 22336 6848 22342 6860
rect 22833 6851 22891 6857
rect 22833 6848 22845 6851
rect 22336 6820 22845 6848
rect 22336 6808 22342 6820
rect 22833 6817 22845 6820
rect 22879 6817 22891 6851
rect 22833 6811 22891 6817
rect 24118 6808 24124 6860
rect 24176 6848 24182 6860
rect 24397 6851 24455 6857
rect 24397 6848 24409 6851
rect 24176 6820 24409 6848
rect 24176 6808 24182 6820
rect 24397 6817 24409 6820
rect 24443 6817 24455 6851
rect 24397 6811 24455 6817
rect 24489 6851 24547 6857
rect 24489 6817 24501 6851
rect 24535 6848 24547 6851
rect 24854 6848 24860 6860
rect 24535 6820 24860 6848
rect 24535 6817 24547 6820
rect 24489 6811 24547 6817
rect 2682 6780 2688 6792
rect 2643 6752 2688 6780
rect 2682 6740 2688 6752
rect 2740 6740 2746 6792
rect 2774 6740 2780 6792
rect 2832 6780 2838 6792
rect 2832 6752 2877 6780
rect 2832 6740 2838 6752
rect 5166 6740 5172 6792
rect 5224 6780 5230 6792
rect 5721 6783 5779 6789
rect 5721 6780 5733 6783
rect 5224 6752 5733 6780
rect 5224 6740 5230 6752
rect 5721 6749 5733 6752
rect 5767 6749 5779 6783
rect 5721 6743 5779 6749
rect 5905 6783 5963 6789
rect 5905 6749 5917 6783
rect 5951 6780 5963 6783
rect 5994 6780 6000 6792
rect 5951 6752 6000 6780
rect 5951 6749 5963 6752
rect 5905 6743 5963 6749
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 6457 6783 6515 6789
rect 6457 6749 6469 6783
rect 6503 6780 6515 6783
rect 7098 6780 7104 6792
rect 6503 6752 7104 6780
rect 6503 6749 6515 6752
rect 6457 6743 6515 6749
rect 7098 6740 7104 6752
rect 7156 6740 7162 6792
rect 8478 6780 8484 6792
rect 8439 6752 8484 6780
rect 8478 6740 8484 6752
rect 8536 6740 8542 6792
rect 8662 6780 8668 6792
rect 8623 6752 8668 6780
rect 8662 6740 8668 6752
rect 8720 6740 8726 6792
rect 9493 6783 9551 6789
rect 9493 6749 9505 6783
rect 9539 6780 9551 6783
rect 10134 6780 10140 6792
rect 9539 6752 10140 6780
rect 9539 6749 9551 6752
rect 9493 6743 9551 6749
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 10321 6783 10379 6789
rect 10321 6749 10333 6783
rect 10367 6749 10379 6783
rect 10321 6743 10379 6749
rect 2225 6715 2283 6721
rect 2225 6681 2237 6715
rect 2271 6712 2283 6715
rect 7190 6712 7196 6724
rect 2271 6684 7196 6712
rect 2271 6681 2283 6684
rect 2225 6675 2283 6681
rect 7190 6672 7196 6684
rect 7248 6672 7254 6724
rect 7558 6712 7564 6724
rect 7519 6684 7564 6712
rect 7558 6672 7564 6684
rect 7616 6672 7622 6724
rect 7929 6715 7987 6721
rect 7929 6681 7941 6715
rect 7975 6712 7987 6715
rect 8202 6712 8208 6724
rect 7975 6684 8208 6712
rect 7975 6681 7987 6684
rect 7929 6675 7987 6681
rect 8202 6672 8208 6684
rect 8260 6672 8266 6724
rect 10336 6712 10364 6743
rect 11882 6740 11888 6792
rect 11940 6780 11946 6792
rect 12805 6783 12863 6789
rect 11940 6752 11985 6780
rect 11940 6740 11946 6752
rect 12805 6749 12817 6783
rect 12851 6780 12863 6783
rect 13446 6780 13452 6792
rect 12851 6752 13452 6780
rect 12851 6749 12863 6752
rect 12805 6743 12863 6749
rect 13446 6740 13452 6752
rect 13504 6740 13510 6792
rect 14642 6740 14648 6792
rect 14700 6780 14706 6792
rect 15841 6783 15899 6789
rect 14700 6752 15700 6780
rect 14700 6740 14706 6752
rect 10778 6712 10784 6724
rect 10336 6684 10784 6712
rect 10778 6672 10784 6684
rect 10836 6672 10842 6724
rect 15102 6712 15108 6724
rect 14200 6684 15108 6712
rect 14200 6656 14228 6684
rect 15102 6672 15108 6684
rect 15160 6672 15166 6724
rect 15286 6712 15292 6724
rect 15247 6684 15292 6712
rect 15286 6672 15292 6684
rect 15344 6672 15350 6724
rect 15672 6712 15700 6752
rect 15841 6749 15853 6783
rect 15887 6749 15899 6783
rect 18046 6780 18052 6792
rect 17959 6752 18052 6780
rect 15841 6743 15899 6749
rect 15856 6712 15884 6743
rect 18046 6740 18052 6752
rect 18104 6780 18110 6792
rect 18966 6780 18972 6792
rect 18104 6752 18972 6780
rect 18104 6740 18110 6752
rect 18966 6740 18972 6752
rect 19024 6740 19030 6792
rect 19518 6780 19524 6792
rect 19479 6752 19524 6780
rect 19518 6740 19524 6752
rect 19576 6740 19582 6792
rect 19705 6783 19763 6789
rect 19705 6749 19717 6783
rect 19751 6780 19763 6783
rect 20070 6780 20076 6792
rect 19751 6752 20076 6780
rect 19751 6749 19763 6752
rect 19705 6743 19763 6749
rect 20070 6740 20076 6752
rect 20128 6740 20134 6792
rect 21358 6780 21364 6792
rect 21319 6752 21364 6780
rect 21358 6740 21364 6752
rect 21416 6740 21422 6792
rect 21542 6780 21548 6792
rect 21503 6752 21548 6780
rect 21542 6740 21548 6752
rect 21600 6740 21606 6792
rect 22094 6740 22100 6792
rect 22152 6780 22158 6792
rect 22922 6780 22928 6792
rect 22152 6752 22784 6780
rect 22883 6752 22928 6780
rect 22152 6740 22158 6752
rect 16482 6712 16488 6724
rect 15672 6684 16488 6712
rect 16482 6672 16488 6684
rect 16540 6672 16546 6724
rect 19061 6715 19119 6721
rect 19061 6681 19073 6715
rect 19107 6712 19119 6715
rect 19150 6712 19156 6724
rect 19107 6684 19156 6712
rect 19107 6681 19119 6684
rect 19061 6675 19119 6681
rect 19150 6672 19156 6684
rect 19208 6672 19214 6724
rect 22278 6712 22284 6724
rect 22239 6684 22284 6712
rect 22278 6672 22284 6684
rect 22336 6672 22342 6724
rect 22462 6712 22468 6724
rect 22423 6684 22468 6712
rect 22462 6672 22468 6684
rect 22520 6672 22526 6724
rect 22756 6712 22784 6752
rect 22922 6740 22928 6752
rect 22980 6740 22986 6792
rect 23017 6783 23075 6789
rect 23017 6749 23029 6783
rect 23063 6749 23075 6783
rect 23017 6743 23075 6749
rect 23032 6712 23060 6743
rect 23198 6740 23204 6792
rect 23256 6780 23262 6792
rect 24504 6780 24532 6811
rect 24854 6808 24860 6820
rect 24912 6808 24918 6860
rect 23256 6752 24532 6780
rect 24581 6783 24639 6789
rect 23256 6740 23262 6752
rect 24581 6749 24593 6783
rect 24627 6749 24639 6783
rect 24581 6743 24639 6749
rect 24026 6712 24032 6724
rect 22756 6684 23060 6712
rect 23987 6684 24032 6712
rect 24026 6672 24032 6684
rect 24084 6672 24090 6724
rect 24596 6712 24624 6743
rect 25041 6715 25099 6721
rect 25041 6712 25053 6715
rect 24504 6684 25053 6712
rect 1946 6604 1952 6656
rect 2004 6644 2010 6656
rect 2041 6647 2099 6653
rect 2041 6644 2053 6647
rect 2004 6616 2053 6644
rect 2004 6604 2010 6616
rect 2041 6613 2053 6616
rect 2087 6613 2099 6647
rect 5258 6644 5264 6656
rect 5219 6616 5264 6644
rect 2041 6607 2099 6613
rect 5258 6604 5264 6616
rect 5316 6604 5322 6656
rect 7098 6644 7104 6656
rect 7059 6616 7104 6644
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 8018 6644 8024 6656
rect 7979 6616 8024 6644
rect 8018 6604 8024 6616
rect 8076 6604 8082 6656
rect 8570 6604 8576 6656
rect 8628 6644 8634 6656
rect 9677 6647 9735 6653
rect 9677 6644 9689 6647
rect 8628 6616 9689 6644
rect 8628 6604 8634 6616
rect 9677 6613 9689 6616
rect 9723 6613 9735 6647
rect 9677 6607 9735 6613
rect 11882 6604 11888 6656
rect 11940 6644 11946 6656
rect 12066 6644 12072 6656
rect 11940 6616 12072 6644
rect 11940 6604 11946 6616
rect 12066 6604 12072 6616
rect 12124 6604 12130 6656
rect 12437 6647 12495 6653
rect 12437 6613 12449 6647
rect 12483 6644 12495 6647
rect 12710 6644 12716 6656
rect 12483 6616 12716 6644
rect 12483 6613 12495 6616
rect 12437 6607 12495 6613
rect 12710 6604 12716 6616
rect 12768 6604 12774 6656
rect 12897 6647 12955 6653
rect 12897 6613 12909 6647
rect 12943 6644 12955 6647
rect 13078 6644 13084 6656
rect 12943 6616 13084 6644
rect 12943 6613 12955 6616
rect 12897 6607 12955 6613
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 14001 6647 14059 6653
rect 14001 6613 14013 6647
rect 14047 6644 14059 6647
rect 14182 6644 14188 6656
rect 14047 6616 14188 6644
rect 14047 6613 14059 6616
rect 14001 6607 14059 6613
rect 14182 6604 14188 6616
rect 14240 6604 14246 6656
rect 14274 6604 14280 6656
rect 14332 6644 14338 6656
rect 14829 6647 14887 6653
rect 14829 6644 14841 6647
rect 14332 6616 14841 6644
rect 14332 6604 14338 6616
rect 14829 6613 14841 6616
rect 14875 6613 14887 6647
rect 14829 6607 14887 6613
rect 14921 6647 14979 6653
rect 14921 6613 14933 6647
rect 14967 6644 14979 6647
rect 16298 6644 16304 6656
rect 14967 6616 16304 6644
rect 14967 6613 14979 6616
rect 14921 6607 14979 6613
rect 16298 6604 16304 6616
rect 16356 6604 16362 6656
rect 17402 6644 17408 6656
rect 17363 6616 17408 6644
rect 17402 6604 17408 6616
rect 17460 6604 17466 6656
rect 18506 6644 18512 6656
rect 18467 6616 18512 6644
rect 18506 6604 18512 6616
rect 18564 6604 18570 6656
rect 18782 6644 18788 6656
rect 18743 6616 18788 6644
rect 18782 6604 18788 6616
rect 18840 6604 18846 6656
rect 19978 6604 19984 6656
rect 20036 6644 20042 6656
rect 20073 6647 20131 6653
rect 20073 6644 20085 6647
rect 20036 6616 20085 6644
rect 20036 6604 20042 6616
rect 20073 6613 20085 6616
rect 20119 6613 20131 6647
rect 20073 6607 20131 6613
rect 20533 6647 20591 6653
rect 20533 6613 20545 6647
rect 20579 6644 20591 6647
rect 20622 6644 20628 6656
rect 20579 6616 20628 6644
rect 20579 6613 20591 6616
rect 20533 6607 20591 6613
rect 20622 6604 20628 6616
rect 20680 6604 20686 6656
rect 20901 6647 20959 6653
rect 20901 6613 20913 6647
rect 20947 6644 20959 6647
rect 20990 6644 20996 6656
rect 20947 6616 20996 6644
rect 20947 6613 20959 6616
rect 20901 6607 20959 6613
rect 20990 6604 20996 6616
rect 21048 6604 21054 6656
rect 21910 6644 21916 6656
rect 21871 6616 21916 6644
rect 21910 6604 21916 6616
rect 21968 6604 21974 6656
rect 22186 6604 22192 6656
rect 22244 6644 22250 6656
rect 24504 6644 24532 6684
rect 25041 6681 25053 6684
rect 25087 6712 25099 6715
rect 25130 6712 25136 6724
rect 25087 6684 25136 6712
rect 25087 6681 25099 6684
rect 25041 6675 25099 6681
rect 25130 6672 25136 6684
rect 25188 6672 25194 6724
rect 25406 6644 25412 6656
rect 22244 6616 24532 6644
rect 25367 6616 25412 6644
rect 22244 6604 22250 6616
rect 25406 6604 25412 6616
rect 25464 6604 25470 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 1949 6443 2007 6449
rect 1949 6409 1961 6443
rect 1995 6440 2007 6443
rect 2590 6440 2596 6452
rect 1995 6412 2596 6440
rect 1995 6409 2007 6412
rect 1949 6403 2007 6409
rect 2590 6400 2596 6412
rect 2648 6400 2654 6452
rect 4154 6400 4160 6452
rect 4212 6440 4218 6452
rect 4433 6443 4491 6449
rect 4433 6440 4445 6443
rect 4212 6412 4445 6440
rect 4212 6400 4218 6412
rect 4433 6409 4445 6412
rect 4479 6440 4491 6443
rect 6641 6443 6699 6449
rect 4479 6412 5488 6440
rect 4479 6409 4491 6412
rect 4433 6403 4491 6409
rect 2317 6375 2375 6381
rect 2317 6341 2329 6375
rect 2363 6372 2375 6375
rect 2685 6375 2743 6381
rect 2685 6372 2697 6375
rect 2363 6344 2697 6372
rect 2363 6341 2375 6344
rect 2317 6335 2375 6341
rect 2685 6341 2697 6344
rect 2731 6372 2743 6375
rect 2774 6372 2780 6384
rect 2731 6344 2780 6372
rect 2731 6341 2743 6344
rect 2685 6335 2743 6341
rect 2774 6332 2780 6344
rect 2832 6332 2838 6384
rect 5460 6313 5488 6412
rect 6641 6409 6653 6443
rect 6687 6440 6699 6443
rect 7006 6440 7012 6452
rect 6687 6412 7012 6440
rect 6687 6409 6699 6412
rect 6641 6403 6699 6409
rect 7006 6400 7012 6412
rect 7064 6400 7070 6452
rect 9674 6440 9680 6452
rect 9635 6412 9680 6440
rect 9674 6400 9680 6412
rect 9732 6400 9738 6452
rect 11514 6440 11520 6452
rect 11475 6412 11520 6440
rect 11514 6400 11520 6412
rect 11572 6400 11578 6452
rect 11698 6400 11704 6452
rect 11756 6440 11762 6452
rect 11885 6443 11943 6449
rect 11885 6440 11897 6443
rect 11756 6412 11897 6440
rect 11756 6400 11762 6412
rect 11885 6409 11897 6412
rect 11931 6409 11943 6443
rect 13354 6440 13360 6452
rect 13315 6412 13360 6440
rect 11885 6403 11943 6409
rect 13354 6400 13360 6412
rect 13412 6400 13418 6452
rect 13722 6400 13728 6452
rect 13780 6440 13786 6452
rect 13817 6443 13875 6449
rect 13817 6440 13829 6443
rect 13780 6412 13829 6440
rect 13780 6400 13786 6412
rect 13817 6409 13829 6412
rect 13863 6440 13875 6443
rect 14274 6440 14280 6452
rect 13863 6412 14280 6440
rect 13863 6409 13875 6412
rect 13817 6403 13875 6409
rect 14274 6400 14280 6412
rect 14332 6400 14338 6452
rect 15562 6400 15568 6452
rect 15620 6440 15626 6452
rect 16117 6443 16175 6449
rect 16117 6440 16129 6443
rect 15620 6412 16129 6440
rect 15620 6400 15626 6412
rect 16117 6409 16129 6412
rect 16163 6409 16175 6443
rect 16117 6403 16175 6409
rect 17497 6443 17555 6449
rect 17497 6409 17509 6443
rect 17543 6440 17555 6443
rect 17862 6440 17868 6452
rect 17543 6412 17868 6440
rect 17543 6409 17555 6412
rect 17497 6403 17555 6409
rect 17862 6400 17868 6412
rect 17920 6400 17926 6452
rect 19150 6440 19156 6452
rect 19111 6412 19156 6440
rect 19150 6400 19156 6412
rect 19208 6400 19214 6452
rect 21361 6443 21419 6449
rect 21361 6409 21373 6443
rect 21407 6440 21419 6443
rect 21634 6440 21640 6452
rect 21407 6412 21640 6440
rect 21407 6409 21419 6412
rect 21361 6403 21419 6409
rect 21634 6400 21640 6412
rect 21692 6400 21698 6452
rect 21729 6443 21787 6449
rect 21729 6409 21741 6443
rect 21775 6440 21787 6443
rect 22002 6440 22008 6452
rect 21775 6412 22008 6440
rect 21775 6409 21787 6412
rect 21729 6403 21787 6409
rect 22002 6400 22008 6412
rect 22060 6440 22066 6452
rect 23661 6443 23719 6449
rect 22060 6412 22324 6440
rect 22060 6400 22066 6412
rect 11241 6375 11299 6381
rect 11241 6341 11253 6375
rect 11287 6372 11299 6375
rect 11330 6372 11336 6384
rect 11287 6344 11336 6372
rect 11287 6341 11299 6344
rect 11241 6335 11299 6341
rect 11330 6332 11336 6344
rect 11388 6372 11394 6384
rect 11790 6372 11796 6384
rect 11388 6344 11796 6372
rect 11388 6332 11394 6344
rect 11790 6332 11796 6344
rect 11848 6332 11854 6384
rect 15010 6332 15016 6384
rect 15068 6372 15074 6384
rect 15657 6375 15715 6381
rect 15657 6372 15669 6375
rect 15068 6344 15669 6372
rect 15068 6332 15074 6344
rect 15657 6341 15669 6344
rect 15703 6372 15715 6375
rect 15930 6372 15936 6384
rect 15703 6344 15936 6372
rect 15703 6341 15715 6344
rect 15657 6335 15715 6341
rect 15930 6332 15936 6344
rect 15988 6332 15994 6384
rect 17126 6332 17132 6384
rect 17184 6372 17190 6384
rect 18049 6375 18107 6381
rect 18049 6372 18061 6375
rect 17184 6344 18061 6372
rect 17184 6332 17190 6344
rect 18049 6341 18061 6344
rect 18095 6372 18107 6375
rect 19242 6372 19248 6384
rect 18095 6344 19248 6372
rect 18095 6341 18107 6344
rect 18049 6335 18107 6341
rect 19242 6332 19248 6344
rect 19300 6332 19306 6384
rect 5445 6307 5503 6313
rect 5445 6273 5457 6307
rect 5491 6273 5503 6307
rect 5445 6267 5503 6273
rect 5629 6307 5687 6313
rect 5629 6273 5641 6307
rect 5675 6304 5687 6307
rect 5994 6304 6000 6316
rect 5675 6276 6000 6304
rect 5675 6273 5687 6276
rect 5629 6267 5687 6273
rect 5994 6264 6000 6276
rect 6052 6264 6058 6316
rect 8570 6304 8576 6316
rect 8531 6276 8576 6304
rect 8570 6264 8576 6276
rect 8628 6264 8634 6316
rect 8662 6264 8668 6316
rect 8720 6304 8726 6316
rect 8720 6276 8813 6304
rect 8720 6264 8726 6276
rect 1762 6196 1768 6248
rect 1820 6236 1826 6248
rect 2777 6239 2835 6245
rect 2777 6236 2789 6239
rect 1820 6208 2789 6236
rect 1820 6196 1826 6208
rect 2777 6205 2789 6208
rect 2823 6236 2835 6239
rect 3602 6236 3608 6248
rect 2823 6208 3608 6236
rect 2823 6205 2835 6208
rect 2777 6199 2835 6205
rect 3602 6196 3608 6208
rect 3660 6196 3666 6248
rect 4982 6236 4988 6248
rect 4172 6208 4988 6236
rect 2958 6128 2964 6180
rect 3016 6177 3022 6180
rect 3016 6171 3080 6177
rect 3016 6137 3034 6171
rect 3068 6137 3080 6171
rect 3016 6131 3080 6137
rect 3016 6128 3022 6131
rect 4172 6109 4200 6208
rect 4982 6196 4988 6208
rect 5040 6196 5046 6248
rect 5350 6236 5356 6248
rect 5311 6208 5356 6236
rect 5350 6196 5356 6208
rect 5408 6196 5414 6248
rect 7009 6239 7067 6245
rect 7009 6205 7021 6239
rect 7055 6236 7067 6239
rect 7558 6236 7564 6248
rect 7055 6208 7564 6236
rect 7055 6205 7067 6208
rect 7009 6199 7067 6205
rect 7558 6196 7564 6208
rect 7616 6196 7622 6248
rect 8386 6196 8392 6248
rect 8444 6236 8450 6248
rect 8481 6239 8539 6245
rect 8481 6236 8493 6239
rect 8444 6208 8493 6236
rect 8444 6196 8450 6208
rect 8481 6205 8493 6208
rect 8527 6205 8539 6239
rect 8680 6236 8708 6264
rect 8481 6199 8539 6205
rect 8588 6208 8708 6236
rect 8588 6168 8616 6208
rect 9674 6196 9680 6248
rect 9732 6236 9738 6248
rect 9861 6239 9919 6245
rect 9861 6236 9873 6239
rect 9732 6208 9873 6236
rect 9732 6196 9738 6208
rect 9861 6205 9873 6208
rect 9907 6236 9919 6239
rect 10870 6236 10876 6248
rect 9907 6208 10876 6236
rect 9907 6205 9919 6208
rect 9861 6199 9919 6205
rect 10870 6196 10876 6208
rect 10928 6196 10934 6248
rect 12621 6239 12679 6245
rect 12621 6205 12633 6239
rect 12667 6236 12679 6239
rect 12710 6236 12716 6248
rect 12667 6208 12716 6236
rect 12667 6205 12679 6208
rect 12621 6199 12679 6205
rect 12710 6196 12716 6208
rect 12768 6196 12774 6248
rect 14182 6245 14188 6248
rect 13909 6239 13967 6245
rect 13909 6205 13921 6239
rect 13955 6205 13967 6239
rect 14176 6236 14188 6245
rect 14143 6208 14188 6236
rect 13909 6199 13967 6205
rect 14176 6199 14188 6208
rect 7944 6140 8616 6168
rect 9401 6171 9459 6177
rect 4157 6103 4215 6109
rect 4157 6069 4169 6103
rect 4203 6069 4215 6103
rect 4798 6100 4804 6112
rect 4759 6072 4804 6100
rect 4157 6063 4215 6069
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 4982 6100 4988 6112
rect 4943 6072 4988 6100
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 5994 6100 6000 6112
rect 5955 6072 6000 6100
rect 5994 6060 6000 6072
rect 6052 6060 6058 6112
rect 7190 6100 7196 6112
rect 7151 6072 7196 6100
rect 7190 6060 7196 6072
rect 7248 6060 7254 6112
rect 7650 6100 7656 6112
rect 7611 6072 7656 6100
rect 7650 6060 7656 6072
rect 7708 6100 7714 6112
rect 7944 6109 7972 6140
rect 9401 6137 9413 6171
rect 9447 6168 9459 6171
rect 10106 6171 10164 6177
rect 10106 6168 10118 6171
rect 9447 6140 10118 6168
rect 9447 6137 9459 6140
rect 9401 6131 9459 6137
rect 9876 6112 9904 6140
rect 10106 6137 10118 6140
rect 10152 6168 10164 6171
rect 11054 6168 11060 6180
rect 10152 6140 11060 6168
rect 10152 6137 10164 6140
rect 10106 6131 10164 6137
rect 11054 6128 11060 6140
rect 11112 6128 11118 6180
rect 12894 6168 12900 6180
rect 12855 6140 12900 6168
rect 12894 6128 12900 6140
rect 12952 6128 12958 6180
rect 13924 6168 13952 6199
rect 14182 6196 14188 6199
rect 14240 6196 14246 6248
rect 15948 6236 15976 6332
rect 16298 6264 16304 6316
rect 16356 6304 16362 6316
rect 16669 6307 16727 6313
rect 16669 6304 16681 6307
rect 16356 6276 16681 6304
rect 16356 6264 16362 6276
rect 16669 6273 16681 6276
rect 16715 6273 16727 6307
rect 16669 6267 16727 6273
rect 18506 6264 18512 6316
rect 18564 6304 18570 6316
rect 18693 6307 18751 6313
rect 18693 6304 18705 6307
rect 18564 6276 18705 6304
rect 18564 6264 18570 6276
rect 18693 6273 18705 6276
rect 18739 6304 18751 6307
rect 19150 6304 19156 6316
rect 18739 6276 19156 6304
rect 18739 6273 18751 6276
rect 18693 6267 18751 6273
rect 19150 6264 19156 6276
rect 19208 6264 19214 6316
rect 22296 6313 22324 6412
rect 23661 6409 23673 6443
rect 23707 6440 23719 6443
rect 24670 6440 24676 6452
rect 23707 6412 24676 6440
rect 23707 6409 23719 6412
rect 23661 6403 23719 6409
rect 24670 6400 24676 6412
rect 24728 6440 24734 6452
rect 25406 6440 25412 6452
rect 24728 6412 25412 6440
rect 24728 6400 24734 6412
rect 25406 6400 25412 6412
rect 25464 6400 25470 6452
rect 25590 6400 25596 6452
rect 25648 6440 25654 6452
rect 26145 6443 26203 6449
rect 26145 6440 26157 6443
rect 25648 6412 26157 6440
rect 25648 6400 25654 6412
rect 26145 6409 26157 6412
rect 26191 6409 26203 6443
rect 26145 6403 26203 6409
rect 24765 6375 24823 6381
rect 24765 6341 24777 6375
rect 24811 6372 24823 6375
rect 24854 6372 24860 6384
rect 24811 6344 24860 6372
rect 24811 6341 24823 6344
rect 24765 6335 24823 6341
rect 24854 6332 24860 6344
rect 24912 6372 24918 6384
rect 26234 6372 26240 6384
rect 24912 6344 26240 6372
rect 24912 6332 24918 6344
rect 26234 6332 26240 6344
rect 26292 6332 26298 6384
rect 22281 6307 22339 6313
rect 22281 6273 22293 6307
rect 22327 6273 22339 6307
rect 22281 6267 22339 6273
rect 22465 6307 22523 6313
rect 22465 6273 22477 6307
rect 22511 6273 22523 6307
rect 22465 6267 22523 6273
rect 16577 6239 16635 6245
rect 16577 6236 16589 6239
rect 15948 6208 16589 6236
rect 16577 6205 16589 6208
rect 16623 6205 16635 6239
rect 16577 6199 16635 6205
rect 19613 6239 19671 6245
rect 19613 6205 19625 6239
rect 19659 6236 19671 6239
rect 20254 6236 20260 6248
rect 19659 6208 20260 6236
rect 19659 6205 19671 6208
rect 19613 6199 19671 6205
rect 20254 6196 20260 6208
rect 20312 6196 20318 6248
rect 21910 6196 21916 6248
rect 21968 6236 21974 6248
rect 21968 6208 22324 6236
rect 21968 6196 21974 6208
rect 14826 6168 14832 6180
rect 13924 6140 14832 6168
rect 14826 6128 14832 6140
rect 14884 6128 14890 6180
rect 16022 6168 16028 6180
rect 14936 6140 16028 6168
rect 7929 6103 7987 6109
rect 7929 6100 7941 6103
rect 7708 6072 7941 6100
rect 7708 6060 7714 6072
rect 7929 6069 7941 6072
rect 7975 6069 7987 6103
rect 8110 6100 8116 6112
rect 8071 6072 8116 6100
rect 7929 6063 7987 6069
rect 8110 6060 8116 6072
rect 8168 6060 8174 6112
rect 9858 6060 9864 6112
rect 9916 6060 9922 6112
rect 13630 6060 13636 6112
rect 13688 6100 13694 6112
rect 14936 6100 14964 6140
rect 16022 6128 16028 6140
rect 16080 6168 16086 6180
rect 16080 6140 17908 6168
rect 16080 6128 16086 6140
rect 15286 6100 15292 6112
rect 13688 6072 14964 6100
rect 15247 6072 15292 6100
rect 13688 6060 13694 6072
rect 15286 6060 15292 6072
rect 15344 6060 15350 6112
rect 15930 6100 15936 6112
rect 15891 6072 15936 6100
rect 15930 6060 15936 6072
rect 15988 6100 15994 6112
rect 17880 6109 17908 6140
rect 17954 6128 17960 6180
rect 18012 6168 18018 6180
rect 18509 6171 18567 6177
rect 18509 6168 18521 6171
rect 18012 6140 18521 6168
rect 18012 6128 18018 6140
rect 18509 6137 18521 6140
rect 18555 6168 18567 6171
rect 18782 6168 18788 6180
rect 18555 6140 18788 6168
rect 18555 6137 18567 6140
rect 18509 6131 18567 6137
rect 18782 6128 18788 6140
rect 18840 6128 18846 6180
rect 19858 6171 19916 6177
rect 19858 6168 19870 6171
rect 19536 6140 19870 6168
rect 19536 6112 19564 6140
rect 19858 6137 19870 6140
rect 19904 6137 19916 6171
rect 19858 6131 19916 6137
rect 21634 6128 21640 6180
rect 21692 6168 21698 6180
rect 22189 6171 22247 6177
rect 22189 6168 22201 6171
rect 21692 6140 22201 6168
rect 21692 6128 21698 6140
rect 22189 6137 22201 6140
rect 22235 6137 22247 6171
rect 22296 6168 22324 6208
rect 22370 6168 22376 6180
rect 22283 6140 22376 6168
rect 22189 6131 22247 6137
rect 22370 6128 22376 6140
rect 22428 6168 22434 6180
rect 22480 6168 22508 6267
rect 23750 6264 23756 6316
rect 23808 6304 23814 6316
rect 24213 6307 24271 6313
rect 24213 6304 24225 6307
rect 23808 6276 24225 6304
rect 23808 6264 23814 6276
rect 24213 6273 24225 6276
rect 24259 6304 24271 6307
rect 25041 6307 25099 6313
rect 25041 6304 25053 6307
rect 24259 6276 25053 6304
rect 24259 6273 24271 6276
rect 24213 6267 24271 6273
rect 25041 6273 25053 6276
rect 25087 6273 25099 6307
rect 25041 6267 25099 6273
rect 23658 6196 23664 6248
rect 23716 6236 23722 6248
rect 24029 6239 24087 6245
rect 24029 6236 24041 6239
rect 23716 6208 24041 6236
rect 23716 6196 23722 6208
rect 24029 6205 24041 6208
rect 24075 6205 24087 6239
rect 24029 6199 24087 6205
rect 24854 6196 24860 6248
rect 24912 6236 24918 6248
rect 25225 6239 25283 6245
rect 25225 6236 25237 6239
rect 24912 6208 25237 6236
rect 24912 6196 24918 6208
rect 25225 6205 25237 6208
rect 25271 6236 25283 6239
rect 25777 6239 25835 6245
rect 25777 6236 25789 6239
rect 25271 6208 25789 6236
rect 25271 6205 25283 6208
rect 25225 6199 25283 6205
rect 25777 6205 25789 6208
rect 25823 6205 25835 6239
rect 25777 6199 25835 6205
rect 23474 6168 23480 6180
rect 22428 6140 22508 6168
rect 23387 6140 23480 6168
rect 22428 6128 22434 6140
rect 23474 6128 23480 6140
rect 23532 6168 23538 6180
rect 24121 6171 24179 6177
rect 24121 6168 24133 6171
rect 23532 6140 24133 6168
rect 23532 6128 23538 6140
rect 24121 6137 24133 6140
rect 24167 6168 24179 6171
rect 24762 6168 24768 6180
rect 24167 6140 24768 6168
rect 24167 6137 24179 6140
rect 24121 6131 24179 6137
rect 24762 6128 24768 6140
rect 24820 6128 24826 6180
rect 16485 6103 16543 6109
rect 16485 6100 16497 6103
rect 15988 6072 16497 6100
rect 15988 6060 15994 6072
rect 16485 6069 16497 6072
rect 16531 6069 16543 6103
rect 16485 6063 16543 6069
rect 17865 6103 17923 6109
rect 17865 6069 17877 6103
rect 17911 6100 17923 6103
rect 18417 6103 18475 6109
rect 18417 6100 18429 6103
rect 17911 6072 18429 6100
rect 17911 6069 17923 6072
rect 17865 6063 17923 6069
rect 18417 6069 18429 6072
rect 18463 6100 18475 6103
rect 18966 6100 18972 6112
rect 18463 6072 18972 6100
rect 18463 6069 18475 6072
rect 18417 6063 18475 6069
rect 18966 6060 18972 6072
rect 19024 6060 19030 6112
rect 19518 6100 19524 6112
rect 19479 6072 19524 6100
rect 19518 6060 19524 6072
rect 19576 6060 19582 6112
rect 20714 6060 20720 6112
rect 20772 6100 20778 6112
rect 20993 6103 21051 6109
rect 20993 6100 21005 6103
rect 20772 6072 21005 6100
rect 20772 6060 20778 6072
rect 20993 6069 21005 6072
rect 21039 6069 21051 6103
rect 21818 6100 21824 6112
rect 21779 6072 21824 6100
rect 20993 6063 21051 6069
rect 21818 6060 21824 6072
rect 21876 6060 21882 6112
rect 22922 6100 22928 6112
rect 22883 6072 22928 6100
rect 22922 6060 22928 6072
rect 22980 6060 22986 6112
rect 25406 6100 25412 6112
rect 25367 6072 25412 6100
rect 25406 6060 25412 6072
rect 25464 6060 25470 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1673 5899 1731 5905
rect 1673 5865 1685 5899
rect 1719 5896 1731 5899
rect 2682 5896 2688 5908
rect 1719 5868 2688 5896
rect 1719 5865 1731 5868
rect 1673 5859 1731 5865
rect 2682 5856 2688 5868
rect 2740 5856 2746 5908
rect 2774 5856 2780 5908
rect 2832 5896 2838 5908
rect 3145 5899 3203 5905
rect 3145 5896 3157 5899
rect 2832 5868 3157 5896
rect 2832 5856 2838 5868
rect 3145 5865 3157 5868
rect 3191 5865 3203 5899
rect 3145 5859 3203 5865
rect 4525 5899 4583 5905
rect 4525 5865 4537 5899
rect 4571 5896 4583 5899
rect 5166 5896 5172 5908
rect 4571 5868 5172 5896
rect 4571 5865 4583 5868
rect 4525 5859 4583 5865
rect 5166 5856 5172 5868
rect 5224 5856 5230 5908
rect 6362 5896 6368 5908
rect 6323 5868 6368 5896
rect 6362 5856 6368 5868
rect 6420 5856 6426 5908
rect 6822 5896 6828 5908
rect 6783 5868 6828 5896
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 7929 5899 7987 5905
rect 7929 5865 7941 5899
rect 7975 5896 7987 5899
rect 8570 5896 8576 5908
rect 7975 5868 8576 5896
rect 7975 5865 7987 5868
rect 7929 5859 7987 5865
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 11054 5896 11060 5908
rect 11015 5868 11060 5896
rect 11054 5856 11060 5868
rect 11112 5856 11118 5908
rect 11330 5896 11336 5908
rect 11291 5868 11336 5896
rect 11330 5856 11336 5868
rect 11388 5856 11394 5908
rect 14642 5896 14648 5908
rect 14603 5868 14648 5896
rect 14642 5856 14648 5868
rect 14700 5856 14706 5908
rect 15010 5896 15016 5908
rect 14971 5868 15016 5896
rect 15010 5856 15016 5868
rect 15068 5856 15074 5908
rect 16666 5896 16672 5908
rect 15120 5868 16672 5896
rect 5442 5828 5448 5840
rect 4632 5800 5448 5828
rect 1762 5760 1768 5772
rect 1723 5732 1768 5760
rect 1762 5720 1768 5732
rect 1820 5720 1826 5772
rect 2038 5769 2044 5772
rect 2032 5760 2044 5769
rect 1999 5732 2044 5760
rect 2032 5723 2044 5732
rect 2038 5720 2044 5723
rect 2096 5720 2102 5772
rect 3513 5763 3571 5769
rect 3513 5729 3525 5763
rect 3559 5760 3571 5763
rect 3602 5760 3608 5772
rect 3559 5732 3608 5760
rect 3559 5729 3571 5732
rect 3513 5723 3571 5729
rect 3602 5720 3608 5732
rect 3660 5760 3666 5772
rect 4632 5769 4660 5800
rect 5442 5788 5448 5800
rect 5500 5788 5506 5840
rect 7558 5828 7564 5840
rect 7519 5800 7564 5828
rect 7558 5788 7564 5800
rect 7616 5788 7622 5840
rect 8478 5788 8484 5840
rect 8536 5828 8542 5840
rect 9033 5831 9091 5837
rect 9033 5828 9045 5831
rect 8536 5800 9045 5828
rect 8536 5788 8542 5800
rect 9033 5797 9045 5800
rect 9079 5797 9091 5831
rect 9033 5791 9091 5797
rect 9766 5788 9772 5840
rect 9824 5828 9830 5840
rect 9922 5831 9980 5837
rect 9922 5828 9934 5831
rect 9824 5800 9934 5828
rect 9824 5788 9830 5800
rect 9922 5797 9934 5800
rect 9968 5797 9980 5831
rect 9922 5791 9980 5797
rect 10870 5788 10876 5840
rect 10928 5828 10934 5840
rect 11422 5828 11428 5840
rect 10928 5800 11428 5828
rect 10928 5788 10934 5800
rect 11422 5788 11428 5800
rect 11480 5828 11486 5840
rect 11701 5831 11759 5837
rect 11701 5828 11713 5831
rect 11480 5800 11713 5828
rect 11480 5788 11486 5800
rect 11701 5797 11713 5800
rect 11747 5797 11759 5831
rect 11701 5791 11759 5797
rect 12253 5831 12311 5837
rect 12253 5797 12265 5831
rect 12299 5828 12311 5831
rect 12434 5828 12440 5840
rect 12299 5800 12440 5828
rect 12299 5797 12311 5800
rect 12253 5791 12311 5797
rect 4890 5769 4896 5772
rect 3881 5763 3939 5769
rect 3881 5760 3893 5763
rect 3660 5732 3893 5760
rect 3660 5720 3666 5732
rect 3881 5729 3893 5732
rect 3927 5760 3939 5763
rect 4617 5763 4675 5769
rect 4617 5760 4629 5763
rect 3927 5732 4629 5760
rect 3927 5729 3939 5732
rect 3881 5723 3939 5729
rect 4617 5729 4629 5732
rect 4663 5729 4675 5763
rect 4884 5760 4896 5769
rect 4851 5732 4896 5760
rect 4617 5723 4675 5729
rect 4884 5723 4896 5732
rect 4890 5720 4896 5723
rect 4948 5720 4954 5772
rect 6914 5760 6920 5772
rect 6875 5732 6920 5760
rect 6914 5720 6920 5732
rect 6972 5720 6978 5772
rect 8294 5720 8300 5772
rect 8352 5760 8358 5772
rect 8389 5763 8447 5769
rect 8389 5760 8401 5763
rect 8352 5732 8401 5760
rect 8352 5720 8358 5732
rect 8389 5729 8401 5732
rect 8435 5760 8447 5763
rect 9582 5760 9588 5772
rect 8435 5732 9588 5760
rect 8435 5729 8447 5732
rect 8389 5723 8447 5729
rect 9582 5720 9588 5732
rect 9640 5720 9646 5772
rect 9674 5720 9680 5772
rect 9732 5760 9738 5772
rect 9732 5732 9777 5760
rect 9732 5720 9738 5732
rect 7742 5652 7748 5704
rect 7800 5692 7806 5704
rect 8110 5692 8116 5704
rect 7800 5664 8116 5692
rect 7800 5652 7806 5664
rect 8110 5652 8116 5664
rect 8168 5692 8174 5704
rect 8481 5695 8539 5701
rect 8481 5692 8493 5695
rect 8168 5664 8493 5692
rect 8168 5652 8174 5664
rect 8481 5661 8493 5664
rect 8527 5661 8539 5695
rect 8662 5692 8668 5704
rect 8623 5664 8668 5692
rect 8481 5655 8539 5661
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 11716 5692 11744 5791
rect 12434 5788 12440 5800
rect 12492 5788 12498 5840
rect 14093 5831 14151 5837
rect 14093 5797 14105 5831
rect 14139 5828 14151 5831
rect 14182 5828 14188 5840
rect 14139 5800 14188 5828
rect 14139 5797 14151 5800
rect 14093 5791 14151 5797
rect 14182 5788 14188 5800
rect 14240 5828 14246 5840
rect 15120 5828 15148 5868
rect 16666 5856 16672 5868
rect 16724 5856 16730 5908
rect 17126 5896 17132 5908
rect 17087 5868 17132 5896
rect 17126 5856 17132 5868
rect 17184 5856 17190 5908
rect 17497 5899 17555 5905
rect 17497 5865 17509 5899
rect 17543 5896 17555 5899
rect 17770 5896 17776 5908
rect 17543 5868 17776 5896
rect 17543 5865 17555 5868
rect 17497 5859 17555 5865
rect 17770 5856 17776 5868
rect 17828 5856 17834 5908
rect 19521 5899 19579 5905
rect 19521 5865 19533 5899
rect 19567 5896 19579 5899
rect 20070 5896 20076 5908
rect 19567 5868 20076 5896
rect 19567 5865 19579 5868
rect 19521 5859 19579 5865
rect 20070 5856 20076 5868
rect 20128 5856 20134 5908
rect 20898 5896 20904 5908
rect 20859 5868 20904 5896
rect 20898 5856 20904 5868
rect 20956 5856 20962 5908
rect 21358 5856 21364 5908
rect 21416 5896 21422 5908
rect 21729 5899 21787 5905
rect 21729 5896 21741 5899
rect 21416 5868 21741 5896
rect 21416 5856 21422 5868
rect 21729 5865 21741 5868
rect 21775 5865 21787 5899
rect 21729 5859 21787 5865
rect 22186 5856 22192 5908
rect 22244 5896 22250 5908
rect 23293 5899 23351 5905
rect 23293 5896 23305 5899
rect 22244 5868 23305 5896
rect 22244 5856 22250 5868
rect 23293 5865 23305 5868
rect 23339 5865 23351 5899
rect 23658 5896 23664 5908
rect 23619 5868 23664 5896
rect 23293 5859 23351 5865
rect 23658 5856 23664 5868
rect 23716 5856 23722 5908
rect 24118 5896 24124 5908
rect 24079 5868 24124 5896
rect 24118 5856 24124 5868
rect 24176 5856 24182 5908
rect 24397 5899 24455 5905
rect 24397 5865 24409 5899
rect 24443 5896 24455 5899
rect 24670 5896 24676 5908
rect 24443 5868 24676 5896
rect 24443 5865 24455 5868
rect 24397 5859 24455 5865
rect 24670 5856 24676 5868
rect 24728 5856 24734 5908
rect 25501 5899 25559 5905
rect 25501 5865 25513 5899
rect 25547 5896 25559 5899
rect 25590 5896 25596 5908
rect 25547 5868 25596 5896
rect 25547 5865 25559 5868
rect 25501 5859 25559 5865
rect 25590 5856 25596 5868
rect 25648 5856 25654 5908
rect 14240 5800 15148 5828
rect 15556 5831 15614 5837
rect 14240 5788 14246 5800
rect 15556 5797 15568 5831
rect 15602 5828 15614 5831
rect 15746 5828 15752 5840
rect 15602 5800 15752 5828
rect 15602 5797 15614 5800
rect 15556 5791 15614 5797
rect 15746 5788 15752 5800
rect 15804 5788 15810 5840
rect 17862 5788 17868 5840
rect 17920 5828 17926 5840
rect 18046 5837 18052 5840
rect 18040 5828 18052 5837
rect 17920 5800 18052 5828
rect 17920 5788 17926 5800
rect 18040 5791 18052 5800
rect 18046 5788 18052 5791
rect 18104 5788 18110 5840
rect 20717 5831 20775 5837
rect 20717 5797 20729 5831
rect 20763 5828 20775 5831
rect 21818 5828 21824 5840
rect 20763 5800 21824 5828
rect 20763 5797 20775 5800
rect 20717 5791 20775 5797
rect 21818 5788 21824 5800
rect 21876 5788 21882 5840
rect 25869 5831 25927 5837
rect 25869 5797 25881 5831
rect 25915 5828 25927 5831
rect 26142 5828 26148 5840
rect 25915 5800 26148 5828
rect 25915 5797 25927 5800
rect 25869 5791 25927 5797
rect 26142 5788 26148 5800
rect 26200 5828 26206 5840
rect 26326 5828 26332 5840
rect 26200 5800 26332 5828
rect 26200 5788 26206 5800
rect 26326 5788 26332 5800
rect 26384 5788 26390 5840
rect 11790 5720 11796 5772
rect 11848 5760 11854 5772
rect 12612 5763 12670 5769
rect 12612 5760 12624 5763
rect 11848 5732 12624 5760
rect 11848 5720 11854 5732
rect 12612 5729 12624 5732
rect 12658 5760 12670 5763
rect 13170 5760 13176 5772
rect 12658 5732 13176 5760
rect 12658 5729 12670 5732
rect 12612 5723 12670 5729
rect 13170 5720 13176 5732
rect 13228 5720 13234 5772
rect 14826 5720 14832 5772
rect 14884 5760 14890 5772
rect 15289 5763 15347 5769
rect 15289 5760 15301 5763
rect 14884 5732 15301 5760
rect 14884 5720 14890 5732
rect 15289 5729 15301 5732
rect 15335 5760 15347 5763
rect 17773 5763 17831 5769
rect 17773 5760 17785 5763
rect 15335 5732 17785 5760
rect 15335 5729 15347 5732
rect 15289 5723 15347 5729
rect 17773 5729 17785 5732
rect 17819 5760 17831 5763
rect 18322 5760 18328 5772
rect 17819 5732 18328 5760
rect 17819 5729 17831 5732
rect 17773 5723 17831 5729
rect 18322 5720 18328 5732
rect 18380 5760 18386 5772
rect 18598 5760 18604 5772
rect 18380 5732 18604 5760
rect 18380 5720 18386 5732
rect 18598 5720 18604 5732
rect 18656 5720 18662 5772
rect 21453 5763 21511 5769
rect 21453 5729 21465 5763
rect 21499 5760 21511 5763
rect 21542 5760 21548 5772
rect 21499 5732 21548 5760
rect 21499 5729 21511 5732
rect 21453 5723 21511 5729
rect 21542 5720 21548 5732
rect 21600 5720 21606 5772
rect 22186 5769 22192 5772
rect 22180 5760 22192 5769
rect 22147 5732 22192 5760
rect 22180 5723 22192 5732
rect 22186 5720 22192 5723
rect 22244 5720 22250 5772
rect 22922 5720 22928 5772
rect 22980 5760 22986 5772
rect 24765 5763 24823 5769
rect 24765 5760 24777 5763
rect 22980 5732 24777 5760
rect 22980 5720 22986 5732
rect 24765 5729 24777 5732
rect 24811 5760 24823 5763
rect 25038 5760 25044 5772
rect 24811 5732 25044 5760
rect 24811 5729 24823 5732
rect 24765 5723 24823 5729
rect 25038 5720 25044 5732
rect 25096 5720 25102 5772
rect 12345 5695 12403 5701
rect 12345 5692 12357 5695
rect 11716 5664 12357 5692
rect 12345 5661 12357 5664
rect 12391 5661 12403 5695
rect 12345 5655 12403 5661
rect 13814 5652 13820 5704
rect 13872 5692 13878 5704
rect 15010 5692 15016 5704
rect 13872 5664 15016 5692
rect 13872 5652 13878 5664
rect 15010 5652 15016 5664
rect 15068 5652 15074 5704
rect 20254 5652 20260 5704
rect 20312 5692 20318 5704
rect 21726 5692 21732 5704
rect 20312 5664 21732 5692
rect 20312 5652 20318 5664
rect 21726 5652 21732 5664
rect 21784 5692 21790 5704
rect 21913 5695 21971 5701
rect 21913 5692 21925 5695
rect 21784 5664 21925 5692
rect 21784 5652 21790 5664
rect 21913 5661 21925 5664
rect 21959 5661 21971 5695
rect 21913 5655 21971 5661
rect 23382 5652 23388 5704
rect 23440 5692 23446 5704
rect 24857 5695 24915 5701
rect 24857 5692 24869 5695
rect 23440 5664 24869 5692
rect 23440 5652 23446 5664
rect 24857 5661 24869 5664
rect 24903 5661 24915 5695
rect 24857 5655 24915 5661
rect 24949 5695 25007 5701
rect 24949 5661 24961 5695
rect 24995 5692 25007 5695
rect 25130 5692 25136 5704
rect 24995 5664 25136 5692
rect 24995 5661 25007 5664
rect 24949 5655 25007 5661
rect 7101 5627 7159 5633
rect 7101 5593 7113 5627
rect 7147 5624 7159 5627
rect 7558 5624 7564 5636
rect 7147 5596 7564 5624
rect 7147 5593 7159 5596
rect 7101 5587 7159 5593
rect 7558 5584 7564 5596
rect 7616 5584 7622 5636
rect 8018 5624 8024 5636
rect 7979 5596 8024 5624
rect 8018 5584 8024 5596
rect 8076 5584 8082 5636
rect 19334 5584 19340 5636
rect 19392 5624 19398 5636
rect 19889 5627 19947 5633
rect 19889 5624 19901 5627
rect 19392 5596 19901 5624
rect 19392 5584 19398 5596
rect 19889 5593 19901 5596
rect 19935 5593 19947 5627
rect 19889 5587 19947 5593
rect 5994 5556 6000 5568
rect 5955 5528 6000 5556
rect 5994 5516 6000 5528
rect 6052 5516 6058 5568
rect 8202 5516 8208 5568
rect 8260 5556 8266 5568
rect 9493 5559 9551 5565
rect 9493 5556 9505 5559
rect 8260 5528 9505 5556
rect 8260 5516 8266 5528
rect 9493 5525 9505 5528
rect 9539 5556 9551 5559
rect 10778 5556 10784 5568
rect 9539 5528 10784 5556
rect 9539 5525 9551 5528
rect 9493 5519 9551 5525
rect 10778 5516 10784 5528
rect 10836 5516 10842 5568
rect 12526 5516 12532 5568
rect 12584 5556 12590 5568
rect 13725 5559 13783 5565
rect 13725 5556 13737 5559
rect 12584 5528 13737 5556
rect 12584 5516 12590 5528
rect 13725 5525 13737 5528
rect 13771 5525 13783 5559
rect 19150 5556 19156 5568
rect 19111 5528 19156 5556
rect 13725 5519 13783 5525
rect 19150 5516 19156 5528
rect 19208 5516 19214 5568
rect 20349 5559 20407 5565
rect 20349 5525 20361 5559
rect 20395 5556 20407 5559
rect 20990 5556 20996 5568
rect 20395 5528 20996 5556
rect 20395 5525 20407 5528
rect 20349 5519 20407 5525
rect 20990 5516 20996 5528
rect 21048 5516 21054 5568
rect 21634 5516 21640 5568
rect 21692 5556 21698 5568
rect 23566 5556 23572 5568
rect 21692 5528 23572 5556
rect 21692 5516 21698 5528
rect 23566 5516 23572 5528
rect 23624 5556 23630 5568
rect 24118 5556 24124 5568
rect 23624 5528 24124 5556
rect 23624 5516 23630 5528
rect 24118 5516 24124 5528
rect 24176 5516 24182 5568
rect 24872 5556 24900 5655
rect 25130 5652 25136 5664
rect 25188 5652 25194 5704
rect 25222 5556 25228 5568
rect 24872 5528 25228 5556
rect 25222 5516 25228 5528
rect 25280 5516 25286 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 2501 5355 2559 5361
rect 2501 5321 2513 5355
rect 2547 5352 2559 5355
rect 4249 5355 4307 5361
rect 4249 5352 4261 5355
rect 2547 5324 4261 5352
rect 2547 5321 2559 5324
rect 2501 5315 2559 5321
rect 4249 5321 4261 5324
rect 4295 5321 4307 5355
rect 4249 5315 4307 5321
rect 4614 5312 4620 5364
rect 4672 5352 4678 5364
rect 4985 5355 5043 5361
rect 4985 5352 4997 5355
rect 4672 5324 4997 5352
rect 4672 5312 4678 5324
rect 4985 5321 4997 5324
rect 5031 5352 5043 5355
rect 5074 5352 5080 5364
rect 5031 5324 5080 5352
rect 5031 5321 5043 5324
rect 4985 5315 5043 5321
rect 5074 5312 5080 5324
rect 5132 5312 5138 5364
rect 7285 5355 7343 5361
rect 7285 5321 7297 5355
rect 7331 5352 7343 5355
rect 8110 5352 8116 5364
rect 7331 5324 8116 5352
rect 7331 5321 7343 5324
rect 7285 5315 7343 5321
rect 8110 5312 8116 5324
rect 8168 5312 8174 5364
rect 11422 5352 11428 5364
rect 11383 5324 11428 5352
rect 11422 5312 11428 5324
rect 11480 5312 11486 5364
rect 11790 5312 11796 5364
rect 11848 5352 11854 5364
rect 12161 5355 12219 5361
rect 12161 5352 12173 5355
rect 11848 5324 12173 5352
rect 11848 5312 11854 5324
rect 12161 5321 12173 5324
rect 12207 5321 12219 5355
rect 12161 5315 12219 5321
rect 13449 5355 13507 5361
rect 13449 5321 13461 5355
rect 13495 5352 13507 5355
rect 14090 5352 14096 5364
rect 13495 5324 14096 5352
rect 13495 5321 13507 5324
rect 13449 5315 13507 5321
rect 2866 5284 2872 5296
rect 1872 5256 2872 5284
rect 1872 5225 1900 5256
rect 2866 5244 2872 5256
rect 2924 5244 2930 5296
rect 12066 5244 12072 5296
rect 12124 5284 12130 5296
rect 12526 5284 12532 5296
rect 12124 5256 12532 5284
rect 12124 5244 12130 5256
rect 12526 5244 12532 5256
rect 12584 5244 12590 5296
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5185 1915 5219
rect 1857 5179 1915 5185
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5216 4675 5219
rect 4890 5216 4896 5228
rect 4663 5188 4896 5216
rect 4663 5185 4675 5188
rect 4617 5179 4675 5185
rect 4890 5176 4896 5188
rect 4948 5176 4954 5228
rect 5629 5219 5687 5225
rect 5629 5216 5641 5219
rect 5000 5188 5641 5216
rect 2869 5151 2927 5157
rect 2869 5117 2881 5151
rect 2915 5148 2927 5151
rect 3602 5148 3608 5160
rect 2915 5120 3608 5148
rect 2915 5117 2927 5120
rect 2869 5111 2927 5117
rect 3602 5108 3608 5120
rect 3660 5108 3666 5160
rect 4798 5108 4804 5160
rect 4856 5148 4862 5160
rect 5000 5148 5028 5188
rect 5629 5185 5641 5188
rect 5675 5216 5687 5219
rect 5994 5216 6000 5228
rect 5675 5188 6000 5216
rect 5675 5185 5687 5188
rect 5629 5179 5687 5185
rect 5994 5176 6000 5188
rect 6052 5176 6058 5228
rect 9674 5176 9680 5228
rect 9732 5176 9738 5228
rect 9766 5176 9772 5228
rect 9824 5216 9830 5228
rect 14016 5225 14044 5324
rect 14090 5312 14096 5324
rect 14148 5312 14154 5364
rect 15013 5355 15071 5361
rect 15013 5321 15025 5355
rect 15059 5352 15071 5355
rect 15746 5352 15752 5364
rect 15059 5324 15752 5352
rect 15059 5321 15071 5324
rect 15013 5315 15071 5321
rect 15746 5312 15752 5324
rect 15804 5312 15810 5364
rect 16482 5352 16488 5364
rect 16443 5324 16488 5352
rect 16482 5312 16488 5324
rect 16540 5312 16546 5364
rect 16850 5352 16856 5364
rect 16811 5324 16856 5352
rect 16850 5312 16856 5324
rect 16908 5312 16914 5364
rect 17862 5352 17868 5364
rect 17823 5324 17868 5352
rect 17862 5312 17868 5324
rect 17920 5312 17926 5364
rect 20714 5352 20720 5364
rect 20675 5324 20720 5352
rect 20714 5312 20720 5324
rect 20772 5312 20778 5364
rect 21082 5312 21088 5364
rect 21140 5352 21146 5364
rect 22186 5352 22192 5364
rect 21140 5324 22192 5352
rect 21140 5312 21146 5324
rect 22186 5312 22192 5324
rect 22244 5312 22250 5364
rect 23474 5352 23480 5364
rect 23435 5324 23480 5352
rect 23474 5312 23480 5324
rect 23532 5312 23538 5364
rect 25682 5312 25688 5364
rect 25740 5352 25746 5364
rect 26142 5352 26148 5364
rect 25740 5324 26148 5352
rect 25740 5312 25746 5324
rect 26142 5312 26148 5324
rect 26200 5312 26206 5364
rect 10505 5219 10563 5225
rect 10505 5216 10517 5219
rect 9824 5188 10517 5216
rect 9824 5176 9830 5188
rect 10505 5185 10517 5188
rect 10551 5185 10563 5219
rect 10505 5179 10563 5185
rect 14001 5219 14059 5225
rect 14001 5185 14013 5219
rect 14047 5185 14059 5219
rect 14182 5216 14188 5228
rect 14143 5188 14188 5216
rect 14001 5179 14059 5185
rect 14182 5176 14188 5188
rect 14240 5176 14246 5228
rect 14826 5176 14832 5228
rect 14884 5216 14890 5228
rect 15105 5219 15163 5225
rect 15105 5216 15117 5219
rect 14884 5188 15117 5216
rect 14884 5176 14890 5188
rect 15105 5185 15117 5188
rect 15151 5185 15163 5219
rect 15105 5179 15163 5185
rect 20530 5176 20536 5228
rect 20588 5216 20594 5228
rect 20732 5216 20760 5312
rect 22094 5244 22100 5296
rect 22152 5284 22158 5296
rect 22465 5287 22523 5293
rect 22465 5284 22477 5287
rect 22152 5256 22477 5284
rect 22152 5244 22158 5256
rect 22465 5253 22477 5256
rect 22511 5253 22523 5287
rect 22465 5247 22523 5253
rect 23492 5216 23520 5312
rect 23658 5244 23664 5296
rect 23716 5284 23722 5296
rect 24302 5284 24308 5296
rect 23716 5256 24308 5284
rect 23716 5244 23722 5256
rect 24302 5244 24308 5256
rect 24360 5244 24366 5296
rect 25222 5244 25228 5296
rect 25280 5244 25286 5296
rect 25590 5244 25596 5296
rect 25648 5284 25654 5296
rect 25866 5284 25872 5296
rect 25648 5256 25872 5284
rect 25648 5244 25654 5256
rect 25866 5244 25872 5256
rect 25924 5244 25930 5296
rect 24213 5219 24271 5225
rect 24213 5216 24225 5219
rect 20588 5188 20944 5216
rect 23492 5188 24225 5216
rect 20588 5176 20594 5188
rect 4856 5120 5028 5148
rect 4856 5108 4862 5120
rect 5442 5108 5448 5160
rect 5500 5148 5506 5160
rect 5537 5151 5595 5157
rect 5537 5148 5549 5151
rect 5500 5120 5549 5148
rect 5500 5108 5506 5120
rect 5537 5117 5549 5120
rect 5583 5117 5595 5151
rect 5537 5111 5595 5117
rect 7745 5151 7803 5157
rect 7745 5117 7757 5151
rect 7791 5148 7803 5151
rect 8386 5148 8392 5160
rect 7791 5120 8392 5148
rect 7791 5117 7803 5120
rect 7745 5111 7803 5117
rect 8386 5108 8392 5120
rect 8444 5148 8450 5160
rect 9692 5148 9720 5176
rect 8444 5120 9720 5148
rect 8444 5108 8450 5120
rect 10042 5108 10048 5160
rect 10100 5148 10106 5160
rect 10321 5151 10379 5157
rect 10321 5148 10333 5151
rect 10100 5120 10333 5148
rect 10100 5108 10106 5120
rect 10321 5117 10333 5120
rect 10367 5117 10379 5151
rect 10321 5111 10379 5117
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5117 12495 5151
rect 12437 5111 12495 5117
rect 18233 5151 18291 5157
rect 18233 5117 18245 5151
rect 18279 5148 18291 5151
rect 18322 5148 18328 5160
rect 18279 5120 18328 5148
rect 18279 5117 18291 5120
rect 18233 5111 18291 5117
rect 3114 5083 3172 5089
rect 3114 5080 3126 5083
rect 2700 5052 3126 5080
rect 2700 5024 2728 5052
rect 3114 5049 3126 5052
rect 3160 5049 3172 5083
rect 7650 5080 7656 5092
rect 7563 5052 7656 5080
rect 3114 5043 3172 5049
rect 7650 5040 7656 5052
rect 7708 5080 7714 5092
rect 8012 5083 8070 5089
rect 8012 5080 8024 5083
rect 7708 5052 8024 5080
rect 7708 5040 7714 5052
rect 8012 5049 8024 5052
rect 8058 5080 8070 5083
rect 8846 5080 8852 5092
rect 8058 5052 8852 5080
rect 8058 5049 8070 5052
rect 8012 5043 8070 5049
rect 8846 5040 8852 5052
rect 8904 5040 8910 5092
rect 9674 5040 9680 5092
rect 9732 5080 9738 5092
rect 12452 5080 12480 5111
rect 18322 5108 18328 5120
rect 18380 5108 18386 5160
rect 20254 5108 20260 5160
rect 20312 5148 20318 5160
rect 20809 5151 20867 5157
rect 20809 5148 20821 5151
rect 20312 5120 20821 5148
rect 20312 5108 20318 5120
rect 20809 5117 20821 5120
rect 20855 5117 20867 5151
rect 20916 5148 20944 5188
rect 24213 5185 24225 5188
rect 24259 5185 24271 5219
rect 24213 5179 24271 5185
rect 24765 5219 24823 5225
rect 24765 5185 24777 5219
rect 24811 5216 24823 5219
rect 25240 5216 25268 5244
rect 27154 5216 27160 5228
rect 24811 5188 27160 5216
rect 24811 5185 24823 5188
rect 24765 5179 24823 5185
rect 27154 5176 27160 5188
rect 27212 5176 27218 5228
rect 21065 5151 21123 5157
rect 21065 5148 21077 5151
rect 20916 5120 21077 5148
rect 20809 5111 20867 5117
rect 21065 5117 21077 5120
rect 21111 5117 21123 5151
rect 21065 5111 21123 5117
rect 24029 5151 24087 5157
rect 24029 5117 24041 5151
rect 24075 5148 24087 5151
rect 24486 5148 24492 5160
rect 24075 5120 24492 5148
rect 24075 5117 24087 5120
rect 24029 5111 24087 5117
rect 24486 5108 24492 5120
rect 24544 5108 24550 5160
rect 25225 5151 25283 5157
rect 25225 5117 25237 5151
rect 25271 5148 25283 5151
rect 25777 5151 25835 5157
rect 25777 5148 25789 5151
rect 25271 5120 25789 5148
rect 25271 5117 25283 5120
rect 25225 5111 25283 5117
rect 25777 5117 25789 5120
rect 25823 5148 25835 5151
rect 26050 5148 26056 5160
rect 25823 5120 26056 5148
rect 25823 5117 25835 5120
rect 25777 5111 25835 5117
rect 26050 5108 26056 5120
rect 26108 5108 26114 5160
rect 13909 5083 13967 5089
rect 13909 5080 13921 5083
rect 9732 5052 10456 5080
rect 9732 5040 9738 5052
rect 1762 5012 1768 5024
rect 1723 4984 1768 5012
rect 1762 4972 1768 4984
rect 1820 4972 1826 5024
rect 2038 4972 2044 5024
rect 2096 5012 2102 5024
rect 2317 5015 2375 5021
rect 2317 5012 2329 5015
rect 2096 4984 2329 5012
rect 2096 4972 2102 4984
rect 2317 4981 2329 4984
rect 2363 5012 2375 5015
rect 2501 5015 2559 5021
rect 2501 5012 2513 5015
rect 2363 4984 2513 5012
rect 2363 4981 2375 4984
rect 2317 4975 2375 4981
rect 2501 4981 2513 4984
rect 2547 4981 2559 5015
rect 2682 5012 2688 5024
rect 2643 4984 2688 5012
rect 2501 4975 2559 4981
rect 2682 4972 2688 4984
rect 2740 4972 2746 5024
rect 5074 5012 5080 5024
rect 5035 4984 5080 5012
rect 5074 4972 5080 4984
rect 5132 4972 5138 5024
rect 5166 4972 5172 5024
rect 5224 5012 5230 5024
rect 5445 5015 5503 5021
rect 5445 5012 5457 5015
rect 5224 4984 5457 5012
rect 5224 4972 5230 4984
rect 5445 4981 5457 4984
rect 5491 4981 5503 5015
rect 5445 4975 5503 4981
rect 6181 5015 6239 5021
rect 6181 4981 6193 5015
rect 6227 5012 6239 5015
rect 6454 5012 6460 5024
rect 6227 4984 6460 5012
rect 6227 4981 6239 4984
rect 6181 4975 6239 4981
rect 6454 4972 6460 4984
rect 6512 4972 6518 5024
rect 6641 5015 6699 5021
rect 6641 4981 6653 5015
rect 6687 5012 6699 5015
rect 6822 5012 6828 5024
rect 6687 4984 6828 5012
rect 6687 4981 6699 4984
rect 6641 4975 6699 4981
rect 6822 4972 6828 4984
rect 6880 4972 6886 5024
rect 9122 5012 9128 5024
rect 9083 4984 9128 5012
rect 9122 4972 9128 4984
rect 9180 5012 9186 5024
rect 9401 5015 9459 5021
rect 9401 5012 9413 5015
rect 9180 4984 9413 5012
rect 9180 4972 9186 4984
rect 9401 4981 9413 4984
rect 9447 5012 9459 5015
rect 9766 5012 9772 5024
rect 9447 4984 9772 5012
rect 9447 4981 9459 4984
rect 9401 4975 9459 4981
rect 9766 4972 9772 4984
rect 9824 4972 9830 5024
rect 9950 5012 9956 5024
rect 9911 4984 9956 5012
rect 9950 4972 9956 4984
rect 10008 4972 10014 5024
rect 10428 5021 10456 5052
rect 11808 5052 12480 5080
rect 13004 5052 13921 5080
rect 10413 5015 10471 5021
rect 10413 4981 10425 5015
rect 10459 5012 10471 5015
rect 10965 5015 11023 5021
rect 10965 5012 10977 5015
rect 10459 4984 10977 5012
rect 10459 4981 10471 4984
rect 10413 4975 10471 4981
rect 10965 4981 10977 4984
rect 11011 4981 11023 5015
rect 10965 4975 11023 4981
rect 11330 4972 11336 5024
rect 11388 5012 11394 5024
rect 11808 5021 11836 5052
rect 13004 5024 13032 5052
rect 13909 5049 13921 5052
rect 13955 5049 13967 5083
rect 13909 5043 13967 5049
rect 14645 5083 14703 5089
rect 14645 5049 14657 5083
rect 14691 5080 14703 5083
rect 14826 5080 14832 5092
rect 14691 5052 14832 5080
rect 14691 5049 14703 5052
rect 14645 5043 14703 5049
rect 14826 5040 14832 5052
rect 14884 5080 14890 5092
rect 15350 5083 15408 5089
rect 15350 5080 15362 5083
rect 14884 5052 15362 5080
rect 14884 5040 14890 5052
rect 15350 5049 15362 5052
rect 15396 5049 15408 5083
rect 15350 5043 15408 5049
rect 17497 5083 17555 5089
rect 17497 5049 17509 5083
rect 17543 5080 17555 5083
rect 18500 5083 18558 5089
rect 18500 5080 18512 5083
rect 17543 5052 18512 5080
rect 17543 5049 17555 5052
rect 17497 5043 17555 5049
rect 18500 5049 18512 5052
rect 18546 5080 18558 5083
rect 19150 5080 19156 5092
rect 18546 5052 19156 5080
rect 18546 5049 18558 5052
rect 18500 5043 18558 5049
rect 19150 5040 19156 5052
rect 19208 5040 19214 5092
rect 24121 5083 24179 5089
rect 24121 5080 24133 5083
rect 23032 5052 24133 5080
rect 23032 5024 23060 5052
rect 24121 5049 24133 5052
rect 24167 5049 24179 5083
rect 24121 5043 24179 5049
rect 25038 5040 25044 5092
rect 25096 5080 25102 5092
rect 25133 5083 25191 5089
rect 25133 5080 25145 5083
rect 25096 5052 25145 5080
rect 25096 5040 25102 5052
rect 25133 5049 25145 5052
rect 25179 5080 25191 5083
rect 25866 5080 25872 5092
rect 25179 5052 25872 5080
rect 25179 5049 25191 5052
rect 25133 5043 25191 5049
rect 25866 5040 25872 5052
rect 25924 5040 25930 5092
rect 11793 5015 11851 5021
rect 11793 5012 11805 5015
rect 11388 4984 11805 5012
rect 11388 4972 11394 4984
rect 11793 4981 11805 4984
rect 11839 4981 11851 5015
rect 12618 5012 12624 5024
rect 12579 4984 12624 5012
rect 11793 4975 11851 4981
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 12986 5012 12992 5024
rect 12947 4984 12992 5012
rect 12986 4972 12992 4984
rect 13044 4972 13050 5024
rect 13538 5012 13544 5024
rect 13499 4984 13544 5012
rect 13538 4972 13544 4984
rect 13596 4972 13602 5024
rect 19518 4972 19524 5024
rect 19576 5012 19582 5024
rect 19613 5015 19671 5021
rect 19613 5012 19625 5015
rect 19576 4984 19625 5012
rect 19576 4972 19582 4984
rect 19613 4981 19625 4984
rect 19659 4981 19671 5015
rect 19613 4975 19671 4981
rect 19981 5015 20039 5021
rect 19981 4981 19993 5015
rect 20027 5012 20039 5015
rect 20070 5012 20076 5024
rect 20027 4984 20076 5012
rect 20027 4981 20039 4984
rect 19981 4975 20039 4981
rect 20070 4972 20076 4984
rect 20128 4972 20134 5024
rect 20254 5012 20260 5024
rect 20215 4984 20260 5012
rect 20254 4972 20260 4984
rect 20312 4972 20318 5024
rect 23014 5012 23020 5024
rect 22975 4984 23020 5012
rect 23014 4972 23020 4984
rect 23072 4972 23078 5024
rect 23658 5012 23664 5024
rect 23619 4984 23664 5012
rect 23658 4972 23664 4984
rect 23716 4972 23722 5024
rect 25409 5015 25467 5021
rect 25409 4981 25421 5015
rect 25455 5012 25467 5015
rect 25682 5012 25688 5024
rect 25455 4984 25688 5012
rect 25455 4981 25467 4984
rect 25409 4975 25467 4981
rect 25682 4972 25688 4984
rect 25740 4972 25746 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1210 4768 1216 4820
rect 1268 4808 1274 4820
rect 1581 4811 1639 4817
rect 1581 4808 1593 4811
rect 1268 4780 1593 4808
rect 1268 4768 1274 4780
rect 1581 4777 1593 4780
rect 1627 4777 1639 4811
rect 1581 4771 1639 4777
rect 1596 4740 1624 4771
rect 1762 4768 1768 4820
rect 1820 4808 1826 4820
rect 2869 4811 2927 4817
rect 2869 4808 2881 4811
rect 1820 4780 2881 4808
rect 1820 4768 1826 4780
rect 2869 4777 2881 4780
rect 2915 4808 2927 4811
rect 5074 4808 5080 4820
rect 2915 4780 5080 4808
rect 2915 4777 2927 4780
rect 2869 4771 2927 4777
rect 5074 4768 5080 4780
rect 5132 4768 5138 4820
rect 7282 4808 7288 4820
rect 7243 4780 7288 4808
rect 7282 4768 7288 4780
rect 7340 4768 7346 4820
rect 7742 4808 7748 4820
rect 7703 4780 7748 4808
rect 7742 4768 7748 4780
rect 7800 4768 7806 4820
rect 8113 4811 8171 4817
rect 8113 4777 8125 4811
rect 8159 4808 8171 4811
rect 8662 4808 8668 4820
rect 8159 4780 8668 4808
rect 8159 4777 8171 4780
rect 8113 4771 8171 4777
rect 8662 4768 8668 4780
rect 8720 4808 8726 4820
rect 9122 4808 9128 4820
rect 8720 4780 9128 4808
rect 8720 4768 8726 4780
rect 9122 4768 9128 4780
rect 9180 4768 9186 4820
rect 9674 4808 9680 4820
rect 9635 4780 9680 4808
rect 9674 4768 9680 4780
rect 9732 4768 9738 4820
rect 10042 4768 10048 4820
rect 10100 4808 10106 4820
rect 10689 4811 10747 4817
rect 10689 4808 10701 4811
rect 10100 4780 10701 4808
rect 10100 4768 10106 4780
rect 10689 4777 10701 4780
rect 10735 4777 10747 4811
rect 13078 4808 13084 4820
rect 13039 4780 13084 4808
rect 10689 4771 10747 4777
rect 13078 4768 13084 4780
rect 13136 4808 13142 4820
rect 14001 4811 14059 4817
rect 14001 4808 14013 4811
rect 13136 4780 14013 4808
rect 13136 4768 13142 4780
rect 14001 4777 14013 4780
rect 14047 4777 14059 4811
rect 15010 4808 15016 4820
rect 14971 4780 15016 4808
rect 14001 4771 14059 4777
rect 15010 4768 15016 4780
rect 15068 4768 15074 4820
rect 15654 4808 15660 4820
rect 15615 4780 15660 4808
rect 15654 4768 15660 4780
rect 15712 4768 15718 4820
rect 17497 4811 17555 4817
rect 17497 4777 17509 4811
rect 17543 4808 17555 4811
rect 17954 4808 17960 4820
rect 17543 4780 17960 4808
rect 17543 4777 17555 4780
rect 17497 4771 17555 4777
rect 17954 4768 17960 4780
rect 18012 4768 18018 4820
rect 19061 4811 19119 4817
rect 19061 4777 19073 4811
rect 19107 4808 19119 4811
rect 19242 4808 19248 4820
rect 19107 4780 19248 4808
rect 19107 4777 19119 4780
rect 19061 4771 19119 4777
rect 19242 4768 19248 4780
rect 19300 4768 19306 4820
rect 19426 4768 19432 4820
rect 19484 4808 19490 4820
rect 19521 4811 19579 4817
rect 19521 4808 19533 4811
rect 19484 4780 19533 4808
rect 19484 4768 19490 4780
rect 19521 4777 19533 4780
rect 19567 4777 19579 4811
rect 20346 4808 20352 4820
rect 20307 4780 20352 4808
rect 19521 4771 19579 4777
rect 20346 4768 20352 4780
rect 20404 4768 20410 4820
rect 20714 4768 20720 4820
rect 20772 4808 20778 4820
rect 20901 4811 20959 4817
rect 20901 4808 20913 4811
rect 20772 4780 20913 4808
rect 20772 4768 20778 4780
rect 20901 4777 20913 4780
rect 20947 4777 20959 4811
rect 20901 4771 20959 4777
rect 20990 4768 20996 4820
rect 21048 4808 21054 4820
rect 21361 4811 21419 4817
rect 21361 4808 21373 4811
rect 21048 4780 21373 4808
rect 21048 4768 21054 4780
rect 21361 4777 21373 4780
rect 21407 4777 21419 4811
rect 21361 4771 21419 4777
rect 22005 4811 22063 4817
rect 22005 4777 22017 4811
rect 22051 4808 22063 4811
rect 22186 4808 22192 4820
rect 22051 4780 22192 4808
rect 22051 4777 22063 4780
rect 22005 4771 22063 4777
rect 22186 4768 22192 4780
rect 22244 4768 22250 4820
rect 22922 4808 22928 4820
rect 22883 4780 22928 4808
rect 22922 4768 22928 4780
rect 22980 4768 22986 4820
rect 24029 4811 24087 4817
rect 24029 4777 24041 4811
rect 24075 4777 24087 4811
rect 24029 4771 24087 4777
rect 1949 4743 2007 4749
rect 1949 4740 1961 4743
rect 1596 4712 1961 4740
rect 1949 4709 1961 4712
rect 1995 4740 2007 4743
rect 2222 4740 2228 4752
rect 1995 4712 2228 4740
rect 1995 4709 2007 4712
rect 1949 4703 2007 4709
rect 2222 4700 2228 4712
rect 2280 4700 2286 4752
rect 3881 4743 3939 4749
rect 3881 4709 3893 4743
rect 3927 4740 3939 4743
rect 4525 4743 4583 4749
rect 4525 4740 4537 4743
rect 3927 4712 4537 4740
rect 3927 4709 3939 4712
rect 3881 4703 3939 4709
rect 4525 4709 4537 4712
rect 4571 4740 4583 4743
rect 4982 4740 4988 4752
rect 4571 4712 4988 4740
rect 4571 4709 4583 4712
rect 4525 4703 4583 4709
rect 4982 4700 4988 4712
rect 5040 4700 5046 4752
rect 5534 4700 5540 4752
rect 5592 4740 5598 4752
rect 6454 4740 6460 4752
rect 5592 4712 6460 4740
rect 5592 4700 5598 4712
rect 2777 4675 2835 4681
rect 2777 4641 2789 4675
rect 2823 4672 2835 4675
rect 2866 4672 2872 4684
rect 2823 4644 2872 4672
rect 2823 4641 2835 4644
rect 2777 4635 2835 4641
rect 2866 4632 2872 4644
rect 2924 4632 2930 4684
rect 3513 4675 3571 4681
rect 3513 4641 3525 4675
rect 3559 4672 3571 4675
rect 4433 4675 4491 4681
rect 4433 4672 4445 4675
rect 3559 4644 4445 4672
rect 3559 4641 3571 4644
rect 3513 4635 3571 4641
rect 4433 4641 4445 4644
rect 4479 4672 4491 4675
rect 5258 4672 5264 4684
rect 4479 4644 5264 4672
rect 4479 4641 4491 4644
rect 4433 4635 4491 4641
rect 5258 4632 5264 4644
rect 5316 4632 5322 4684
rect 5920 4681 5948 4712
rect 6454 4700 6460 4712
rect 6512 4700 6518 4752
rect 11514 4700 11520 4752
rect 11572 4740 11578 4752
rect 11692 4743 11750 4749
rect 11692 4740 11704 4743
rect 11572 4712 11704 4740
rect 11572 4700 11578 4712
rect 11692 4709 11704 4712
rect 11738 4740 11750 4743
rect 12066 4740 12072 4752
rect 11738 4712 12072 4740
rect 11738 4709 11750 4712
rect 11692 4703 11750 4709
rect 12066 4700 12072 4712
rect 12124 4700 12130 4752
rect 15028 4740 15056 4768
rect 15749 4743 15807 4749
rect 15749 4740 15761 4743
rect 15028 4712 15761 4740
rect 15749 4709 15761 4712
rect 15795 4709 15807 4743
rect 15749 4703 15807 4709
rect 17310 4700 17316 4752
rect 17368 4740 17374 4752
rect 17865 4743 17923 4749
rect 17865 4740 17877 4743
rect 17368 4712 17877 4740
rect 17368 4700 17374 4712
rect 17865 4709 17877 4712
rect 17911 4709 17923 4743
rect 17865 4703 17923 4709
rect 22833 4743 22891 4749
rect 22833 4709 22845 4743
rect 22879 4740 22891 4743
rect 23106 4740 23112 4752
rect 22879 4712 23112 4740
rect 22879 4709 22891 4712
rect 22833 4703 22891 4709
rect 23106 4700 23112 4712
rect 23164 4700 23170 4752
rect 24044 4740 24072 4771
rect 24118 4768 24124 4820
rect 24176 4808 24182 4820
rect 24397 4811 24455 4817
rect 24397 4808 24409 4811
rect 24176 4780 24409 4808
rect 24176 4768 24182 4780
rect 24397 4777 24409 4780
rect 24443 4808 24455 4811
rect 24670 4808 24676 4820
rect 24443 4780 24676 4808
rect 24443 4777 24455 4780
rect 24397 4771 24455 4777
rect 24670 4768 24676 4780
rect 24728 4768 24734 4820
rect 25130 4808 25136 4820
rect 25091 4780 25136 4808
rect 25130 4768 25136 4780
rect 25188 4768 25194 4820
rect 26237 4811 26295 4817
rect 26237 4777 26249 4811
rect 26283 4808 26295 4811
rect 26326 4808 26332 4820
rect 26283 4780 26332 4808
rect 26283 4777 26295 4780
rect 26237 4771 26295 4777
rect 26326 4768 26332 4780
rect 26384 4768 26390 4820
rect 25498 4740 25504 4752
rect 24044 4712 25504 4740
rect 25498 4700 25504 4712
rect 25556 4700 25562 4752
rect 5905 4675 5963 4681
rect 5905 4641 5917 4675
rect 5951 4641 5963 4675
rect 5905 4635 5963 4641
rect 5994 4632 6000 4684
rect 6052 4672 6058 4684
rect 6161 4675 6219 4681
rect 6161 4672 6173 4675
rect 6052 4644 6173 4672
rect 6052 4632 6058 4644
rect 6161 4641 6173 4644
rect 6207 4641 6219 4675
rect 8478 4672 8484 4684
rect 8439 4644 8484 4672
rect 6161 4635 6219 4641
rect 8478 4632 8484 4644
rect 8536 4632 8542 4684
rect 9125 4675 9183 4681
rect 9125 4641 9137 4675
rect 9171 4672 9183 4675
rect 10045 4675 10103 4681
rect 10045 4672 10057 4675
rect 9171 4644 10057 4672
rect 9171 4641 9183 4644
rect 9125 4635 9183 4641
rect 10045 4641 10057 4644
rect 10091 4672 10103 4675
rect 10962 4672 10968 4684
rect 10091 4644 10968 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 10962 4632 10968 4644
rect 11020 4632 11026 4684
rect 11422 4672 11428 4684
rect 11383 4644 11428 4672
rect 11422 4632 11428 4644
rect 11480 4632 11486 4684
rect 12250 4672 12256 4684
rect 11532 4644 12256 4672
rect 2038 4564 2044 4616
rect 2096 4604 2102 4616
rect 3053 4607 3111 4613
rect 3053 4604 3065 4607
rect 2096 4576 3065 4604
rect 2096 4564 2102 4576
rect 3053 4573 3065 4576
rect 3099 4604 3111 4607
rect 3786 4604 3792 4616
rect 3099 4576 3792 4604
rect 3099 4573 3111 4576
rect 3053 4567 3111 4573
rect 3786 4564 3792 4576
rect 3844 4604 3850 4616
rect 4617 4607 4675 4613
rect 4617 4604 4629 4607
rect 3844 4576 4629 4604
rect 3844 4564 3850 4576
rect 4617 4573 4629 4576
rect 4663 4573 4675 4607
rect 10137 4607 10195 4613
rect 10137 4604 10149 4607
rect 4617 4567 4675 4573
rect 9416 4576 10149 4604
rect 2409 4539 2467 4545
rect 2409 4505 2421 4539
rect 2455 4536 2467 4539
rect 2590 4536 2596 4548
rect 2455 4508 2596 4536
rect 2455 4505 2467 4508
rect 2409 4499 2467 4505
rect 2590 4496 2596 4508
rect 2648 4496 2654 4548
rect 2774 4496 2780 4548
rect 2832 4536 2838 4548
rect 4065 4539 4123 4545
rect 4065 4536 4077 4539
rect 2832 4508 4077 4536
rect 2832 4496 2838 4508
rect 4065 4505 4077 4508
rect 4111 4505 4123 4539
rect 8662 4536 8668 4548
rect 8623 4508 8668 4536
rect 4065 4499 4123 4505
rect 8662 4496 8668 4508
rect 8720 4496 8726 4548
rect 4798 4428 4804 4480
rect 4856 4468 4862 4480
rect 5077 4471 5135 4477
rect 5077 4468 5089 4471
rect 4856 4440 5089 4468
rect 4856 4428 4862 4440
rect 5077 4437 5089 4440
rect 5123 4437 5135 4471
rect 5442 4468 5448 4480
rect 5403 4440 5448 4468
rect 5077 4431 5135 4437
rect 5442 4428 5448 4440
rect 5500 4428 5506 4480
rect 8294 4428 8300 4480
rect 8352 4468 8358 4480
rect 9416 4477 9444 4576
rect 10137 4573 10149 4576
rect 10183 4573 10195 4607
rect 10137 4567 10195 4573
rect 10226 4564 10232 4616
rect 10284 4604 10290 4616
rect 11532 4604 11560 4644
rect 12250 4632 12256 4644
rect 12308 4672 12314 4684
rect 16206 4672 16212 4684
rect 12308 4644 16212 4672
rect 12308 4632 12314 4644
rect 16206 4632 16212 4644
rect 16264 4632 16270 4684
rect 16482 4632 16488 4684
rect 16540 4672 16546 4684
rect 16577 4675 16635 4681
rect 16577 4672 16589 4675
rect 16540 4644 16589 4672
rect 16540 4632 16546 4644
rect 16577 4641 16589 4644
rect 16623 4672 16635 4675
rect 17770 4672 17776 4684
rect 16623 4644 17776 4672
rect 16623 4641 16635 4644
rect 16577 4635 16635 4641
rect 17770 4632 17776 4644
rect 17828 4632 17834 4684
rect 19426 4672 19432 4684
rect 19339 4644 19432 4672
rect 19426 4632 19432 4644
rect 19484 4672 19490 4684
rect 19978 4672 19984 4684
rect 19484 4644 19984 4672
rect 19484 4632 19490 4644
rect 19978 4632 19984 4644
rect 20036 4632 20042 4684
rect 20898 4632 20904 4684
rect 20956 4672 20962 4684
rect 21269 4675 21327 4681
rect 21269 4672 21281 4675
rect 20956 4644 21281 4672
rect 20956 4632 20962 4644
rect 21269 4641 21281 4644
rect 21315 4641 21327 4675
rect 21269 4635 21327 4641
rect 23290 4632 23296 4684
rect 23348 4672 23354 4684
rect 24489 4675 24547 4681
rect 24489 4672 24501 4675
rect 23348 4644 24501 4672
rect 23348 4632 23354 4644
rect 24489 4641 24501 4644
rect 24535 4672 24547 4675
rect 25777 4675 25835 4681
rect 25777 4672 25789 4675
rect 24535 4644 25789 4672
rect 24535 4641 24547 4644
rect 24489 4635 24547 4641
rect 25777 4641 25789 4644
rect 25823 4641 25835 4675
rect 25777 4635 25835 4641
rect 10284 4576 10329 4604
rect 11440 4576 11560 4604
rect 13541 4607 13599 4613
rect 10284 4564 10290 4576
rect 11440 4548 11468 4576
rect 13541 4573 13553 4607
rect 13587 4604 13599 4607
rect 14090 4604 14096 4616
rect 13587 4576 14096 4604
rect 13587 4573 13599 4576
rect 13541 4567 13599 4573
rect 14090 4564 14096 4576
rect 14148 4564 14154 4616
rect 14182 4564 14188 4616
rect 14240 4604 14246 4616
rect 15930 4604 15936 4616
rect 14240 4576 14285 4604
rect 15891 4576 15936 4604
rect 14240 4564 14246 4576
rect 15930 4564 15936 4576
rect 15988 4564 15994 4616
rect 17402 4564 17408 4616
rect 17460 4604 17466 4616
rect 17957 4607 18015 4613
rect 17957 4604 17969 4607
rect 17460 4576 17969 4604
rect 17460 4564 17466 4576
rect 17957 4573 17969 4576
rect 18003 4573 18015 4607
rect 17957 4567 18015 4573
rect 18049 4607 18107 4613
rect 18049 4573 18061 4607
rect 18095 4573 18107 4607
rect 18049 4567 18107 4573
rect 18969 4607 19027 4613
rect 18969 4573 18981 4607
rect 19015 4604 19027 4607
rect 19518 4604 19524 4616
rect 19015 4576 19524 4604
rect 19015 4573 19027 4576
rect 18969 4567 19027 4573
rect 11422 4496 11428 4548
rect 11480 4496 11486 4548
rect 13630 4536 13636 4548
rect 13591 4508 13636 4536
rect 13630 4496 13636 4508
rect 13688 4496 13694 4548
rect 14737 4539 14795 4545
rect 14737 4505 14749 4539
rect 14783 4536 14795 4539
rect 15286 4536 15292 4548
rect 14783 4508 15292 4536
rect 14783 4505 14795 4508
rect 14737 4499 14795 4505
rect 15286 4496 15292 4508
rect 15344 4496 15350 4548
rect 17313 4539 17371 4545
rect 17313 4505 17325 4539
rect 17359 4536 17371 4539
rect 17862 4536 17868 4548
rect 17359 4508 17868 4536
rect 17359 4505 17371 4508
rect 17313 4499 17371 4505
rect 17862 4496 17868 4508
rect 17920 4536 17926 4548
rect 18064 4536 18092 4567
rect 19518 4564 19524 4576
rect 19576 4604 19582 4616
rect 19705 4607 19763 4613
rect 19705 4604 19717 4607
rect 19576 4576 19717 4604
rect 19576 4564 19582 4576
rect 19705 4573 19717 4576
rect 19751 4604 19763 4607
rect 20717 4607 20775 4613
rect 20717 4604 20729 4607
rect 19751 4576 20729 4604
rect 19751 4573 19763 4576
rect 19705 4567 19763 4573
rect 20717 4573 20729 4576
rect 20763 4604 20775 4607
rect 21453 4607 21511 4613
rect 21453 4604 21465 4607
rect 20763 4576 21465 4604
rect 20763 4573 20775 4576
rect 20717 4567 20775 4573
rect 21453 4573 21465 4576
rect 21499 4573 21511 4607
rect 21453 4567 21511 4573
rect 22370 4564 22376 4616
rect 22428 4604 22434 4616
rect 23017 4607 23075 4613
rect 23017 4604 23029 4607
rect 22428 4576 23029 4604
rect 22428 4564 22434 4576
rect 23017 4573 23029 4576
rect 23063 4573 23075 4607
rect 23017 4567 23075 4573
rect 24673 4607 24731 4613
rect 24673 4573 24685 4607
rect 24719 4604 24731 4607
rect 25130 4604 25136 4616
rect 24719 4576 25136 4604
rect 24719 4573 24731 4576
rect 24673 4567 24731 4573
rect 25130 4564 25136 4576
rect 25188 4564 25194 4616
rect 17920 4508 18092 4536
rect 17920 4496 17926 4508
rect 24486 4496 24492 4548
rect 24544 4496 24550 4548
rect 9401 4471 9459 4477
rect 9401 4468 9413 4471
rect 8352 4440 9413 4468
rect 8352 4428 8358 4440
rect 9401 4437 9413 4440
rect 9447 4437 9459 4471
rect 9401 4431 9459 4437
rect 11333 4471 11391 4477
rect 11333 4437 11345 4471
rect 11379 4468 11391 4471
rect 12342 4468 12348 4480
rect 11379 4440 12348 4468
rect 11379 4437 11391 4440
rect 11333 4431 11391 4437
rect 12342 4428 12348 4440
rect 12400 4428 12406 4480
rect 12805 4471 12863 4477
rect 12805 4437 12817 4471
rect 12851 4468 12863 4471
rect 12986 4468 12992 4480
rect 12851 4440 12992 4468
rect 12851 4437 12863 4440
rect 12805 4431 12863 4437
rect 12986 4428 12992 4440
rect 13044 4428 13050 4480
rect 17034 4468 17040 4480
rect 16995 4440 17040 4468
rect 17034 4428 17040 4440
rect 17092 4428 17098 4480
rect 18506 4468 18512 4480
rect 18467 4440 18512 4468
rect 18506 4428 18512 4440
rect 18564 4428 18570 4480
rect 22094 4428 22100 4480
rect 22152 4468 22158 4480
rect 22373 4471 22431 4477
rect 22373 4468 22385 4471
rect 22152 4440 22385 4468
rect 22152 4428 22158 4440
rect 22373 4437 22385 4440
rect 22419 4468 22431 4471
rect 22465 4471 22523 4477
rect 22465 4468 22477 4471
rect 22419 4440 22477 4468
rect 22419 4437 22431 4440
rect 22373 4431 22431 4437
rect 22465 4437 22477 4440
rect 22511 4437 22523 4471
rect 23658 4468 23664 4480
rect 23619 4440 23664 4468
rect 22465 4431 22523 4437
rect 23658 4428 23664 4440
rect 23716 4468 23722 4480
rect 24504 4468 24532 4496
rect 23716 4440 24532 4468
rect 23716 4428 23722 4440
rect 24854 4428 24860 4480
rect 24912 4468 24918 4480
rect 25409 4471 25467 4477
rect 25409 4468 25421 4471
rect 24912 4440 25421 4468
rect 24912 4428 24918 4440
rect 25409 4437 25421 4440
rect 25455 4437 25467 4471
rect 25409 4431 25467 4437
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 2038 4264 2044 4276
rect 1999 4236 2044 4264
rect 2038 4224 2044 4236
rect 2096 4224 2102 4276
rect 4433 4267 4491 4273
rect 4433 4233 4445 4267
rect 4479 4264 4491 4267
rect 5442 4264 5448 4276
rect 4479 4236 5448 4264
rect 4479 4233 4491 4236
rect 4433 4227 4491 4233
rect 5442 4224 5448 4236
rect 5500 4224 5506 4276
rect 9858 4264 9864 4276
rect 9819 4236 9864 4264
rect 9858 4224 9864 4236
rect 9916 4224 9922 4276
rect 11514 4264 11520 4276
rect 11475 4236 11520 4264
rect 11514 4224 11520 4236
rect 11572 4224 11578 4276
rect 13725 4267 13783 4273
rect 13725 4233 13737 4267
rect 13771 4264 13783 4267
rect 14182 4264 14188 4276
rect 13771 4236 14188 4264
rect 13771 4233 13783 4236
rect 13725 4227 13783 4233
rect 2409 4199 2467 4205
rect 2409 4165 2421 4199
rect 2455 4196 2467 4199
rect 2682 4196 2688 4208
rect 2455 4168 2688 4196
rect 2455 4165 2467 4168
rect 2409 4159 2467 4165
rect 2682 4156 2688 4168
rect 2740 4196 2746 4208
rect 4798 4196 4804 4208
rect 2740 4168 4804 4196
rect 2740 4156 2746 4168
rect 2038 4088 2044 4140
rect 2096 4128 2102 4140
rect 2314 4128 2320 4140
rect 2096 4100 2320 4128
rect 2096 4088 2102 4100
rect 2314 4088 2320 4100
rect 2372 4088 2378 4140
rect 3326 4128 3332 4140
rect 2884 4100 3332 4128
rect 2777 4063 2835 4069
rect 2777 4029 2789 4063
rect 2823 4060 2835 4063
rect 2884 4060 2912 4100
rect 3326 4088 3332 4100
rect 3384 4088 3390 4140
rect 3436 4137 3464 4168
rect 4798 4156 4804 4168
rect 4856 4156 4862 4208
rect 4982 4156 4988 4208
rect 5040 4196 5046 4208
rect 5040 4168 5488 4196
rect 5040 4156 5046 4168
rect 5092 4137 5120 4168
rect 3421 4131 3479 4137
rect 3421 4097 3433 4131
rect 3467 4097 3479 4131
rect 3421 4091 3479 4097
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 5460 4128 5488 4168
rect 8846 4156 8852 4208
rect 8904 4196 8910 4208
rect 9217 4199 9275 4205
rect 9217 4196 9229 4199
rect 8904 4168 9229 4196
rect 8904 4156 8910 4168
rect 9217 4165 9229 4168
rect 9263 4196 9275 4199
rect 9398 4196 9404 4208
rect 9263 4168 9404 4196
rect 9263 4165 9275 4168
rect 9217 4159 9275 4165
rect 9398 4156 9404 4168
rect 9456 4156 9462 4208
rect 5537 4131 5595 4137
rect 5537 4128 5549 4131
rect 5123 4100 5157 4128
rect 5460 4100 5549 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 5537 4097 5549 4100
rect 5583 4097 5595 4131
rect 6822 4128 6828 4140
rect 6783 4100 6828 4128
rect 5537 4091 5595 4097
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 9876 4128 9904 4224
rect 10045 4199 10103 4205
rect 10045 4165 10057 4199
rect 10091 4196 10103 4199
rect 12710 4196 12716 4208
rect 10091 4168 12716 4196
rect 10091 4165 10103 4168
rect 10045 4159 10103 4165
rect 12710 4156 12716 4168
rect 12768 4156 12774 4208
rect 10597 4131 10655 4137
rect 10597 4128 10609 4131
rect 9876 4100 10609 4128
rect 10597 4097 10609 4100
rect 10643 4097 10655 4131
rect 10597 4091 10655 4097
rect 11146 4088 11152 4140
rect 11204 4128 11210 4140
rect 11606 4128 11612 4140
rect 11204 4100 11612 4128
rect 11204 4088 11210 4100
rect 11606 4088 11612 4100
rect 11664 4088 11670 4140
rect 13081 4131 13139 4137
rect 13081 4128 13093 4131
rect 12176 4100 13093 4128
rect 2823 4032 2912 4060
rect 2823 4029 2835 4032
rect 2777 4023 2835 4029
rect 2958 4020 2964 4072
rect 3016 4060 3022 4072
rect 3237 4063 3295 4069
rect 3237 4060 3249 4063
rect 3016 4032 3249 4060
rect 3016 4020 3022 4032
rect 3237 4029 3249 4032
rect 3283 4029 3295 4063
rect 7742 4060 7748 4072
rect 3237 4023 3295 4029
rect 3344 4032 7748 4060
rect 1854 3952 1860 4004
rect 1912 3992 1918 4004
rect 3344 3992 3372 4032
rect 7742 4020 7748 4032
rect 7800 4020 7806 4072
rect 7837 4063 7895 4069
rect 7837 4029 7849 4063
rect 7883 4060 7895 4063
rect 8386 4060 8392 4072
rect 7883 4032 8392 4060
rect 7883 4029 7895 4032
rect 7837 4023 7895 4029
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 9950 4020 9956 4072
rect 10008 4060 10014 4072
rect 10413 4063 10471 4069
rect 10413 4060 10425 4063
rect 10008 4032 10425 4060
rect 10008 4020 10014 4032
rect 10413 4029 10425 4032
rect 10459 4060 10471 4063
rect 11793 4063 11851 4069
rect 11793 4060 11805 4063
rect 10459 4032 11805 4060
rect 10459 4029 10471 4032
rect 10413 4023 10471 4029
rect 11793 4029 11805 4032
rect 11839 4029 11851 4063
rect 11793 4023 11851 4029
rect 11974 4020 11980 4072
rect 12032 4020 12038 4072
rect 1912 3964 3372 3992
rect 1912 3952 1918 3964
rect 3418 3952 3424 4004
rect 3476 3992 3482 4004
rect 3878 3992 3884 4004
rect 3476 3964 3884 3992
rect 3476 3952 3482 3964
rect 3878 3952 3884 3964
rect 3936 3992 3942 4004
rect 4801 3995 4859 4001
rect 4801 3992 4813 3995
rect 3936 3964 4813 3992
rect 3936 3952 3942 3964
rect 4801 3961 4813 3964
rect 4847 3961 4859 3995
rect 4801 3955 4859 3961
rect 5166 3952 5172 4004
rect 5224 3992 5230 4004
rect 5905 3995 5963 4001
rect 5905 3992 5917 3995
rect 5224 3964 5917 3992
rect 5224 3952 5230 3964
rect 5905 3961 5917 3964
rect 5951 3992 5963 3995
rect 5994 3992 6000 4004
rect 5951 3964 6000 3992
rect 5951 3961 5963 3964
rect 5905 3955 5963 3961
rect 5994 3952 6000 3964
rect 6052 3952 6058 4004
rect 8082 3995 8140 4001
rect 8082 3992 8094 3995
rect 7668 3964 8094 3992
rect 7668 3936 7696 3964
rect 8082 3961 8094 3964
rect 8128 3961 8140 3995
rect 8082 3955 8140 3961
rect 9398 3952 9404 4004
rect 9456 3992 9462 4004
rect 9493 3995 9551 4001
rect 9493 3992 9505 3995
rect 9456 3964 9505 3992
rect 9456 3952 9462 3964
rect 9493 3961 9505 3964
rect 9539 3992 9551 3995
rect 10226 3992 10232 4004
rect 9539 3964 10232 3992
rect 9539 3961 9551 3964
rect 9493 3955 9551 3961
rect 10226 3952 10232 3964
rect 10284 3952 10290 4004
rect 10505 3995 10563 4001
rect 10505 3961 10517 3995
rect 10551 3992 10563 3995
rect 10686 3992 10692 4004
rect 10551 3964 10692 3992
rect 10551 3961 10563 3964
rect 10505 3955 10563 3961
rect 10686 3952 10692 3964
rect 10744 3992 10750 4004
rect 11057 3995 11115 4001
rect 11057 3992 11069 3995
rect 10744 3964 11069 3992
rect 10744 3952 10750 3964
rect 11057 3961 11069 3964
rect 11103 3961 11115 3995
rect 11057 3955 11115 3961
rect 11330 3952 11336 4004
rect 11388 3992 11394 4004
rect 11992 3992 12020 4020
rect 11388 3964 12020 3992
rect 11388 3952 11394 3964
rect 1670 3924 1676 3936
rect 1631 3896 1676 3924
rect 1670 3884 1676 3896
rect 1728 3884 1734 3936
rect 2866 3924 2872 3936
rect 2827 3896 2872 3924
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 4246 3924 4252 3936
rect 4207 3896 4252 3924
rect 4246 3884 4252 3896
rect 4304 3924 4310 3936
rect 4706 3924 4712 3936
rect 4304 3896 4712 3924
rect 4304 3884 4310 3896
rect 4706 3884 4712 3896
rect 4764 3924 4770 3936
rect 4893 3927 4951 3933
rect 4893 3924 4905 3927
rect 4764 3896 4905 3924
rect 4764 3884 4770 3896
rect 4893 3893 4905 3896
rect 4939 3893 4951 3927
rect 4893 3887 4951 3893
rect 6365 3927 6423 3933
rect 6365 3893 6377 3927
rect 6411 3924 6423 3927
rect 6454 3924 6460 3936
rect 6411 3896 6460 3924
rect 6411 3893 6423 3896
rect 6365 3887 6423 3893
rect 6454 3884 6460 3896
rect 6512 3924 6518 3936
rect 7374 3924 7380 3936
rect 6512 3896 7380 3924
rect 6512 3884 6518 3896
rect 7374 3884 7380 3896
rect 7432 3884 7438 3936
rect 7650 3924 7656 3936
rect 7611 3896 7656 3924
rect 7650 3884 7656 3896
rect 7708 3884 7714 3936
rect 10042 3884 10048 3936
rect 10100 3924 10106 3936
rect 10962 3924 10968 3936
rect 10100 3896 10968 3924
rect 10100 3884 10106 3896
rect 10962 3884 10968 3896
rect 11020 3884 11026 3936
rect 12066 3884 12072 3936
rect 12124 3924 12130 3936
rect 12176 3933 12204 4100
rect 13081 4097 13093 4100
rect 13127 4128 13139 4131
rect 13740 4128 13768 4227
rect 14182 4224 14188 4236
rect 14240 4224 14246 4276
rect 17402 4264 17408 4276
rect 17363 4236 17408 4264
rect 17402 4224 17408 4236
rect 17460 4224 17466 4276
rect 19242 4264 19248 4276
rect 19076 4236 19248 4264
rect 15565 4199 15623 4205
rect 15565 4165 15577 4199
rect 15611 4196 15623 4199
rect 15930 4196 15936 4208
rect 15611 4168 15936 4196
rect 15611 4165 15623 4168
rect 15565 4159 15623 4165
rect 15930 4156 15936 4168
rect 15988 4196 15994 4208
rect 16301 4199 16359 4205
rect 16301 4196 16313 4199
rect 15988 4168 16313 4196
rect 15988 4156 15994 4168
rect 16301 4165 16313 4168
rect 16347 4196 16359 4199
rect 19076 4196 19104 4236
rect 19242 4224 19248 4236
rect 19300 4224 19306 4276
rect 22557 4267 22615 4273
rect 22557 4233 22569 4267
rect 22603 4264 22615 4267
rect 22922 4264 22928 4276
rect 22603 4236 22928 4264
rect 22603 4233 22615 4236
rect 22557 4227 22615 4233
rect 22922 4224 22928 4236
rect 22980 4224 22986 4276
rect 24670 4264 24676 4276
rect 24631 4236 24676 4264
rect 24670 4224 24676 4236
rect 24728 4224 24734 4276
rect 25130 4264 25136 4276
rect 25091 4236 25136 4264
rect 25130 4224 25136 4236
rect 25188 4224 25194 4276
rect 19426 4196 19432 4208
rect 16347 4168 16988 4196
rect 16347 4165 16359 4168
rect 16301 4159 16359 4165
rect 16850 4128 16856 4140
rect 13127 4100 13768 4128
rect 16811 4100 16856 4128
rect 13127 4097 13139 4100
rect 13081 4091 13139 4097
rect 16850 4088 16856 4100
rect 16908 4088 16914 4140
rect 16960 4137 16988 4168
rect 18984 4168 19104 4196
rect 19260 4168 19432 4196
rect 18984 4137 19012 4168
rect 16945 4131 17003 4137
rect 16945 4097 16957 4131
rect 16991 4097 17003 4131
rect 16945 4091 17003 4097
rect 18969 4131 19027 4137
rect 18969 4097 18981 4131
rect 19015 4097 19027 4131
rect 18969 4091 19027 4097
rect 12618 4020 12624 4072
rect 12676 4060 12682 4072
rect 12805 4063 12863 4069
rect 12805 4060 12817 4063
rect 12676 4032 12817 4060
rect 12676 4020 12682 4032
rect 12805 4029 12817 4032
rect 12851 4060 12863 4063
rect 13722 4060 13728 4072
rect 12851 4032 13728 4060
rect 12851 4029 12863 4032
rect 12805 4023 12863 4029
rect 13722 4020 13728 4032
rect 13780 4020 13786 4072
rect 14185 4063 14243 4069
rect 14185 4029 14197 4063
rect 14231 4060 14243 4063
rect 14734 4060 14740 4072
rect 14231 4032 14740 4060
rect 14231 4029 14243 4032
rect 14185 4023 14243 4029
rect 14734 4020 14740 4032
rect 14792 4020 14798 4072
rect 18782 4060 18788 4072
rect 17788 4032 18788 4060
rect 12342 3952 12348 4004
rect 12400 3992 12406 4004
rect 14093 3995 14151 4001
rect 12400 3964 12940 3992
rect 12400 3952 12406 3964
rect 12161 3927 12219 3933
rect 12161 3924 12173 3927
rect 12124 3896 12173 3924
rect 12124 3884 12130 3896
rect 12161 3893 12173 3896
rect 12207 3893 12219 3927
rect 12161 3887 12219 3893
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 12912 3933 12940 3964
rect 14093 3961 14105 3995
rect 14139 3992 14151 3995
rect 14274 3992 14280 4004
rect 14139 3964 14280 3992
rect 14139 3961 14151 3964
rect 14093 3955 14151 3961
rect 14274 3952 14280 3964
rect 14332 3992 14338 4004
rect 14430 3995 14488 4001
rect 14430 3992 14442 3995
rect 14332 3964 14442 3992
rect 14332 3952 14338 3964
rect 14430 3961 14442 3964
rect 14476 3961 14488 3995
rect 17494 3992 17500 4004
rect 14430 3955 14488 3961
rect 14559 3964 17500 3992
rect 12897 3927 12955 3933
rect 12492 3896 12537 3924
rect 12492 3884 12498 3896
rect 12897 3893 12909 3927
rect 12943 3924 12955 3927
rect 14559 3924 14587 3964
rect 17494 3952 17500 3964
rect 17552 3952 17558 4004
rect 17788 3936 17816 4032
rect 18782 4020 18788 4032
rect 18840 4020 18846 4072
rect 19260 3992 19288 4168
rect 19426 4156 19432 4168
rect 19484 4156 19490 4208
rect 20993 4199 21051 4205
rect 20993 4165 21005 4199
rect 21039 4196 21051 4199
rect 22278 4196 22284 4208
rect 21039 4168 22284 4196
rect 21039 4165 21051 4168
rect 20993 4159 21051 4165
rect 19797 4131 19855 4137
rect 19797 4097 19809 4131
rect 19843 4128 19855 4131
rect 20530 4128 20536 4140
rect 19843 4100 20536 4128
rect 19843 4097 19855 4100
rect 19797 4091 19855 4097
rect 20530 4088 20536 4100
rect 20588 4088 20594 4140
rect 21928 4137 21956 4168
rect 22278 4156 22284 4168
rect 22336 4196 22342 4208
rect 25038 4196 25044 4208
rect 22336 4168 25044 4196
rect 22336 4156 22342 4168
rect 25038 4156 25044 4168
rect 25096 4156 25102 4208
rect 21913 4131 21971 4137
rect 21913 4097 21925 4131
rect 21959 4097 21971 4131
rect 21913 4091 21971 4097
rect 22097 4131 22155 4137
rect 22097 4097 22109 4131
rect 22143 4128 22155 4131
rect 22370 4128 22376 4140
rect 22143 4100 22376 4128
rect 22143 4097 22155 4100
rect 22097 4091 22155 4097
rect 22370 4088 22376 4100
rect 22428 4088 22434 4140
rect 22925 4131 22983 4137
rect 22925 4097 22937 4131
rect 22971 4128 22983 4131
rect 23106 4128 23112 4140
rect 22971 4100 23112 4128
rect 22971 4097 22983 4100
rect 22925 4091 22983 4097
rect 23106 4088 23112 4100
rect 23164 4088 23170 4140
rect 23474 4088 23480 4140
rect 23532 4128 23538 4140
rect 24213 4131 24271 4137
rect 24213 4128 24225 4131
rect 23532 4100 24225 4128
rect 23532 4088 23538 4100
rect 24213 4097 24225 4100
rect 24259 4097 24271 4131
rect 24213 4091 24271 4097
rect 19334 4020 19340 4072
rect 19392 4060 19398 4072
rect 20257 4063 20315 4069
rect 20257 4060 20269 4063
rect 19392 4032 20269 4060
rect 19392 4020 19398 4032
rect 20257 4029 20269 4032
rect 20303 4029 20315 4063
rect 20257 4023 20315 4029
rect 20349 4063 20407 4069
rect 20349 4029 20361 4063
rect 20395 4060 20407 4063
rect 20622 4060 20628 4072
rect 20395 4032 20628 4060
rect 20395 4029 20407 4032
rect 20349 4023 20407 4029
rect 20622 4020 20628 4032
rect 20680 4020 20686 4072
rect 24118 4060 24124 4072
rect 24079 4032 24124 4060
rect 24118 4020 24124 4032
rect 24176 4020 24182 4072
rect 25222 4060 25228 4072
rect 25183 4032 25228 4060
rect 25222 4020 25228 4032
rect 25280 4060 25286 4072
rect 25961 4063 26019 4069
rect 25961 4060 25973 4063
rect 25280 4032 25973 4060
rect 25280 4020 25286 4032
rect 25961 4029 25973 4032
rect 26007 4029 26019 4063
rect 26326 4060 26332 4072
rect 26287 4032 26332 4060
rect 25961 4023 26019 4029
rect 26326 4020 26332 4032
rect 26384 4020 26390 4072
rect 18340 3964 19288 3992
rect 19429 3995 19487 4001
rect 12943 3896 14587 3924
rect 12943 3893 12955 3896
rect 12897 3887 12955 3893
rect 16298 3884 16304 3936
rect 16356 3924 16362 3936
rect 16393 3927 16451 3933
rect 16393 3924 16405 3927
rect 16356 3896 16405 3924
rect 16356 3884 16362 3896
rect 16393 3893 16405 3896
rect 16439 3893 16451 3927
rect 16758 3924 16764 3936
rect 16719 3896 16764 3924
rect 16393 3887 16451 3893
rect 16758 3884 16764 3896
rect 16816 3884 16822 3936
rect 17770 3924 17776 3936
rect 17731 3896 17776 3924
rect 17770 3884 17776 3896
rect 17828 3884 17834 3936
rect 18340 3933 18368 3964
rect 19429 3961 19441 3995
rect 19475 3992 19487 3995
rect 20714 3992 20720 4004
rect 19475 3964 20720 3992
rect 19475 3961 19487 3964
rect 19429 3955 19487 3961
rect 18325 3927 18383 3933
rect 18325 3893 18337 3927
rect 18371 3893 18383 3927
rect 18325 3887 18383 3893
rect 18506 3884 18512 3936
rect 18564 3924 18570 3936
rect 18693 3927 18751 3933
rect 18693 3924 18705 3927
rect 18564 3896 18705 3924
rect 18564 3884 18570 3896
rect 18693 3893 18705 3896
rect 18739 3893 18751 3927
rect 18693 3887 18751 3893
rect 19334 3884 19340 3936
rect 19392 3924 19398 3936
rect 19444 3924 19472 3955
rect 20714 3952 20720 3964
rect 20772 3952 20778 4004
rect 21821 3995 21879 4001
rect 21821 3992 21833 3995
rect 21284 3964 21833 3992
rect 19392 3896 19472 3924
rect 19889 3927 19947 3933
rect 19392 3884 19398 3896
rect 19889 3893 19901 3927
rect 19935 3924 19947 3927
rect 19978 3924 19984 3936
rect 19935 3896 19984 3924
rect 19935 3893 19947 3896
rect 19889 3887 19947 3893
rect 19978 3884 19984 3896
rect 20036 3884 20042 3936
rect 21082 3884 21088 3936
rect 21140 3924 21146 3936
rect 21284 3933 21312 3964
rect 21821 3961 21833 3964
rect 21867 3961 21879 3995
rect 24026 3992 24032 4004
rect 23987 3964 24032 3992
rect 21821 3955 21879 3961
rect 24026 3952 24032 3964
rect 24084 3992 24090 4004
rect 24762 3992 24768 4004
rect 24084 3964 24768 3992
rect 24084 3952 24090 3964
rect 24762 3952 24768 3964
rect 24820 3952 24826 4004
rect 24946 3952 24952 4004
rect 25004 3992 25010 4004
rect 25501 3995 25559 4001
rect 25501 3992 25513 3995
rect 25004 3964 25513 3992
rect 25004 3952 25010 3964
rect 25501 3961 25513 3964
rect 25547 3961 25559 3995
rect 25501 3955 25559 3961
rect 21269 3927 21327 3933
rect 21269 3924 21281 3927
rect 21140 3896 21281 3924
rect 21140 3884 21146 3896
rect 21269 3893 21281 3896
rect 21315 3893 21327 3927
rect 21269 3887 21327 3893
rect 21358 3884 21364 3936
rect 21416 3924 21422 3936
rect 21453 3927 21511 3933
rect 21453 3924 21465 3927
rect 21416 3896 21465 3924
rect 21416 3884 21422 3896
rect 21453 3893 21465 3896
rect 21499 3893 21511 3927
rect 23474 3924 23480 3936
rect 23435 3896 23480 3924
rect 21453 3887 21511 3893
rect 23474 3884 23480 3896
rect 23532 3884 23538 3936
rect 23566 3884 23572 3936
rect 23624 3924 23630 3936
rect 23661 3927 23719 3933
rect 23661 3924 23673 3927
rect 23624 3896 23673 3924
rect 23624 3884 23630 3896
rect 23661 3893 23673 3896
rect 23707 3893 23719 3927
rect 23661 3887 23719 3893
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1394 3720 1400 3732
rect 1355 3692 1400 3720
rect 1394 3680 1400 3692
rect 1452 3680 1458 3732
rect 1670 3680 1676 3732
rect 1728 3720 1734 3732
rect 2958 3720 2964 3732
rect 1728 3692 1900 3720
rect 2919 3692 2964 3720
rect 1728 3680 1734 3692
rect 1578 3612 1584 3664
rect 1636 3652 1642 3664
rect 1765 3655 1823 3661
rect 1765 3652 1777 3655
rect 1636 3624 1777 3652
rect 1636 3612 1642 3624
rect 1765 3621 1777 3624
rect 1811 3621 1823 3655
rect 1765 3615 1823 3621
rect 1780 3448 1808 3615
rect 1872 3593 1900 3692
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 3786 3720 3792 3732
rect 3747 3692 3792 3720
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 4062 3720 4068 3732
rect 4023 3692 4068 3720
rect 4062 3680 4068 3692
rect 4120 3680 4126 3732
rect 4433 3723 4491 3729
rect 4433 3689 4445 3723
rect 4479 3720 4491 3723
rect 5534 3720 5540 3732
rect 4479 3692 5540 3720
rect 4479 3689 4491 3692
rect 4433 3683 4491 3689
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 7374 3680 7380 3732
rect 7432 3720 7438 3732
rect 7561 3723 7619 3729
rect 7561 3720 7573 3723
rect 7432 3692 7573 3720
rect 7432 3680 7438 3692
rect 7561 3689 7573 3692
rect 7607 3689 7619 3723
rect 7561 3683 7619 3689
rect 8205 3723 8263 3729
rect 8205 3689 8217 3723
rect 8251 3720 8263 3723
rect 8386 3720 8392 3732
rect 8251 3692 8392 3720
rect 8251 3689 8263 3692
rect 8205 3683 8263 3689
rect 8386 3680 8392 3692
rect 8444 3680 8450 3732
rect 8478 3680 8484 3732
rect 8536 3720 8542 3732
rect 9033 3723 9091 3729
rect 9033 3720 9045 3723
rect 8536 3692 9045 3720
rect 8536 3680 8542 3692
rect 9033 3689 9045 3692
rect 9079 3720 9091 3723
rect 9122 3720 9128 3732
rect 9079 3692 9128 3720
rect 9079 3689 9091 3692
rect 9033 3683 9091 3689
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 9493 3723 9551 3729
rect 9493 3689 9505 3723
rect 9539 3720 9551 3723
rect 10137 3723 10195 3729
rect 10137 3720 10149 3723
rect 9539 3692 10149 3720
rect 9539 3689 9551 3692
rect 9493 3683 9551 3689
rect 10137 3689 10149 3692
rect 10183 3720 10195 3723
rect 12805 3723 12863 3729
rect 12805 3720 12817 3723
rect 10183 3692 12817 3720
rect 10183 3689 10195 3692
rect 10137 3683 10195 3689
rect 12805 3689 12817 3692
rect 12851 3689 12863 3723
rect 12805 3683 12863 3689
rect 13173 3723 13231 3729
rect 13173 3689 13185 3723
rect 13219 3720 13231 3723
rect 14366 3720 14372 3732
rect 13219 3692 14372 3720
rect 13219 3689 13231 3692
rect 13173 3683 13231 3689
rect 2866 3612 2872 3664
rect 2924 3652 2930 3664
rect 5077 3655 5135 3661
rect 5077 3652 5089 3655
rect 2924 3624 5089 3652
rect 2924 3612 2930 3624
rect 5077 3621 5089 3624
rect 5123 3621 5135 3655
rect 5077 3615 5135 3621
rect 6086 3612 6092 3664
rect 6144 3661 6150 3664
rect 6144 3655 6208 3661
rect 6144 3621 6162 3655
rect 6196 3621 6208 3655
rect 6144 3615 6208 3621
rect 8573 3655 8631 3661
rect 8573 3621 8585 3655
rect 8619 3652 8631 3655
rect 9582 3652 9588 3664
rect 8619 3624 9588 3652
rect 8619 3621 8631 3624
rect 8573 3615 8631 3621
rect 6144 3612 6150 3615
rect 9582 3612 9588 3624
rect 9640 3612 9646 3664
rect 9858 3612 9864 3664
rect 9916 3652 9922 3664
rect 11330 3652 11336 3664
rect 9916 3624 11336 3652
rect 9916 3612 9922 3624
rect 11330 3612 11336 3624
rect 11388 3612 11394 3664
rect 11514 3612 11520 3664
rect 11572 3652 11578 3664
rect 11701 3655 11759 3661
rect 11701 3652 11713 3655
rect 11572 3624 11713 3652
rect 11572 3612 11578 3624
rect 11701 3621 11713 3624
rect 11747 3621 11759 3655
rect 11701 3615 11759 3621
rect 11790 3612 11796 3664
rect 11848 3612 11854 3664
rect 12710 3612 12716 3664
rect 12768 3652 12774 3664
rect 13188 3652 13216 3683
rect 14366 3680 14372 3692
rect 14424 3680 14430 3732
rect 14642 3720 14648 3732
rect 14603 3692 14648 3720
rect 14642 3680 14648 3692
rect 14700 3680 14706 3732
rect 15105 3723 15163 3729
rect 15105 3689 15117 3723
rect 15151 3720 15163 3723
rect 16758 3720 16764 3732
rect 15151 3692 16764 3720
rect 15151 3689 15163 3692
rect 15105 3683 15163 3689
rect 16758 3680 16764 3692
rect 16816 3720 16822 3732
rect 19061 3723 19119 3729
rect 19061 3720 19073 3723
rect 16816 3692 19073 3720
rect 16816 3680 16822 3692
rect 19061 3689 19073 3692
rect 19107 3689 19119 3723
rect 19518 3720 19524 3732
rect 19431 3692 19524 3720
rect 19061 3683 19119 3689
rect 19518 3680 19524 3692
rect 19576 3720 19582 3732
rect 20162 3720 20168 3732
rect 19576 3692 20168 3720
rect 19576 3680 19582 3692
rect 20162 3680 20168 3692
rect 20220 3680 20226 3732
rect 20898 3720 20904 3732
rect 20859 3692 20904 3720
rect 20898 3680 20904 3692
rect 20956 3680 20962 3732
rect 21361 3723 21419 3729
rect 21361 3689 21373 3723
rect 21407 3720 21419 3723
rect 21910 3720 21916 3732
rect 21407 3692 21916 3720
rect 21407 3689 21419 3692
rect 21361 3683 21419 3689
rect 21910 3680 21916 3692
rect 21968 3680 21974 3732
rect 22005 3723 22063 3729
rect 22005 3689 22017 3723
rect 22051 3720 22063 3723
rect 22370 3720 22376 3732
rect 22051 3692 22376 3720
rect 22051 3689 22063 3692
rect 22005 3683 22063 3689
rect 22370 3680 22376 3692
rect 22428 3680 22434 3732
rect 22465 3723 22523 3729
rect 22465 3689 22477 3723
rect 22511 3720 22523 3723
rect 23014 3720 23020 3732
rect 22511 3692 23020 3720
rect 22511 3689 22523 3692
rect 22465 3683 22523 3689
rect 23014 3680 23020 3692
rect 23072 3680 23078 3732
rect 24118 3680 24124 3732
rect 24176 3720 24182 3732
rect 25409 3723 25467 3729
rect 25409 3720 25421 3723
rect 24176 3692 25421 3720
rect 24176 3680 24182 3692
rect 25409 3689 25421 3692
rect 25455 3689 25467 3723
rect 25774 3720 25780 3732
rect 25735 3692 25780 3720
rect 25409 3683 25467 3689
rect 25774 3680 25780 3692
rect 25832 3680 25838 3732
rect 26142 3720 26148 3732
rect 26103 3692 26148 3720
rect 26142 3680 26148 3692
rect 26200 3680 26206 3732
rect 12768 3624 13216 3652
rect 13265 3655 13323 3661
rect 12768 3612 12774 3624
rect 13265 3621 13277 3655
rect 13311 3652 13323 3655
rect 13446 3652 13452 3664
rect 13311 3624 13452 3652
rect 13311 3621 13323 3624
rect 13265 3615 13323 3621
rect 13446 3612 13452 3624
rect 13504 3612 13510 3664
rect 15556 3655 15614 3661
rect 15556 3621 15568 3655
rect 15602 3652 15614 3655
rect 15930 3652 15936 3664
rect 15602 3624 15936 3652
rect 15602 3621 15614 3624
rect 15556 3615 15614 3621
rect 15930 3612 15936 3624
rect 15988 3612 15994 3664
rect 17310 3652 17316 3664
rect 17271 3624 17316 3652
rect 17310 3612 17316 3624
rect 17368 3612 17374 3664
rect 18601 3655 18659 3661
rect 18601 3621 18613 3655
rect 18647 3652 18659 3655
rect 18874 3652 18880 3664
rect 18647 3624 18880 3652
rect 18647 3621 18659 3624
rect 18601 3615 18659 3621
rect 18874 3612 18880 3624
rect 18932 3612 18938 3664
rect 19334 3612 19340 3664
rect 19392 3652 19398 3664
rect 20257 3655 20315 3661
rect 20257 3652 20269 3655
rect 19392 3624 20269 3652
rect 19392 3612 19398 3624
rect 20257 3621 20269 3624
rect 20303 3652 20315 3655
rect 21634 3652 21640 3664
rect 20303 3624 21640 3652
rect 20303 3621 20315 3624
rect 20257 3615 20315 3621
rect 21634 3612 21640 3624
rect 21692 3612 21698 3664
rect 22922 3652 22928 3664
rect 22883 3624 22928 3652
rect 22922 3612 22928 3624
rect 22980 3612 22986 3664
rect 24486 3652 24492 3664
rect 24447 3624 24492 3652
rect 24486 3612 24492 3624
rect 24544 3652 24550 3664
rect 24762 3652 24768 3664
rect 24544 3624 24768 3652
rect 24544 3612 24550 3624
rect 24762 3612 24768 3624
rect 24820 3612 24826 3664
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3584 1915 3587
rect 3142 3584 3148 3596
rect 1903 3556 3148 3584
rect 1903 3553 1915 3556
rect 1857 3547 1915 3553
rect 3142 3544 3148 3556
rect 3200 3584 3206 3596
rect 4525 3587 4583 3593
rect 3200 3556 3372 3584
rect 3200 3544 3206 3556
rect 2041 3519 2099 3525
rect 2041 3485 2053 3519
rect 2087 3516 2099 3519
rect 2222 3516 2228 3528
rect 2087 3488 2228 3516
rect 2087 3485 2099 3488
rect 2041 3479 2099 3485
rect 2222 3476 2228 3488
rect 2280 3516 2286 3528
rect 3237 3519 3295 3525
rect 3237 3516 3249 3519
rect 2280 3488 3249 3516
rect 2280 3476 2286 3488
rect 3237 3485 3249 3488
rect 3283 3485 3295 3519
rect 3237 3479 3295 3485
rect 2409 3451 2467 3457
rect 2409 3448 2421 3451
rect 1780 3420 2421 3448
rect 2409 3417 2421 3420
rect 2455 3417 2467 3451
rect 2409 3411 2467 3417
rect 1394 3340 1400 3392
rect 1452 3380 1458 3392
rect 1946 3380 1952 3392
rect 1452 3352 1952 3380
rect 1452 3340 1458 3352
rect 1946 3340 1952 3352
rect 2004 3340 2010 3392
rect 3344 3380 3372 3556
rect 4525 3553 4537 3587
rect 4571 3584 4583 3587
rect 5258 3584 5264 3596
rect 4571 3556 5264 3584
rect 4571 3553 4583 3556
rect 4525 3547 4583 3553
rect 5258 3544 5264 3556
rect 5316 3544 5322 3596
rect 5905 3587 5963 3593
rect 5905 3553 5917 3587
rect 5951 3584 5963 3587
rect 5994 3584 6000 3596
rect 5951 3556 6000 3584
rect 5951 3553 5963 3556
rect 5905 3547 5963 3553
rect 5994 3544 6000 3556
rect 6052 3584 6058 3596
rect 6454 3584 6460 3596
rect 6052 3556 6460 3584
rect 6052 3544 6058 3556
rect 6454 3544 6460 3556
rect 6512 3544 6518 3596
rect 8018 3544 8024 3596
rect 8076 3584 8082 3596
rect 8297 3587 8355 3593
rect 8297 3584 8309 3587
rect 8076 3556 8309 3584
rect 8076 3544 8082 3556
rect 8297 3553 8309 3556
rect 8343 3553 8355 3587
rect 8297 3547 8355 3553
rect 9766 3544 9772 3596
rect 9824 3584 9830 3596
rect 10045 3587 10103 3593
rect 10045 3584 10057 3587
rect 9824 3556 10057 3584
rect 9824 3544 9830 3556
rect 10045 3553 10057 3556
rect 10091 3553 10103 3587
rect 10045 3547 10103 3553
rect 10781 3587 10839 3593
rect 10781 3553 10793 3587
rect 10827 3584 10839 3587
rect 10962 3584 10968 3596
rect 10827 3556 10968 3584
rect 10827 3553 10839 3556
rect 10781 3547 10839 3553
rect 10962 3544 10968 3556
rect 11020 3584 11026 3596
rect 11422 3584 11428 3596
rect 11020 3556 11428 3584
rect 11020 3544 11026 3556
rect 11422 3544 11428 3556
rect 11480 3544 11486 3596
rect 11609 3587 11667 3593
rect 11609 3553 11621 3587
rect 11655 3584 11667 3587
rect 11808 3584 11836 3612
rect 13078 3584 13084 3596
rect 11655 3556 13084 3584
rect 11655 3553 11667 3556
rect 11609 3547 11667 3553
rect 13078 3544 13084 3556
rect 13136 3544 13142 3596
rect 14734 3544 14740 3596
rect 14792 3584 14798 3596
rect 15289 3587 15347 3593
rect 15289 3584 15301 3587
rect 14792 3556 15301 3584
rect 14792 3544 14798 3556
rect 15289 3553 15301 3556
rect 15335 3553 15347 3587
rect 15289 3547 15347 3553
rect 16390 3544 16396 3596
rect 16448 3584 16454 3596
rect 16758 3584 16764 3596
rect 16448 3556 16764 3584
rect 16448 3544 16454 3556
rect 16758 3544 16764 3556
rect 16816 3544 16822 3596
rect 17586 3544 17592 3596
rect 17644 3584 17650 3596
rect 17865 3587 17923 3593
rect 17865 3584 17877 3587
rect 17644 3556 17877 3584
rect 17644 3544 17650 3556
rect 17865 3553 17877 3556
rect 17911 3553 17923 3587
rect 17865 3547 17923 3553
rect 19058 3544 19064 3596
rect 19116 3584 19122 3596
rect 19429 3587 19487 3593
rect 19429 3584 19441 3587
rect 19116 3556 19441 3584
rect 19116 3544 19122 3556
rect 19429 3553 19441 3556
rect 19475 3553 19487 3587
rect 21266 3584 21272 3596
rect 21227 3556 21272 3584
rect 19429 3547 19487 3553
rect 21266 3544 21272 3556
rect 21324 3544 21330 3596
rect 22462 3544 22468 3596
rect 22520 3584 22526 3596
rect 22833 3587 22891 3593
rect 22833 3584 22845 3587
rect 22520 3556 22845 3584
rect 22520 3544 22526 3556
rect 22833 3553 22845 3556
rect 22879 3553 22891 3587
rect 22833 3547 22891 3553
rect 24397 3587 24455 3593
rect 24397 3553 24409 3587
rect 24443 3584 24455 3587
rect 25792 3584 25820 3680
rect 24443 3556 25820 3584
rect 24443 3553 24455 3556
rect 24397 3547 24455 3553
rect 4706 3516 4712 3528
rect 4619 3488 4712 3516
rect 4706 3476 4712 3488
rect 4764 3516 4770 3528
rect 5442 3516 5448 3528
rect 4764 3488 5448 3516
rect 4764 3476 4770 3488
rect 5442 3476 5448 3488
rect 5500 3476 5506 3528
rect 9398 3476 9404 3528
rect 9456 3516 9462 3528
rect 10229 3519 10287 3525
rect 10229 3516 10241 3519
rect 9456 3488 10241 3516
rect 9456 3476 9462 3488
rect 10229 3485 10241 3488
rect 10275 3485 10287 3519
rect 10229 3479 10287 3485
rect 11054 3476 11060 3528
rect 11112 3516 11118 3528
rect 11793 3519 11851 3525
rect 11112 3488 11284 3516
rect 11112 3476 11118 3488
rect 7282 3448 7288 3460
rect 7243 3420 7288 3448
rect 7282 3408 7288 3420
rect 7340 3408 7346 3460
rect 9674 3448 9680 3460
rect 9635 3420 9680 3448
rect 9674 3408 9680 3420
rect 9732 3408 9738 3460
rect 10042 3408 10048 3460
rect 10100 3448 10106 3460
rect 10870 3448 10876 3460
rect 10100 3420 10876 3448
rect 10100 3408 10106 3420
rect 10870 3408 10876 3420
rect 10928 3408 10934 3460
rect 11256 3457 11284 3488
rect 11793 3485 11805 3519
rect 11839 3516 11851 3519
rect 13449 3519 13507 3525
rect 13449 3516 13461 3519
rect 11839 3488 13461 3516
rect 11839 3485 11851 3488
rect 11793 3479 11851 3485
rect 13449 3485 13461 3488
rect 13495 3516 13507 3519
rect 13817 3519 13875 3525
rect 13817 3516 13829 3519
rect 13495 3488 13829 3516
rect 13495 3485 13507 3488
rect 13449 3479 13507 3485
rect 13817 3485 13829 3488
rect 13863 3485 13875 3519
rect 13817 3479 13875 3485
rect 11241 3451 11299 3457
rect 11241 3417 11253 3451
rect 11287 3417 11299 3451
rect 11808 3448 11836 3479
rect 16850 3476 16856 3528
rect 16908 3516 16914 3528
rect 16945 3519 17003 3525
rect 16945 3516 16957 3519
rect 16908 3488 16957 3516
rect 16908 3476 16914 3488
rect 16945 3485 16957 3488
rect 16991 3516 17003 3519
rect 16991 3488 17724 3516
rect 16991 3485 17003 3488
rect 16945 3479 17003 3485
rect 11241 3411 11299 3417
rect 11716 3420 11836 3448
rect 12529 3451 12587 3457
rect 6822 3380 6828 3392
rect 3344 3352 6828 3380
rect 6822 3340 6828 3352
rect 6880 3340 6886 3392
rect 10778 3340 10784 3392
rect 10836 3380 10842 3392
rect 11054 3380 11060 3392
rect 10836 3352 11060 3380
rect 10836 3340 10842 3352
rect 11054 3340 11060 3352
rect 11112 3380 11118 3392
rect 11716 3380 11744 3420
rect 12529 3417 12541 3451
rect 12575 3448 12587 3451
rect 12802 3448 12808 3460
rect 12575 3420 12808 3448
rect 12575 3417 12587 3420
rect 12529 3411 12587 3417
rect 12802 3408 12808 3420
rect 12860 3408 12866 3460
rect 17494 3448 17500 3460
rect 17455 3420 17500 3448
rect 17494 3408 17500 3420
rect 17552 3408 17558 3460
rect 17696 3448 17724 3488
rect 17770 3476 17776 3528
rect 17828 3516 17834 3528
rect 17957 3519 18015 3525
rect 17957 3516 17969 3519
rect 17828 3488 17969 3516
rect 17828 3476 17834 3488
rect 17957 3485 17969 3488
rect 18003 3485 18015 3519
rect 17957 3479 18015 3485
rect 18049 3519 18107 3525
rect 18049 3485 18061 3519
rect 18095 3485 18107 3519
rect 18049 3479 18107 3485
rect 18064 3448 18092 3479
rect 18322 3476 18328 3528
rect 18380 3516 18386 3528
rect 19613 3519 19671 3525
rect 19613 3516 19625 3519
rect 18380 3488 19625 3516
rect 18380 3476 18386 3488
rect 19613 3485 19625 3488
rect 19659 3516 19671 3519
rect 20530 3516 20536 3528
rect 19659 3488 20536 3516
rect 19659 3485 19671 3488
rect 19613 3479 19671 3485
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 20714 3516 20720 3528
rect 20627 3488 20720 3516
rect 20714 3476 20720 3488
rect 20772 3516 20778 3528
rect 21542 3516 21548 3528
rect 20772 3488 21548 3516
rect 20772 3476 20778 3488
rect 21542 3476 21548 3488
rect 21600 3476 21606 3528
rect 18598 3448 18604 3460
rect 17696 3420 18604 3448
rect 18598 3408 18604 3420
rect 18656 3448 18662 3460
rect 18877 3451 18935 3457
rect 18877 3448 18889 3451
rect 18656 3420 18889 3448
rect 18656 3408 18662 3420
rect 18877 3417 18889 3420
rect 18923 3417 18935 3451
rect 22848 3448 22876 3547
rect 22922 3476 22928 3528
rect 22980 3516 22986 3528
rect 23017 3519 23075 3525
rect 23017 3516 23029 3519
rect 22980 3488 23029 3516
rect 22980 3476 22986 3488
rect 23017 3485 23029 3488
rect 23063 3485 23075 3519
rect 24670 3516 24676 3528
rect 24631 3488 24676 3516
rect 23017 3479 23075 3485
rect 24670 3476 24676 3488
rect 24728 3476 24734 3528
rect 25041 3451 25099 3457
rect 25041 3448 25053 3451
rect 22848 3420 25053 3448
rect 18877 3411 18935 3417
rect 25041 3417 25053 3420
rect 25087 3417 25099 3451
rect 25041 3411 25099 3417
rect 14366 3380 14372 3392
rect 11112 3352 11744 3380
rect 14327 3352 14372 3380
rect 11112 3340 11118 3352
rect 14366 3340 14372 3352
rect 14424 3340 14430 3392
rect 15654 3340 15660 3392
rect 15712 3380 15718 3392
rect 16669 3383 16727 3389
rect 16669 3380 16681 3383
rect 15712 3352 16681 3380
rect 15712 3340 15718 3352
rect 16669 3349 16681 3352
rect 16715 3349 16727 3383
rect 23750 3380 23756 3392
rect 23711 3352 23756 3380
rect 16669 3343 16727 3349
rect 23750 3340 23756 3352
rect 23808 3340 23814 3392
rect 24026 3380 24032 3392
rect 23987 3352 24032 3380
rect 24026 3340 24032 3352
rect 24084 3340 24090 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1397 3179 1455 3185
rect 1397 3145 1409 3179
rect 1443 3176 1455 3179
rect 1486 3176 1492 3188
rect 1443 3148 1492 3176
rect 1443 3145 1455 3148
rect 1397 3139 1455 3145
rect 1486 3136 1492 3148
rect 1544 3136 1550 3188
rect 2869 3179 2927 3185
rect 2869 3145 2881 3179
rect 2915 3176 2927 3179
rect 3326 3176 3332 3188
rect 2915 3148 3332 3176
rect 2915 3145 2927 3148
rect 2869 3139 2927 3145
rect 2409 3111 2467 3117
rect 2409 3108 2421 3111
rect 1872 3080 2421 3108
rect 1670 3000 1676 3052
rect 1728 3040 1734 3052
rect 1872 3049 1900 3080
rect 2409 3077 2421 3080
rect 2455 3077 2467 3111
rect 2409 3071 2467 3077
rect 1857 3043 1915 3049
rect 1857 3040 1869 3043
rect 1728 3012 1869 3040
rect 1728 3000 1734 3012
rect 1857 3009 1869 3012
rect 1903 3009 1915 3043
rect 1857 3003 1915 3009
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3040 2099 3043
rect 2222 3040 2228 3052
rect 2087 3012 2228 3040
rect 2087 3009 2099 3012
rect 2041 3003 2099 3009
rect 2222 3000 2228 3012
rect 2280 3000 2286 3052
rect 1762 2972 1768 2984
rect 1675 2944 1768 2972
rect 1762 2932 1768 2944
rect 1820 2972 1826 2984
rect 2884 2972 2912 3139
rect 3326 3136 3332 3148
rect 3384 3136 3390 3188
rect 3421 3179 3479 3185
rect 3421 3145 3433 3179
rect 3467 3176 3479 3179
rect 4706 3176 4712 3188
rect 3467 3148 4712 3176
rect 3467 3145 3479 3148
rect 3421 3139 3479 3145
rect 4706 3136 4712 3148
rect 4764 3136 4770 3188
rect 5258 3176 5264 3188
rect 5219 3148 5264 3176
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 5629 3179 5687 3185
rect 5629 3145 5641 3179
rect 5675 3176 5687 3179
rect 6086 3176 6092 3188
rect 5675 3148 6092 3176
rect 5675 3145 5687 3148
rect 5629 3139 5687 3145
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 6917 3179 6975 3185
rect 6917 3145 6929 3179
rect 6963 3176 6975 3179
rect 8202 3176 8208 3188
rect 6963 3148 8208 3176
rect 6963 3145 6975 3148
rect 6917 3139 6975 3145
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 9858 3176 9864 3188
rect 9771 3148 9864 3176
rect 9858 3136 9864 3148
rect 9916 3176 9922 3188
rect 12434 3176 12440 3188
rect 9916 3148 11836 3176
rect 12395 3148 12440 3176
rect 9916 3136 9922 3148
rect 7742 3068 7748 3120
rect 7800 3108 7806 3120
rect 8297 3111 8355 3117
rect 8297 3108 8309 3111
rect 7800 3080 8309 3108
rect 7800 3068 7806 3080
rect 8297 3077 8309 3080
rect 8343 3077 8355 3111
rect 8297 3071 8355 3077
rect 6273 3043 6331 3049
rect 6273 3009 6285 3043
rect 6319 3040 6331 3043
rect 7469 3043 7527 3049
rect 7469 3040 7481 3043
rect 6319 3012 7481 3040
rect 6319 3009 6331 3012
rect 6273 3003 6331 3009
rect 7469 3009 7481 3012
rect 7515 3040 7527 3043
rect 7650 3040 7656 3052
rect 7515 3012 7656 3040
rect 7515 3009 7527 3012
rect 7469 3003 7527 3009
rect 7650 3000 7656 3012
rect 7708 3000 7714 3052
rect 8312 3040 8340 3071
rect 9766 3068 9772 3120
rect 9824 3108 9830 3120
rect 10689 3111 10747 3117
rect 10689 3108 10701 3111
rect 9824 3080 10701 3108
rect 9824 3068 9830 3080
rect 10689 3077 10701 3080
rect 10735 3077 10747 3111
rect 11330 3108 11336 3120
rect 10689 3071 10747 3077
rect 11164 3080 11336 3108
rect 11164 3049 11192 3080
rect 11330 3068 11336 3080
rect 11388 3068 11394 3120
rect 11514 3068 11520 3120
rect 11572 3108 11578 3120
rect 11701 3111 11759 3117
rect 11701 3108 11713 3111
rect 11572 3080 11713 3108
rect 11572 3068 11578 3080
rect 11701 3077 11713 3080
rect 11747 3077 11759 3111
rect 11701 3071 11759 3077
rect 10597 3043 10655 3049
rect 8312 3012 8616 3040
rect 1820 2944 2912 2972
rect 1820 2932 1826 2944
rect 3142 2932 3148 2984
rect 3200 2972 3206 2984
rect 3513 2975 3571 2981
rect 3513 2972 3525 2975
rect 3200 2944 3525 2972
rect 3200 2932 3206 2944
rect 3513 2941 3525 2944
rect 3559 2972 3571 2975
rect 3602 2972 3608 2984
rect 3559 2944 3608 2972
rect 3559 2941 3571 2944
rect 3513 2935 3571 2941
rect 3602 2932 3608 2944
rect 3660 2932 3666 2984
rect 3786 2981 3792 2984
rect 3780 2972 3792 2981
rect 3747 2944 3792 2972
rect 3780 2935 3792 2944
rect 3786 2932 3792 2935
rect 3844 2932 3850 2984
rect 7190 2932 7196 2984
rect 7248 2972 7254 2984
rect 7285 2975 7343 2981
rect 7285 2972 7297 2975
rect 7248 2944 7297 2972
rect 7248 2932 7254 2944
rect 7285 2941 7297 2944
rect 7331 2941 7343 2975
rect 8018 2972 8024 2984
rect 7979 2944 8024 2972
rect 7285 2935 7343 2941
rect 8018 2932 8024 2944
rect 8076 2932 8082 2984
rect 8386 2932 8392 2984
rect 8444 2972 8450 2984
rect 8481 2975 8539 2981
rect 8481 2972 8493 2975
rect 8444 2944 8493 2972
rect 8444 2932 8450 2944
rect 8481 2941 8493 2944
rect 8527 2941 8539 2975
rect 8588 2972 8616 3012
rect 10597 3009 10609 3043
rect 10643 3040 10655 3043
rect 11149 3043 11207 3049
rect 11149 3040 11161 3043
rect 10643 3012 11161 3040
rect 10643 3009 10655 3012
rect 10597 3003 10655 3009
rect 11149 3009 11161 3012
rect 11195 3009 11207 3043
rect 11149 3003 11207 3009
rect 11241 3043 11299 3049
rect 11241 3009 11253 3043
rect 11287 3009 11299 3043
rect 11808 3040 11836 3148
rect 12434 3136 12440 3148
rect 12492 3136 12498 3188
rect 14826 3176 14832 3188
rect 14787 3148 14832 3176
rect 14826 3136 14832 3148
rect 14884 3176 14890 3188
rect 15654 3176 15660 3188
rect 14884 3148 15660 3176
rect 14884 3136 14890 3148
rect 13081 3043 13139 3049
rect 13081 3040 13093 3043
rect 11808 3012 13093 3040
rect 11241 3003 11299 3009
rect 13081 3009 13093 3012
rect 13127 3040 13139 3043
rect 14185 3043 14243 3049
rect 14185 3040 14197 3043
rect 13127 3012 14197 3040
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 14185 3009 14197 3012
rect 14231 3009 14243 3043
rect 14185 3003 14243 3009
rect 8754 2981 8760 2984
rect 8737 2975 8760 2981
rect 8737 2972 8749 2975
rect 8588 2944 8749 2972
rect 8481 2935 8539 2941
rect 8737 2941 8749 2944
rect 8812 2972 8818 2984
rect 8812 2944 8885 2972
rect 8737 2935 8760 2941
rect 1578 2864 1584 2916
rect 1636 2904 1642 2916
rect 2498 2904 2504 2916
rect 1636 2876 2504 2904
rect 1636 2864 1642 2876
rect 2498 2864 2504 2876
rect 2556 2864 2562 2916
rect 5721 2907 5779 2913
rect 4724 2876 5212 2904
rect 658 2796 664 2848
rect 716 2836 722 2848
rect 4724 2836 4752 2876
rect 716 2808 4752 2836
rect 4893 2839 4951 2845
rect 716 2796 722 2808
rect 4893 2805 4905 2839
rect 4939 2836 4951 2839
rect 5074 2836 5080 2848
rect 4939 2808 5080 2836
rect 4939 2805 4951 2808
rect 4893 2799 4951 2805
rect 5074 2796 5080 2808
rect 5132 2796 5138 2848
rect 5184 2836 5212 2876
rect 5721 2873 5733 2907
rect 5767 2904 5779 2907
rect 6270 2904 6276 2916
rect 5767 2876 6276 2904
rect 5767 2873 5779 2876
rect 5721 2867 5779 2873
rect 6270 2864 6276 2876
rect 6328 2864 6334 2916
rect 6638 2904 6644 2916
rect 6551 2876 6644 2904
rect 6638 2864 6644 2876
rect 6696 2904 6702 2916
rect 7377 2907 7435 2913
rect 7377 2904 7389 2907
rect 6696 2876 7389 2904
rect 6696 2864 6702 2876
rect 7377 2873 7389 2876
rect 7423 2904 7435 2907
rect 7926 2904 7932 2916
rect 7423 2876 7932 2904
rect 7423 2873 7435 2876
rect 7377 2867 7435 2873
rect 7926 2864 7932 2876
rect 7984 2864 7990 2916
rect 8496 2904 8524 2935
rect 8754 2932 8760 2935
rect 8812 2932 8818 2944
rect 9950 2932 9956 2984
rect 10008 2972 10014 2984
rect 10137 2975 10195 2981
rect 10137 2972 10149 2975
rect 10008 2944 10149 2972
rect 10008 2932 10014 2944
rect 10137 2941 10149 2944
rect 10183 2972 10195 2975
rect 11054 2972 11060 2984
rect 10183 2944 11060 2972
rect 10183 2941 10195 2944
rect 10137 2935 10195 2941
rect 11054 2932 11060 2944
rect 11112 2972 11118 2984
rect 11256 2972 11284 3003
rect 14366 3000 14372 3052
rect 14424 3040 14430 3052
rect 15580 3049 15608 3148
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 15930 3176 15936 3188
rect 15891 3148 15936 3176
rect 15930 3136 15936 3148
rect 15988 3136 15994 3188
rect 18046 3176 18052 3188
rect 18007 3148 18052 3176
rect 18046 3136 18052 3148
rect 18104 3136 18110 3188
rect 19518 3176 19524 3188
rect 19479 3148 19524 3176
rect 19518 3136 19524 3148
rect 19576 3136 19582 3188
rect 20530 3136 20536 3188
rect 20588 3176 20594 3188
rect 20625 3179 20683 3185
rect 20625 3176 20637 3179
rect 20588 3148 20637 3176
rect 20588 3136 20594 3148
rect 20625 3145 20637 3148
rect 20671 3145 20683 3179
rect 21174 3176 21180 3188
rect 21135 3148 21180 3176
rect 20625 3139 20683 3145
rect 21174 3136 21180 3148
rect 21232 3136 21238 3188
rect 25038 3176 25044 3188
rect 24999 3148 25044 3176
rect 25038 3136 25044 3148
rect 25096 3136 25102 3188
rect 26326 3176 26332 3188
rect 26287 3148 26332 3176
rect 26326 3136 26332 3148
rect 26384 3136 26390 3188
rect 16206 3068 16212 3120
rect 16264 3108 16270 3120
rect 19058 3108 19064 3120
rect 16264 3080 19064 3108
rect 16264 3068 16270 3080
rect 19058 3068 19064 3080
rect 19116 3068 19122 3120
rect 19610 3108 19616 3120
rect 19571 3080 19616 3108
rect 19610 3068 19616 3080
rect 19668 3068 19674 3120
rect 15565 3043 15623 3049
rect 14424 3012 15424 3040
rect 14424 3000 14430 3012
rect 12802 2972 12808 2984
rect 11112 2944 11284 2972
rect 12763 2944 12808 2972
rect 11112 2932 11118 2944
rect 12802 2932 12808 2944
rect 12860 2932 12866 2984
rect 12897 2975 12955 2981
rect 12897 2941 12909 2975
rect 12943 2972 12955 2975
rect 13817 2975 13875 2981
rect 13817 2972 13829 2975
rect 12943 2944 13829 2972
rect 12943 2941 12955 2944
rect 12897 2935 12955 2941
rect 13817 2941 13829 2944
rect 13863 2972 13875 2975
rect 13906 2972 13912 2984
rect 13863 2944 13912 2972
rect 13863 2941 13875 2944
rect 13817 2935 13875 2941
rect 13906 2932 13912 2944
rect 13964 2932 13970 2984
rect 15286 2972 15292 2984
rect 15247 2944 15292 2972
rect 15286 2932 15292 2944
rect 15344 2932 15350 2984
rect 15396 2981 15424 3012
rect 15565 3009 15577 3043
rect 15611 3009 15623 3043
rect 15565 3003 15623 3009
rect 16393 3043 16451 3049
rect 16393 3009 16405 3043
rect 16439 3040 16451 3043
rect 16669 3043 16727 3049
rect 16669 3040 16681 3043
rect 16439 3012 16681 3040
rect 16439 3009 16451 3012
rect 16393 3003 16451 3009
rect 16669 3009 16681 3012
rect 16715 3040 16727 3043
rect 16758 3040 16764 3052
rect 16715 3012 16764 3040
rect 16715 3009 16727 3012
rect 16669 3003 16727 3009
rect 16758 3000 16764 3012
rect 16816 3000 16822 3052
rect 18598 3040 18604 3052
rect 18559 3012 18604 3040
rect 18598 3000 18604 3012
rect 18656 3000 18662 3052
rect 20162 3040 20168 3052
rect 20123 3012 20168 3040
rect 20162 3000 20168 3012
rect 20220 3000 20226 3052
rect 20806 3000 20812 3052
rect 20864 3040 20870 3052
rect 20993 3043 21051 3049
rect 20993 3040 21005 3043
rect 20864 3012 21005 3040
rect 20864 3000 20870 3012
rect 20993 3009 21005 3012
rect 21039 3009 21051 3043
rect 21634 3040 21640 3052
rect 21595 3012 21640 3040
rect 20993 3003 21051 3009
rect 15381 2975 15439 2981
rect 15381 2941 15393 2975
rect 15427 2972 15439 2975
rect 16298 2972 16304 2984
rect 15427 2944 16304 2972
rect 15427 2941 15439 2944
rect 15381 2935 15439 2941
rect 16298 2932 16304 2944
rect 16356 2932 16362 2984
rect 16482 2972 16488 2984
rect 16443 2944 16488 2972
rect 16482 2932 16488 2944
rect 16540 2932 16546 2984
rect 18509 2975 18567 2981
rect 18509 2941 18521 2975
rect 18555 2972 18567 2975
rect 18874 2972 18880 2984
rect 18555 2944 18880 2972
rect 18555 2941 18567 2944
rect 18509 2935 18567 2941
rect 18874 2932 18880 2944
rect 18932 2932 18938 2984
rect 20070 2972 20076 2984
rect 20031 2944 20076 2972
rect 20070 2932 20076 2944
rect 20128 2972 20134 2984
rect 20714 2972 20720 2984
rect 20128 2944 20720 2972
rect 20128 2932 20134 2944
rect 20714 2932 20720 2944
rect 20772 2932 20778 2984
rect 9582 2904 9588 2916
rect 8496 2876 9588 2904
rect 9582 2864 9588 2876
rect 9640 2864 9646 2916
rect 12253 2907 12311 2913
rect 12253 2904 12265 2907
rect 10612 2876 12265 2904
rect 10612 2836 10640 2876
rect 12253 2873 12265 2876
rect 12299 2904 12311 2907
rect 12710 2904 12716 2916
rect 12299 2876 12716 2904
rect 12299 2873 12311 2876
rect 12253 2867 12311 2873
rect 12710 2864 12716 2876
rect 12768 2864 12774 2916
rect 13630 2904 13636 2916
rect 12820 2876 13636 2904
rect 12820 2848 12848 2876
rect 13630 2864 13636 2876
rect 13688 2864 13694 2916
rect 15562 2864 15568 2916
rect 15620 2904 15626 2916
rect 18230 2904 18236 2916
rect 15620 2876 18236 2904
rect 15620 2864 15626 2876
rect 18230 2864 18236 2876
rect 18288 2864 18294 2916
rect 21008 2904 21036 3003
rect 21634 3000 21640 3012
rect 21692 3000 21698 3052
rect 21729 3043 21787 3049
rect 21729 3009 21741 3043
rect 21775 3040 21787 3043
rect 22465 3043 22523 3049
rect 22465 3040 22477 3043
rect 21775 3012 22477 3040
rect 21775 3009 21787 3012
rect 21729 3003 21787 3009
rect 22465 3009 22477 3012
rect 22511 3040 22523 3043
rect 22922 3040 22928 3052
rect 22511 3012 22928 3040
rect 22511 3009 22523 3012
rect 22465 3003 22523 3009
rect 21450 2932 21456 2984
rect 21508 2972 21514 2984
rect 21545 2975 21603 2981
rect 21545 2972 21557 2975
rect 21508 2944 21557 2972
rect 21508 2932 21514 2944
rect 21545 2941 21557 2944
rect 21591 2941 21603 2975
rect 21744 2972 21772 3003
rect 22922 3000 22928 3012
rect 22980 3000 22986 3052
rect 23014 3000 23020 3052
rect 23072 3040 23078 3052
rect 23474 3040 23480 3052
rect 23072 3012 23480 3040
rect 23072 3000 23078 3012
rect 23474 3000 23480 3012
rect 23532 3040 23538 3052
rect 24213 3043 24271 3049
rect 24213 3040 24225 3043
rect 23532 3012 24225 3040
rect 23532 3000 23538 3012
rect 24213 3009 24225 3012
rect 24259 3040 24271 3043
rect 24670 3040 24676 3052
rect 24259 3012 24676 3040
rect 24259 3009 24271 3012
rect 24213 3003 24271 3009
rect 24670 3000 24676 3012
rect 24728 3000 24734 3052
rect 21545 2935 21603 2941
rect 21652 2944 21772 2972
rect 21652 2904 21680 2944
rect 23750 2932 23756 2984
rect 23808 2972 23814 2984
rect 24026 2972 24032 2984
rect 23808 2944 24032 2972
rect 23808 2932 23814 2944
rect 24026 2932 24032 2944
rect 24084 2932 24090 2984
rect 25225 2975 25283 2981
rect 25225 2941 25237 2975
rect 25271 2972 25283 2975
rect 25314 2972 25320 2984
rect 25271 2944 25320 2972
rect 25271 2941 25283 2944
rect 25225 2935 25283 2941
rect 25314 2932 25320 2944
rect 25372 2972 25378 2984
rect 25961 2975 26019 2981
rect 25961 2972 25973 2975
rect 25372 2944 25973 2972
rect 25372 2932 25378 2944
rect 25961 2941 25973 2944
rect 26007 2941 26019 2975
rect 25961 2935 26019 2941
rect 21008 2876 21680 2904
rect 23477 2907 23535 2913
rect 23477 2873 23489 2907
rect 23523 2904 23535 2907
rect 23934 2904 23940 2916
rect 23523 2876 23940 2904
rect 23523 2873 23535 2876
rect 23477 2867 23535 2873
rect 23934 2864 23940 2876
rect 23992 2904 23998 2916
rect 24121 2907 24179 2913
rect 24121 2904 24133 2907
rect 23992 2876 24133 2904
rect 23992 2864 23998 2876
rect 24121 2873 24133 2876
rect 24167 2873 24179 2907
rect 25498 2904 25504 2916
rect 25459 2876 25504 2904
rect 24121 2867 24179 2873
rect 25498 2864 25504 2876
rect 25556 2864 25562 2916
rect 5184 2808 10640 2836
rect 10962 2796 10968 2848
rect 11020 2836 11026 2848
rect 11057 2839 11115 2845
rect 11057 2836 11069 2839
rect 11020 2808 11069 2836
rect 11020 2796 11026 2808
rect 11057 2805 11069 2808
rect 11103 2805 11115 2839
rect 11057 2799 11115 2805
rect 12802 2796 12808 2848
rect 12860 2796 12866 2848
rect 13446 2836 13452 2848
rect 13407 2808 13452 2836
rect 13446 2796 13452 2808
rect 13504 2796 13510 2848
rect 14918 2836 14924 2848
rect 14879 2808 14924 2836
rect 14918 2796 14924 2808
rect 14976 2796 14982 2848
rect 17494 2836 17500 2848
rect 17455 2808 17500 2836
rect 17494 2796 17500 2808
rect 17552 2836 17558 2848
rect 17770 2836 17776 2848
rect 17552 2808 17776 2836
rect 17552 2796 17558 2808
rect 17770 2796 17776 2808
rect 17828 2796 17834 2848
rect 18138 2796 18144 2848
rect 18196 2836 18202 2848
rect 18414 2836 18420 2848
rect 18196 2808 18420 2836
rect 18196 2796 18202 2808
rect 18414 2796 18420 2808
rect 18472 2796 18478 2848
rect 19981 2839 20039 2845
rect 19981 2805 19993 2839
rect 20027 2836 20039 2839
rect 20070 2836 20076 2848
rect 20027 2808 20076 2836
rect 20027 2805 20039 2808
rect 19981 2799 20039 2805
rect 20070 2796 20076 2808
rect 20128 2836 20134 2848
rect 20254 2836 20260 2848
rect 20128 2808 20260 2836
rect 20128 2796 20134 2808
rect 20254 2796 20260 2808
rect 20312 2796 20318 2848
rect 23014 2836 23020 2848
rect 22975 2808 23020 2836
rect 23014 2796 23020 2808
rect 23072 2796 23078 2848
rect 23658 2836 23664 2848
rect 23619 2808 23664 2836
rect 23658 2796 23664 2808
rect 23716 2796 23722 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1397 2635 1455 2641
rect 1397 2601 1409 2635
rect 1443 2632 1455 2635
rect 2130 2632 2136 2644
rect 1443 2604 2136 2632
rect 1443 2601 1455 2604
rect 1397 2595 1455 2601
rect 2130 2592 2136 2604
rect 2188 2592 2194 2644
rect 3605 2635 3663 2641
rect 3605 2601 3617 2635
rect 3651 2632 3663 2635
rect 3786 2632 3792 2644
rect 3651 2604 3792 2632
rect 3651 2601 3663 2604
rect 3605 2595 3663 2601
rect 3786 2592 3792 2604
rect 3844 2592 3850 2644
rect 5994 2592 6000 2644
rect 6052 2632 6058 2644
rect 6089 2635 6147 2641
rect 6089 2632 6101 2635
rect 6052 2604 6101 2632
rect 6052 2592 6058 2604
rect 6089 2601 6101 2604
rect 6135 2601 6147 2635
rect 7190 2632 7196 2644
rect 7151 2604 7196 2632
rect 6089 2595 6147 2601
rect 7190 2592 7196 2604
rect 7248 2592 7254 2644
rect 8846 2632 8852 2644
rect 8807 2604 8852 2632
rect 8846 2592 8852 2604
rect 8904 2592 8910 2644
rect 9398 2592 9404 2644
rect 9456 2632 9462 2644
rect 9493 2635 9551 2641
rect 9493 2632 9505 2635
rect 9456 2604 9505 2632
rect 9456 2592 9462 2604
rect 9493 2601 9505 2604
rect 9539 2601 9551 2635
rect 9493 2595 9551 2601
rect 9582 2592 9588 2644
rect 9640 2632 9646 2644
rect 11701 2635 11759 2641
rect 9640 2604 10180 2632
rect 9640 2592 9646 2604
rect 1670 2524 1676 2576
rect 1728 2564 1734 2576
rect 1765 2567 1823 2573
rect 1765 2564 1777 2567
rect 1728 2536 1777 2564
rect 1728 2524 1734 2536
rect 1765 2533 1777 2536
rect 1811 2564 1823 2567
rect 2869 2567 2927 2573
rect 2869 2564 2881 2567
rect 1811 2536 2881 2564
rect 1811 2533 1823 2536
rect 1765 2527 1823 2533
rect 2869 2533 2881 2536
rect 2915 2564 2927 2567
rect 4614 2564 4620 2576
rect 2915 2536 4620 2564
rect 2915 2533 2927 2536
rect 2869 2527 2927 2533
rect 4614 2524 4620 2536
rect 4672 2524 4678 2576
rect 5074 2524 5080 2576
rect 5132 2564 5138 2576
rect 5721 2567 5779 2573
rect 5721 2564 5733 2567
rect 5132 2536 5733 2564
rect 5132 2524 5138 2536
rect 5721 2533 5733 2536
rect 5767 2533 5779 2567
rect 8386 2564 8392 2576
rect 5721 2527 5779 2533
rect 7484 2536 8392 2564
rect 1394 2456 1400 2508
rect 1452 2496 1458 2508
rect 1857 2499 1915 2505
rect 1857 2496 1869 2499
rect 1452 2468 1869 2496
rect 1452 2456 1458 2468
rect 1857 2465 1869 2468
rect 1903 2496 1915 2499
rect 2409 2499 2467 2505
rect 2409 2496 2421 2499
rect 1903 2468 2421 2496
rect 1903 2465 1915 2468
rect 1857 2459 1915 2465
rect 2409 2465 2421 2468
rect 2455 2465 2467 2499
rect 2409 2459 2467 2465
rect 3142 2456 3148 2508
rect 3200 2496 3206 2508
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 3200 2468 4077 2496
rect 3200 2456 3206 2468
rect 4065 2465 4077 2468
rect 4111 2465 4123 2499
rect 4065 2459 4123 2465
rect 4332 2499 4390 2505
rect 4332 2465 4344 2499
rect 4378 2496 4390 2499
rect 5092 2496 5120 2524
rect 7484 2505 7512 2536
rect 8386 2524 8392 2536
rect 8444 2524 8450 2576
rect 9217 2567 9275 2573
rect 9217 2533 9229 2567
rect 9263 2564 9275 2567
rect 9766 2564 9772 2576
rect 9263 2536 9772 2564
rect 9263 2533 9275 2536
rect 9217 2527 9275 2533
rect 9766 2524 9772 2536
rect 9824 2524 9830 2576
rect 7742 2505 7748 2508
rect 4378 2468 5120 2496
rect 7469 2499 7527 2505
rect 4378 2465 4390 2468
rect 4332 2459 4390 2465
rect 7469 2465 7481 2499
rect 7515 2465 7527 2499
rect 7736 2496 7748 2505
rect 7469 2459 7527 2465
rect 7576 2468 7748 2496
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2428 2099 2431
rect 2222 2428 2228 2440
rect 2087 2400 2228 2428
rect 2087 2397 2099 2400
rect 2041 2391 2099 2397
rect 2222 2388 2228 2400
rect 2280 2388 2286 2440
rect 2958 2428 2964 2440
rect 2919 2400 2964 2428
rect 2958 2388 2964 2400
rect 3016 2388 3022 2440
rect 6733 2431 6791 2437
rect 6733 2397 6745 2431
rect 6779 2428 6791 2431
rect 7576 2428 7604 2468
rect 7736 2459 7748 2468
rect 7742 2456 7748 2459
rect 7800 2456 7806 2508
rect 6779 2400 7604 2428
rect 10152 2428 10180 2604
rect 11701 2601 11713 2635
rect 11747 2632 11759 2635
rect 13998 2632 14004 2644
rect 11747 2604 12388 2632
rect 13959 2604 14004 2632
rect 11747 2601 11759 2604
rect 11701 2595 11759 2601
rect 11790 2524 11796 2576
rect 11848 2564 11854 2576
rect 11977 2567 12035 2573
rect 11977 2564 11989 2567
rect 11848 2536 11989 2564
rect 11848 2524 11854 2536
rect 11977 2533 11989 2536
rect 12023 2533 12035 2567
rect 12360 2564 12388 2604
rect 13998 2592 14004 2604
rect 14056 2592 14062 2644
rect 16390 2592 16396 2644
rect 16448 2632 16454 2644
rect 16485 2635 16543 2641
rect 16485 2632 16497 2635
rect 16448 2604 16497 2632
rect 16448 2592 16454 2604
rect 16485 2601 16497 2604
rect 16531 2601 16543 2635
rect 18138 2632 18144 2644
rect 18099 2604 18144 2632
rect 16485 2595 16543 2601
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 18690 2632 18696 2644
rect 18651 2604 18696 2632
rect 18690 2592 18696 2604
rect 18748 2592 18754 2644
rect 19705 2635 19763 2641
rect 19705 2601 19717 2635
rect 19751 2632 19763 2635
rect 20162 2632 20168 2644
rect 19751 2604 20168 2632
rect 19751 2601 19763 2604
rect 19705 2595 19763 2601
rect 14550 2564 14556 2576
rect 12360 2536 12572 2564
rect 14511 2536 14556 2564
rect 11977 2527 12035 2533
rect 10594 2505 10600 2508
rect 10229 2499 10287 2505
rect 10229 2465 10241 2499
rect 10275 2496 10287 2499
rect 10588 2496 10600 2505
rect 10275 2468 10600 2496
rect 10275 2465 10287 2468
rect 10229 2459 10287 2465
rect 10588 2459 10600 2468
rect 10594 2456 10600 2459
rect 10652 2456 10658 2508
rect 12544 2496 12572 2536
rect 14550 2524 14556 2536
rect 14608 2524 14614 2576
rect 14752 2536 16712 2564
rect 12888 2499 12946 2505
rect 12888 2496 12900 2499
rect 12544 2468 12900 2496
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 10152 2400 10333 2428
rect 6779 2397 6791 2400
rect 6733 2391 6791 2397
rect 10321 2397 10333 2400
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 12437 2431 12495 2437
rect 12437 2397 12449 2431
rect 12483 2428 12495 2431
rect 12544 2428 12572 2468
rect 12888 2465 12900 2468
rect 12934 2496 12946 2499
rect 14752 2496 14780 2536
rect 12934 2468 14780 2496
rect 15841 2499 15899 2505
rect 12934 2465 12946 2468
rect 12888 2459 12946 2465
rect 15841 2465 15853 2499
rect 15887 2465 15899 2499
rect 15841 2459 15899 2465
rect 12483 2400 12572 2428
rect 12621 2431 12679 2437
rect 12483 2397 12495 2400
rect 12437 2391 12495 2397
rect 12621 2397 12633 2431
rect 12667 2397 12679 2431
rect 12621 2391 12679 2397
rect 5442 2292 5448 2304
rect 5403 2264 5448 2292
rect 5442 2252 5448 2264
rect 5500 2252 5506 2304
rect 10336 2292 10364 2391
rect 12636 2292 12664 2391
rect 14458 2388 14464 2440
rect 14516 2428 14522 2440
rect 14829 2431 14887 2437
rect 14829 2428 14841 2431
rect 14516 2400 14841 2428
rect 14516 2388 14522 2400
rect 14829 2397 14841 2400
rect 14875 2428 14887 2431
rect 15856 2428 15884 2459
rect 14875 2400 15884 2428
rect 15933 2431 15991 2437
rect 14875 2397 14887 2400
rect 14829 2391 14887 2397
rect 15933 2397 15945 2431
rect 15979 2397 15991 2431
rect 15933 2391 15991 2397
rect 16117 2431 16175 2437
rect 16117 2397 16129 2431
rect 16163 2428 16175 2431
rect 16390 2428 16396 2440
rect 16163 2400 16396 2428
rect 16163 2397 16175 2400
rect 16117 2391 16175 2397
rect 13722 2320 13728 2372
rect 13780 2360 13786 2372
rect 15473 2363 15531 2369
rect 15473 2360 15485 2363
rect 13780 2332 15485 2360
rect 13780 2320 13786 2332
rect 15473 2329 15485 2332
rect 15519 2329 15531 2363
rect 15473 2323 15531 2329
rect 15286 2292 15292 2304
rect 10336 2264 12664 2292
rect 15247 2264 15292 2292
rect 15286 2252 15292 2264
rect 15344 2292 15350 2304
rect 15948 2292 15976 2391
rect 16390 2388 16396 2400
rect 16448 2388 16454 2440
rect 16684 2428 16712 2536
rect 16758 2456 16764 2508
rect 16816 2496 16822 2508
rect 17037 2499 17095 2505
rect 17037 2496 17049 2499
rect 16816 2468 17049 2496
rect 16816 2456 16822 2468
rect 17037 2465 17049 2468
rect 17083 2465 17095 2499
rect 17037 2459 17095 2465
rect 18322 2456 18328 2508
rect 18380 2496 18386 2508
rect 18785 2499 18843 2505
rect 18785 2496 18797 2499
rect 18380 2468 18797 2496
rect 18380 2456 18386 2468
rect 18785 2465 18797 2468
rect 18831 2465 18843 2499
rect 18785 2459 18843 2465
rect 16945 2431 17003 2437
rect 16945 2428 16957 2431
rect 16684 2400 16957 2428
rect 16945 2397 16957 2400
rect 16991 2428 17003 2431
rect 18969 2431 19027 2437
rect 18969 2428 18981 2431
rect 16991 2400 18981 2428
rect 16991 2397 17003 2400
rect 16945 2391 17003 2397
rect 18969 2397 18981 2400
rect 19015 2428 19027 2431
rect 19720 2428 19748 2595
rect 20162 2592 20168 2604
rect 20220 2592 20226 2644
rect 20714 2592 20720 2644
rect 20772 2632 20778 2644
rect 21177 2635 21235 2641
rect 21177 2632 21189 2635
rect 20772 2604 21189 2632
rect 20772 2592 20778 2604
rect 21177 2601 21189 2604
rect 21223 2601 21235 2635
rect 21634 2632 21640 2644
rect 21595 2604 21640 2632
rect 21177 2595 21235 2601
rect 21634 2592 21640 2604
rect 21692 2592 21698 2644
rect 22738 2632 22744 2644
rect 22699 2604 22744 2632
rect 22738 2592 22744 2604
rect 22796 2592 22802 2644
rect 23934 2592 23940 2644
rect 23992 2632 23998 2644
rect 24029 2635 24087 2641
rect 24029 2632 24041 2635
rect 23992 2604 24041 2632
rect 23992 2592 23998 2604
rect 24029 2601 24041 2604
rect 24075 2601 24087 2635
rect 24029 2595 24087 2601
rect 20898 2564 20904 2576
rect 20859 2536 20904 2564
rect 20898 2524 20904 2536
rect 20956 2564 20962 2576
rect 21545 2567 21603 2573
rect 21545 2564 21557 2567
rect 20956 2536 21557 2564
rect 20956 2524 20962 2536
rect 21545 2533 21557 2536
rect 21591 2533 21603 2567
rect 21545 2527 21603 2533
rect 19978 2496 19984 2508
rect 19939 2468 19984 2496
rect 19978 2456 19984 2468
rect 20036 2496 20042 2508
rect 20533 2499 20591 2505
rect 20533 2496 20545 2499
rect 20036 2468 20545 2496
rect 20036 2456 20042 2468
rect 20533 2465 20545 2468
rect 20579 2465 20591 2499
rect 22756 2496 22784 2592
rect 24044 2564 24072 2595
rect 24762 2592 24768 2644
rect 24820 2632 24826 2644
rect 25409 2635 25467 2641
rect 25409 2632 25421 2635
rect 24820 2604 25421 2632
rect 24820 2592 24826 2604
rect 25409 2601 25421 2604
rect 25455 2601 25467 2635
rect 26418 2632 26424 2644
rect 26379 2604 26424 2632
rect 25409 2595 25467 2601
rect 26418 2592 26424 2604
rect 26476 2592 26482 2644
rect 26053 2567 26111 2573
rect 26053 2564 26065 2567
rect 24044 2536 26065 2564
rect 26053 2533 26065 2536
rect 26099 2533 26111 2567
rect 26053 2527 26111 2533
rect 22833 2499 22891 2505
rect 22833 2496 22845 2499
rect 22756 2468 22845 2496
rect 20533 2459 20591 2465
rect 22833 2465 22845 2468
rect 22879 2465 22891 2499
rect 22833 2459 22891 2465
rect 23474 2456 23480 2508
rect 23532 2496 23538 2508
rect 24397 2499 24455 2505
rect 24397 2496 24409 2499
rect 23532 2468 24409 2496
rect 23532 2456 23538 2468
rect 24397 2465 24409 2468
rect 24443 2465 24455 2499
rect 24397 2459 24455 2465
rect 21726 2428 21732 2440
rect 19015 2400 19748 2428
rect 21687 2400 21732 2428
rect 19015 2397 19027 2400
rect 18969 2391 19027 2397
rect 21726 2388 21732 2400
rect 21784 2428 21790 2440
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 21784 2400 22201 2428
rect 21784 2388 21790 2400
rect 22189 2397 22201 2400
rect 22235 2428 22247 2431
rect 23014 2428 23020 2440
rect 22235 2400 23020 2428
rect 22235 2397 22247 2400
rect 22189 2391 22247 2397
rect 23014 2388 23020 2400
rect 23072 2388 23078 2440
rect 23658 2388 23664 2440
rect 23716 2428 23722 2440
rect 23753 2431 23811 2437
rect 23753 2428 23765 2431
rect 23716 2400 23765 2428
rect 23716 2388 23722 2400
rect 23753 2397 23765 2400
rect 23799 2428 23811 2431
rect 24489 2431 24547 2437
rect 24489 2428 24501 2431
rect 23799 2400 24501 2428
rect 23799 2397 23811 2400
rect 23753 2391 23811 2397
rect 24489 2397 24501 2400
rect 24535 2397 24547 2431
rect 24670 2428 24676 2440
rect 24631 2400 24676 2428
rect 24489 2391 24547 2397
rect 24670 2388 24676 2400
rect 24728 2428 24734 2440
rect 25041 2431 25099 2437
rect 25041 2428 25053 2431
rect 24728 2400 25053 2428
rect 24728 2388 24734 2400
rect 25041 2397 25053 2400
rect 25087 2397 25099 2431
rect 25590 2428 25596 2440
rect 25551 2400 25596 2428
rect 25041 2391 25099 2397
rect 25590 2388 25596 2400
rect 25648 2388 25654 2440
rect 15344 2264 15976 2292
rect 15344 2252 15350 2264
rect 17126 2252 17132 2304
rect 17184 2292 17190 2304
rect 17221 2295 17279 2301
rect 17221 2292 17233 2295
rect 17184 2264 17233 2292
rect 17184 2252 17190 2264
rect 17221 2261 17233 2264
rect 17267 2261 17279 2295
rect 17586 2292 17592 2304
rect 17547 2264 17592 2292
rect 17221 2255 17279 2261
rect 17586 2252 17592 2264
rect 17644 2252 17650 2304
rect 18322 2292 18328 2304
rect 18283 2264 18328 2292
rect 18322 2252 18328 2264
rect 18380 2252 18386 2304
rect 20162 2292 20168 2304
rect 20123 2264 20168 2292
rect 20162 2252 20168 2264
rect 20220 2252 20226 2304
rect 23014 2292 23020 2304
rect 22975 2264 23020 2292
rect 23014 2252 23020 2264
rect 23072 2252 23078 2304
rect 23474 2292 23480 2304
rect 23435 2264 23480 2292
rect 23474 2252 23480 2264
rect 23532 2252 23538 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 11514 2048 11520 2100
rect 11572 2088 11578 2100
rect 13446 2088 13452 2100
rect 11572 2060 13452 2088
rect 11572 2048 11578 2060
rect 13446 2048 13452 2060
rect 13504 2048 13510 2100
rect 12526 1912 12532 1964
rect 12584 1952 12590 1964
rect 18782 1952 18788 1964
rect 12584 1924 18788 1952
rect 12584 1912 12590 1924
rect 18782 1912 18788 1924
rect 18840 1912 18846 1964
rect 22646 552 22652 604
rect 22704 592 22710 604
rect 22738 592 22744 604
rect 22704 564 22744 592
rect 22704 552 22710 564
rect 22738 552 22744 564
rect 22796 552 22802 604
rect 23750 552 23756 604
rect 23808 592 23814 604
rect 25682 592 25688 604
rect 23808 564 25688 592
rect 23808 552 23814 564
rect 25682 552 25688 564
rect 25740 552 25746 604
<< via1 >>
rect 3516 27548 3568 27600
rect 9128 27548 9180 27600
rect 3332 26188 3384 26240
rect 11152 26256 11204 26308
rect 10784 26188 10836 26240
rect 14464 26256 14516 26308
rect 16120 26256 16172 26308
rect 12348 26188 12400 26240
rect 19524 26188 19576 26240
rect 5540 26120 5592 26172
rect 18144 26120 18196 26172
rect 6736 26052 6788 26104
rect 11888 26052 11940 26104
rect 13452 26052 13504 26104
rect 18880 26052 18932 26104
rect 9220 25984 9272 26036
rect 16580 25984 16632 26036
rect 4620 25916 4672 25968
rect 11796 25916 11848 25968
rect 11888 25916 11940 25968
rect 25136 25916 25188 25968
rect 9956 25848 10008 25900
rect 12164 25848 12216 25900
rect 13544 25848 13596 25900
rect 21272 25848 21324 25900
rect 8024 25780 8076 25832
rect 17132 25780 17184 25832
rect 19524 25780 19576 25832
rect 8944 25712 8996 25764
rect 13820 25712 13872 25764
rect 17224 25712 17276 25764
rect 19156 25712 19208 25764
rect 10692 25644 10744 25696
rect 18328 25644 18380 25696
rect 21916 25644 21968 25696
rect 26516 25644 26568 25696
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 2228 25440 2280 25492
rect 10692 25440 10744 25492
rect 12256 25440 12308 25492
rect 12348 25440 12400 25492
rect 13728 25440 13780 25492
rect 13820 25440 13872 25492
rect 10876 25304 10928 25356
rect 11612 25304 11664 25356
rect 12716 25304 12768 25356
rect 9864 25236 9916 25288
rect 14096 25440 14148 25492
rect 16212 25440 16264 25492
rect 16580 25372 16632 25424
rect 21364 25440 21416 25492
rect 21916 25483 21968 25492
rect 21916 25449 21925 25483
rect 21925 25449 21959 25483
rect 21959 25449 21968 25483
rect 21916 25440 21968 25449
rect 22928 25440 22980 25492
rect 25872 25440 25924 25492
rect 23020 25372 23072 25424
rect 15292 25304 15344 25356
rect 16120 25304 16172 25356
rect 16304 25304 16356 25356
rect 14372 25279 14424 25288
rect 14372 25245 14381 25279
rect 14381 25245 14415 25279
rect 14415 25245 14424 25279
rect 14372 25236 14424 25245
rect 14648 25236 14700 25288
rect 16488 25236 16540 25288
rect 17316 25304 17368 25356
rect 19064 25304 19116 25356
rect 19984 25347 20036 25356
rect 19984 25313 19993 25347
rect 19993 25313 20027 25347
rect 20027 25313 20036 25347
rect 19984 25304 20036 25313
rect 22008 25304 22060 25356
rect 22744 25304 22796 25356
rect 24768 25372 24820 25424
rect 24032 25304 24084 25356
rect 14556 25168 14608 25220
rect 8852 25100 8904 25152
rect 13360 25100 13412 25152
rect 14740 25100 14792 25152
rect 15292 25168 15344 25220
rect 18420 25168 18472 25220
rect 23848 25236 23900 25288
rect 24768 25236 24820 25288
rect 22928 25168 22980 25220
rect 27068 25168 27120 25220
rect 16764 25100 16816 25152
rect 17868 25100 17920 25152
rect 23296 25100 23348 25152
rect 23848 25143 23900 25152
rect 23848 25109 23857 25143
rect 23857 25109 23891 25143
rect 23891 25109 23900 25143
rect 23848 25100 23900 25109
rect 24216 25100 24268 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 1584 24939 1636 24948
rect 1584 24905 1593 24939
rect 1593 24905 1627 24939
rect 1627 24905 1636 24939
rect 1584 24896 1636 24905
rect 9220 24939 9272 24948
rect 9220 24905 9229 24939
rect 9229 24905 9263 24939
rect 9263 24905 9272 24939
rect 9220 24896 9272 24905
rect 9312 24896 9364 24948
rect 14372 24896 14424 24948
rect 14648 24939 14700 24948
rect 14648 24905 14657 24939
rect 14657 24905 14691 24939
rect 14691 24905 14700 24939
rect 14648 24896 14700 24905
rect 14740 24896 14792 24948
rect 15292 24896 15344 24948
rect 9864 24828 9916 24880
rect 13452 24828 13504 24880
rect 13728 24828 13780 24880
rect 14004 24760 14056 24812
rect 14280 24760 14332 24812
rect 14832 24760 14884 24812
rect 15108 24828 15160 24880
rect 24676 24896 24728 24948
rect 25596 24939 25648 24948
rect 25596 24905 25605 24939
rect 25605 24905 25639 24939
rect 25639 24905 25648 24939
rect 25596 24896 25648 24905
rect 15476 24760 15528 24812
rect 16396 24760 16448 24812
rect 20720 24828 20772 24880
rect 23848 24828 23900 24880
rect 23388 24760 23440 24812
rect 14464 24692 14516 24744
rect 16304 24692 16356 24744
rect 16580 24692 16632 24744
rect 17592 24692 17644 24744
rect 13176 24624 13228 24676
rect 14832 24624 14884 24676
rect 16212 24624 16264 24676
rect 16672 24667 16724 24676
rect 16672 24633 16681 24667
rect 16681 24633 16715 24667
rect 16715 24633 16724 24667
rect 16672 24624 16724 24633
rect 20168 24735 20220 24744
rect 20168 24701 20177 24735
rect 20177 24701 20211 24735
rect 20211 24701 20220 24735
rect 20168 24692 20220 24701
rect 24124 24624 24176 24676
rect 2228 24556 2280 24608
rect 8852 24556 8904 24608
rect 10048 24599 10100 24608
rect 10048 24565 10057 24599
rect 10057 24565 10091 24599
rect 10091 24565 10100 24599
rect 10048 24556 10100 24565
rect 10876 24556 10928 24608
rect 11244 24556 11296 24608
rect 11428 24599 11480 24608
rect 11428 24565 11437 24599
rect 11437 24565 11471 24599
rect 11471 24565 11480 24599
rect 11428 24556 11480 24565
rect 11612 24556 11664 24608
rect 12256 24556 12308 24608
rect 12992 24599 13044 24608
rect 12992 24565 13001 24599
rect 13001 24565 13035 24599
rect 13035 24565 13044 24599
rect 12992 24556 13044 24565
rect 13360 24599 13412 24608
rect 13360 24565 13369 24599
rect 13369 24565 13403 24599
rect 13403 24565 13412 24599
rect 13360 24556 13412 24565
rect 14924 24556 14976 24608
rect 15108 24599 15160 24608
rect 15108 24565 15117 24599
rect 15117 24565 15151 24599
rect 15151 24565 15160 24599
rect 15108 24556 15160 24565
rect 16120 24599 16172 24608
rect 16120 24565 16129 24599
rect 16129 24565 16163 24599
rect 16163 24565 16172 24599
rect 16120 24556 16172 24565
rect 16304 24599 16356 24608
rect 16304 24565 16313 24599
rect 16313 24565 16347 24599
rect 16347 24565 16356 24599
rect 16304 24556 16356 24565
rect 16764 24599 16816 24608
rect 16764 24565 16773 24599
rect 16773 24565 16807 24599
rect 16807 24565 16816 24599
rect 16764 24556 16816 24565
rect 17316 24599 17368 24608
rect 17316 24565 17325 24599
rect 17325 24565 17359 24599
rect 17359 24565 17368 24599
rect 17316 24556 17368 24565
rect 17776 24599 17828 24608
rect 17776 24565 17785 24599
rect 17785 24565 17819 24599
rect 17819 24565 17828 24599
rect 17776 24556 17828 24565
rect 19064 24599 19116 24608
rect 19064 24565 19073 24599
rect 19073 24565 19107 24599
rect 19107 24565 19116 24599
rect 19064 24556 19116 24565
rect 19984 24599 20036 24608
rect 19984 24565 19993 24599
rect 19993 24565 20027 24599
rect 20027 24565 20036 24599
rect 19984 24556 20036 24565
rect 21088 24599 21140 24608
rect 21088 24565 21097 24599
rect 21097 24565 21131 24599
rect 21131 24565 21140 24599
rect 21088 24556 21140 24565
rect 21732 24556 21784 24608
rect 22008 24556 22060 24608
rect 22836 24556 22888 24608
rect 23480 24599 23532 24608
rect 23480 24565 23489 24599
rect 23489 24565 23523 24599
rect 23523 24565 23532 24599
rect 23480 24556 23532 24565
rect 23756 24556 23808 24608
rect 24860 24599 24912 24608
rect 24860 24565 24869 24599
rect 24869 24565 24903 24599
rect 24903 24565 24912 24599
rect 24860 24556 24912 24565
rect 25320 24599 25372 24608
rect 25320 24565 25329 24599
rect 25329 24565 25363 24599
rect 25363 24565 25372 24599
rect 25320 24556 25372 24565
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 1492 24352 1544 24404
rect 7932 24352 7984 24404
rect 8668 24395 8720 24404
rect 8668 24361 8677 24395
rect 8677 24361 8711 24395
rect 8711 24361 8720 24395
rect 8668 24352 8720 24361
rect 11520 24352 11572 24404
rect 13452 24395 13504 24404
rect 13452 24361 13461 24395
rect 13461 24361 13495 24395
rect 13495 24361 13504 24395
rect 13452 24352 13504 24361
rect 13820 24395 13872 24404
rect 13820 24361 13829 24395
rect 13829 24361 13863 24395
rect 13863 24361 13872 24395
rect 13820 24352 13872 24361
rect 14096 24352 14148 24404
rect 15476 24352 15528 24404
rect 15568 24352 15620 24404
rect 15844 24352 15896 24404
rect 16856 24395 16908 24404
rect 16856 24361 16865 24395
rect 16865 24361 16899 24395
rect 16899 24361 16908 24395
rect 16856 24352 16908 24361
rect 18052 24395 18104 24404
rect 18052 24361 18061 24395
rect 18061 24361 18095 24395
rect 18095 24361 18104 24395
rect 18052 24352 18104 24361
rect 18512 24352 18564 24404
rect 19156 24352 19208 24404
rect 19340 24352 19392 24404
rect 21364 24395 21416 24404
rect 15292 24284 15344 24336
rect 2044 24216 2096 24268
rect 7564 24216 7616 24268
rect 8300 24216 8352 24268
rect 10232 24259 10284 24268
rect 10232 24225 10241 24259
rect 10241 24225 10275 24259
rect 10275 24225 10284 24259
rect 10232 24216 10284 24225
rect 11612 24216 11664 24268
rect 12348 24216 12400 24268
rect 14648 24216 14700 24268
rect 17408 24284 17460 24336
rect 21364 24361 21373 24395
rect 21373 24361 21407 24395
rect 21407 24361 21416 24395
rect 21364 24352 21416 24361
rect 21180 24284 21232 24336
rect 16948 24216 17000 24268
rect 19156 24216 19208 24268
rect 23848 24216 23900 24268
rect 25044 24259 25096 24268
rect 25044 24225 25053 24259
rect 25053 24225 25087 24259
rect 25087 24225 25096 24259
rect 25044 24216 25096 24225
rect 13912 24191 13964 24200
rect 10416 24123 10468 24132
rect 10416 24089 10425 24123
rect 10425 24089 10459 24123
rect 10459 24089 10468 24123
rect 10416 24080 10468 24089
rect 11704 24080 11756 24132
rect 11796 24080 11848 24132
rect 13912 24157 13921 24191
rect 13921 24157 13955 24191
rect 13955 24157 13964 24191
rect 13912 24148 13964 24157
rect 14096 24191 14148 24200
rect 14096 24157 14105 24191
rect 14105 24157 14139 24191
rect 14139 24157 14148 24191
rect 14096 24148 14148 24157
rect 15292 24148 15344 24200
rect 16488 24148 16540 24200
rect 18604 24148 18656 24200
rect 19064 24191 19116 24200
rect 19064 24157 19073 24191
rect 19073 24157 19107 24191
rect 19107 24157 19116 24191
rect 19064 24148 19116 24157
rect 21548 24191 21600 24200
rect 21548 24157 21557 24191
rect 21557 24157 21591 24191
rect 21591 24157 21600 24191
rect 21548 24148 21600 24157
rect 23112 24148 23164 24200
rect 23480 24080 23532 24132
rect 24952 24148 25004 24200
rect 8852 24012 8904 24064
rect 10784 24055 10836 24064
rect 10784 24021 10793 24055
rect 10793 24021 10827 24055
rect 10827 24021 10836 24055
rect 10784 24012 10836 24021
rect 12808 24012 12860 24064
rect 13360 24012 13412 24064
rect 15660 24012 15712 24064
rect 15752 24012 15804 24064
rect 16028 24012 16080 24064
rect 16396 24012 16448 24064
rect 16672 24012 16724 24064
rect 16856 24012 16908 24064
rect 19616 24055 19668 24064
rect 19616 24021 19625 24055
rect 19625 24021 19659 24055
rect 19659 24021 19668 24055
rect 19616 24012 19668 24021
rect 22560 24012 22612 24064
rect 22744 24012 22796 24064
rect 23296 24012 23348 24064
rect 23572 24012 23624 24064
rect 24032 24080 24084 24132
rect 24860 24080 24912 24132
rect 25320 24148 25372 24200
rect 24124 24055 24176 24064
rect 24124 24021 24133 24055
rect 24133 24021 24167 24055
rect 24167 24021 24176 24055
rect 24124 24012 24176 24021
rect 24676 24055 24728 24064
rect 24676 24021 24685 24055
rect 24685 24021 24719 24055
rect 24719 24021 24728 24055
rect 24676 24012 24728 24021
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1676 23808 1728 23860
rect 2688 23851 2740 23860
rect 2688 23817 2697 23851
rect 2697 23817 2731 23851
rect 2731 23817 2740 23851
rect 2688 23808 2740 23817
rect 8024 23851 8076 23860
rect 8024 23817 8033 23851
rect 8033 23817 8067 23851
rect 8067 23817 8076 23851
rect 8024 23808 8076 23817
rect 9128 23851 9180 23860
rect 9128 23817 9137 23851
rect 9137 23817 9171 23851
rect 9171 23817 9180 23851
rect 9128 23808 9180 23817
rect 9496 23851 9548 23860
rect 9496 23817 9505 23851
rect 9505 23817 9539 23851
rect 9539 23817 9548 23851
rect 9496 23808 9548 23817
rect 10232 23851 10284 23860
rect 10232 23817 10241 23851
rect 10241 23817 10275 23851
rect 10275 23817 10284 23851
rect 10232 23808 10284 23817
rect 10692 23808 10744 23860
rect 13820 23808 13872 23860
rect 15476 23808 15528 23860
rect 15844 23808 15896 23860
rect 16764 23808 16816 23860
rect 20352 23851 20404 23860
rect 20352 23817 20361 23851
rect 20361 23817 20395 23851
rect 20395 23817 20404 23851
rect 20352 23808 20404 23817
rect 20720 23851 20772 23860
rect 20720 23817 20729 23851
rect 20729 23817 20763 23851
rect 20763 23817 20772 23851
rect 20720 23808 20772 23817
rect 7288 23740 7340 23792
rect 7840 23740 7892 23792
rect 1676 23604 1728 23656
rect 2320 23604 2372 23656
rect 9312 23740 9364 23792
rect 17040 23783 17092 23792
rect 11704 23672 11756 23724
rect 13728 23672 13780 23724
rect 9496 23604 9548 23656
rect 10784 23604 10836 23656
rect 13544 23604 13596 23656
rect 8300 23536 8352 23588
rect 11980 23536 12032 23588
rect 14096 23536 14148 23588
rect 2044 23511 2096 23520
rect 2044 23477 2053 23511
rect 2053 23477 2087 23511
rect 2087 23477 2096 23511
rect 2044 23468 2096 23477
rect 4436 23468 4488 23520
rect 4896 23468 4948 23520
rect 7564 23468 7616 23520
rect 8944 23468 8996 23520
rect 11612 23468 11664 23520
rect 12348 23468 12400 23520
rect 12808 23468 12860 23520
rect 15200 23672 15252 23724
rect 16488 23672 16540 23724
rect 17040 23749 17049 23783
rect 17049 23749 17083 23783
rect 17083 23749 17092 23783
rect 17040 23740 17092 23749
rect 17408 23783 17460 23792
rect 17408 23749 17417 23783
rect 17417 23749 17451 23783
rect 17451 23749 17460 23783
rect 17408 23740 17460 23749
rect 17592 23740 17644 23792
rect 18328 23740 18380 23792
rect 17960 23672 18012 23724
rect 18604 23715 18656 23724
rect 18604 23681 18613 23715
rect 18613 23681 18647 23715
rect 18647 23681 18656 23715
rect 18604 23672 18656 23681
rect 20168 23672 20220 23724
rect 21456 23808 21508 23860
rect 23204 23808 23256 23860
rect 24216 23808 24268 23860
rect 24860 23808 24912 23860
rect 25412 23851 25464 23860
rect 25412 23817 25421 23851
rect 25421 23817 25455 23851
rect 25455 23817 25464 23851
rect 25412 23808 25464 23817
rect 22928 23740 22980 23792
rect 24952 23740 25004 23792
rect 15936 23604 15988 23656
rect 16212 23604 16264 23656
rect 16396 23604 16448 23656
rect 17132 23604 17184 23656
rect 18144 23604 18196 23656
rect 18512 23647 18564 23656
rect 18512 23613 18521 23647
rect 18521 23613 18555 23647
rect 18555 23613 18564 23647
rect 18512 23604 18564 23613
rect 18788 23604 18840 23656
rect 19616 23647 19668 23656
rect 19616 23613 19625 23647
rect 19625 23613 19659 23647
rect 19659 23613 19668 23647
rect 19616 23604 19668 23613
rect 20352 23604 20404 23656
rect 16304 23536 16356 23588
rect 14648 23468 14700 23520
rect 16948 23468 17000 23520
rect 19156 23468 19208 23520
rect 20168 23468 20220 23520
rect 21364 23468 21416 23520
rect 24308 23715 24360 23724
rect 24308 23681 24317 23715
rect 24317 23681 24351 23715
rect 24351 23681 24360 23715
rect 24308 23672 24360 23681
rect 25044 23672 25096 23724
rect 25872 23672 25924 23724
rect 24124 23579 24176 23588
rect 24124 23545 24133 23579
rect 24133 23545 24167 23579
rect 24167 23545 24176 23579
rect 24124 23536 24176 23545
rect 22468 23468 22520 23520
rect 23020 23511 23072 23520
rect 23020 23477 23029 23511
rect 23029 23477 23063 23511
rect 23063 23477 23072 23511
rect 23020 23468 23072 23477
rect 23664 23511 23716 23520
rect 23664 23477 23673 23511
rect 23673 23477 23707 23511
rect 23707 23477 23716 23511
rect 23664 23468 23716 23477
rect 24308 23468 24360 23520
rect 26148 23468 26200 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 7196 23307 7248 23316
rect 7196 23273 7205 23307
rect 7205 23273 7239 23307
rect 7239 23273 7248 23307
rect 7196 23264 7248 23273
rect 11888 23264 11940 23316
rect 15108 23307 15160 23316
rect 15108 23273 15117 23307
rect 15117 23273 15151 23307
rect 15151 23273 15160 23307
rect 15108 23264 15160 23273
rect 16580 23264 16632 23316
rect 17224 23264 17276 23316
rect 18144 23307 18196 23316
rect 18144 23273 18153 23307
rect 18153 23273 18187 23307
rect 18187 23273 18196 23307
rect 18144 23264 18196 23273
rect 18420 23307 18472 23316
rect 18420 23273 18429 23307
rect 18429 23273 18463 23307
rect 18463 23273 18472 23307
rect 18420 23264 18472 23273
rect 18696 23264 18748 23316
rect 21180 23307 21232 23316
rect 21180 23273 21189 23307
rect 21189 23273 21223 23307
rect 21223 23273 21232 23307
rect 21180 23264 21232 23273
rect 25228 23307 25280 23316
rect 8208 23196 8260 23248
rect 11152 23196 11204 23248
rect 2412 23128 2464 23180
rect 7472 23128 7524 23180
rect 9312 23128 9364 23180
rect 10692 23128 10744 23180
rect 11888 23128 11940 23180
rect 13268 23128 13320 23180
rect 15016 23196 15068 23248
rect 15844 23196 15896 23248
rect 17868 23196 17920 23248
rect 25228 23273 25237 23307
rect 25237 23273 25271 23307
rect 25271 23273 25280 23307
rect 25228 23264 25280 23273
rect 17132 23128 17184 23180
rect 18696 23128 18748 23180
rect 24308 23196 24360 23248
rect 1676 23103 1728 23112
rect 1676 23069 1685 23103
rect 1685 23069 1719 23103
rect 1719 23069 1728 23103
rect 1676 23060 1728 23069
rect 2320 23103 2372 23112
rect 2320 23069 2329 23103
rect 2329 23069 2363 23103
rect 2363 23069 2372 23103
rect 2320 23060 2372 23069
rect 10600 23103 10652 23112
rect 10600 23069 10609 23103
rect 10609 23069 10643 23103
rect 10643 23069 10652 23103
rect 12072 23103 12124 23112
rect 10600 23060 10652 23069
rect 12072 23069 12081 23103
rect 12081 23069 12115 23103
rect 12115 23069 12124 23103
rect 12072 23060 12124 23069
rect 9496 22992 9548 23044
rect 11796 22992 11848 23044
rect 13452 23060 13504 23112
rect 13728 23103 13780 23112
rect 13728 23069 13737 23103
rect 13737 23069 13771 23103
rect 13771 23069 13780 23103
rect 13728 23060 13780 23069
rect 15660 23060 15712 23112
rect 15936 23103 15988 23112
rect 15936 23069 15945 23103
rect 15945 23069 15979 23103
rect 15979 23069 15988 23103
rect 15936 23060 15988 23069
rect 17408 23103 17460 23112
rect 13360 22992 13412 23044
rect 13544 22992 13596 23044
rect 14004 22992 14056 23044
rect 17408 23069 17417 23103
rect 17417 23069 17451 23103
rect 17451 23069 17460 23103
rect 17408 23060 17460 23069
rect 18880 23103 18932 23112
rect 18880 23069 18889 23103
rect 18889 23069 18923 23103
rect 18923 23069 18932 23103
rect 18880 23060 18932 23069
rect 20076 23128 20128 23180
rect 21180 23128 21232 23180
rect 23848 23171 23900 23180
rect 23848 23137 23857 23171
rect 23857 23137 23891 23171
rect 23891 23137 23900 23171
rect 23848 23128 23900 23137
rect 25044 23171 25096 23180
rect 25044 23137 25053 23171
rect 25053 23137 25087 23171
rect 25087 23137 25096 23171
rect 25044 23128 25096 23137
rect 21548 23060 21600 23112
rect 22468 23103 22520 23112
rect 22468 23069 22477 23103
rect 22477 23069 22511 23103
rect 22511 23069 22520 23103
rect 23940 23103 23992 23112
rect 22468 23060 22520 23069
rect 23940 23069 23949 23103
rect 23949 23069 23983 23103
rect 23983 23069 23992 23103
rect 23940 23060 23992 23069
rect 24124 23103 24176 23112
rect 24124 23069 24133 23103
rect 24133 23069 24167 23103
rect 24167 23069 24176 23103
rect 24124 23060 24176 23069
rect 24768 22992 24820 23044
rect 7012 22924 7064 22976
rect 8944 22924 8996 22976
rect 10968 22924 11020 22976
rect 12900 22924 12952 22976
rect 13912 22924 13964 22976
rect 16212 22924 16264 22976
rect 17592 22924 17644 22976
rect 20352 22967 20404 22976
rect 20352 22933 20361 22967
rect 20361 22933 20395 22967
rect 20395 22933 20404 22967
rect 20352 22924 20404 22933
rect 20720 22967 20772 22976
rect 20720 22933 20729 22967
rect 20729 22933 20763 22967
rect 20763 22933 20772 22967
rect 20720 22924 20772 22933
rect 21456 22967 21508 22976
rect 21456 22933 21465 22967
rect 21465 22933 21499 22967
rect 21499 22933 21508 22967
rect 21456 22924 21508 22933
rect 21916 22967 21968 22976
rect 21916 22933 21925 22967
rect 21925 22933 21959 22967
rect 21959 22933 21968 22967
rect 21916 22924 21968 22933
rect 23388 22924 23440 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 1584 22763 1636 22772
rect 1584 22729 1593 22763
rect 1593 22729 1627 22763
rect 1627 22729 1636 22763
rect 1584 22720 1636 22729
rect 4068 22720 4120 22772
rect 9036 22763 9088 22772
rect 9036 22729 9045 22763
rect 9045 22729 9079 22763
rect 9079 22729 9088 22763
rect 9036 22720 9088 22729
rect 10048 22720 10100 22772
rect 10600 22720 10652 22772
rect 11612 22720 11664 22772
rect 12072 22720 12124 22772
rect 13268 22763 13320 22772
rect 13268 22729 13277 22763
rect 13277 22729 13311 22763
rect 13311 22729 13320 22763
rect 13268 22720 13320 22729
rect 15660 22720 15712 22772
rect 17224 22720 17276 22772
rect 17684 22720 17736 22772
rect 19616 22763 19668 22772
rect 19616 22729 19625 22763
rect 19625 22729 19659 22763
rect 19659 22729 19668 22763
rect 19616 22720 19668 22729
rect 21824 22763 21876 22772
rect 21824 22729 21833 22763
rect 21833 22729 21867 22763
rect 21867 22729 21876 22763
rect 21824 22720 21876 22729
rect 25044 22763 25096 22772
rect 25044 22729 25053 22763
rect 25053 22729 25087 22763
rect 25087 22729 25096 22763
rect 25044 22720 25096 22729
rect 25596 22763 25648 22772
rect 25596 22729 25605 22763
rect 25605 22729 25639 22763
rect 25639 22729 25648 22763
rect 25596 22720 25648 22729
rect 9404 22652 9456 22704
rect 6644 22584 6696 22636
rect 8116 22584 8168 22636
rect 9496 22627 9548 22636
rect 9496 22593 9505 22627
rect 9505 22593 9539 22627
rect 9539 22593 9548 22627
rect 9496 22584 9548 22593
rect 18144 22652 18196 22704
rect 5356 22516 5408 22568
rect 7104 22559 7156 22568
rect 7104 22525 7113 22559
rect 7113 22525 7147 22559
rect 7147 22525 7156 22559
rect 7656 22559 7708 22568
rect 7104 22516 7156 22525
rect 7656 22525 7665 22559
rect 7665 22525 7699 22559
rect 7699 22525 7708 22559
rect 7656 22516 7708 22525
rect 9036 22516 9088 22568
rect 4804 22448 4856 22500
rect 7012 22448 7064 22500
rect 7288 22448 7340 22500
rect 2136 22380 2188 22432
rect 2412 22423 2464 22432
rect 2412 22389 2421 22423
rect 2421 22389 2455 22423
rect 2455 22389 2464 22423
rect 2412 22380 2464 22389
rect 6644 22423 6696 22432
rect 6644 22389 6653 22423
rect 6653 22389 6687 22423
rect 6687 22389 6696 22423
rect 6644 22380 6696 22389
rect 7196 22423 7248 22432
rect 7196 22389 7205 22423
rect 7205 22389 7239 22423
rect 7239 22389 7248 22423
rect 7196 22380 7248 22389
rect 8208 22423 8260 22432
rect 8208 22389 8217 22423
rect 8217 22389 8251 22423
rect 8251 22389 8260 22423
rect 8208 22380 8260 22389
rect 9956 22380 10008 22432
rect 12900 22584 12952 22636
rect 10968 22516 11020 22568
rect 12440 22516 12492 22568
rect 13820 22516 13872 22568
rect 14372 22584 14424 22636
rect 14556 22516 14608 22568
rect 13728 22448 13780 22500
rect 15936 22584 15988 22636
rect 17224 22584 17276 22636
rect 18236 22584 18288 22636
rect 18328 22584 18380 22636
rect 23848 22695 23900 22704
rect 23848 22661 23857 22695
rect 23857 22661 23891 22695
rect 23891 22661 23900 22695
rect 23848 22652 23900 22661
rect 24768 22652 24820 22704
rect 20076 22584 20128 22636
rect 23204 22584 23256 22636
rect 24124 22584 24176 22636
rect 24492 22627 24544 22636
rect 24492 22593 24501 22627
rect 24501 22593 24535 22627
rect 24535 22593 24544 22627
rect 24492 22584 24544 22593
rect 18144 22516 18196 22568
rect 18696 22516 18748 22568
rect 25412 22559 25464 22568
rect 25412 22525 25421 22559
rect 25421 22525 25455 22559
rect 25455 22525 25464 22559
rect 25412 22516 25464 22525
rect 10692 22380 10744 22432
rect 11060 22380 11112 22432
rect 11888 22380 11940 22432
rect 14740 22423 14792 22432
rect 14740 22389 14749 22423
rect 14749 22389 14783 22423
rect 14783 22389 14792 22423
rect 14740 22380 14792 22389
rect 15108 22423 15160 22432
rect 15108 22389 15117 22423
rect 15117 22389 15151 22423
rect 15151 22389 15160 22423
rect 15108 22380 15160 22389
rect 15844 22423 15896 22432
rect 15844 22389 15853 22423
rect 15853 22389 15887 22423
rect 15887 22389 15896 22423
rect 15844 22380 15896 22389
rect 16580 22448 16632 22500
rect 16396 22423 16448 22432
rect 16396 22389 16405 22423
rect 16405 22389 16439 22423
rect 16439 22389 16448 22423
rect 16396 22380 16448 22389
rect 17132 22423 17184 22432
rect 17132 22389 17141 22423
rect 17141 22389 17175 22423
rect 17175 22389 17184 22423
rect 17132 22380 17184 22389
rect 17500 22380 17552 22432
rect 20352 22448 20404 22500
rect 24400 22448 24452 22500
rect 18328 22380 18380 22432
rect 19432 22423 19484 22432
rect 19432 22389 19441 22423
rect 19441 22389 19475 22423
rect 19475 22389 19484 22423
rect 19432 22380 19484 22389
rect 20076 22423 20128 22432
rect 20076 22389 20085 22423
rect 20085 22389 20119 22423
rect 20119 22389 20128 22423
rect 20076 22380 20128 22389
rect 21180 22380 21232 22432
rect 21548 22380 21600 22432
rect 22284 22423 22336 22432
rect 22284 22389 22293 22423
rect 22293 22389 22327 22423
rect 22327 22389 22336 22423
rect 22284 22380 22336 22389
rect 23480 22423 23532 22432
rect 23480 22389 23489 22423
rect 23489 22389 23523 22423
rect 23523 22389 23532 22423
rect 23480 22380 23532 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 4804 22219 4856 22228
rect 4804 22185 4813 22219
rect 4813 22185 4847 22219
rect 4847 22185 4856 22219
rect 4804 22176 4856 22185
rect 13452 22219 13504 22228
rect 13452 22185 13461 22219
rect 13461 22185 13495 22219
rect 13495 22185 13504 22219
rect 13452 22176 13504 22185
rect 13912 22176 13964 22228
rect 16396 22176 16448 22228
rect 5356 22151 5408 22160
rect 5356 22117 5365 22151
rect 5365 22117 5399 22151
rect 5399 22117 5408 22151
rect 5356 22108 5408 22117
rect 2320 22040 2372 22092
rect 4988 22040 5040 22092
rect 7380 22083 7432 22092
rect 7380 22049 7414 22083
rect 7414 22049 7432 22083
rect 9404 22108 9456 22160
rect 7380 22040 7432 22049
rect 10692 22108 10744 22160
rect 11520 22108 11572 22160
rect 9956 22083 10008 22092
rect 9956 22049 9990 22083
rect 9990 22049 10008 22083
rect 9956 22040 10008 22049
rect 11796 22040 11848 22092
rect 14004 22108 14056 22160
rect 15844 22108 15896 22160
rect 16028 22108 16080 22160
rect 16120 22108 16172 22160
rect 20260 22176 20312 22228
rect 20720 22176 20772 22228
rect 22284 22176 22336 22228
rect 23940 22176 23992 22228
rect 14832 22040 14884 22092
rect 7104 22015 7156 22024
rect 7104 21981 7113 22015
rect 7113 21981 7147 22015
rect 7147 21981 7156 22015
rect 7104 21972 7156 21981
rect 8944 21972 8996 22024
rect 12348 22015 12400 22024
rect 12348 21981 12357 22015
rect 12357 21981 12391 22015
rect 12391 21981 12400 22015
rect 12348 21972 12400 21981
rect 12716 21972 12768 22024
rect 12808 21972 12860 22024
rect 13912 22015 13964 22024
rect 13912 21981 13921 22015
rect 13921 21981 13955 22015
rect 13955 21981 13964 22015
rect 13912 21972 13964 21981
rect 14556 21972 14608 22024
rect 15844 21972 15896 22024
rect 16764 22040 16816 22092
rect 16856 22040 16908 22092
rect 17684 22040 17736 22092
rect 1400 21904 1452 21956
rect 8116 21904 8168 21956
rect 11152 21904 11204 21956
rect 12072 21904 12124 21956
rect 14648 21904 14700 21956
rect 17684 21904 17736 21956
rect 17868 22108 17920 22160
rect 18420 22108 18472 22160
rect 18604 22151 18656 22160
rect 18604 22117 18613 22151
rect 18613 22117 18647 22151
rect 18647 22117 18656 22151
rect 18604 22108 18656 22117
rect 21548 22108 21600 22160
rect 21732 22108 21784 22160
rect 21824 22108 21876 22160
rect 22100 22108 22152 22160
rect 17868 21972 17920 22024
rect 18696 22015 18748 22024
rect 18696 21981 18705 22015
rect 18705 21981 18739 22015
rect 18739 21981 18748 22015
rect 18696 21972 18748 21981
rect 19524 22040 19576 22092
rect 20628 22040 20680 22092
rect 22008 22083 22060 22092
rect 22008 22049 22017 22083
rect 22017 22049 22051 22083
rect 22051 22049 22060 22083
rect 22008 22040 22060 22049
rect 24124 22108 24176 22160
rect 23204 22040 23256 22092
rect 23940 22040 23992 22092
rect 20076 21972 20128 22024
rect 20444 21972 20496 22024
rect 20996 21972 21048 22024
rect 22284 22015 22336 22024
rect 22284 21981 22293 22015
rect 22293 21981 22327 22015
rect 22327 21981 22336 22015
rect 22284 21972 22336 21981
rect 23480 21972 23532 22024
rect 18236 21947 18288 21956
rect 18236 21913 18245 21947
rect 18245 21913 18279 21947
rect 18279 21913 18288 21947
rect 18236 21904 18288 21913
rect 18972 21904 19024 21956
rect 21088 21904 21140 21956
rect 23204 21904 23256 21956
rect 24400 22015 24452 22024
rect 24400 21981 24409 22015
rect 24409 21981 24443 22015
rect 24443 21981 24452 22015
rect 24860 22040 24912 22092
rect 24400 21972 24452 21981
rect 6276 21836 6328 21888
rect 6552 21879 6604 21888
rect 6552 21845 6561 21879
rect 6561 21845 6595 21879
rect 6595 21845 6604 21879
rect 6552 21836 6604 21845
rect 6920 21879 6972 21888
rect 6920 21845 6929 21879
rect 6929 21845 6963 21879
rect 6963 21845 6972 21879
rect 6920 21836 6972 21845
rect 9036 21879 9088 21888
rect 9036 21845 9045 21879
rect 9045 21845 9079 21879
rect 9079 21845 9088 21879
rect 9036 21836 9088 21845
rect 9128 21836 9180 21888
rect 9588 21836 9640 21888
rect 10048 21836 10100 21888
rect 13268 21879 13320 21888
rect 13268 21845 13277 21879
rect 13277 21845 13311 21879
rect 13311 21845 13320 21879
rect 13268 21836 13320 21845
rect 15936 21879 15988 21888
rect 15936 21845 15945 21879
rect 15945 21845 15979 21879
rect 15979 21845 15988 21879
rect 15936 21836 15988 21845
rect 18052 21836 18104 21888
rect 18420 21836 18472 21888
rect 18880 21836 18932 21888
rect 19248 21879 19300 21888
rect 19248 21845 19257 21879
rect 19257 21845 19291 21879
rect 19291 21845 19300 21879
rect 19248 21836 19300 21845
rect 20904 21836 20956 21888
rect 22468 21836 22520 21888
rect 24216 21836 24268 21888
rect 24676 21836 24728 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1492 21632 1544 21684
rect 3516 21632 3568 21684
rect 4804 21632 4856 21684
rect 4896 21632 4948 21684
rect 6644 21675 6696 21684
rect 6644 21641 6653 21675
rect 6653 21641 6687 21675
rect 6687 21641 6696 21675
rect 6644 21632 6696 21641
rect 7380 21632 7432 21684
rect 10692 21632 10744 21684
rect 12808 21632 12860 21684
rect 14096 21632 14148 21684
rect 3792 21564 3844 21616
rect 5540 21564 5592 21616
rect 2044 21539 2096 21548
rect 2044 21505 2053 21539
rect 2053 21505 2087 21539
rect 2087 21505 2096 21539
rect 2044 21496 2096 21505
rect 5816 21539 5868 21548
rect 5816 21505 5825 21539
rect 5825 21505 5859 21539
rect 5859 21505 5868 21539
rect 5816 21496 5868 21505
rect 3056 21471 3108 21480
rect 3056 21437 3065 21471
rect 3065 21437 3099 21471
rect 3099 21437 3108 21471
rect 3056 21428 3108 21437
rect 4988 21428 5040 21480
rect 4896 21360 4948 21412
rect 6828 21360 6880 21412
rect 2320 21335 2372 21344
rect 2320 21301 2329 21335
rect 2329 21301 2363 21335
rect 2363 21301 2372 21335
rect 2320 21292 2372 21301
rect 2780 21292 2832 21344
rect 5172 21335 5224 21344
rect 5172 21301 5181 21335
rect 5181 21301 5215 21335
rect 5215 21301 5224 21335
rect 5172 21292 5224 21301
rect 5540 21335 5592 21344
rect 5540 21301 5549 21335
rect 5549 21301 5583 21335
rect 5583 21301 5592 21335
rect 5540 21292 5592 21301
rect 7104 21428 7156 21480
rect 8944 21496 8996 21548
rect 12348 21496 12400 21548
rect 18604 21632 18656 21684
rect 20076 21632 20128 21684
rect 16764 21564 16816 21616
rect 17132 21564 17184 21616
rect 18696 21564 18748 21616
rect 8208 21428 8260 21480
rect 10692 21428 10744 21480
rect 12992 21428 13044 21480
rect 14832 21428 14884 21480
rect 18880 21496 18932 21548
rect 19064 21428 19116 21480
rect 20352 21632 20404 21684
rect 21640 21632 21692 21684
rect 22008 21675 22060 21684
rect 22008 21641 22017 21675
rect 22017 21641 22051 21675
rect 22051 21641 22060 21675
rect 22008 21632 22060 21641
rect 22100 21632 22152 21684
rect 23204 21632 23256 21684
rect 23756 21632 23808 21684
rect 24676 21632 24728 21684
rect 25688 21632 25740 21684
rect 20904 21539 20956 21548
rect 20904 21505 20913 21539
rect 20913 21505 20947 21539
rect 20947 21505 20956 21539
rect 20904 21496 20956 21505
rect 22284 21564 22336 21616
rect 22376 21496 22428 21548
rect 23388 21496 23440 21548
rect 25044 21496 25096 21548
rect 22008 21428 22060 21480
rect 22100 21428 22152 21480
rect 24216 21471 24268 21480
rect 24216 21437 24225 21471
rect 24225 21437 24259 21471
rect 24259 21437 24268 21471
rect 24216 21428 24268 21437
rect 25228 21428 25280 21480
rect 9496 21360 9548 21412
rect 10048 21360 10100 21412
rect 13728 21360 13780 21412
rect 13912 21360 13964 21412
rect 16764 21360 16816 21412
rect 17500 21360 17552 21412
rect 7656 21292 7708 21344
rect 8852 21335 8904 21344
rect 8852 21301 8861 21335
rect 8861 21301 8895 21335
rect 8895 21301 8904 21335
rect 8852 21292 8904 21301
rect 9404 21292 9456 21344
rect 9956 21292 10008 21344
rect 11060 21335 11112 21344
rect 11060 21301 11069 21335
rect 11069 21301 11103 21335
rect 11103 21301 11112 21335
rect 11060 21292 11112 21301
rect 11244 21292 11296 21344
rect 13268 21335 13320 21344
rect 13268 21301 13277 21335
rect 13277 21301 13311 21335
rect 13311 21301 13320 21335
rect 13268 21292 13320 21301
rect 14280 21292 14332 21344
rect 14556 21292 14608 21344
rect 16672 21292 16724 21344
rect 17132 21292 17184 21344
rect 17868 21292 17920 21344
rect 18052 21335 18104 21344
rect 18052 21301 18061 21335
rect 18061 21301 18095 21335
rect 18095 21301 18104 21335
rect 18052 21292 18104 21301
rect 18420 21335 18472 21344
rect 18420 21301 18429 21335
rect 18429 21301 18463 21335
rect 18463 21301 18472 21335
rect 18420 21292 18472 21301
rect 22744 21292 22796 21344
rect 23480 21335 23532 21344
rect 23480 21301 23489 21335
rect 23489 21301 23523 21335
rect 23523 21301 23532 21335
rect 23480 21292 23532 21301
rect 23940 21292 23992 21344
rect 25044 21292 25096 21344
rect 25688 21292 25740 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1584 21131 1636 21140
rect 1584 21097 1593 21131
rect 1593 21097 1627 21131
rect 1627 21097 1636 21131
rect 1584 21088 1636 21097
rect 2596 21088 2648 21140
rect 3516 21131 3568 21140
rect 3516 21097 3525 21131
rect 3525 21097 3559 21131
rect 3559 21097 3568 21131
rect 3516 21088 3568 21097
rect 4896 21131 4948 21140
rect 4896 21097 4905 21131
rect 4905 21097 4939 21131
rect 4939 21097 4948 21131
rect 4896 21088 4948 21097
rect 5540 21088 5592 21140
rect 5448 21020 5500 21072
rect 6552 21088 6604 21140
rect 9036 21088 9088 21140
rect 9680 21088 9732 21140
rect 10140 21088 10192 21140
rect 11152 21088 11204 21140
rect 16396 21131 16448 21140
rect 16396 21097 16405 21131
rect 16405 21097 16439 21131
rect 16439 21097 16448 21131
rect 16396 21088 16448 21097
rect 17776 21088 17828 21140
rect 18144 21131 18196 21140
rect 18144 21097 18153 21131
rect 18153 21097 18187 21131
rect 18187 21097 18196 21131
rect 18144 21088 18196 21097
rect 19524 21131 19576 21140
rect 19524 21097 19533 21131
rect 19533 21097 19567 21131
rect 19567 21097 19576 21131
rect 19524 21088 19576 21097
rect 20996 21131 21048 21140
rect 20996 21097 21005 21131
rect 21005 21097 21039 21131
rect 21039 21097 21048 21131
rect 20996 21088 21048 21097
rect 23388 21131 23440 21140
rect 23388 21097 23397 21131
rect 23397 21097 23431 21131
rect 23431 21097 23440 21131
rect 23388 21088 23440 21097
rect 24860 21088 24912 21140
rect 8668 21020 8720 21072
rect 10600 21020 10652 21072
rect 11244 21020 11296 21072
rect 12716 21020 12768 21072
rect 14096 21063 14148 21072
rect 14096 21029 14105 21063
rect 14105 21029 14139 21063
rect 14139 21029 14148 21063
rect 14096 21020 14148 21029
rect 14280 21020 14332 21072
rect 2044 20952 2096 21004
rect 3148 20952 3200 21004
rect 5540 20952 5592 21004
rect 8024 20952 8076 21004
rect 4988 20884 5040 20936
rect 5080 20884 5132 20936
rect 5816 20884 5868 20936
rect 6000 20884 6052 20936
rect 9588 20952 9640 21004
rect 9864 20952 9916 21004
rect 10692 20952 10744 21004
rect 13820 20952 13872 21004
rect 15292 20995 15344 21004
rect 15292 20961 15301 20995
rect 15301 20961 15335 20995
rect 15335 20961 15344 20995
rect 15292 20952 15344 20961
rect 15476 21020 15528 21072
rect 22284 21020 22336 21072
rect 23664 21020 23716 21072
rect 16580 20952 16632 21004
rect 18696 20952 18748 21004
rect 19248 20952 19300 21004
rect 19708 20995 19760 21004
rect 19708 20961 19717 20995
rect 19717 20961 19751 20995
rect 19751 20961 19760 20995
rect 19708 20952 19760 20961
rect 20720 20952 20772 21004
rect 23756 20995 23808 21004
rect 23756 20961 23765 20995
rect 23765 20961 23799 20995
rect 23799 20961 23808 20995
rect 23756 20952 23808 20961
rect 24032 20952 24084 21004
rect 24952 20995 25004 21004
rect 24952 20961 24961 20995
rect 24961 20961 24995 20995
rect 24995 20961 25004 20995
rect 24952 20952 25004 20961
rect 25136 20952 25188 21004
rect 5540 20816 5592 20868
rect 8300 20816 8352 20868
rect 9496 20884 9548 20936
rect 15936 20884 15988 20936
rect 17040 20927 17092 20936
rect 17040 20893 17049 20927
rect 17049 20893 17083 20927
rect 17083 20893 17092 20927
rect 17040 20884 17092 20893
rect 17408 20884 17460 20936
rect 18144 20884 18196 20936
rect 8852 20816 8904 20868
rect 9956 20816 10008 20868
rect 13728 20816 13780 20868
rect 14832 20816 14884 20868
rect 18880 20884 18932 20936
rect 20996 20884 21048 20936
rect 22376 20884 22428 20936
rect 23664 20884 23716 20936
rect 24860 20884 24912 20936
rect 19892 20859 19944 20868
rect 19892 20825 19901 20859
rect 19901 20825 19935 20859
rect 19935 20825 19944 20859
rect 19892 20816 19944 20825
rect 22744 20816 22796 20868
rect 24124 20816 24176 20868
rect 5172 20748 5224 20800
rect 6184 20748 6236 20800
rect 9496 20748 9548 20800
rect 10324 20791 10376 20800
rect 10324 20757 10333 20791
rect 10333 20757 10367 20791
rect 10367 20757 10376 20791
rect 10324 20748 10376 20757
rect 10692 20748 10744 20800
rect 15384 20748 15436 20800
rect 17316 20748 17368 20800
rect 19064 20748 19116 20800
rect 22284 20748 22336 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 2688 20587 2740 20596
rect 2688 20553 2697 20587
rect 2697 20553 2731 20587
rect 2731 20553 2740 20587
rect 2688 20544 2740 20553
rect 5264 20544 5316 20596
rect 6552 20544 6604 20596
rect 8300 20544 8352 20596
rect 9312 20544 9364 20596
rect 9680 20544 9732 20596
rect 13820 20544 13872 20596
rect 14188 20587 14240 20596
rect 14188 20553 14197 20587
rect 14197 20553 14231 20587
rect 14231 20553 14240 20587
rect 14188 20544 14240 20553
rect 14372 20587 14424 20596
rect 14372 20553 14381 20587
rect 14381 20553 14415 20587
rect 14415 20553 14424 20587
rect 14372 20544 14424 20553
rect 15384 20544 15436 20596
rect 16488 20544 16540 20596
rect 20996 20587 21048 20596
rect 20996 20553 21005 20587
rect 21005 20553 21039 20587
rect 21039 20553 21048 20587
rect 20996 20544 21048 20553
rect 21824 20544 21876 20596
rect 24952 20587 25004 20596
rect 24952 20553 24961 20587
rect 24961 20553 24995 20587
rect 24995 20553 25004 20587
rect 24952 20544 25004 20553
rect 25412 20587 25464 20596
rect 25412 20553 25421 20587
rect 25421 20553 25455 20587
rect 25455 20553 25464 20587
rect 25412 20544 25464 20553
rect 2044 20519 2096 20528
rect 2044 20485 2053 20519
rect 2053 20485 2087 20519
rect 2087 20485 2096 20519
rect 2044 20476 2096 20485
rect 3884 20476 3936 20528
rect 8392 20476 8444 20528
rect 5540 20408 5592 20460
rect 5724 20451 5776 20460
rect 5724 20417 5733 20451
rect 5733 20417 5767 20451
rect 5767 20417 5776 20451
rect 5724 20408 5776 20417
rect 6920 20408 6972 20460
rect 2504 20383 2556 20392
rect 2504 20349 2513 20383
rect 2513 20349 2547 20383
rect 2547 20349 2556 20383
rect 2504 20340 2556 20349
rect 3608 20383 3660 20392
rect 3608 20349 3617 20383
rect 3617 20349 3651 20383
rect 3651 20349 3660 20383
rect 3608 20340 3660 20349
rect 6644 20383 6696 20392
rect 6644 20349 6653 20383
rect 6653 20349 6687 20383
rect 6687 20349 6696 20383
rect 8668 20408 8720 20460
rect 9404 20408 9456 20460
rect 10692 20451 10744 20460
rect 10692 20417 10701 20451
rect 10701 20417 10735 20451
rect 10735 20417 10744 20451
rect 10692 20408 10744 20417
rect 12716 20408 12768 20460
rect 15936 20476 15988 20528
rect 17868 20476 17920 20528
rect 18144 20476 18196 20528
rect 14924 20451 14976 20460
rect 14924 20417 14933 20451
rect 14933 20417 14967 20451
rect 14967 20417 14976 20451
rect 14924 20408 14976 20417
rect 15844 20408 15896 20460
rect 17316 20408 17368 20460
rect 20076 20408 20128 20460
rect 6644 20340 6696 20349
rect 10324 20340 10376 20392
rect 10784 20340 10836 20392
rect 15936 20340 15988 20392
rect 16396 20340 16448 20392
rect 18420 20383 18472 20392
rect 18420 20349 18429 20383
rect 18429 20349 18463 20383
rect 18463 20349 18472 20383
rect 18420 20340 18472 20349
rect 18512 20383 18564 20392
rect 18512 20349 18521 20383
rect 18521 20349 18555 20383
rect 18555 20349 18564 20383
rect 18512 20340 18564 20349
rect 19432 20340 19484 20392
rect 3148 20315 3200 20324
rect 3148 20281 3157 20315
rect 3157 20281 3191 20315
rect 3191 20281 3200 20315
rect 3148 20272 3200 20281
rect 5080 20272 5132 20324
rect 5540 20315 5592 20324
rect 5540 20281 5549 20315
rect 5549 20281 5583 20315
rect 5583 20281 5592 20315
rect 5540 20272 5592 20281
rect 8944 20315 8996 20324
rect 8944 20281 8953 20315
rect 8953 20281 8987 20315
rect 8987 20281 8996 20315
rect 8944 20272 8996 20281
rect 13176 20272 13228 20324
rect 1400 20204 1452 20256
rect 2412 20247 2464 20256
rect 2412 20213 2421 20247
rect 2421 20213 2455 20247
rect 2455 20213 2464 20247
rect 2412 20204 2464 20213
rect 3792 20247 3844 20256
rect 3792 20213 3801 20247
rect 3801 20213 3835 20247
rect 3835 20213 3844 20247
rect 3792 20204 3844 20213
rect 4988 20247 5040 20256
rect 4988 20213 4997 20247
rect 4997 20213 5031 20247
rect 5031 20213 5040 20247
rect 4988 20204 5040 20213
rect 5264 20204 5316 20256
rect 6000 20204 6052 20256
rect 7196 20247 7248 20256
rect 7196 20213 7205 20247
rect 7205 20213 7239 20247
rect 7239 20213 7248 20247
rect 7196 20204 7248 20213
rect 9128 20204 9180 20256
rect 9588 20204 9640 20256
rect 11244 20247 11296 20256
rect 11244 20213 11253 20247
rect 11253 20213 11287 20247
rect 11287 20213 11296 20247
rect 11244 20204 11296 20213
rect 12440 20247 12492 20256
rect 12440 20213 12449 20247
rect 12449 20213 12483 20247
rect 12483 20213 12492 20247
rect 12808 20247 12860 20256
rect 12440 20204 12492 20213
rect 12808 20213 12817 20247
rect 12817 20213 12851 20247
rect 12851 20213 12860 20247
rect 12808 20204 12860 20213
rect 14648 20204 14700 20256
rect 15936 20247 15988 20256
rect 15936 20213 15945 20247
rect 15945 20213 15979 20247
rect 15979 20213 15988 20247
rect 15936 20204 15988 20213
rect 16764 20247 16816 20256
rect 16764 20213 16773 20247
rect 16773 20213 16807 20247
rect 16807 20213 16816 20247
rect 16764 20204 16816 20213
rect 17408 20247 17460 20256
rect 17408 20213 17417 20247
rect 17417 20213 17451 20247
rect 17451 20213 17460 20247
rect 17408 20204 17460 20213
rect 17868 20247 17920 20256
rect 17868 20213 17877 20247
rect 17877 20213 17911 20247
rect 17911 20213 17920 20247
rect 17868 20204 17920 20213
rect 19248 20204 19300 20256
rect 19708 20272 19760 20324
rect 19524 20204 19576 20256
rect 20720 20451 20772 20460
rect 20720 20417 20729 20451
rect 20729 20417 20763 20451
rect 20763 20417 20772 20451
rect 20720 20408 20772 20417
rect 21640 20408 21692 20460
rect 22376 20408 22428 20460
rect 23204 20408 23256 20460
rect 24216 20476 24268 20528
rect 24584 20476 24636 20528
rect 24860 20476 24912 20528
rect 24124 20451 24176 20460
rect 24124 20417 24133 20451
rect 24133 20417 24167 20451
rect 24167 20417 24176 20451
rect 24124 20408 24176 20417
rect 24768 20408 24820 20460
rect 23664 20340 23716 20392
rect 21364 20272 21416 20324
rect 22284 20272 22336 20324
rect 22376 20272 22428 20324
rect 22836 20272 22888 20324
rect 24952 20340 25004 20392
rect 20812 20204 20864 20256
rect 21180 20247 21232 20256
rect 21180 20213 21189 20247
rect 21189 20213 21223 20247
rect 21223 20213 21232 20247
rect 21180 20204 21232 20213
rect 21640 20247 21692 20256
rect 21640 20213 21649 20247
rect 21649 20213 21683 20247
rect 21683 20213 21692 20247
rect 21640 20204 21692 20213
rect 23112 20204 23164 20256
rect 23480 20247 23532 20256
rect 23480 20213 23489 20247
rect 23489 20213 23523 20247
rect 23523 20213 23532 20247
rect 23480 20204 23532 20213
rect 23756 20204 23808 20256
rect 24216 20204 24268 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 4252 20043 4304 20052
rect 4252 20009 4261 20043
rect 4261 20009 4295 20043
rect 4295 20009 4304 20043
rect 4252 20000 4304 20009
rect 4712 20043 4764 20052
rect 4712 20009 4721 20043
rect 4721 20009 4755 20043
rect 4755 20009 4764 20043
rect 4712 20000 4764 20009
rect 6092 20000 6144 20052
rect 7656 20000 7708 20052
rect 8024 20043 8076 20052
rect 8024 20009 8033 20043
rect 8033 20009 8067 20043
rect 8067 20009 8076 20043
rect 8024 20000 8076 20009
rect 9864 20043 9916 20052
rect 9864 20009 9873 20043
rect 9873 20009 9907 20043
rect 9907 20009 9916 20043
rect 9864 20000 9916 20009
rect 11060 20043 11112 20052
rect 11060 20009 11069 20043
rect 11069 20009 11103 20043
rect 11103 20009 11112 20043
rect 11060 20000 11112 20009
rect 11520 20043 11572 20052
rect 11520 20009 11529 20043
rect 11529 20009 11563 20043
rect 11563 20009 11572 20043
rect 11520 20000 11572 20009
rect 12808 20000 12860 20052
rect 13728 20000 13780 20052
rect 15108 20043 15160 20052
rect 15108 20009 15117 20043
rect 15117 20009 15151 20043
rect 15151 20009 15160 20043
rect 15108 20000 15160 20009
rect 16580 20000 16632 20052
rect 18236 20000 18288 20052
rect 18972 20043 19024 20052
rect 18972 20009 18981 20043
rect 18981 20009 19015 20043
rect 19015 20009 19024 20043
rect 18972 20000 19024 20009
rect 20076 20043 20128 20052
rect 20076 20009 20085 20043
rect 20085 20009 20119 20043
rect 20119 20009 20128 20043
rect 20076 20000 20128 20009
rect 22100 20000 22152 20052
rect 24032 20043 24084 20052
rect 24032 20009 24041 20043
rect 24041 20009 24075 20043
rect 24075 20009 24084 20043
rect 24032 20000 24084 20009
rect 24216 20000 24268 20052
rect 2504 19932 2556 19984
rect 2596 19932 2648 19984
rect 4804 19932 4856 19984
rect 2320 19660 2372 19712
rect 2872 19703 2924 19712
rect 2872 19669 2881 19703
rect 2881 19669 2915 19703
rect 2915 19669 2924 19703
rect 2872 19660 2924 19669
rect 4988 19864 5040 19916
rect 5724 19864 5776 19916
rect 6828 19932 6880 19984
rect 7196 19932 7248 19984
rect 11152 19932 11204 19984
rect 12348 19932 12400 19984
rect 12992 19932 13044 19984
rect 14648 19975 14700 19984
rect 6092 19907 6144 19916
rect 6092 19873 6126 19907
rect 6126 19873 6144 19907
rect 6092 19864 6144 19873
rect 6644 19864 6696 19916
rect 8392 19907 8444 19916
rect 8392 19873 8401 19907
rect 8401 19873 8435 19907
rect 8435 19873 8444 19907
rect 8392 19864 8444 19873
rect 4804 19796 4856 19848
rect 5080 19796 5132 19848
rect 8024 19796 8076 19848
rect 8668 19839 8720 19848
rect 8668 19805 8677 19839
rect 8677 19805 8711 19839
rect 8711 19805 8720 19839
rect 8668 19796 8720 19805
rect 9864 19796 9916 19848
rect 11704 19864 11756 19916
rect 12716 19864 12768 19916
rect 13268 19907 13320 19916
rect 13268 19873 13302 19907
rect 13302 19873 13320 19907
rect 13268 19864 13320 19873
rect 13728 19864 13780 19916
rect 14648 19941 14657 19975
rect 14657 19941 14691 19975
rect 14691 19941 14700 19975
rect 14648 19932 14700 19941
rect 16764 19932 16816 19984
rect 15384 19864 15436 19916
rect 16396 19864 16448 19916
rect 18512 19864 18564 19916
rect 22008 19864 22060 19916
rect 11244 19796 11296 19848
rect 12992 19839 13044 19848
rect 12992 19805 13001 19839
rect 13001 19805 13035 19839
rect 13035 19805 13044 19839
rect 12992 19796 13044 19805
rect 19064 19839 19116 19848
rect 19064 19805 19073 19839
rect 19073 19805 19107 19839
rect 19107 19805 19116 19839
rect 21548 19839 21600 19848
rect 19064 19796 19116 19805
rect 21548 19805 21557 19839
rect 21557 19805 21591 19839
rect 21591 19805 21600 19839
rect 21548 19796 21600 19805
rect 9588 19728 9640 19780
rect 12256 19728 12308 19780
rect 23940 19932 23992 19984
rect 24860 19932 24912 19984
rect 22836 19907 22888 19916
rect 22836 19873 22845 19907
rect 22845 19873 22879 19907
rect 22879 19873 22888 19907
rect 22836 19864 22888 19873
rect 23480 19864 23532 19916
rect 24032 19864 24084 19916
rect 24584 19864 24636 19916
rect 25044 19864 25096 19916
rect 22928 19839 22980 19848
rect 22928 19805 22937 19839
rect 22937 19805 22971 19839
rect 22971 19805 22980 19839
rect 22928 19796 22980 19805
rect 23204 19796 23256 19848
rect 23296 19796 23348 19848
rect 24492 19839 24544 19848
rect 24492 19805 24501 19839
rect 24501 19805 24535 19839
rect 24535 19805 24544 19839
rect 24492 19796 24544 19805
rect 23388 19728 23440 19780
rect 24768 19796 24820 19848
rect 4252 19660 4304 19712
rect 7196 19703 7248 19712
rect 7196 19669 7205 19703
rect 7205 19669 7239 19703
rect 7239 19669 7248 19703
rect 7196 19660 7248 19669
rect 9128 19703 9180 19712
rect 9128 19669 9137 19703
rect 9137 19669 9171 19703
rect 9171 19669 9180 19703
rect 9128 19660 9180 19669
rect 11244 19660 11296 19712
rect 15844 19703 15896 19712
rect 15844 19669 15853 19703
rect 15853 19669 15887 19703
rect 15887 19669 15896 19703
rect 15844 19660 15896 19669
rect 18236 19703 18288 19712
rect 18236 19669 18245 19703
rect 18245 19669 18279 19703
rect 18279 19669 18288 19703
rect 18236 19660 18288 19669
rect 19432 19660 19484 19712
rect 19708 19703 19760 19712
rect 19708 19669 19717 19703
rect 19717 19669 19751 19703
rect 19751 19669 19760 19703
rect 19708 19660 19760 19669
rect 20352 19703 20404 19712
rect 20352 19669 20361 19703
rect 20361 19669 20395 19703
rect 20395 19669 20404 19703
rect 20352 19660 20404 19669
rect 20904 19703 20956 19712
rect 20904 19669 20913 19703
rect 20913 19669 20947 19703
rect 20947 19669 20956 19703
rect 20904 19660 20956 19669
rect 21088 19660 21140 19712
rect 21640 19660 21692 19712
rect 25228 19660 25280 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 2044 19456 2096 19508
rect 2228 19456 2280 19508
rect 4712 19499 4764 19508
rect 4712 19465 4721 19499
rect 4721 19465 4755 19499
rect 4755 19465 4764 19499
rect 4712 19456 4764 19465
rect 8392 19499 8444 19508
rect 8392 19465 8401 19499
rect 8401 19465 8435 19499
rect 8435 19465 8444 19499
rect 8392 19456 8444 19465
rect 10784 19499 10836 19508
rect 10784 19465 10793 19499
rect 10793 19465 10827 19499
rect 10827 19465 10836 19499
rect 10784 19456 10836 19465
rect 11520 19456 11572 19508
rect 12532 19456 12584 19508
rect 12900 19456 12952 19508
rect 4804 19388 4856 19440
rect 6460 19388 6512 19440
rect 7104 19388 7156 19440
rect 12256 19388 12308 19440
rect 14188 19456 14240 19508
rect 14556 19456 14608 19508
rect 16396 19456 16448 19508
rect 6092 19320 6144 19372
rect 7656 19320 7708 19372
rect 3608 19252 3660 19304
rect 3976 19252 4028 19304
rect 4344 19252 4396 19304
rect 5172 19252 5224 19304
rect 7012 19252 7064 19304
rect 8208 19252 8260 19304
rect 9404 19252 9456 19304
rect 10232 19295 10284 19304
rect 10232 19261 10241 19295
rect 10241 19261 10275 19295
rect 10275 19261 10284 19295
rect 11152 19320 11204 19372
rect 11244 19320 11296 19372
rect 10232 19252 10284 19261
rect 10784 19252 10836 19304
rect 10968 19252 11020 19304
rect 12072 19320 12124 19372
rect 2780 19184 2832 19236
rect 2320 19116 2372 19168
rect 2872 19116 2924 19168
rect 3056 19159 3108 19168
rect 3056 19125 3065 19159
rect 3065 19125 3099 19159
rect 3099 19125 3108 19159
rect 3056 19116 3108 19125
rect 6276 19184 6328 19236
rect 8300 19184 8352 19236
rect 3976 19159 4028 19168
rect 3976 19125 3985 19159
rect 3985 19125 4019 19159
rect 4019 19125 4028 19159
rect 3976 19116 4028 19125
rect 4988 19159 5040 19168
rect 4988 19125 4997 19159
rect 4997 19125 5031 19159
rect 5031 19125 5040 19159
rect 4988 19116 5040 19125
rect 5356 19116 5408 19168
rect 6368 19116 6420 19168
rect 6644 19116 6696 19168
rect 8024 19159 8076 19168
rect 8024 19125 8033 19159
rect 8033 19125 8067 19159
rect 8067 19125 8076 19159
rect 8024 19116 8076 19125
rect 10968 19116 11020 19168
rect 11244 19227 11296 19236
rect 11244 19193 11253 19227
rect 11253 19193 11287 19227
rect 11287 19193 11296 19227
rect 11244 19184 11296 19193
rect 11704 19184 11756 19236
rect 12072 19184 12124 19236
rect 11796 19116 11848 19168
rect 11980 19116 12032 19168
rect 15200 19388 15252 19440
rect 16764 19456 16816 19508
rect 20628 19456 20680 19508
rect 22836 19456 22888 19508
rect 23664 19499 23716 19508
rect 23664 19465 23673 19499
rect 23673 19465 23707 19499
rect 23707 19465 23716 19499
rect 23664 19456 23716 19465
rect 14556 19363 14608 19372
rect 14556 19329 14565 19363
rect 14565 19329 14599 19363
rect 14599 19329 14608 19363
rect 14556 19320 14608 19329
rect 15384 19320 15436 19372
rect 20076 19388 20128 19440
rect 13452 19252 13504 19304
rect 13820 19252 13872 19304
rect 14096 19252 14148 19304
rect 15292 19295 15344 19304
rect 15292 19261 15301 19295
rect 15301 19261 15335 19295
rect 15335 19261 15344 19295
rect 15292 19252 15344 19261
rect 12624 19116 12676 19168
rect 13452 19159 13504 19168
rect 13452 19125 13461 19159
rect 13461 19125 13495 19159
rect 13495 19125 13504 19159
rect 13452 19116 13504 19125
rect 13912 19116 13964 19168
rect 20352 19320 20404 19372
rect 21824 19320 21876 19372
rect 22284 19320 22336 19372
rect 23940 19320 23992 19372
rect 24584 19388 24636 19440
rect 15844 19252 15896 19304
rect 16580 19252 16632 19304
rect 18972 19252 19024 19304
rect 19340 19252 19392 19304
rect 20260 19252 20312 19304
rect 20628 19252 20680 19304
rect 22744 19252 22796 19304
rect 22928 19295 22980 19304
rect 22928 19261 22937 19295
rect 22937 19261 22971 19295
rect 22971 19261 22980 19295
rect 22928 19252 22980 19261
rect 24676 19252 24728 19304
rect 24860 19252 24912 19304
rect 25504 19252 25556 19304
rect 26240 19295 26292 19304
rect 26240 19261 26249 19295
rect 26249 19261 26283 19295
rect 26283 19261 26292 19295
rect 26240 19252 26292 19261
rect 18236 19184 18288 19236
rect 15844 19116 15896 19168
rect 16856 19116 16908 19168
rect 17408 19116 17460 19168
rect 17684 19116 17736 19168
rect 18604 19116 18656 19168
rect 19340 19116 19392 19168
rect 20260 19116 20312 19168
rect 20720 19159 20772 19168
rect 20720 19125 20729 19159
rect 20729 19125 20763 19159
rect 20763 19125 20772 19159
rect 20720 19116 20772 19125
rect 21180 19159 21232 19168
rect 21180 19125 21189 19159
rect 21189 19125 21223 19159
rect 21223 19125 21232 19159
rect 21180 19116 21232 19125
rect 23296 19116 23348 19168
rect 24768 19159 24820 19168
rect 24768 19125 24777 19159
rect 24777 19125 24811 19159
rect 24811 19125 24820 19159
rect 24768 19116 24820 19125
rect 25044 19116 25096 19168
rect 25596 19116 25648 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1860 18912 1912 18964
rect 2964 18912 3016 18964
rect 3700 18955 3752 18964
rect 3700 18921 3709 18955
rect 3709 18921 3743 18955
rect 3743 18921 3752 18955
rect 3700 18912 3752 18921
rect 4712 18955 4764 18964
rect 1952 18844 2004 18896
rect 4712 18921 4721 18955
rect 4721 18921 4755 18955
rect 4755 18921 4764 18955
rect 4712 18912 4764 18921
rect 5448 18912 5500 18964
rect 5264 18844 5316 18896
rect 6184 18912 6236 18964
rect 6092 18844 6144 18896
rect 6368 18887 6420 18896
rect 6368 18853 6377 18887
rect 6377 18853 6411 18887
rect 6411 18853 6420 18887
rect 6368 18844 6420 18853
rect 4620 18776 4672 18828
rect 5080 18776 5132 18828
rect 3056 18751 3108 18760
rect 3056 18717 3065 18751
rect 3065 18717 3099 18751
rect 3099 18717 3108 18751
rect 3056 18708 3108 18717
rect 5540 18708 5592 18760
rect 6000 18751 6052 18760
rect 6000 18717 6009 18751
rect 6009 18717 6043 18751
rect 6043 18717 6052 18751
rect 6000 18708 6052 18717
rect 1124 18640 1176 18692
rect 7012 18912 7064 18964
rect 8300 18955 8352 18964
rect 8300 18921 8309 18955
rect 8309 18921 8343 18955
rect 8343 18921 8352 18955
rect 8300 18912 8352 18921
rect 11060 18912 11112 18964
rect 13728 18912 13780 18964
rect 8484 18844 8536 18896
rect 9864 18844 9916 18896
rect 11520 18887 11572 18896
rect 11520 18853 11529 18887
rect 11529 18853 11563 18887
rect 11563 18853 11572 18887
rect 11520 18844 11572 18853
rect 11796 18844 11848 18896
rect 6828 18776 6880 18828
rect 7196 18819 7248 18828
rect 7196 18785 7230 18819
rect 7230 18785 7248 18819
rect 7196 18776 7248 18785
rect 9956 18776 10008 18828
rect 10324 18776 10376 18828
rect 10876 18776 10928 18828
rect 12808 18819 12860 18828
rect 12808 18785 12817 18819
rect 12817 18785 12851 18819
rect 12851 18785 12860 18819
rect 12808 18776 12860 18785
rect 12992 18844 13044 18896
rect 14556 18844 14608 18896
rect 16304 18912 16356 18964
rect 16396 18912 16448 18964
rect 16764 18912 16816 18964
rect 17684 18912 17736 18964
rect 20628 18912 20680 18964
rect 21824 18912 21876 18964
rect 22192 18912 22244 18964
rect 23480 18912 23532 18964
rect 23664 18955 23716 18964
rect 23664 18921 23673 18955
rect 23673 18921 23707 18955
rect 23707 18921 23716 18955
rect 23664 18912 23716 18921
rect 24124 18912 24176 18964
rect 24492 18955 24544 18964
rect 24492 18921 24501 18955
rect 24501 18921 24535 18955
rect 24535 18921 24544 18955
rect 24492 18912 24544 18921
rect 19064 18844 19116 18896
rect 15384 18776 15436 18828
rect 15844 18776 15896 18828
rect 11152 18708 11204 18760
rect 11520 18708 11572 18760
rect 11704 18751 11756 18760
rect 11704 18717 11713 18751
rect 11713 18717 11747 18751
rect 11747 18717 11756 18751
rect 11704 18708 11756 18717
rect 11888 18708 11940 18760
rect 12532 18708 12584 18760
rect 13820 18640 13872 18692
rect 16488 18708 16540 18760
rect 1952 18615 2004 18624
rect 1952 18581 1961 18615
rect 1961 18581 1995 18615
rect 1995 18581 2004 18615
rect 1952 18572 2004 18581
rect 2504 18572 2556 18624
rect 6828 18615 6880 18624
rect 6828 18581 6837 18615
rect 6837 18581 6871 18615
rect 6871 18581 6880 18615
rect 6828 18572 6880 18581
rect 7564 18572 7616 18624
rect 9864 18615 9916 18624
rect 9864 18581 9873 18615
rect 9873 18581 9907 18615
rect 9907 18581 9916 18615
rect 9864 18572 9916 18581
rect 10324 18615 10376 18624
rect 10324 18581 10333 18615
rect 10333 18581 10367 18615
rect 10367 18581 10376 18615
rect 10324 18572 10376 18581
rect 10968 18572 11020 18624
rect 11612 18572 11664 18624
rect 12532 18615 12584 18624
rect 12532 18581 12541 18615
rect 12541 18581 12575 18615
rect 12575 18581 12584 18615
rect 12532 18572 12584 18581
rect 14832 18615 14884 18624
rect 14832 18581 14841 18615
rect 14841 18581 14875 18615
rect 14875 18581 14884 18615
rect 14832 18572 14884 18581
rect 16304 18615 16356 18624
rect 16304 18581 16313 18615
rect 16313 18581 16347 18615
rect 16347 18581 16356 18615
rect 16304 18572 16356 18581
rect 16856 18776 16908 18828
rect 23204 18844 23256 18896
rect 23940 18844 23992 18896
rect 19432 18819 19484 18828
rect 19432 18785 19441 18819
rect 19441 18785 19475 18819
rect 19475 18785 19484 18819
rect 19432 18776 19484 18785
rect 21824 18776 21876 18828
rect 22100 18776 22152 18828
rect 19524 18751 19576 18760
rect 19524 18717 19533 18751
rect 19533 18717 19567 18751
rect 19567 18717 19576 18751
rect 19524 18708 19576 18717
rect 21364 18751 21416 18760
rect 21364 18717 21373 18751
rect 21373 18717 21407 18751
rect 21407 18717 21416 18751
rect 21364 18708 21416 18717
rect 21640 18708 21692 18760
rect 19432 18640 19484 18692
rect 21916 18640 21968 18692
rect 23480 18776 23532 18828
rect 24676 18844 24728 18896
rect 25044 18776 25096 18828
rect 23112 18751 23164 18760
rect 23112 18717 23121 18751
rect 23121 18717 23155 18751
rect 23155 18717 23164 18751
rect 23112 18708 23164 18717
rect 23296 18708 23348 18760
rect 24676 18708 24728 18760
rect 17408 18572 17460 18624
rect 18144 18615 18196 18624
rect 18144 18581 18153 18615
rect 18153 18581 18187 18615
rect 18187 18581 18196 18615
rect 18144 18572 18196 18581
rect 18512 18615 18564 18624
rect 18512 18581 18521 18615
rect 18521 18581 18555 18615
rect 18555 18581 18564 18615
rect 18512 18572 18564 18581
rect 18972 18615 19024 18624
rect 18972 18581 18981 18615
rect 18981 18581 19015 18615
rect 19015 18581 19024 18615
rect 18972 18572 19024 18581
rect 20260 18572 20312 18624
rect 20812 18572 20864 18624
rect 21548 18572 21600 18624
rect 22284 18572 22336 18624
rect 24952 18572 25004 18624
rect 25228 18572 25280 18624
rect 26240 18572 26292 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 2964 18368 3016 18420
rect 4620 18411 4672 18420
rect 4620 18377 4629 18411
rect 4629 18377 4663 18411
rect 4663 18377 4672 18411
rect 4620 18368 4672 18377
rect 5080 18411 5132 18420
rect 5080 18377 5089 18411
rect 5089 18377 5123 18411
rect 5123 18377 5132 18411
rect 5080 18368 5132 18377
rect 6000 18368 6052 18420
rect 7196 18368 7248 18420
rect 9312 18368 9364 18420
rect 848 18300 900 18352
rect 1952 18232 2004 18284
rect 2596 18275 2648 18284
rect 2596 18241 2605 18275
rect 2605 18241 2639 18275
rect 2639 18241 2648 18275
rect 2596 18232 2648 18241
rect 1584 18164 1636 18216
rect 4344 18232 4396 18284
rect 4712 18232 4764 18284
rect 7012 18343 7064 18352
rect 7012 18309 7021 18343
rect 7021 18309 7055 18343
rect 7055 18309 7064 18343
rect 7012 18300 7064 18309
rect 7932 18300 7984 18352
rect 8300 18300 8352 18352
rect 12992 18368 13044 18420
rect 13452 18411 13504 18420
rect 13452 18377 13461 18411
rect 13461 18377 13495 18411
rect 13495 18377 13504 18411
rect 13452 18368 13504 18377
rect 14004 18411 14056 18420
rect 14004 18377 14013 18411
rect 14013 18377 14047 18411
rect 14047 18377 14056 18411
rect 14004 18368 14056 18377
rect 15384 18368 15436 18420
rect 15936 18368 15988 18420
rect 6828 18232 6880 18284
rect 7472 18275 7524 18284
rect 7472 18241 7481 18275
rect 7481 18241 7515 18275
rect 7515 18241 7524 18275
rect 7472 18232 7524 18241
rect 9036 18275 9088 18284
rect 1492 18028 1544 18080
rect 3884 18164 3936 18216
rect 4068 18207 4120 18216
rect 4068 18173 4077 18207
rect 4077 18173 4111 18207
rect 4111 18173 4120 18207
rect 4068 18164 4120 18173
rect 4528 18164 4580 18216
rect 9036 18241 9045 18275
rect 9045 18241 9079 18275
rect 9079 18241 9088 18275
rect 9036 18232 9088 18241
rect 12256 18300 12308 18352
rect 13728 18300 13780 18352
rect 17684 18368 17736 18420
rect 17960 18368 18012 18420
rect 21364 18368 21416 18420
rect 23388 18368 23440 18420
rect 23756 18368 23808 18420
rect 24952 18368 25004 18420
rect 16580 18300 16632 18352
rect 22100 18300 22152 18352
rect 22284 18300 22336 18352
rect 23112 18300 23164 18352
rect 24676 18343 24728 18352
rect 8208 18164 8260 18216
rect 8576 18164 8628 18216
rect 9404 18164 9456 18216
rect 12808 18232 12860 18284
rect 14556 18275 14608 18284
rect 14556 18241 14565 18275
rect 14565 18241 14599 18275
rect 14599 18241 14608 18275
rect 14556 18232 14608 18241
rect 16764 18275 16816 18284
rect 16764 18241 16773 18275
rect 16773 18241 16807 18275
rect 16807 18241 16816 18275
rect 16764 18232 16816 18241
rect 19064 18232 19116 18284
rect 19616 18232 19668 18284
rect 20352 18232 20404 18284
rect 11244 18164 11296 18216
rect 11520 18164 11572 18216
rect 13912 18164 13964 18216
rect 2044 18071 2096 18080
rect 2044 18037 2053 18071
rect 2053 18037 2087 18071
rect 2087 18037 2096 18071
rect 2044 18028 2096 18037
rect 2228 18028 2280 18080
rect 2688 18028 2740 18080
rect 3884 18028 3936 18080
rect 5448 18028 5500 18080
rect 5632 18071 5684 18080
rect 5632 18037 5641 18071
rect 5641 18037 5675 18071
rect 5675 18037 5684 18071
rect 5632 18028 5684 18037
rect 7564 18028 7616 18080
rect 7932 18028 7984 18080
rect 8576 18071 8628 18080
rect 8576 18037 8585 18071
rect 8585 18037 8619 18071
rect 8619 18037 8628 18071
rect 8576 18028 8628 18037
rect 10692 18096 10744 18148
rect 10784 18096 10836 18148
rect 9772 18028 9824 18080
rect 11060 18096 11112 18148
rect 10968 18028 11020 18080
rect 11704 18028 11756 18080
rect 12164 18071 12216 18080
rect 12164 18037 12173 18071
rect 12173 18037 12207 18071
rect 12207 18037 12216 18071
rect 12164 18028 12216 18037
rect 12440 18071 12492 18080
rect 12440 18037 12449 18071
rect 12449 18037 12483 18071
rect 12483 18037 12492 18071
rect 12440 18028 12492 18037
rect 15384 18096 15436 18148
rect 17316 18096 17368 18148
rect 13176 18028 13228 18080
rect 14372 18071 14424 18080
rect 14372 18037 14381 18071
rect 14381 18037 14415 18071
rect 14415 18037 14424 18071
rect 14372 18028 14424 18037
rect 15108 18071 15160 18080
rect 15108 18037 15117 18071
rect 15117 18037 15151 18071
rect 15151 18037 15160 18071
rect 15108 18028 15160 18037
rect 15844 18071 15896 18080
rect 15844 18037 15853 18071
rect 15853 18037 15887 18071
rect 15887 18037 15896 18071
rect 15844 18028 15896 18037
rect 16580 18071 16632 18080
rect 16580 18037 16589 18071
rect 16589 18037 16623 18071
rect 16623 18037 16632 18071
rect 16580 18028 16632 18037
rect 17132 18028 17184 18080
rect 19248 18164 19300 18216
rect 20904 18164 20956 18216
rect 20720 18139 20772 18148
rect 20720 18105 20729 18139
rect 20729 18105 20763 18139
rect 20763 18105 20772 18139
rect 23664 18232 23716 18284
rect 24676 18309 24685 18343
rect 24685 18309 24719 18343
rect 24719 18309 24728 18343
rect 24676 18300 24728 18309
rect 25504 18275 25556 18284
rect 25504 18241 25513 18275
rect 25513 18241 25547 18275
rect 25547 18241 25556 18275
rect 25504 18232 25556 18241
rect 26332 18275 26384 18284
rect 26332 18241 26341 18275
rect 26341 18241 26375 18275
rect 26375 18241 26384 18275
rect 26332 18232 26384 18241
rect 23848 18164 23900 18216
rect 25228 18207 25280 18216
rect 25228 18173 25237 18207
rect 25237 18173 25271 18207
rect 25271 18173 25280 18207
rect 25228 18164 25280 18173
rect 20720 18096 20772 18105
rect 23756 18096 23808 18148
rect 19064 18071 19116 18080
rect 19064 18037 19073 18071
rect 19073 18037 19107 18071
rect 19107 18037 19116 18071
rect 19064 18028 19116 18037
rect 19248 18071 19300 18080
rect 19248 18037 19257 18071
rect 19257 18037 19291 18071
rect 19291 18037 19300 18071
rect 19248 18028 19300 18037
rect 20904 18028 20956 18080
rect 21364 18028 21416 18080
rect 23112 18028 23164 18080
rect 25228 18028 25280 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 2412 17867 2464 17876
rect 2412 17833 2421 17867
rect 2421 17833 2455 17867
rect 2455 17833 2464 17867
rect 2412 17824 2464 17833
rect 4344 17867 4396 17876
rect 4344 17833 4353 17867
rect 4353 17833 4387 17867
rect 4387 17833 4396 17867
rect 4344 17824 4396 17833
rect 5264 17824 5316 17876
rect 6000 17824 6052 17876
rect 6920 17824 6972 17876
rect 7196 17824 7248 17876
rect 8484 17867 8536 17876
rect 8484 17833 8493 17867
rect 8493 17833 8527 17867
rect 8527 17833 8536 17867
rect 8484 17824 8536 17833
rect 8852 17867 8904 17876
rect 8852 17833 8861 17867
rect 8861 17833 8895 17867
rect 8895 17833 8904 17867
rect 8852 17824 8904 17833
rect 13084 17824 13136 17876
rect 13452 17824 13504 17876
rect 14188 17867 14240 17876
rect 14188 17833 14197 17867
rect 14197 17833 14231 17867
rect 14231 17833 14240 17867
rect 14188 17824 14240 17833
rect 15108 17867 15160 17876
rect 15108 17833 15117 17867
rect 15117 17833 15151 17867
rect 15151 17833 15160 17867
rect 15108 17824 15160 17833
rect 15292 17867 15344 17876
rect 15292 17833 15301 17867
rect 15301 17833 15335 17867
rect 15335 17833 15344 17867
rect 15292 17824 15344 17833
rect 15936 17824 15988 17876
rect 16396 17867 16448 17876
rect 16396 17833 16405 17867
rect 16405 17833 16439 17867
rect 16439 17833 16448 17867
rect 16396 17824 16448 17833
rect 16856 17867 16908 17876
rect 16856 17833 16865 17867
rect 16865 17833 16899 17867
rect 16899 17833 16908 17867
rect 16856 17824 16908 17833
rect 17408 17824 17460 17876
rect 17960 17824 18012 17876
rect 19524 17824 19576 17876
rect 1952 17756 2004 17808
rect 2596 17756 2648 17808
rect 6644 17756 6696 17808
rect 9680 17799 9732 17808
rect 9680 17765 9689 17799
rect 9689 17765 9723 17799
rect 9723 17765 9732 17799
rect 9680 17756 9732 17765
rect 10968 17756 11020 17808
rect 2872 17663 2924 17672
rect 2872 17629 2881 17663
rect 2881 17629 2915 17663
rect 2915 17629 2924 17663
rect 2872 17620 2924 17629
rect 6184 17688 6236 17740
rect 7564 17688 7616 17740
rect 8392 17688 8444 17740
rect 11060 17731 11112 17740
rect 11060 17697 11069 17731
rect 11069 17697 11103 17731
rect 11103 17697 11112 17731
rect 11060 17688 11112 17697
rect 3884 17620 3936 17672
rect 4988 17663 5040 17672
rect 4988 17629 4997 17663
rect 4997 17629 5031 17663
rect 5031 17629 5040 17663
rect 4988 17620 5040 17629
rect 5080 17663 5132 17672
rect 5080 17629 5089 17663
rect 5089 17629 5123 17663
rect 5123 17629 5132 17663
rect 5080 17620 5132 17629
rect 5540 17620 5592 17672
rect 6000 17620 6052 17672
rect 10968 17620 11020 17672
rect 11336 17756 11388 17808
rect 11888 17756 11940 17808
rect 12808 17756 12860 17808
rect 14556 17756 14608 17808
rect 12900 17688 12952 17740
rect 14648 17688 14700 17740
rect 11336 17663 11388 17672
rect 11336 17629 11345 17663
rect 11345 17629 11379 17663
rect 11379 17629 11388 17663
rect 11336 17620 11388 17629
rect 13084 17663 13136 17672
rect 13084 17629 13093 17663
rect 13093 17629 13127 17663
rect 13127 17629 13136 17663
rect 13084 17620 13136 17629
rect 14372 17620 14424 17672
rect 14740 17620 14792 17672
rect 13452 17552 13504 17604
rect 14924 17552 14976 17604
rect 18512 17756 18564 17808
rect 19984 17824 20036 17876
rect 20076 17756 20128 17808
rect 20352 17824 20404 17876
rect 22008 17824 22060 17876
rect 22192 17824 22244 17876
rect 23296 17867 23348 17876
rect 23296 17833 23305 17867
rect 23305 17833 23339 17867
rect 23339 17833 23348 17867
rect 23296 17824 23348 17833
rect 23848 17824 23900 17876
rect 24308 17824 24360 17876
rect 21548 17756 21600 17808
rect 21824 17756 21876 17808
rect 24032 17756 24084 17808
rect 17408 17731 17460 17740
rect 17408 17697 17442 17731
rect 17442 17697 17460 17731
rect 17408 17688 17460 17697
rect 19984 17688 20036 17740
rect 20352 17688 20404 17740
rect 21364 17688 21416 17740
rect 22376 17688 22428 17740
rect 23204 17731 23256 17740
rect 23204 17697 23213 17731
rect 23213 17697 23247 17731
rect 23247 17697 23256 17731
rect 23204 17688 23256 17697
rect 24676 17688 24728 17740
rect 20904 17620 20956 17672
rect 23388 17663 23440 17672
rect 16488 17552 16540 17604
rect 21180 17552 21232 17604
rect 23388 17629 23397 17663
rect 23397 17629 23431 17663
rect 23431 17629 23440 17663
rect 23388 17620 23440 17629
rect 23940 17620 23992 17672
rect 25044 17824 25096 17876
rect 22008 17552 22060 17604
rect 23480 17552 23532 17604
rect 25044 17620 25096 17672
rect 1676 17527 1728 17536
rect 1676 17493 1685 17527
rect 1685 17493 1719 17527
rect 1719 17493 1728 17527
rect 1676 17484 1728 17493
rect 2688 17484 2740 17536
rect 3056 17484 3108 17536
rect 4068 17484 4120 17536
rect 6000 17484 6052 17536
rect 6368 17484 6420 17536
rect 8116 17527 8168 17536
rect 8116 17493 8125 17527
rect 8125 17493 8159 17527
rect 8159 17493 8168 17527
rect 8116 17484 8168 17493
rect 9772 17484 9824 17536
rect 13820 17484 13872 17536
rect 13912 17484 13964 17536
rect 14740 17527 14792 17536
rect 14740 17493 14749 17527
rect 14749 17493 14783 17527
rect 14783 17493 14792 17527
rect 14740 17484 14792 17493
rect 16764 17484 16816 17536
rect 18880 17484 18932 17536
rect 21640 17484 21692 17536
rect 24216 17484 24268 17536
rect 25228 17484 25280 17536
rect 26240 17527 26292 17536
rect 26240 17493 26249 17527
rect 26249 17493 26283 17527
rect 26283 17493 26292 17527
rect 26240 17484 26292 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 1584 17323 1636 17332
rect 1584 17289 1593 17323
rect 1593 17289 1627 17323
rect 1627 17289 1636 17323
rect 1584 17280 1636 17289
rect 2596 17323 2648 17332
rect 2596 17289 2605 17323
rect 2605 17289 2639 17323
rect 2639 17289 2648 17323
rect 2596 17280 2648 17289
rect 6368 17280 6420 17332
rect 6736 17280 6788 17332
rect 7472 17280 7524 17332
rect 8300 17280 8352 17332
rect 2228 17187 2280 17196
rect 2228 17153 2237 17187
rect 2237 17153 2271 17187
rect 2271 17153 2280 17187
rect 2228 17144 2280 17153
rect 3424 17144 3476 17196
rect 5080 17212 5132 17264
rect 6184 17255 6236 17264
rect 6184 17221 6193 17255
rect 6193 17221 6227 17255
rect 6227 17221 6236 17255
rect 6184 17212 6236 17221
rect 5172 17187 5224 17196
rect 5172 17153 5181 17187
rect 5181 17153 5215 17187
rect 5215 17153 5224 17187
rect 5172 17144 5224 17153
rect 5264 17187 5316 17196
rect 5264 17153 5273 17187
rect 5273 17153 5307 17187
rect 5307 17153 5316 17187
rect 5264 17144 5316 17153
rect 6092 17144 6144 17196
rect 8944 17212 8996 17264
rect 8760 17187 8812 17196
rect 8760 17153 8769 17187
rect 8769 17153 8803 17187
rect 8803 17153 8812 17187
rect 8760 17144 8812 17153
rect 9312 17144 9364 17196
rect 10048 17280 10100 17332
rect 10784 17280 10836 17332
rect 11244 17280 11296 17332
rect 14004 17280 14056 17332
rect 14464 17280 14516 17332
rect 14832 17323 14884 17332
rect 14832 17289 14841 17323
rect 14841 17289 14875 17323
rect 14875 17289 14884 17323
rect 14832 17280 14884 17289
rect 18052 17323 18104 17332
rect 18052 17289 18061 17323
rect 18061 17289 18095 17323
rect 18095 17289 18104 17323
rect 18052 17280 18104 17289
rect 19248 17280 19300 17332
rect 19432 17280 19484 17332
rect 22376 17280 22428 17332
rect 22652 17280 22704 17332
rect 23756 17280 23808 17332
rect 24676 17280 24728 17332
rect 26332 17323 26384 17332
rect 26332 17289 26341 17323
rect 26341 17289 26375 17323
rect 26375 17289 26384 17323
rect 26332 17280 26384 17289
rect 10968 17212 11020 17264
rect 12256 17212 12308 17264
rect 2872 17076 2924 17128
rect 3608 17076 3660 17128
rect 5080 17119 5132 17128
rect 5080 17085 5089 17119
rect 5089 17085 5123 17119
rect 5123 17085 5132 17119
rect 5080 17076 5132 17085
rect 7104 17076 7156 17128
rect 8576 17076 8628 17128
rect 9588 17076 9640 17128
rect 11060 17144 11112 17196
rect 1676 17008 1728 17060
rect 2688 17008 2740 17060
rect 4988 17008 5040 17060
rect 7564 17008 7616 17060
rect 9312 17008 9364 17060
rect 10140 17008 10192 17060
rect 13176 17076 13228 17128
rect 12716 17008 12768 17060
rect 2412 16940 2464 16992
rect 3148 16983 3200 16992
rect 3148 16949 3157 16983
rect 3157 16949 3191 16983
rect 3191 16949 3200 16983
rect 3148 16940 3200 16949
rect 3516 16983 3568 16992
rect 3516 16949 3525 16983
rect 3525 16949 3559 16983
rect 3559 16949 3568 16983
rect 3516 16940 3568 16949
rect 3976 16940 4028 16992
rect 4712 16983 4764 16992
rect 4712 16949 4721 16983
rect 4721 16949 4755 16983
rect 4755 16949 4764 16983
rect 4712 16940 4764 16949
rect 6460 16940 6512 16992
rect 8116 16940 8168 16992
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 13636 16940 13688 16992
rect 14648 17212 14700 17264
rect 24032 17212 24084 17264
rect 25320 17212 25372 17264
rect 25872 17212 25924 17264
rect 17408 17144 17460 17196
rect 18696 17187 18748 17196
rect 18696 17153 18705 17187
rect 18705 17153 18739 17187
rect 18739 17153 18748 17187
rect 18696 17144 18748 17153
rect 19432 17144 19484 17196
rect 21548 17144 21600 17196
rect 23112 17144 23164 17196
rect 23664 17144 23716 17196
rect 24216 17144 24268 17196
rect 25412 17187 25464 17196
rect 14464 17119 14516 17128
rect 14464 17085 14473 17119
rect 14473 17085 14507 17119
rect 14507 17085 14516 17119
rect 14464 17076 14516 17085
rect 14648 17119 14700 17128
rect 14648 17085 14657 17119
rect 14657 17085 14691 17119
rect 14691 17085 14700 17119
rect 14648 17076 14700 17085
rect 15200 17076 15252 17128
rect 18052 17076 18104 17128
rect 18512 17119 18564 17128
rect 18512 17085 18521 17119
rect 18521 17085 18555 17119
rect 18555 17085 18564 17119
rect 18512 17076 18564 17085
rect 19248 17076 19300 17128
rect 21824 17076 21876 17128
rect 25412 17153 25421 17187
rect 25421 17153 25455 17187
rect 25455 17153 25464 17187
rect 25412 17144 25464 17153
rect 24768 17076 24820 17128
rect 24952 17076 25004 17128
rect 16580 17008 16632 17060
rect 17684 17008 17736 17060
rect 18604 17008 18656 17060
rect 20352 17008 20404 17060
rect 14096 16940 14148 16992
rect 15108 16940 15160 16992
rect 15936 16940 15988 16992
rect 19340 16940 19392 16992
rect 20076 16983 20128 16992
rect 20076 16949 20085 16983
rect 20085 16949 20119 16983
rect 20119 16949 20128 16983
rect 20076 16940 20128 16949
rect 20904 16983 20956 16992
rect 20904 16949 20913 16983
rect 20913 16949 20947 16983
rect 20947 16949 20956 16983
rect 20904 16940 20956 16949
rect 21180 16940 21232 16992
rect 21548 16940 21600 16992
rect 22008 16940 22060 16992
rect 23480 17008 23532 17060
rect 23296 16940 23348 16992
rect 23756 16940 23808 16992
rect 24032 16983 24084 16992
rect 24032 16949 24041 16983
rect 24041 16949 24075 16983
rect 24075 16949 24084 16983
rect 24032 16940 24084 16949
rect 24216 16940 24268 16992
rect 24676 16940 24728 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 2228 16736 2280 16788
rect 2964 16779 3016 16788
rect 1676 16668 1728 16720
rect 2412 16711 2464 16720
rect 2412 16677 2421 16711
rect 2421 16677 2455 16711
rect 2455 16677 2464 16711
rect 2412 16668 2464 16677
rect 2964 16745 2973 16779
rect 2973 16745 3007 16779
rect 3007 16745 3016 16779
rect 2964 16736 3016 16745
rect 4344 16736 4396 16788
rect 4160 16600 4212 16652
rect 4712 16668 4764 16720
rect 6092 16736 6144 16788
rect 7196 16779 7248 16788
rect 1952 16532 2004 16584
rect 2136 16532 2188 16584
rect 3424 16532 3476 16584
rect 6092 16575 6144 16584
rect 6092 16541 6101 16575
rect 6101 16541 6135 16575
rect 6135 16541 6144 16575
rect 6092 16532 6144 16541
rect 6184 16575 6236 16584
rect 6184 16541 6193 16575
rect 6193 16541 6227 16575
rect 6227 16541 6236 16575
rect 6184 16532 6236 16541
rect 7196 16745 7205 16779
rect 7205 16745 7239 16779
rect 7239 16745 7248 16779
rect 7196 16736 7248 16745
rect 7748 16736 7800 16788
rect 8392 16779 8444 16788
rect 8392 16745 8401 16779
rect 8401 16745 8435 16779
rect 8435 16745 8444 16779
rect 8392 16736 8444 16745
rect 8576 16736 8628 16788
rect 9036 16779 9088 16788
rect 9036 16745 9045 16779
rect 9045 16745 9079 16779
rect 9079 16745 9088 16779
rect 9036 16736 9088 16745
rect 9404 16779 9456 16788
rect 9404 16745 9413 16779
rect 9413 16745 9447 16779
rect 9447 16745 9456 16779
rect 9404 16736 9456 16745
rect 9956 16736 10008 16788
rect 10140 16736 10192 16788
rect 11336 16779 11388 16788
rect 11336 16745 11345 16779
rect 11345 16745 11379 16779
rect 11379 16745 11388 16779
rect 11336 16736 11388 16745
rect 12900 16736 12952 16788
rect 14372 16779 14424 16788
rect 14372 16745 14381 16779
rect 14381 16745 14415 16779
rect 14415 16745 14424 16779
rect 14372 16736 14424 16745
rect 14648 16779 14700 16788
rect 14648 16745 14657 16779
rect 14657 16745 14691 16779
rect 14691 16745 14700 16779
rect 14648 16736 14700 16745
rect 16580 16736 16632 16788
rect 17408 16736 17460 16788
rect 17868 16736 17920 16788
rect 19524 16736 19576 16788
rect 20352 16779 20404 16788
rect 20352 16745 20361 16779
rect 20361 16745 20395 16779
rect 20395 16745 20404 16779
rect 20352 16736 20404 16745
rect 21364 16736 21416 16788
rect 22376 16736 22428 16788
rect 23388 16736 23440 16788
rect 23664 16736 23716 16788
rect 24860 16736 24912 16788
rect 10232 16668 10284 16720
rect 12072 16668 12124 16720
rect 14096 16668 14148 16720
rect 14556 16668 14608 16720
rect 6644 16643 6696 16652
rect 6644 16609 6653 16643
rect 6653 16609 6687 16643
rect 6687 16609 6696 16643
rect 6644 16600 6696 16609
rect 6552 16532 6604 16584
rect 7656 16600 7708 16652
rect 8760 16600 8812 16652
rect 9956 16643 10008 16652
rect 9956 16609 9990 16643
rect 9990 16609 10008 16643
rect 9956 16600 10008 16609
rect 11888 16600 11940 16652
rect 7472 16532 7524 16584
rect 9588 16532 9640 16584
rect 6644 16464 6696 16516
rect 1860 16396 1912 16448
rect 2044 16396 2096 16448
rect 3424 16439 3476 16448
rect 3424 16405 3433 16439
rect 3433 16405 3467 16439
rect 3467 16405 3476 16439
rect 3424 16396 3476 16405
rect 4068 16439 4120 16448
rect 4068 16405 4077 16439
rect 4077 16405 4111 16439
rect 4111 16405 4120 16439
rect 4068 16396 4120 16405
rect 5172 16439 5224 16448
rect 5172 16405 5181 16439
rect 5181 16405 5215 16439
rect 5215 16405 5224 16439
rect 5172 16396 5224 16405
rect 8300 16396 8352 16448
rect 8576 16396 8628 16448
rect 11336 16464 11388 16516
rect 11796 16396 11848 16448
rect 12440 16396 12492 16448
rect 13268 16600 13320 16652
rect 13636 16600 13688 16652
rect 15200 16600 15252 16652
rect 16304 16600 16356 16652
rect 17040 16600 17092 16652
rect 18052 16600 18104 16652
rect 18880 16668 18932 16720
rect 18972 16668 19024 16720
rect 19156 16668 19208 16720
rect 21548 16668 21600 16720
rect 19616 16600 19668 16652
rect 13912 16532 13964 16584
rect 14280 16532 14332 16584
rect 14372 16532 14424 16584
rect 25044 16668 25096 16720
rect 26240 16668 26292 16720
rect 22744 16600 22796 16652
rect 24676 16600 24728 16652
rect 25136 16643 25188 16652
rect 25136 16609 25145 16643
rect 25145 16609 25179 16643
rect 25179 16609 25188 16643
rect 25136 16600 25188 16609
rect 25412 16643 25464 16652
rect 25412 16609 25421 16643
rect 25421 16609 25455 16643
rect 25455 16609 25464 16643
rect 25412 16600 25464 16609
rect 25504 16600 25556 16652
rect 25780 16600 25832 16652
rect 20536 16532 20588 16584
rect 22376 16532 22428 16584
rect 23848 16532 23900 16584
rect 26332 16532 26384 16584
rect 13452 16507 13504 16516
rect 13452 16473 13461 16507
rect 13461 16473 13495 16507
rect 13495 16473 13504 16507
rect 13452 16464 13504 16473
rect 13636 16464 13688 16516
rect 15108 16464 15160 16516
rect 16764 16396 16816 16448
rect 18420 16396 18472 16448
rect 23296 16464 23348 16516
rect 23940 16464 23992 16516
rect 25136 16464 25188 16516
rect 22468 16396 22520 16448
rect 23848 16396 23900 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 940 16192 992 16244
rect 3332 16192 3384 16244
rect 3424 16192 3476 16244
rect 6644 16192 6696 16244
rect 7748 16192 7800 16244
rect 10140 16192 10192 16244
rect 10508 16235 10560 16244
rect 6460 16124 6512 16176
rect 2044 16099 2096 16108
rect 2044 16065 2053 16099
rect 2053 16065 2087 16099
rect 2087 16065 2096 16099
rect 2044 16056 2096 16065
rect 5356 16056 5408 16108
rect 1768 16031 1820 16040
rect 1768 15997 1777 16031
rect 1777 15997 1811 16031
rect 1811 15997 1820 16031
rect 1768 15988 1820 15997
rect 2228 15988 2280 16040
rect 2964 16031 3016 16040
rect 2964 15997 2973 16031
rect 2973 15997 3007 16031
rect 3007 15997 3016 16031
rect 2964 15988 3016 15997
rect 5448 15988 5500 16040
rect 7104 16099 7156 16108
rect 7104 16065 7113 16099
rect 7113 16065 7147 16099
rect 7147 16065 7156 16099
rect 7104 16056 7156 16065
rect 8300 16099 8352 16108
rect 8300 16065 8309 16099
rect 8309 16065 8343 16099
rect 8343 16065 8352 16099
rect 8300 16056 8352 16065
rect 8392 15988 8444 16040
rect 10508 16201 10517 16235
rect 10517 16201 10551 16235
rect 10551 16201 10560 16235
rect 10508 16192 10560 16201
rect 11796 16192 11848 16244
rect 12072 16235 12124 16244
rect 12072 16201 12081 16235
rect 12081 16201 12115 16235
rect 12115 16201 12124 16235
rect 12072 16192 12124 16201
rect 13084 16192 13136 16244
rect 11612 16056 11664 16108
rect 11796 16056 11848 16108
rect 13636 16056 13688 16108
rect 14372 16192 14424 16244
rect 15660 16192 15712 16244
rect 16304 16192 16356 16244
rect 17040 16235 17092 16244
rect 16212 16124 16264 16176
rect 17040 16201 17049 16235
rect 17049 16201 17083 16235
rect 17083 16201 17092 16235
rect 17040 16192 17092 16201
rect 17868 16192 17920 16244
rect 18880 16192 18932 16244
rect 18052 16124 18104 16176
rect 18604 16124 18656 16176
rect 20536 16192 20588 16244
rect 21916 16192 21968 16244
rect 22100 16192 22152 16244
rect 23388 16235 23440 16244
rect 18696 16099 18748 16108
rect 1676 15920 1728 15972
rect 3240 15963 3292 15972
rect 1400 15895 1452 15904
rect 1400 15861 1409 15895
rect 1409 15861 1443 15895
rect 1443 15861 1452 15895
rect 1400 15852 1452 15861
rect 1860 15895 1912 15904
rect 1860 15861 1869 15895
rect 1869 15861 1903 15895
rect 1903 15861 1912 15895
rect 1860 15852 1912 15861
rect 1952 15852 2004 15904
rect 2688 15852 2740 15904
rect 3240 15929 3249 15963
rect 3249 15929 3283 15963
rect 3283 15929 3292 15963
rect 3240 15920 3292 15929
rect 6092 15920 6144 15972
rect 7196 15920 7248 15972
rect 3700 15852 3752 15904
rect 5540 15852 5592 15904
rect 6276 15852 6328 15904
rect 7472 15852 7524 15904
rect 7656 15895 7708 15904
rect 7656 15861 7665 15895
rect 7665 15861 7699 15895
rect 7699 15861 7708 15895
rect 7656 15852 7708 15861
rect 9956 15920 10008 15972
rect 10876 15895 10928 15904
rect 10876 15861 10885 15895
rect 10885 15861 10919 15895
rect 10919 15861 10928 15895
rect 10876 15852 10928 15861
rect 12808 15852 12860 15904
rect 14372 15920 14424 15972
rect 15660 15920 15712 15972
rect 16212 15920 16264 15972
rect 18696 16065 18705 16099
rect 18705 16065 18739 16099
rect 18739 16065 18748 16099
rect 18696 16056 18748 16065
rect 21548 16124 21600 16176
rect 22744 16124 22796 16176
rect 22468 16099 22520 16108
rect 17592 15988 17644 16040
rect 18420 16031 18472 16040
rect 18420 15997 18429 16031
rect 18429 15997 18463 16031
rect 18463 15997 18472 16031
rect 18420 15988 18472 15997
rect 15936 15895 15988 15904
rect 15936 15861 15945 15895
rect 15945 15861 15979 15895
rect 15979 15861 15988 15895
rect 15936 15852 15988 15861
rect 17132 15852 17184 15904
rect 19064 15920 19116 15972
rect 22468 16065 22477 16099
rect 22477 16065 22511 16099
rect 22511 16065 22520 16099
rect 22468 16056 22520 16065
rect 23388 16201 23397 16235
rect 23397 16201 23431 16235
rect 23431 16201 23440 16235
rect 23388 16192 23440 16201
rect 23480 16192 23532 16244
rect 24676 16192 24728 16244
rect 23388 16056 23440 16108
rect 24032 16056 24084 16108
rect 24676 16056 24728 16108
rect 26056 16192 26108 16244
rect 26240 16235 26292 16244
rect 26240 16201 26249 16235
rect 26249 16201 26283 16235
rect 26283 16201 26292 16235
rect 26240 16192 26292 16201
rect 26332 16056 26384 16108
rect 23480 15988 23532 16040
rect 25228 16031 25280 16040
rect 25228 15997 25237 16031
rect 25237 15997 25271 16031
rect 25271 15997 25280 16031
rect 25228 15988 25280 15997
rect 22100 15920 22152 15972
rect 23572 15920 23624 15972
rect 18052 15895 18104 15904
rect 18052 15861 18061 15895
rect 18061 15861 18095 15895
rect 18095 15861 18104 15895
rect 18052 15852 18104 15861
rect 20996 15895 21048 15904
rect 20996 15861 21005 15895
rect 21005 15861 21039 15895
rect 21039 15861 21048 15895
rect 20996 15852 21048 15861
rect 22008 15852 22060 15904
rect 22192 15895 22244 15904
rect 22192 15861 22201 15895
rect 22201 15861 22235 15895
rect 22235 15861 22244 15895
rect 22192 15852 22244 15861
rect 23848 15852 23900 15904
rect 25044 15895 25096 15904
rect 25044 15861 25053 15895
rect 25053 15861 25087 15895
rect 25087 15861 25096 15895
rect 25044 15852 25096 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2136 15648 2188 15700
rect 5172 15648 5224 15700
rect 6184 15648 6236 15700
rect 6552 15691 6604 15700
rect 6552 15657 6561 15691
rect 6561 15657 6595 15691
rect 6595 15657 6604 15691
rect 6552 15648 6604 15657
rect 6920 15648 6972 15700
rect 9404 15691 9456 15700
rect 9404 15657 9413 15691
rect 9413 15657 9447 15691
rect 9447 15657 9456 15691
rect 9404 15648 9456 15657
rect 9680 15648 9732 15700
rect 12900 15648 12952 15700
rect 14372 15648 14424 15700
rect 14464 15648 14516 15700
rect 15476 15648 15528 15700
rect 15936 15648 15988 15700
rect 16212 15648 16264 15700
rect 22100 15648 22152 15700
rect 22192 15648 22244 15700
rect 23572 15691 23624 15700
rect 23572 15657 23581 15691
rect 23581 15657 23615 15691
rect 23615 15657 23624 15691
rect 23572 15648 23624 15657
rect 24032 15691 24084 15700
rect 24032 15657 24041 15691
rect 24041 15657 24075 15691
rect 24075 15657 24084 15691
rect 24032 15648 24084 15657
rect 25136 15648 25188 15700
rect 25320 15691 25372 15700
rect 25320 15657 25329 15691
rect 25329 15657 25363 15691
rect 25363 15657 25372 15691
rect 25320 15648 25372 15657
rect 4712 15580 4764 15632
rect 5632 15580 5684 15632
rect 8668 15580 8720 15632
rect 3516 15512 3568 15564
rect 4620 15555 4672 15564
rect 4620 15521 4654 15555
rect 4654 15521 4672 15555
rect 4620 15512 4672 15521
rect 8116 15555 8168 15564
rect 1676 15444 1728 15496
rect 1768 15308 1820 15360
rect 1952 15308 2004 15360
rect 3148 15376 3200 15428
rect 2964 15351 3016 15360
rect 2964 15317 2973 15351
rect 2973 15317 3007 15351
rect 3007 15317 3016 15351
rect 2964 15308 3016 15317
rect 3424 15351 3476 15360
rect 3424 15317 3433 15351
rect 3433 15317 3467 15351
rect 3467 15317 3476 15351
rect 3424 15308 3476 15317
rect 6092 15376 6144 15428
rect 7104 15487 7156 15496
rect 7104 15453 7113 15487
rect 7113 15453 7147 15487
rect 7147 15453 7156 15487
rect 8116 15521 8125 15555
rect 8125 15521 8159 15555
rect 8159 15521 8168 15555
rect 8116 15512 8168 15521
rect 10416 15580 10468 15632
rect 11060 15580 11112 15632
rect 13452 15580 13504 15632
rect 15844 15580 15896 15632
rect 11244 15555 11296 15564
rect 11244 15521 11253 15555
rect 11253 15521 11287 15555
rect 11287 15521 11296 15555
rect 11244 15512 11296 15521
rect 11612 15512 11664 15564
rect 13636 15512 13688 15564
rect 15292 15512 15344 15564
rect 15476 15512 15528 15564
rect 16212 15512 16264 15564
rect 16580 15512 16632 15564
rect 17868 15512 17920 15564
rect 7104 15444 7156 15453
rect 8208 15444 8260 15496
rect 11060 15444 11112 15496
rect 11428 15487 11480 15496
rect 11428 15453 11437 15487
rect 11437 15453 11471 15487
rect 11471 15453 11480 15487
rect 11428 15444 11480 15453
rect 11888 15444 11940 15496
rect 13912 15444 13964 15496
rect 14372 15376 14424 15428
rect 4528 15308 4580 15360
rect 6552 15308 6604 15360
rect 6828 15308 6880 15360
rect 7656 15351 7708 15360
rect 7656 15317 7665 15351
rect 7665 15317 7699 15351
rect 7699 15317 7708 15351
rect 7656 15308 7708 15317
rect 8392 15308 8444 15360
rect 10324 15351 10376 15360
rect 10324 15317 10333 15351
rect 10333 15317 10367 15351
rect 10367 15317 10376 15351
rect 10324 15308 10376 15317
rect 10692 15351 10744 15360
rect 10692 15317 10701 15351
rect 10701 15317 10735 15351
rect 10735 15317 10744 15351
rect 10692 15308 10744 15317
rect 11428 15308 11480 15360
rect 14832 15308 14884 15360
rect 15660 15376 15712 15428
rect 16396 15444 16448 15496
rect 17684 15487 17736 15496
rect 17684 15453 17693 15487
rect 17693 15453 17727 15487
rect 17727 15453 17736 15487
rect 17684 15444 17736 15453
rect 24676 15580 24728 15632
rect 18696 15512 18748 15564
rect 19156 15512 19208 15564
rect 20628 15512 20680 15564
rect 21180 15512 21232 15564
rect 22008 15512 22060 15564
rect 23940 15555 23992 15564
rect 23940 15521 23949 15555
rect 23949 15521 23983 15555
rect 23983 15521 23992 15555
rect 23940 15512 23992 15521
rect 25136 15555 25188 15564
rect 25136 15521 25145 15555
rect 25145 15521 25179 15555
rect 25179 15521 25188 15555
rect 25136 15512 25188 15521
rect 25320 15512 25372 15564
rect 18604 15487 18656 15496
rect 18604 15453 18613 15487
rect 18613 15453 18647 15487
rect 18647 15453 18656 15487
rect 18604 15444 18656 15453
rect 19984 15444 20036 15496
rect 20352 15444 20404 15496
rect 20536 15444 20588 15496
rect 17960 15376 18012 15428
rect 20076 15376 20128 15428
rect 22744 15419 22796 15428
rect 22744 15385 22753 15419
rect 22753 15385 22787 15419
rect 22787 15385 22796 15419
rect 22744 15376 22796 15385
rect 16948 15308 17000 15360
rect 20352 15308 20404 15360
rect 22928 15308 22980 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 4160 15104 4212 15156
rect 5540 15104 5592 15156
rect 6000 15104 6052 15156
rect 8300 15104 8352 15156
rect 8852 15104 8904 15156
rect 9956 15147 10008 15156
rect 9956 15113 9965 15147
rect 9965 15113 9999 15147
rect 9999 15113 10008 15147
rect 9956 15104 10008 15113
rect 11612 15104 11664 15156
rect 11888 15104 11940 15156
rect 13452 15147 13504 15156
rect 13452 15113 13461 15147
rect 13461 15113 13495 15147
rect 13495 15113 13504 15147
rect 13452 15104 13504 15113
rect 14096 15104 14148 15156
rect 15660 15104 15712 15156
rect 16580 15104 16632 15156
rect 17040 15104 17092 15156
rect 18420 15104 18472 15156
rect 19156 15147 19208 15156
rect 19156 15113 19165 15147
rect 19165 15113 19199 15147
rect 19199 15113 19208 15147
rect 19156 15104 19208 15113
rect 20168 15104 20220 15156
rect 21548 15104 21600 15156
rect 22008 15104 22060 15156
rect 22744 15147 22796 15156
rect 22744 15113 22753 15147
rect 22753 15113 22787 15147
rect 22787 15113 22796 15147
rect 22744 15104 22796 15113
rect 23296 15104 23348 15156
rect 24032 15104 24084 15156
rect 25136 15104 25188 15156
rect 1216 15036 1268 15088
rect 6092 15036 6144 15088
rect 2504 14968 2556 15020
rect 4528 15011 4580 15020
rect 4528 14977 4537 15011
rect 4537 14977 4571 15011
rect 4571 14977 4580 15011
rect 4528 14968 4580 14977
rect 2044 14900 2096 14952
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 4068 14900 4120 14952
rect 4804 14943 4856 14952
rect 3516 14832 3568 14884
rect 4804 14909 4838 14943
rect 4838 14909 4856 14943
rect 6920 14968 6972 15020
rect 11244 15036 11296 15088
rect 15844 15036 15896 15088
rect 16396 15079 16448 15088
rect 16396 15045 16405 15079
rect 16405 15045 16439 15079
rect 16439 15045 16448 15079
rect 16396 15036 16448 15045
rect 17868 15036 17920 15088
rect 19892 15036 19944 15088
rect 20628 15036 20680 15088
rect 21180 15079 21232 15088
rect 21180 15045 21189 15079
rect 21189 15045 21223 15079
rect 21223 15045 21232 15079
rect 21180 15036 21232 15045
rect 7472 14968 7524 15020
rect 10324 14968 10376 15020
rect 14372 15011 14424 15020
rect 14372 14977 14381 15011
rect 14381 14977 14415 15011
rect 14415 14977 14424 15011
rect 14372 14968 14424 14977
rect 14464 15011 14516 15020
rect 14464 14977 14473 15011
rect 14473 14977 14507 15011
rect 14507 14977 14516 15011
rect 14464 14968 14516 14977
rect 16212 14968 16264 15020
rect 16764 14968 16816 15020
rect 17132 14968 17184 15020
rect 17408 14968 17460 15020
rect 17684 14968 17736 15020
rect 4804 14900 4856 14909
rect 6828 14900 6880 14952
rect 8208 14900 8260 14952
rect 8484 14900 8536 14952
rect 11060 14943 11112 14952
rect 11060 14909 11069 14943
rect 11069 14909 11103 14943
rect 11103 14909 11112 14943
rect 11060 14900 11112 14909
rect 11244 14900 11296 14952
rect 13452 14900 13504 14952
rect 13912 14900 13964 14952
rect 7104 14832 7156 14884
rect 8852 14875 8904 14884
rect 8852 14841 8861 14875
rect 8861 14841 8895 14875
rect 8895 14841 8904 14875
rect 8852 14832 8904 14841
rect 10968 14832 11020 14884
rect 15844 14900 15896 14952
rect 18052 14900 18104 14952
rect 19432 14968 19484 15020
rect 22284 15036 22336 15088
rect 22652 15036 22704 15088
rect 23480 15079 23532 15088
rect 23480 15045 23489 15079
rect 23489 15045 23523 15079
rect 23523 15045 23532 15079
rect 23480 15036 23532 15045
rect 18880 14900 18932 14952
rect 20352 14900 20404 14952
rect 22652 14900 22704 14952
rect 23112 14900 23164 14952
rect 23664 14968 23716 15020
rect 24676 14968 24728 15020
rect 25228 14943 25280 14952
rect 25228 14909 25237 14943
rect 25237 14909 25271 14943
rect 25271 14909 25280 14943
rect 25228 14900 25280 14909
rect 16212 14832 16264 14884
rect 16764 14875 16816 14884
rect 16764 14841 16773 14875
rect 16773 14841 16807 14875
rect 16807 14841 16816 14875
rect 16764 14832 16816 14841
rect 17684 14832 17736 14884
rect 17960 14832 18012 14884
rect 20076 14875 20128 14884
rect 20076 14841 20085 14875
rect 20085 14841 20119 14875
rect 20119 14841 20128 14875
rect 20076 14832 20128 14841
rect 20168 14832 20220 14884
rect 23940 14832 23992 14884
rect 1676 14764 1728 14816
rect 1952 14807 2004 14816
rect 1952 14773 1961 14807
rect 1961 14773 1995 14807
rect 1995 14773 2004 14807
rect 1952 14764 2004 14773
rect 3240 14764 3292 14816
rect 4620 14764 4672 14816
rect 5264 14764 5316 14816
rect 5356 14764 5408 14816
rect 6184 14764 6236 14816
rect 11060 14764 11112 14816
rect 13452 14764 13504 14816
rect 14096 14764 14148 14816
rect 15292 14764 15344 14816
rect 17868 14764 17920 14816
rect 19984 14807 20036 14816
rect 19984 14773 19993 14807
rect 19993 14773 20027 14807
rect 20027 14773 20036 14807
rect 19984 14764 20036 14773
rect 20352 14764 20404 14816
rect 21548 14807 21600 14816
rect 21548 14773 21557 14807
rect 21557 14773 21591 14807
rect 21591 14773 21600 14807
rect 21548 14764 21600 14773
rect 23112 14807 23164 14816
rect 23112 14773 23121 14807
rect 23121 14773 23155 14807
rect 23155 14773 23164 14807
rect 23112 14764 23164 14773
rect 24308 14764 24360 14816
rect 26056 14764 26108 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2780 14603 2832 14612
rect 2780 14569 2789 14603
rect 2789 14569 2823 14603
rect 2823 14569 2832 14603
rect 2780 14560 2832 14569
rect 3516 14560 3568 14612
rect 6552 14560 6604 14612
rect 8852 14560 8904 14612
rect 9128 14560 9180 14612
rect 10140 14603 10192 14612
rect 1400 14492 1452 14544
rect 1768 14467 1820 14476
rect 1768 14433 1777 14467
rect 1777 14433 1811 14467
rect 1811 14433 1820 14467
rect 1768 14424 1820 14433
rect 4528 14492 4580 14544
rect 4712 14492 4764 14544
rect 6184 14492 6236 14544
rect 10140 14569 10149 14603
rect 10149 14569 10183 14603
rect 10183 14569 10192 14603
rect 10140 14560 10192 14569
rect 11152 14560 11204 14612
rect 12072 14560 12124 14612
rect 12808 14560 12860 14612
rect 12992 14560 13044 14612
rect 14464 14603 14516 14612
rect 14464 14569 14473 14603
rect 14473 14569 14507 14603
rect 14507 14569 14516 14603
rect 14464 14560 14516 14569
rect 15108 14603 15160 14612
rect 15108 14569 15117 14603
rect 15117 14569 15151 14603
rect 15151 14569 15160 14603
rect 15108 14560 15160 14569
rect 15660 14603 15712 14612
rect 15660 14569 15669 14603
rect 15669 14569 15703 14603
rect 15703 14569 15712 14603
rect 15660 14560 15712 14569
rect 17592 14560 17644 14612
rect 18880 14603 18932 14612
rect 18880 14569 18889 14603
rect 18889 14569 18923 14603
rect 18923 14569 18932 14603
rect 18880 14560 18932 14569
rect 19064 14560 19116 14612
rect 20076 14560 20128 14612
rect 20628 14603 20680 14612
rect 20628 14569 20637 14603
rect 20637 14569 20671 14603
rect 20671 14569 20680 14603
rect 20628 14560 20680 14569
rect 23940 14560 23992 14612
rect 24032 14560 24084 14612
rect 24216 14560 24268 14612
rect 24308 14560 24360 14612
rect 25044 14560 25096 14612
rect 10968 14492 11020 14544
rect 11888 14492 11940 14544
rect 13636 14492 13688 14544
rect 13912 14492 13964 14544
rect 15292 14492 15344 14544
rect 17132 14492 17184 14544
rect 17408 14535 17460 14544
rect 17408 14501 17442 14535
rect 17442 14501 17460 14535
rect 17408 14492 17460 14501
rect 4344 14467 4396 14476
rect 4344 14433 4378 14467
rect 4378 14433 4396 14467
rect 1860 14356 1912 14408
rect 3976 14356 4028 14408
rect 2780 14288 2832 14340
rect 4344 14424 4396 14433
rect 6644 14467 6696 14476
rect 6644 14433 6653 14467
rect 6653 14433 6687 14467
rect 6687 14433 6696 14467
rect 6644 14424 6696 14433
rect 9312 14424 9364 14476
rect 11612 14467 11664 14476
rect 11612 14433 11621 14467
rect 11621 14433 11655 14467
rect 11655 14433 11664 14467
rect 11612 14424 11664 14433
rect 6552 14356 6604 14408
rect 8116 14356 8168 14408
rect 7748 14288 7800 14340
rect 9956 14288 10008 14340
rect 11428 14356 11480 14408
rect 11888 14399 11940 14408
rect 11888 14365 11897 14399
rect 11897 14365 11931 14399
rect 11931 14365 11940 14399
rect 11888 14356 11940 14365
rect 13452 14424 13504 14476
rect 16672 14424 16724 14476
rect 16856 14424 16908 14476
rect 17040 14467 17092 14476
rect 17040 14433 17049 14467
rect 17049 14433 17083 14467
rect 17083 14433 17092 14467
rect 17040 14424 17092 14433
rect 18696 14424 18748 14476
rect 19248 14424 19300 14476
rect 13084 14356 13136 14408
rect 14464 14356 14516 14408
rect 19340 14399 19392 14408
rect 1400 14263 1452 14272
rect 1400 14229 1409 14263
rect 1409 14229 1443 14263
rect 1443 14229 1452 14263
rect 1400 14220 1452 14229
rect 1860 14220 1912 14272
rect 2504 14220 2556 14272
rect 5264 14220 5316 14272
rect 8024 14220 8076 14272
rect 8944 14263 8996 14272
rect 8944 14229 8953 14263
rect 8953 14229 8987 14263
rect 8987 14229 8996 14263
rect 8944 14220 8996 14229
rect 9588 14220 9640 14272
rect 10876 14263 10928 14272
rect 10876 14229 10885 14263
rect 10885 14229 10919 14263
rect 10919 14229 10928 14263
rect 10876 14220 10928 14229
rect 11244 14263 11296 14272
rect 11244 14229 11253 14263
rect 11253 14229 11287 14263
rect 11287 14229 11296 14263
rect 11244 14220 11296 14229
rect 12808 14263 12860 14272
rect 12808 14229 12817 14263
rect 12817 14229 12851 14263
rect 12851 14229 12860 14263
rect 12808 14220 12860 14229
rect 13636 14220 13688 14272
rect 15108 14288 15160 14340
rect 15292 14331 15344 14340
rect 15292 14297 15301 14331
rect 15301 14297 15335 14331
rect 15335 14297 15344 14331
rect 15292 14288 15344 14297
rect 19340 14365 19349 14399
rect 19349 14365 19383 14399
rect 19383 14365 19392 14399
rect 19340 14356 19392 14365
rect 19714 14467 19766 14476
rect 19714 14433 19742 14467
rect 19742 14433 19766 14467
rect 19714 14424 19766 14433
rect 23664 14492 23716 14544
rect 25320 14492 25372 14544
rect 21180 14424 21232 14476
rect 24216 14467 24268 14476
rect 24216 14433 24225 14467
rect 24225 14433 24259 14467
rect 24259 14433 24268 14467
rect 24216 14424 24268 14433
rect 24768 14424 24820 14476
rect 25044 14424 25096 14476
rect 25596 14424 25648 14476
rect 19984 14356 20036 14408
rect 20168 14356 20220 14408
rect 20536 14356 20588 14408
rect 21640 14399 21692 14408
rect 21640 14365 21649 14399
rect 21649 14365 21683 14399
rect 21683 14365 21692 14399
rect 21640 14356 21692 14365
rect 20444 14288 20496 14340
rect 18052 14220 18104 14272
rect 18604 14220 18656 14272
rect 19248 14220 19300 14272
rect 23112 14356 23164 14408
rect 24676 14356 24728 14408
rect 21180 14263 21232 14272
rect 21180 14229 21189 14263
rect 21189 14229 21223 14263
rect 21223 14229 21232 14263
rect 21180 14220 21232 14229
rect 21548 14263 21600 14272
rect 21548 14229 21557 14263
rect 21557 14229 21591 14263
rect 21591 14229 21600 14263
rect 21548 14220 21600 14229
rect 22008 14220 22060 14272
rect 23388 14220 23440 14272
rect 23848 14220 23900 14272
rect 24676 14220 24728 14272
rect 25228 14263 25280 14272
rect 25228 14229 25237 14263
rect 25237 14229 25271 14263
rect 25271 14229 25280 14263
rect 25228 14220 25280 14229
rect 26056 14220 26108 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 4804 14059 4856 14068
rect 4804 14025 4813 14059
rect 4813 14025 4847 14059
rect 4847 14025 4856 14059
rect 4804 14016 4856 14025
rect 5448 14016 5500 14068
rect 6184 14059 6236 14068
rect 6184 14025 6193 14059
rect 6193 14025 6227 14059
rect 6227 14025 6236 14059
rect 6184 14016 6236 14025
rect 6828 14059 6880 14068
rect 6828 14025 6837 14059
rect 6837 14025 6871 14059
rect 6871 14025 6880 14059
rect 6828 14016 6880 14025
rect 8852 14016 8904 14068
rect 10140 14016 10192 14068
rect 11888 14059 11940 14068
rect 2320 13948 2372 14000
rect 2780 13948 2832 14000
rect 1676 13923 1728 13932
rect 1676 13889 1685 13923
rect 1685 13889 1719 13923
rect 1719 13889 1728 13923
rect 1676 13880 1728 13889
rect 1768 13812 1820 13864
rect 2780 13855 2832 13864
rect 2780 13821 2789 13855
rect 2789 13821 2823 13855
rect 2823 13821 2832 13855
rect 7104 13880 7156 13932
rect 8024 13880 8076 13932
rect 2780 13812 2832 13821
rect 4344 13812 4396 13864
rect 2136 13744 2188 13796
rect 2872 13744 2924 13796
rect 6000 13744 6052 13796
rect 6828 13812 6880 13864
rect 8576 13855 8628 13864
rect 8576 13821 8585 13855
rect 8585 13821 8619 13855
rect 8619 13821 8628 13855
rect 8576 13812 8628 13821
rect 9956 13812 10008 13864
rect 11888 14025 11897 14059
rect 11897 14025 11931 14059
rect 11931 14025 11940 14059
rect 11888 14016 11940 14025
rect 12072 14016 12124 14068
rect 12348 14016 12400 14068
rect 12624 14016 12676 14068
rect 13636 14059 13688 14068
rect 13636 14025 13645 14059
rect 13645 14025 13679 14059
rect 13679 14025 13688 14059
rect 13636 14016 13688 14025
rect 14648 14016 14700 14068
rect 15660 14059 15712 14068
rect 15660 14025 15669 14059
rect 15669 14025 15703 14059
rect 15703 14025 15712 14059
rect 15660 14016 15712 14025
rect 16396 14059 16448 14068
rect 16396 14025 16405 14059
rect 16405 14025 16439 14059
rect 16439 14025 16448 14059
rect 16396 14016 16448 14025
rect 17408 14059 17460 14068
rect 17408 14025 17417 14059
rect 17417 14025 17451 14059
rect 17451 14025 17460 14059
rect 17408 14016 17460 14025
rect 19432 14059 19484 14068
rect 19432 14025 19441 14059
rect 19441 14025 19475 14059
rect 19475 14025 19484 14059
rect 19432 14016 19484 14025
rect 19708 14059 19760 14068
rect 19708 14025 19717 14059
rect 19717 14025 19751 14059
rect 19751 14025 19760 14059
rect 19708 14016 19760 14025
rect 20352 14016 20404 14068
rect 20720 14016 20772 14068
rect 20904 14059 20956 14068
rect 20904 14025 20913 14059
rect 20913 14025 20947 14059
rect 20947 14025 20956 14059
rect 20904 14016 20956 14025
rect 22744 14016 22796 14068
rect 23020 14059 23072 14068
rect 23020 14025 23029 14059
rect 23029 14025 23063 14059
rect 23063 14025 23072 14059
rect 23020 14016 23072 14025
rect 23664 14059 23716 14068
rect 23664 14025 23673 14059
rect 23673 14025 23707 14059
rect 23707 14025 23716 14059
rect 23664 14016 23716 14025
rect 24216 14016 24268 14068
rect 10968 13948 11020 14000
rect 11152 13948 11204 14000
rect 13452 13991 13504 14000
rect 10876 13880 10928 13932
rect 12072 13880 12124 13932
rect 8760 13744 8812 13796
rect 9404 13744 9456 13796
rect 9680 13744 9732 13796
rect 10784 13812 10836 13864
rect 13452 13957 13461 13991
rect 13461 13957 13495 13991
rect 13495 13957 13504 13991
rect 13452 13948 13504 13957
rect 13912 13948 13964 14000
rect 21180 13948 21232 14000
rect 12900 13923 12952 13932
rect 12900 13889 12909 13923
rect 12909 13889 12943 13923
rect 12943 13889 12952 13923
rect 12900 13880 12952 13889
rect 12992 13923 13044 13932
rect 12992 13889 13001 13923
rect 13001 13889 13035 13923
rect 13035 13889 13044 13923
rect 14648 13923 14700 13932
rect 12992 13880 13044 13889
rect 14648 13889 14657 13923
rect 14657 13889 14691 13923
rect 14691 13889 14700 13923
rect 14648 13880 14700 13889
rect 17132 13880 17184 13932
rect 22928 13948 22980 14000
rect 10876 13744 10928 13796
rect 11336 13744 11388 13796
rect 14464 13855 14516 13864
rect 14464 13821 14473 13855
rect 14473 13821 14507 13855
rect 14507 13821 14516 13855
rect 14464 13812 14516 13821
rect 16856 13855 16908 13864
rect 16856 13821 16865 13855
rect 16865 13821 16899 13855
rect 16899 13821 16908 13855
rect 16856 13812 16908 13821
rect 17868 13812 17920 13864
rect 18052 13855 18104 13864
rect 18052 13821 18061 13855
rect 18061 13821 18095 13855
rect 18095 13821 18104 13855
rect 18052 13812 18104 13821
rect 18604 13812 18656 13864
rect 20720 13855 20772 13864
rect 20720 13821 20729 13855
rect 20729 13821 20763 13855
rect 20763 13821 20772 13855
rect 20720 13812 20772 13821
rect 21824 13812 21876 13864
rect 23020 13812 23072 13864
rect 1860 13676 1912 13728
rect 5356 13719 5408 13728
rect 5356 13685 5365 13719
rect 5365 13685 5399 13719
rect 5399 13685 5408 13719
rect 5356 13676 5408 13685
rect 5540 13676 5592 13728
rect 8576 13676 8628 13728
rect 11244 13676 11296 13728
rect 12808 13719 12860 13728
rect 12808 13685 12817 13719
rect 12817 13685 12851 13719
rect 12851 13685 12860 13719
rect 12808 13676 12860 13685
rect 12900 13676 12952 13728
rect 16396 13744 16448 13796
rect 16672 13744 16724 13796
rect 16948 13744 17000 13796
rect 17132 13744 17184 13796
rect 23296 13744 23348 13796
rect 25136 13880 25188 13932
rect 25228 13855 25280 13864
rect 25228 13821 25237 13855
rect 25237 13821 25271 13855
rect 25271 13821 25280 13855
rect 25228 13812 25280 13821
rect 18696 13676 18748 13728
rect 22192 13676 22244 13728
rect 22744 13676 22796 13728
rect 23940 13676 23992 13728
rect 26056 13676 26108 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 3148 13472 3200 13524
rect 4160 13472 4212 13524
rect 5632 13472 5684 13524
rect 6828 13472 6880 13524
rect 2596 13404 2648 13456
rect 2780 13447 2832 13456
rect 2780 13413 2789 13447
rect 2789 13413 2823 13447
rect 2823 13413 2832 13447
rect 7012 13472 7064 13524
rect 8024 13515 8076 13524
rect 8024 13481 8033 13515
rect 8033 13481 8067 13515
rect 8067 13481 8076 13515
rect 8024 13472 8076 13481
rect 8668 13472 8720 13524
rect 9772 13472 9824 13524
rect 10784 13472 10836 13524
rect 11336 13472 11388 13524
rect 12256 13472 12308 13524
rect 12440 13472 12492 13524
rect 12808 13472 12860 13524
rect 2780 13404 2832 13413
rect 3148 13336 3200 13388
rect 3884 13336 3936 13388
rect 3976 13336 4028 13388
rect 3516 13311 3568 13320
rect 1768 13132 1820 13184
rect 2044 13132 2096 13184
rect 3516 13277 3525 13311
rect 3525 13277 3559 13311
rect 3559 13277 3568 13311
rect 3516 13268 3568 13277
rect 4528 13311 4580 13320
rect 4528 13277 4537 13311
rect 4537 13277 4571 13311
rect 4571 13277 4580 13311
rect 4528 13268 4580 13277
rect 5264 13336 5316 13388
rect 6460 13268 6512 13320
rect 8300 13404 8352 13456
rect 9588 13404 9640 13456
rect 11520 13404 11572 13456
rect 11704 13447 11756 13456
rect 11704 13413 11716 13447
rect 11716 13413 11756 13447
rect 13084 13447 13136 13456
rect 11704 13404 11756 13413
rect 13084 13413 13093 13447
rect 13093 13413 13127 13447
rect 13127 13413 13136 13447
rect 13084 13404 13136 13413
rect 13452 13447 13504 13456
rect 13452 13413 13461 13447
rect 13461 13413 13495 13447
rect 13495 13413 13504 13447
rect 13452 13404 13504 13413
rect 14096 13404 14148 13456
rect 14280 13404 14332 13456
rect 15936 13472 15988 13524
rect 16856 13472 16908 13524
rect 17040 13472 17092 13524
rect 17408 13472 17460 13524
rect 17592 13472 17644 13524
rect 19984 13472 20036 13524
rect 6736 13336 6788 13388
rect 9128 13336 9180 13388
rect 9496 13336 9548 13388
rect 9680 13336 9732 13388
rect 10324 13336 10376 13388
rect 11244 13336 11296 13388
rect 12440 13336 12492 13388
rect 13912 13336 13964 13388
rect 17960 13404 18012 13456
rect 19432 13404 19484 13456
rect 16396 13336 16448 13388
rect 17132 13336 17184 13388
rect 18052 13336 18104 13388
rect 19248 13336 19300 13388
rect 19340 13336 19392 13388
rect 22008 13472 22060 13524
rect 22928 13472 22980 13524
rect 25964 13472 26016 13524
rect 20996 13404 21048 13456
rect 21640 13404 21692 13456
rect 22468 13404 22520 13456
rect 23296 13404 23348 13456
rect 21548 13336 21600 13388
rect 23112 13336 23164 13388
rect 26056 13404 26108 13456
rect 23480 13379 23532 13388
rect 23480 13345 23514 13379
rect 23514 13345 23532 13379
rect 23480 13336 23532 13345
rect 24032 13336 24084 13388
rect 5356 13200 5408 13252
rect 6000 13200 6052 13252
rect 7472 13268 7524 13320
rect 3240 13132 3292 13184
rect 3516 13132 3568 13184
rect 5540 13132 5592 13184
rect 7472 13175 7524 13184
rect 7472 13141 7481 13175
rect 7481 13141 7515 13175
rect 7515 13141 7524 13175
rect 7472 13132 7524 13141
rect 7932 13175 7984 13184
rect 7932 13141 7941 13175
rect 7941 13141 7975 13175
rect 7975 13141 7984 13175
rect 7932 13132 7984 13141
rect 9956 13200 10008 13252
rect 13820 13268 13872 13320
rect 14556 13268 14608 13320
rect 14648 13268 14700 13320
rect 15292 13311 15344 13320
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 15292 13268 15344 13277
rect 10876 13200 10928 13252
rect 12808 13243 12860 13252
rect 8852 13132 8904 13184
rect 9128 13175 9180 13184
rect 9128 13141 9137 13175
rect 9137 13141 9171 13175
rect 9171 13141 9180 13175
rect 9128 13132 9180 13141
rect 9496 13132 9548 13184
rect 11244 13175 11296 13184
rect 11244 13141 11253 13175
rect 11253 13141 11287 13175
rect 11287 13141 11296 13175
rect 11244 13132 11296 13141
rect 12808 13209 12817 13243
rect 12817 13209 12851 13243
rect 12851 13209 12860 13243
rect 12808 13200 12860 13209
rect 13728 13200 13780 13252
rect 18236 13268 18288 13320
rect 22192 13268 22244 13320
rect 16856 13200 16908 13252
rect 17592 13200 17644 13252
rect 21364 13200 21416 13252
rect 17224 13132 17276 13184
rect 18880 13132 18932 13184
rect 20444 13132 20496 13184
rect 20720 13175 20772 13184
rect 20720 13141 20729 13175
rect 20729 13141 20763 13175
rect 20763 13141 20772 13175
rect 20720 13132 20772 13141
rect 24768 13268 24820 13320
rect 22928 13132 22980 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2964 12928 3016 12980
rect 5540 12928 5592 12980
rect 6000 12928 6052 12980
rect 6736 12928 6788 12980
rect 9036 12971 9088 12980
rect 9036 12937 9045 12971
rect 9045 12937 9079 12971
rect 9079 12937 9088 12971
rect 9036 12928 9088 12937
rect 9772 12928 9824 12980
rect 10140 12928 10192 12980
rect 13360 12928 13412 12980
rect 13636 12928 13688 12980
rect 14556 12928 14608 12980
rect 15752 12928 15804 12980
rect 16948 12928 17000 12980
rect 17132 12928 17184 12980
rect 17684 12928 17736 12980
rect 19432 12971 19484 12980
rect 19432 12937 19441 12971
rect 19441 12937 19475 12971
rect 19475 12937 19484 12971
rect 19432 12928 19484 12937
rect 20260 12971 20312 12980
rect 20260 12937 20269 12971
rect 20269 12937 20303 12971
rect 20303 12937 20312 12971
rect 20260 12928 20312 12937
rect 21180 12971 21232 12980
rect 21180 12937 21189 12971
rect 21189 12937 21223 12971
rect 21223 12937 21232 12971
rect 21180 12928 21232 12937
rect 21916 12928 21968 12980
rect 1124 12860 1176 12912
rect 2780 12860 2832 12912
rect 4068 12860 4120 12912
rect 6460 12903 6512 12912
rect 6460 12869 6469 12903
rect 6469 12869 6503 12903
rect 6503 12869 6512 12903
rect 6460 12860 6512 12869
rect 9128 12860 9180 12912
rect 2136 12835 2188 12844
rect 2136 12801 2145 12835
rect 2145 12801 2179 12835
rect 2179 12801 2188 12835
rect 2136 12792 2188 12801
rect 3424 12792 3476 12844
rect 3792 12835 3844 12844
rect 3792 12801 3801 12835
rect 3801 12801 3835 12835
rect 3835 12801 3844 12835
rect 3792 12792 3844 12801
rect 1216 12724 1268 12776
rect 2596 12724 2648 12776
rect 3516 12767 3568 12776
rect 3516 12733 3525 12767
rect 3525 12733 3559 12767
rect 3559 12733 3568 12767
rect 3516 12724 3568 12733
rect 1400 12588 1452 12640
rect 2504 12588 2556 12640
rect 2780 12588 2832 12640
rect 3148 12588 3200 12640
rect 5172 12835 5224 12844
rect 5172 12801 5181 12835
rect 5181 12801 5215 12835
rect 5215 12801 5224 12835
rect 5172 12792 5224 12801
rect 5264 12835 5316 12844
rect 5264 12801 5273 12835
rect 5273 12801 5307 12835
rect 5307 12801 5316 12835
rect 5264 12792 5316 12801
rect 6552 12792 6604 12844
rect 7932 12792 7984 12844
rect 10048 12860 10100 12912
rect 16212 12860 16264 12912
rect 4712 12724 4764 12776
rect 5080 12767 5132 12776
rect 5080 12733 5089 12767
rect 5089 12733 5123 12767
rect 5123 12733 5132 12767
rect 5080 12724 5132 12733
rect 9128 12724 9180 12776
rect 9404 12767 9456 12776
rect 9404 12733 9413 12767
rect 9413 12733 9447 12767
rect 9447 12733 9456 12767
rect 9404 12724 9456 12733
rect 9680 12724 9732 12776
rect 10324 12792 10376 12844
rect 10692 12792 10744 12844
rect 11244 12835 11296 12844
rect 11244 12801 11253 12835
rect 11253 12801 11287 12835
rect 11287 12801 11296 12835
rect 11244 12792 11296 12801
rect 11704 12792 11756 12844
rect 12440 12835 12492 12844
rect 12440 12801 12449 12835
rect 12449 12801 12483 12835
rect 12483 12801 12492 12835
rect 12440 12792 12492 12801
rect 16580 12792 16632 12844
rect 4528 12656 4580 12708
rect 5264 12656 5316 12708
rect 5356 12656 5408 12708
rect 7472 12656 7524 12708
rect 9864 12656 9916 12708
rect 10232 12656 10284 12708
rect 11152 12656 11204 12708
rect 11612 12724 11664 12776
rect 11980 12724 12032 12776
rect 13820 12724 13872 12776
rect 15292 12724 15344 12776
rect 16396 12724 16448 12776
rect 18880 12835 18932 12844
rect 18880 12801 18889 12835
rect 18889 12801 18923 12835
rect 18923 12801 18932 12835
rect 18880 12792 18932 12801
rect 19064 12835 19116 12844
rect 19064 12801 19073 12835
rect 19073 12801 19107 12835
rect 19107 12801 19116 12835
rect 19064 12792 19116 12801
rect 20168 12860 20220 12912
rect 22928 12928 22980 12980
rect 23480 12928 23532 12980
rect 25320 12971 25372 12980
rect 25320 12937 25329 12971
rect 25329 12937 25363 12971
rect 25363 12937 25372 12971
rect 25320 12928 25372 12937
rect 26056 12971 26108 12980
rect 26056 12937 26065 12971
rect 26065 12937 26099 12971
rect 26099 12937 26108 12971
rect 26056 12928 26108 12937
rect 23020 12792 23072 12844
rect 21640 12767 21692 12776
rect 21640 12733 21649 12767
rect 21649 12733 21683 12767
rect 21683 12733 21692 12767
rect 21640 12724 21692 12733
rect 23112 12724 23164 12776
rect 12808 12656 12860 12708
rect 6552 12588 6604 12640
rect 8024 12588 8076 12640
rect 8852 12588 8904 12640
rect 10876 12588 10928 12640
rect 11520 12588 11572 12640
rect 11980 12588 12032 12640
rect 14924 12699 14976 12708
rect 14924 12665 14958 12699
rect 14958 12665 14976 12699
rect 14924 12656 14976 12665
rect 16580 12656 16632 12708
rect 16672 12656 16724 12708
rect 16948 12656 17000 12708
rect 17684 12656 17736 12708
rect 18420 12656 18472 12708
rect 20996 12699 21048 12708
rect 20996 12665 21005 12699
rect 21005 12665 21039 12699
rect 21039 12665 21048 12699
rect 20996 12656 21048 12665
rect 22652 12656 22704 12708
rect 23020 12656 23072 12708
rect 23296 12656 23348 12708
rect 23572 12656 23624 12708
rect 23848 12656 23900 12708
rect 14464 12588 14516 12640
rect 16212 12588 16264 12640
rect 16396 12588 16448 12640
rect 17316 12588 17368 12640
rect 22468 12588 22520 12640
rect 22836 12588 22888 12640
rect 24768 12588 24820 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1124 12384 1176 12436
rect 3792 12384 3844 12436
rect 3976 12384 4028 12436
rect 4160 12384 4212 12436
rect 4344 12384 4396 12436
rect 5540 12384 5592 12436
rect 8300 12427 8352 12436
rect 8300 12393 8309 12427
rect 8309 12393 8343 12427
rect 8343 12393 8352 12427
rect 8300 12384 8352 12393
rect 8668 12427 8720 12436
rect 8668 12393 8677 12427
rect 8677 12393 8711 12427
rect 8711 12393 8720 12427
rect 8668 12384 8720 12393
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 9864 12384 9916 12436
rect 10784 12384 10836 12436
rect 12256 12384 12308 12436
rect 14096 12384 14148 12436
rect 15844 12384 15896 12436
rect 16212 12384 16264 12436
rect 16580 12384 16632 12436
rect 16948 12427 17000 12436
rect 16948 12393 16957 12427
rect 16957 12393 16991 12427
rect 16991 12393 17000 12427
rect 16948 12384 17000 12393
rect 17316 12427 17368 12436
rect 17316 12393 17325 12427
rect 17325 12393 17359 12427
rect 17359 12393 17368 12427
rect 17316 12384 17368 12393
rect 19064 12384 19116 12436
rect 19156 12384 19208 12436
rect 20996 12384 21048 12436
rect 22284 12384 22336 12436
rect 22468 12384 22520 12436
rect 23848 12384 23900 12436
rect 24124 12427 24176 12436
rect 24124 12393 24133 12427
rect 24133 12393 24167 12427
rect 24167 12393 24176 12427
rect 24124 12384 24176 12393
rect 25412 12384 25464 12436
rect 26056 12427 26108 12436
rect 26056 12393 26065 12427
rect 26065 12393 26099 12427
rect 26099 12393 26108 12427
rect 26056 12384 26108 12393
rect 1400 12316 1452 12368
rect 2320 12316 2372 12368
rect 4712 12359 4764 12368
rect 4712 12325 4721 12359
rect 4721 12325 4755 12359
rect 4755 12325 4764 12359
rect 4712 12316 4764 12325
rect 6552 12316 6604 12368
rect 9588 12316 9640 12368
rect 14004 12316 14056 12368
rect 1860 12248 1912 12300
rect 4160 12248 4212 12300
rect 6184 12248 6236 12300
rect 10324 12248 10376 12300
rect 11520 12291 11572 12300
rect 11520 12257 11529 12291
rect 11529 12257 11563 12291
rect 11563 12257 11572 12291
rect 11520 12248 11572 12257
rect 15292 12291 15344 12300
rect 15292 12257 15301 12291
rect 15301 12257 15335 12291
rect 15335 12257 15344 12291
rect 15292 12248 15344 12257
rect 15752 12316 15804 12368
rect 17040 12316 17092 12368
rect 20812 12316 20864 12368
rect 21916 12316 21968 12368
rect 22652 12316 22704 12368
rect 24952 12316 25004 12368
rect 17500 12291 17552 12300
rect 17500 12257 17509 12291
rect 17509 12257 17543 12291
rect 17543 12257 17552 12291
rect 17500 12248 17552 12257
rect 20904 12291 20956 12300
rect 20904 12257 20913 12291
rect 20913 12257 20947 12291
rect 20947 12257 20956 12291
rect 20904 12248 20956 12257
rect 23020 12248 23072 12300
rect 23388 12248 23440 12300
rect 23848 12248 23900 12300
rect 25228 12248 25280 12300
rect 5448 12223 5500 12232
rect 5448 12189 5457 12223
rect 5457 12189 5491 12223
rect 5491 12189 5500 12223
rect 5448 12180 5500 12189
rect 5080 12112 5132 12164
rect 6460 12180 6512 12232
rect 9956 12180 10008 12232
rect 10508 12180 10560 12232
rect 10784 12180 10836 12232
rect 10968 12180 11020 12232
rect 11336 12180 11388 12232
rect 11704 12223 11756 12232
rect 11704 12189 11713 12223
rect 11713 12189 11747 12223
rect 11747 12189 11756 12223
rect 14464 12223 14516 12232
rect 11704 12180 11756 12189
rect 14464 12189 14473 12223
rect 14473 12189 14507 12223
rect 14507 12189 14516 12223
rect 14464 12180 14516 12189
rect 16580 12180 16632 12232
rect 17592 12180 17644 12232
rect 17776 12180 17828 12232
rect 19340 12180 19392 12232
rect 21916 12180 21968 12232
rect 9680 12112 9732 12164
rect 10140 12112 10192 12164
rect 12256 12112 12308 12164
rect 20260 12155 20312 12164
rect 20260 12121 20269 12155
rect 20269 12121 20303 12155
rect 20303 12121 20312 12155
rect 20260 12112 20312 12121
rect 21088 12155 21140 12164
rect 21088 12121 21097 12155
rect 21097 12121 21131 12155
rect 21131 12121 21140 12155
rect 21088 12112 21140 12121
rect 6092 12087 6144 12096
rect 6092 12053 6101 12087
rect 6101 12053 6135 12087
rect 6135 12053 6144 12087
rect 6092 12044 6144 12053
rect 7932 12087 7984 12096
rect 7932 12053 7941 12087
rect 7941 12053 7975 12087
rect 7975 12053 7984 12087
rect 7932 12044 7984 12053
rect 9404 12044 9456 12096
rect 9956 12044 10008 12096
rect 10692 12087 10744 12096
rect 10692 12053 10701 12087
rect 10701 12053 10735 12087
rect 10735 12053 10744 12087
rect 10692 12044 10744 12053
rect 10784 12044 10836 12096
rect 12532 12087 12584 12096
rect 12532 12053 12541 12087
rect 12541 12053 12575 12087
rect 12575 12053 12584 12087
rect 12532 12044 12584 12053
rect 15292 12044 15344 12096
rect 16396 12044 16448 12096
rect 17592 12044 17644 12096
rect 17960 12044 18012 12096
rect 19984 12044 20036 12096
rect 21640 12087 21692 12096
rect 21640 12053 21649 12087
rect 21649 12053 21683 12087
rect 21683 12053 21692 12087
rect 21640 12044 21692 12053
rect 22008 12044 22060 12096
rect 23940 12044 23992 12096
rect 24676 12044 24728 12096
rect 25596 12087 25648 12096
rect 25596 12053 25605 12087
rect 25605 12053 25639 12087
rect 25639 12053 25648 12087
rect 25596 12044 25648 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2320 11840 2372 11892
rect 2504 11840 2556 11892
rect 5448 11840 5500 11892
rect 6184 11883 6236 11892
rect 6184 11849 6193 11883
rect 6193 11849 6227 11883
rect 6227 11849 6236 11883
rect 6184 11840 6236 11849
rect 6552 11883 6604 11892
rect 6552 11849 6561 11883
rect 6561 11849 6595 11883
rect 6595 11849 6604 11883
rect 6552 11840 6604 11849
rect 7564 11883 7616 11892
rect 7564 11849 7573 11883
rect 7573 11849 7607 11883
rect 7607 11849 7616 11883
rect 7564 11840 7616 11849
rect 9864 11840 9916 11892
rect 10232 11883 10284 11892
rect 10232 11849 10241 11883
rect 10241 11849 10275 11883
rect 10275 11849 10284 11883
rect 10232 11840 10284 11849
rect 10600 11840 10652 11892
rect 11244 11840 11296 11892
rect 13084 11840 13136 11892
rect 13544 11840 13596 11892
rect 13728 11840 13780 11892
rect 16396 11883 16448 11892
rect 16396 11849 16405 11883
rect 16405 11849 16439 11883
rect 16439 11849 16448 11883
rect 16396 11840 16448 11849
rect 17500 11883 17552 11892
rect 17500 11849 17509 11883
rect 17509 11849 17543 11883
rect 17543 11849 17552 11883
rect 17500 11840 17552 11849
rect 20628 11840 20680 11892
rect 21824 11883 21876 11892
rect 21824 11849 21833 11883
rect 21833 11849 21867 11883
rect 21867 11849 21876 11883
rect 21824 11840 21876 11849
rect 23204 11840 23256 11892
rect 23572 11840 23624 11892
rect 24676 11883 24728 11892
rect 24676 11849 24685 11883
rect 24685 11849 24719 11883
rect 24719 11849 24728 11883
rect 24676 11840 24728 11849
rect 26424 11840 26476 11892
rect 5080 11815 5132 11824
rect 5080 11781 5089 11815
rect 5089 11781 5123 11815
rect 5123 11781 5132 11815
rect 5080 11772 5132 11781
rect 7932 11772 7984 11824
rect 9128 11772 9180 11824
rect 9956 11772 10008 11824
rect 10692 11772 10744 11824
rect 14556 11815 14608 11824
rect 6184 11704 6236 11756
rect 6460 11704 6512 11756
rect 9864 11704 9916 11756
rect 10508 11704 10560 11756
rect 14556 11781 14565 11815
rect 14565 11781 14599 11815
rect 14599 11781 14608 11815
rect 14556 11772 14608 11781
rect 25228 11772 25280 11824
rect 10968 11704 11020 11756
rect 12440 11747 12492 11756
rect 12440 11713 12449 11747
rect 12449 11713 12483 11747
rect 12483 11713 12492 11747
rect 12440 11704 12492 11713
rect 13820 11704 13872 11756
rect 16948 11747 17000 11756
rect 16948 11713 16957 11747
rect 16957 11713 16991 11747
rect 16991 11713 17000 11747
rect 16948 11704 17000 11713
rect 17960 11704 18012 11756
rect 6092 11636 6144 11688
rect 7932 11636 7984 11688
rect 11704 11636 11756 11688
rect 13268 11636 13320 11688
rect 13912 11636 13964 11688
rect 14556 11636 14608 11688
rect 20260 11704 20312 11756
rect 2136 11568 2188 11620
rect 2688 11568 2740 11620
rect 5540 11611 5592 11620
rect 5540 11577 5549 11611
rect 5549 11577 5583 11611
rect 5583 11577 5592 11611
rect 5540 11568 5592 11577
rect 10324 11568 10376 11620
rect 12532 11568 12584 11620
rect 13544 11568 13596 11620
rect 15200 11568 15252 11620
rect 17960 11568 18012 11620
rect 19524 11636 19576 11688
rect 20628 11636 20680 11688
rect 22008 11704 22060 11756
rect 22836 11704 22888 11756
rect 23020 11704 23072 11756
rect 24124 11747 24176 11756
rect 24124 11713 24133 11747
rect 24133 11713 24167 11747
rect 24167 11713 24176 11747
rect 24124 11704 24176 11713
rect 23204 11636 23256 11688
rect 25872 11704 25924 11756
rect 25412 11636 25464 11688
rect 19340 11568 19392 11620
rect 21732 11568 21784 11620
rect 22836 11568 22888 11620
rect 24216 11568 24268 11620
rect 24860 11568 24912 11620
rect 1860 11500 1912 11552
rect 2964 11500 3016 11552
rect 3516 11543 3568 11552
rect 3516 11509 3525 11543
rect 3525 11509 3559 11543
rect 3559 11509 3568 11543
rect 3516 11500 3568 11509
rect 5172 11543 5224 11552
rect 5172 11509 5181 11543
rect 5181 11509 5215 11543
rect 5215 11509 5224 11543
rect 5172 11500 5224 11509
rect 6828 11543 6880 11552
rect 6828 11509 6837 11543
rect 6837 11509 6871 11543
rect 6871 11509 6880 11543
rect 6828 11500 6880 11509
rect 9496 11500 9548 11552
rect 10140 11500 10192 11552
rect 10876 11500 10928 11552
rect 11244 11543 11296 11552
rect 11244 11509 11253 11543
rect 11253 11509 11287 11543
rect 11287 11509 11296 11543
rect 11244 11500 11296 11509
rect 11336 11500 11388 11552
rect 12256 11500 12308 11552
rect 13820 11543 13872 11552
rect 13820 11509 13829 11543
rect 13829 11509 13863 11543
rect 13863 11509 13872 11543
rect 13820 11500 13872 11509
rect 14648 11500 14700 11552
rect 15936 11543 15988 11552
rect 15936 11509 15945 11543
rect 15945 11509 15979 11543
rect 15979 11509 15988 11543
rect 15936 11500 15988 11509
rect 17316 11500 17368 11552
rect 19524 11500 19576 11552
rect 20260 11500 20312 11552
rect 21824 11500 21876 11552
rect 26240 11543 26292 11552
rect 26240 11509 26249 11543
rect 26249 11509 26283 11543
rect 26283 11509 26292 11543
rect 26240 11500 26292 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1768 11296 1820 11348
rect 2136 11296 2188 11348
rect 2964 11339 3016 11348
rect 2964 11305 2973 11339
rect 2973 11305 3007 11339
rect 3007 11305 3016 11339
rect 2964 11296 3016 11305
rect 5540 11296 5592 11348
rect 6828 11296 6880 11348
rect 7380 11296 7432 11348
rect 8116 11339 8168 11348
rect 8116 11305 8125 11339
rect 8125 11305 8159 11339
rect 8159 11305 8168 11339
rect 8116 11296 8168 11305
rect 8484 11339 8536 11348
rect 8484 11305 8493 11339
rect 8493 11305 8527 11339
rect 8527 11305 8536 11339
rect 8484 11296 8536 11305
rect 9220 11296 9272 11348
rect 9404 11339 9456 11348
rect 9404 11305 9413 11339
rect 9413 11305 9447 11339
rect 9447 11305 9456 11339
rect 9404 11296 9456 11305
rect 9680 11339 9732 11348
rect 9680 11305 9689 11339
rect 9689 11305 9723 11339
rect 9723 11305 9732 11339
rect 9680 11296 9732 11305
rect 10140 11296 10192 11348
rect 11520 11296 11572 11348
rect 13636 11339 13688 11348
rect 13636 11305 13645 11339
rect 13645 11305 13679 11339
rect 13679 11305 13688 11339
rect 13636 11296 13688 11305
rect 13912 11296 13964 11348
rect 14648 11339 14700 11348
rect 14648 11305 14657 11339
rect 14657 11305 14691 11339
rect 14691 11305 14700 11339
rect 14648 11296 14700 11305
rect 15752 11296 15804 11348
rect 17040 11296 17092 11348
rect 17316 11296 17368 11348
rect 19984 11296 20036 11348
rect 22008 11339 22060 11348
rect 22008 11305 22017 11339
rect 22017 11305 22051 11339
rect 22051 11305 22060 11339
rect 22008 11296 22060 11305
rect 22744 11296 22796 11348
rect 23020 11339 23072 11348
rect 1860 11203 1912 11212
rect 1860 11169 1894 11203
rect 1894 11169 1912 11203
rect 1860 11160 1912 11169
rect 2136 11160 2188 11212
rect 3516 11160 3568 11212
rect 2780 11092 2832 11144
rect 5080 11228 5132 11280
rect 6092 11160 6144 11212
rect 7380 11203 7432 11212
rect 7380 11169 7389 11203
rect 7389 11169 7423 11203
rect 7423 11169 7432 11203
rect 7380 11160 7432 11169
rect 7840 11160 7892 11212
rect 11796 11228 11848 11280
rect 14280 11228 14332 11280
rect 8484 11160 8536 11212
rect 9680 11160 9732 11212
rect 10600 11160 10652 11212
rect 11704 11160 11756 11212
rect 12348 11160 12400 11212
rect 13176 11203 13228 11212
rect 13176 11169 13185 11203
rect 13185 11169 13219 11203
rect 13219 11169 13228 11203
rect 13176 11160 13228 11169
rect 13636 11160 13688 11212
rect 14372 11160 14424 11212
rect 15660 11228 15712 11280
rect 16856 11228 16908 11280
rect 18052 11160 18104 11212
rect 18236 11203 18288 11212
rect 18236 11169 18270 11203
rect 18270 11169 18288 11203
rect 18236 11160 18288 11169
rect 20076 11160 20128 11212
rect 22744 11160 22796 11212
rect 23020 11305 23029 11339
rect 23029 11305 23063 11339
rect 23063 11305 23072 11339
rect 23020 11296 23072 11305
rect 23204 11296 23256 11348
rect 24032 11296 24084 11348
rect 24952 11339 25004 11348
rect 24952 11305 24961 11339
rect 24961 11305 24995 11339
rect 24995 11305 25004 11339
rect 24952 11296 25004 11305
rect 25228 11339 25280 11348
rect 25228 11305 25237 11339
rect 25237 11305 25271 11339
rect 25271 11305 25280 11339
rect 25228 11296 25280 11305
rect 25320 11296 25372 11348
rect 23388 11228 23440 11280
rect 24676 11228 24728 11280
rect 23020 11160 23072 11212
rect 7564 11092 7616 11144
rect 6920 11067 6972 11076
rect 6920 11033 6929 11067
rect 6929 11033 6963 11067
rect 6963 11033 6972 11067
rect 6920 11024 6972 11033
rect 8116 11024 8168 11076
rect 12072 11092 12124 11144
rect 10324 11024 10376 11076
rect 10968 11024 11020 11076
rect 11060 11024 11112 11076
rect 3792 10956 3844 11008
rect 3976 10956 4028 11008
rect 6460 10956 6512 11008
rect 11428 10956 11480 11008
rect 12348 11024 12400 11076
rect 13912 11092 13964 11144
rect 15200 11092 15252 11144
rect 17960 11135 18012 11144
rect 17960 11101 17969 11135
rect 17969 11101 18003 11135
rect 18003 11101 18012 11135
rect 17960 11092 18012 11101
rect 19524 11092 19576 11144
rect 21364 11135 21416 11144
rect 14280 11024 14332 11076
rect 14004 10956 14056 11008
rect 14832 10956 14884 11008
rect 16856 11024 16908 11076
rect 17408 11067 17460 11076
rect 17408 11033 17417 11067
rect 17417 11033 17451 11067
rect 17451 11033 17460 11067
rect 17408 11024 17460 11033
rect 17776 11067 17828 11076
rect 17776 11033 17785 11067
rect 17785 11033 17819 11067
rect 17819 11033 17828 11067
rect 17776 11024 17828 11033
rect 19432 11024 19484 11076
rect 20260 11067 20312 11076
rect 20260 11033 20269 11067
rect 20269 11033 20303 11067
rect 20303 11033 20312 11067
rect 20260 11024 20312 11033
rect 21364 11101 21373 11135
rect 21373 11101 21407 11135
rect 21407 11101 21416 11135
rect 21364 11092 21416 11101
rect 23480 11092 23532 11144
rect 23296 11024 23348 11076
rect 18144 10956 18196 11008
rect 19340 10999 19392 11008
rect 19340 10965 19349 10999
rect 19349 10965 19383 10999
rect 19383 10965 19392 10999
rect 19340 10956 19392 10965
rect 23480 10999 23532 11008
rect 23480 10965 23489 10999
rect 23489 10965 23523 10999
rect 23523 10965 23532 10999
rect 23480 10956 23532 10965
rect 25596 10999 25648 11008
rect 25596 10965 25605 10999
rect 25605 10965 25639 10999
rect 25639 10965 25648 10999
rect 25596 10956 25648 10965
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 2596 10752 2648 10804
rect 1032 10616 1084 10668
rect 1584 10616 1636 10668
rect 5356 10752 5408 10804
rect 6644 10752 6696 10804
rect 8300 10795 8352 10804
rect 8300 10761 8309 10795
rect 8309 10761 8343 10795
rect 8343 10761 8352 10795
rect 8300 10752 8352 10761
rect 10324 10795 10376 10804
rect 10324 10761 10333 10795
rect 10333 10761 10367 10795
rect 10367 10761 10376 10795
rect 10324 10752 10376 10761
rect 13728 10795 13780 10804
rect 13728 10761 13737 10795
rect 13737 10761 13771 10795
rect 13771 10761 13780 10795
rect 13728 10752 13780 10761
rect 5080 10684 5132 10736
rect 6276 10684 6328 10736
rect 7380 10684 7432 10736
rect 7748 10684 7800 10736
rect 11796 10727 11848 10736
rect 11796 10693 11805 10727
rect 11805 10693 11839 10727
rect 11839 10693 11848 10727
rect 11796 10684 11848 10693
rect 13176 10684 13228 10736
rect 16028 10752 16080 10804
rect 16304 10795 16356 10804
rect 16304 10761 16313 10795
rect 16313 10761 16347 10795
rect 16347 10761 16356 10795
rect 16304 10752 16356 10761
rect 14832 10727 14884 10736
rect 14832 10693 14841 10727
rect 14841 10693 14875 10727
rect 14875 10693 14884 10727
rect 14832 10684 14884 10693
rect 15200 10684 15252 10736
rect 15752 10684 15804 10736
rect 7564 10616 7616 10668
rect 8852 10616 8904 10668
rect 10600 10659 10652 10668
rect 10600 10625 10609 10659
rect 10609 10625 10643 10659
rect 10643 10625 10652 10659
rect 10600 10616 10652 10625
rect 11428 10616 11480 10668
rect 15292 10659 15344 10668
rect 15292 10625 15301 10659
rect 15301 10625 15335 10659
rect 15335 10625 15344 10659
rect 15292 10616 15344 10625
rect 18236 10795 18288 10804
rect 17040 10659 17092 10668
rect 2688 10548 2740 10600
rect 3792 10591 3844 10600
rect 3792 10557 3801 10591
rect 3801 10557 3835 10591
rect 3835 10557 3844 10591
rect 3792 10548 3844 10557
rect 6828 10548 6880 10600
rect 7196 10591 7248 10600
rect 7196 10557 7205 10591
rect 7205 10557 7239 10591
rect 7239 10557 7248 10591
rect 7196 10548 7248 10557
rect 8300 10548 8352 10600
rect 8484 10548 8536 10600
rect 9496 10548 9548 10600
rect 11152 10548 11204 10600
rect 14280 10548 14332 10600
rect 17040 10625 17049 10659
rect 17049 10625 17083 10659
rect 17083 10625 17092 10659
rect 18236 10761 18245 10795
rect 18245 10761 18279 10795
rect 18279 10761 18288 10795
rect 18236 10752 18288 10761
rect 18696 10752 18748 10804
rect 20720 10752 20772 10804
rect 21088 10752 21140 10804
rect 20812 10684 20864 10736
rect 17040 10616 17092 10625
rect 21088 10616 21140 10668
rect 17500 10548 17552 10600
rect 18696 10548 18748 10600
rect 20260 10548 20312 10600
rect 20812 10548 20864 10600
rect 21456 10548 21508 10600
rect 23572 10752 23624 10804
rect 24216 10752 24268 10804
rect 24676 10795 24728 10804
rect 24676 10761 24685 10795
rect 24685 10761 24719 10795
rect 24719 10761 24728 10795
rect 24676 10752 24728 10761
rect 24860 10752 24912 10804
rect 25780 10752 25832 10804
rect 22008 10684 22060 10736
rect 22744 10727 22796 10736
rect 22744 10693 22753 10727
rect 22753 10693 22787 10727
rect 22787 10693 22796 10727
rect 22744 10684 22796 10693
rect 23296 10616 23348 10668
rect 25412 10659 25464 10668
rect 25412 10625 25421 10659
rect 25421 10625 25455 10659
rect 25455 10625 25464 10659
rect 25412 10616 25464 10625
rect 23480 10548 23532 10600
rect 25780 10548 25832 10600
rect 4068 10523 4120 10532
rect 4068 10489 4102 10523
rect 4102 10489 4120 10523
rect 4068 10480 4120 10489
rect 7932 10523 7984 10532
rect 7932 10489 7941 10523
rect 7941 10489 7975 10523
rect 7975 10489 7984 10523
rect 7932 10480 7984 10489
rect 15568 10480 15620 10532
rect 15752 10480 15804 10532
rect 2596 10412 2648 10464
rect 3240 10455 3292 10464
rect 3240 10421 3249 10455
rect 3249 10421 3283 10455
rect 3283 10421 3292 10455
rect 3240 10412 3292 10421
rect 6828 10455 6880 10464
rect 6828 10421 6837 10455
rect 6837 10421 6871 10455
rect 6871 10421 6880 10455
rect 6828 10412 6880 10421
rect 8484 10412 8536 10464
rect 11152 10455 11204 10464
rect 11152 10421 11161 10455
rect 11161 10421 11195 10455
rect 11195 10421 11204 10455
rect 11152 10412 11204 10421
rect 11336 10455 11388 10464
rect 11336 10421 11345 10455
rect 11345 10421 11379 10455
rect 11379 10421 11388 10455
rect 11336 10412 11388 10421
rect 12348 10412 12400 10464
rect 14372 10455 14424 10464
rect 14372 10421 14381 10455
rect 14381 10421 14415 10455
rect 14415 10421 14424 10455
rect 14372 10412 14424 10421
rect 15200 10455 15252 10464
rect 15200 10421 15209 10455
rect 15209 10421 15243 10455
rect 15243 10421 15252 10455
rect 15200 10412 15252 10421
rect 15844 10455 15896 10464
rect 15844 10421 15853 10455
rect 15853 10421 15887 10455
rect 15887 10421 15896 10455
rect 15844 10412 15896 10421
rect 16396 10455 16448 10464
rect 16396 10421 16405 10455
rect 16405 10421 16439 10455
rect 16439 10421 16448 10455
rect 16396 10412 16448 10421
rect 16672 10412 16724 10464
rect 16948 10412 17000 10464
rect 18696 10412 18748 10464
rect 19340 10455 19392 10464
rect 19340 10421 19349 10455
rect 19349 10421 19383 10455
rect 19383 10421 19392 10455
rect 19340 10412 19392 10421
rect 22192 10455 22244 10464
rect 22192 10421 22201 10455
rect 22201 10421 22235 10455
rect 22235 10421 22244 10455
rect 22192 10412 22244 10421
rect 24032 10412 24084 10464
rect 25596 10412 25648 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1860 10208 1912 10260
rect 2688 10208 2740 10260
rect 2780 10251 2832 10260
rect 2780 10217 2789 10251
rect 2789 10217 2823 10251
rect 2823 10217 2832 10251
rect 2780 10208 2832 10217
rect 3240 10208 3292 10260
rect 4804 10208 4856 10260
rect 5172 10208 5224 10260
rect 8300 10251 8352 10260
rect 8300 10217 8309 10251
rect 8309 10217 8343 10251
rect 8343 10217 8352 10251
rect 8300 10208 8352 10217
rect 9680 10208 9732 10260
rect 10048 10251 10100 10260
rect 10048 10217 10057 10251
rect 10057 10217 10091 10251
rect 10091 10217 10100 10251
rect 10048 10208 10100 10217
rect 10140 10251 10192 10260
rect 10140 10217 10149 10251
rect 10149 10217 10183 10251
rect 10183 10217 10192 10251
rect 10140 10208 10192 10217
rect 10784 10208 10836 10260
rect 10968 10208 11020 10260
rect 13636 10251 13688 10260
rect 13636 10217 13645 10251
rect 13645 10217 13679 10251
rect 13679 10217 13688 10251
rect 13636 10208 13688 10217
rect 13912 10251 13964 10260
rect 13912 10217 13921 10251
rect 13921 10217 13955 10251
rect 13955 10217 13964 10251
rect 13912 10208 13964 10217
rect 15200 10208 15252 10260
rect 18052 10208 18104 10260
rect 19156 10251 19208 10260
rect 19156 10217 19165 10251
rect 19165 10217 19199 10251
rect 19199 10217 19208 10251
rect 19156 10208 19208 10217
rect 21364 10208 21416 10260
rect 22744 10208 22796 10260
rect 23020 10208 23072 10260
rect 24860 10251 24912 10260
rect 6184 10140 6236 10192
rect 11704 10183 11756 10192
rect 11704 10149 11713 10183
rect 11713 10149 11747 10183
rect 11747 10149 11756 10183
rect 11704 10140 11756 10149
rect 15660 10140 15712 10192
rect 16580 10183 16632 10192
rect 16580 10149 16589 10183
rect 16589 10149 16623 10183
rect 16623 10149 16632 10183
rect 16580 10140 16632 10149
rect 16764 10140 16816 10192
rect 18328 10140 18380 10192
rect 24216 10140 24268 10192
rect 24860 10217 24869 10251
rect 24869 10217 24903 10251
rect 24903 10217 24912 10251
rect 24860 10208 24912 10217
rect 26056 10140 26108 10192
rect 2504 10072 2556 10124
rect 2688 10072 2740 10124
rect 5448 10072 5500 10124
rect 6092 10072 6144 10124
rect 6276 10072 6328 10124
rect 9496 10072 9548 10124
rect 12164 10115 12216 10124
rect 12164 10081 12198 10115
rect 12198 10081 12216 10115
rect 12164 10072 12216 10081
rect 14280 10072 14332 10124
rect 14648 10072 14700 10124
rect 17776 10072 17828 10124
rect 19524 10115 19576 10124
rect 2964 10047 3016 10056
rect 2412 9979 2464 9988
rect 2412 9945 2421 9979
rect 2421 9945 2455 9979
rect 2455 9945 2464 9979
rect 2412 9936 2464 9945
rect 2964 10013 2973 10047
rect 2973 10013 3007 10047
rect 3007 10013 3016 10047
rect 2964 10004 3016 10013
rect 4804 9936 4856 9988
rect 6000 10004 6052 10056
rect 10232 10047 10284 10056
rect 10232 10013 10241 10047
rect 10241 10013 10275 10047
rect 10275 10013 10284 10047
rect 10232 10004 10284 10013
rect 11888 10047 11940 10056
rect 11888 10013 11897 10047
rect 11897 10013 11931 10047
rect 11931 10013 11940 10047
rect 11888 10004 11940 10013
rect 17040 10004 17092 10056
rect 19524 10081 19533 10115
rect 19533 10081 19567 10115
rect 19567 10081 19576 10115
rect 19524 10072 19576 10081
rect 19616 10072 19668 10124
rect 20628 10072 20680 10124
rect 22468 10072 22520 10124
rect 22744 10072 22796 10124
rect 23204 10072 23256 10124
rect 23572 10072 23624 10124
rect 13544 9936 13596 9988
rect 18972 9936 19024 9988
rect 20444 9936 20496 9988
rect 23020 10004 23072 10056
rect 22192 9936 22244 9988
rect 23388 9936 23440 9988
rect 25136 9979 25188 9988
rect 25136 9945 25145 9979
rect 25145 9945 25179 9979
rect 25179 9945 25188 9979
rect 25136 9936 25188 9945
rect 26240 9936 26292 9988
rect 2688 9868 2740 9920
rect 3792 9868 3844 9920
rect 6000 9911 6052 9920
rect 6000 9877 6009 9911
rect 6009 9877 6043 9911
rect 6043 9877 6052 9911
rect 6000 9868 6052 9877
rect 6092 9868 6144 9920
rect 8024 9868 8076 9920
rect 9680 9911 9732 9920
rect 9680 9877 9689 9911
rect 9689 9877 9723 9911
rect 9723 9877 9732 9911
rect 9680 9868 9732 9877
rect 11428 9911 11480 9920
rect 11428 9877 11437 9911
rect 11437 9877 11471 9911
rect 11471 9877 11480 9911
rect 11428 9868 11480 9877
rect 14464 9868 14516 9920
rect 16672 9868 16724 9920
rect 19984 9868 20036 9920
rect 20904 9868 20956 9920
rect 23020 9911 23072 9920
rect 23020 9877 23029 9911
rect 23029 9877 23063 9911
rect 23063 9877 23072 9911
rect 23020 9868 23072 9877
rect 25596 9868 25648 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 1584 9639 1636 9648
rect 1584 9605 1593 9639
rect 1593 9605 1627 9639
rect 1627 9605 1636 9639
rect 1584 9596 1636 9605
rect 1860 9596 1912 9648
rect 4804 9664 4856 9716
rect 6184 9707 6236 9716
rect 6184 9673 6193 9707
rect 6193 9673 6227 9707
rect 6227 9673 6236 9707
rect 6184 9664 6236 9673
rect 4988 9639 5040 9648
rect 4988 9605 4997 9639
rect 4997 9605 5031 9639
rect 5031 9605 5040 9639
rect 4988 9596 5040 9605
rect 10048 9664 10100 9716
rect 6276 9528 6328 9580
rect 1676 9460 1728 9512
rect 2412 9460 2464 9512
rect 3792 9460 3844 9512
rect 6000 9460 6052 9512
rect 8024 9460 8076 9512
rect 10140 9596 10192 9648
rect 11152 9664 11204 9716
rect 12440 9664 12492 9716
rect 14280 9664 14332 9716
rect 11060 9528 11112 9580
rect 11796 9528 11848 9580
rect 14188 9596 14240 9648
rect 10232 9503 10284 9512
rect 10232 9469 10241 9503
rect 10241 9469 10275 9503
rect 10275 9469 10284 9503
rect 10232 9460 10284 9469
rect 2964 9435 3016 9444
rect 2964 9401 2998 9435
rect 2998 9401 3016 9435
rect 2964 9392 3016 9401
rect 4528 9392 4580 9444
rect 6552 9392 6604 9444
rect 8116 9392 8168 9444
rect 11152 9435 11204 9444
rect 11152 9401 11161 9435
rect 11161 9401 11195 9435
rect 11195 9401 11204 9435
rect 11152 9392 11204 9401
rect 12348 9392 12400 9444
rect 12716 9435 12768 9444
rect 12716 9401 12750 9435
rect 12750 9401 12768 9435
rect 12716 9392 12768 9401
rect 14740 9596 14792 9648
rect 16672 9664 16724 9716
rect 16488 9528 16540 9580
rect 16856 9528 16908 9580
rect 17776 9596 17828 9648
rect 18052 9664 18104 9716
rect 18328 9707 18380 9716
rect 18328 9673 18337 9707
rect 18337 9673 18371 9707
rect 18371 9673 18380 9707
rect 18328 9664 18380 9673
rect 21180 9664 21232 9716
rect 22744 9707 22796 9716
rect 22744 9673 22753 9707
rect 22753 9673 22787 9707
rect 22787 9673 22796 9707
rect 22744 9664 22796 9673
rect 24952 9664 25004 9716
rect 19432 9596 19484 9648
rect 20076 9639 20128 9648
rect 20076 9605 20085 9639
rect 20085 9605 20119 9639
rect 20119 9605 20128 9639
rect 20076 9596 20128 9605
rect 21824 9596 21876 9648
rect 21916 9596 21968 9648
rect 18972 9571 19024 9580
rect 18972 9537 18981 9571
rect 18981 9537 19015 9571
rect 19015 9537 19024 9571
rect 18972 9528 19024 9537
rect 14648 9460 14700 9512
rect 15108 9503 15160 9512
rect 15108 9469 15117 9503
rect 15117 9469 15151 9503
rect 15151 9469 15160 9503
rect 15108 9460 15160 9469
rect 16212 9460 16264 9512
rect 18328 9460 18380 9512
rect 18604 9460 18656 9512
rect 19248 9528 19300 9580
rect 20628 9571 20680 9580
rect 20628 9537 20637 9571
rect 20637 9537 20671 9571
rect 20671 9537 20680 9571
rect 20628 9528 20680 9537
rect 21272 9571 21324 9580
rect 21272 9537 21281 9571
rect 21281 9537 21315 9571
rect 21315 9537 21324 9571
rect 21272 9528 21324 9537
rect 22284 9596 22336 9648
rect 19892 9503 19944 9512
rect 19892 9469 19901 9503
rect 19901 9469 19935 9503
rect 19935 9469 19944 9503
rect 19892 9460 19944 9469
rect 22744 9460 22796 9512
rect 23388 9460 23440 9512
rect 23572 9460 23624 9512
rect 23940 9503 23992 9512
rect 23940 9469 23974 9503
rect 23974 9469 23992 9503
rect 15016 9435 15068 9444
rect 15016 9401 15025 9435
rect 15025 9401 15059 9435
rect 15059 9401 15068 9435
rect 15016 9392 15068 9401
rect 16488 9392 16540 9444
rect 18144 9392 18196 9444
rect 19156 9392 19208 9444
rect 20904 9392 20956 9444
rect 23940 9460 23992 9469
rect 3516 9324 3568 9376
rect 4068 9367 4120 9376
rect 4068 9333 4077 9367
rect 4077 9333 4111 9367
rect 4111 9333 4120 9367
rect 4068 9324 4120 9333
rect 5172 9367 5224 9376
rect 5172 9333 5181 9367
rect 5181 9333 5215 9367
rect 5215 9333 5224 9367
rect 5172 9324 5224 9333
rect 6000 9324 6052 9376
rect 10784 9367 10836 9376
rect 10784 9333 10793 9367
rect 10793 9333 10827 9367
rect 10827 9333 10836 9367
rect 10784 9324 10836 9333
rect 12164 9324 12216 9376
rect 13544 9324 13596 9376
rect 16580 9324 16632 9376
rect 19432 9324 19484 9376
rect 20536 9367 20588 9376
rect 20536 9333 20545 9367
rect 20545 9333 20579 9367
rect 20579 9333 20588 9367
rect 20536 9324 20588 9333
rect 20996 9324 21048 9376
rect 21180 9367 21232 9376
rect 21180 9333 21189 9367
rect 21189 9333 21223 9367
rect 21223 9333 21232 9367
rect 21180 9324 21232 9333
rect 21364 9324 21416 9376
rect 25596 9392 25648 9444
rect 22192 9324 22244 9376
rect 24952 9324 25004 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1676 9120 1728 9172
rect 2688 9120 2740 9172
rect 5448 9120 5500 9172
rect 6828 9120 6880 9172
rect 9772 9163 9824 9172
rect 9772 9129 9781 9163
rect 9781 9129 9815 9163
rect 9815 9129 9824 9163
rect 9772 9120 9824 9129
rect 11152 9120 11204 9172
rect 11796 9120 11848 9172
rect 12716 9120 12768 9172
rect 13268 9120 13320 9172
rect 13452 9120 13504 9172
rect 14648 9163 14700 9172
rect 14648 9129 14657 9163
rect 14657 9129 14691 9163
rect 14691 9129 14700 9163
rect 14648 9120 14700 9129
rect 15108 9163 15160 9172
rect 15108 9129 15117 9163
rect 15117 9129 15151 9163
rect 15151 9129 15160 9163
rect 15108 9120 15160 9129
rect 15384 9120 15436 9172
rect 15660 9163 15712 9172
rect 15660 9129 15669 9163
rect 15669 9129 15703 9163
rect 15703 9129 15712 9163
rect 15660 9120 15712 9129
rect 16212 9120 16264 9172
rect 16488 9163 16540 9172
rect 16488 9129 16497 9163
rect 16497 9129 16531 9163
rect 16531 9129 16540 9163
rect 16488 9120 16540 9129
rect 16856 9163 16908 9172
rect 16856 9129 16865 9163
rect 16865 9129 16899 9163
rect 16899 9129 16908 9163
rect 16856 9120 16908 9129
rect 17500 9163 17552 9172
rect 17500 9129 17509 9163
rect 17509 9129 17543 9163
rect 17543 9129 17552 9163
rect 17500 9120 17552 9129
rect 18604 9163 18656 9172
rect 18604 9129 18613 9163
rect 18613 9129 18647 9163
rect 18647 9129 18656 9163
rect 18604 9120 18656 9129
rect 18788 9120 18840 9172
rect 20536 9120 20588 9172
rect 21180 9120 21232 9172
rect 22192 9120 22244 9172
rect 23940 9120 23992 9172
rect 25136 9120 25188 9172
rect 25596 9163 25648 9172
rect 25596 9129 25605 9163
rect 25605 9129 25639 9163
rect 25639 9129 25648 9163
rect 25596 9120 25648 9129
rect 26148 9120 26200 9172
rect 1584 8916 1636 8968
rect 6000 9052 6052 9104
rect 7932 9052 7984 9104
rect 8852 9052 8904 9104
rect 9404 9095 9456 9104
rect 9404 9061 9413 9095
rect 9413 9061 9447 9095
rect 9447 9061 9456 9095
rect 9404 9052 9456 9061
rect 11428 9052 11480 9104
rect 2688 8984 2740 9036
rect 5540 8984 5592 9036
rect 2964 8959 3016 8968
rect 2964 8925 2973 8959
rect 2973 8925 3007 8959
rect 3007 8925 3016 8959
rect 2964 8916 3016 8925
rect 5172 8916 5224 8968
rect 5448 8891 5500 8900
rect 5448 8857 5457 8891
rect 5457 8857 5491 8891
rect 5491 8857 5500 8891
rect 5448 8848 5500 8857
rect 2044 8780 2096 8832
rect 4344 8823 4396 8832
rect 4344 8789 4353 8823
rect 4353 8789 4387 8823
rect 4387 8789 4396 8823
rect 4344 8780 4396 8789
rect 4896 8780 4948 8832
rect 7656 8984 7708 9036
rect 6276 8916 6328 8968
rect 6460 8916 6512 8968
rect 8576 8959 8628 8968
rect 8576 8925 8585 8959
rect 8585 8925 8619 8959
rect 8619 8925 8628 8959
rect 8576 8916 8628 8925
rect 9404 8916 9456 8968
rect 13176 9052 13228 9104
rect 13912 9052 13964 9104
rect 22928 9052 22980 9104
rect 13452 9027 13504 9036
rect 13452 8993 13461 9027
rect 13461 8993 13495 9027
rect 13495 8993 13504 9027
rect 13452 8984 13504 8993
rect 16948 8984 17000 9036
rect 8024 8848 8076 8900
rect 6276 8780 6328 8832
rect 7840 8780 7892 8832
rect 8668 8780 8720 8832
rect 9128 8823 9180 8832
rect 9128 8789 9137 8823
rect 9137 8789 9171 8823
rect 9171 8789 9180 8823
rect 9128 8780 9180 8789
rect 12992 8916 13044 8968
rect 13544 8959 13596 8968
rect 13544 8925 13553 8959
rect 13553 8925 13587 8959
rect 13587 8925 13596 8959
rect 13544 8916 13596 8925
rect 15752 8959 15804 8968
rect 15752 8925 15761 8959
rect 15761 8925 15795 8959
rect 15795 8925 15804 8959
rect 15752 8916 15804 8925
rect 11888 8848 11940 8900
rect 10968 8780 11020 8832
rect 13636 8780 13688 8832
rect 14372 8848 14424 8900
rect 17224 8916 17276 8968
rect 17960 8984 18012 9036
rect 19984 8984 20036 9036
rect 20536 8984 20588 9036
rect 20904 8984 20956 9036
rect 17684 8916 17736 8968
rect 18052 8916 18104 8968
rect 19156 8959 19208 8968
rect 19156 8925 19165 8959
rect 19165 8925 19199 8959
rect 19199 8925 19208 8959
rect 19156 8916 19208 8925
rect 19524 8916 19576 8968
rect 21180 8916 21232 8968
rect 20628 8848 20680 8900
rect 21824 8916 21876 8968
rect 23572 8984 23624 9036
rect 24952 9027 25004 9036
rect 24952 8993 24961 9027
rect 24961 8993 24995 9027
rect 24995 8993 25004 9027
rect 24952 8984 25004 8993
rect 21548 8848 21600 8900
rect 16396 8780 16448 8832
rect 17224 8780 17276 8832
rect 17960 8780 18012 8832
rect 20260 8823 20312 8832
rect 20260 8789 20269 8823
rect 20269 8789 20303 8823
rect 20303 8789 20312 8823
rect 20260 8780 20312 8789
rect 20812 8780 20864 8832
rect 21456 8780 21508 8832
rect 22008 8823 22060 8832
rect 22008 8789 22017 8823
rect 22017 8789 22051 8823
rect 22051 8789 22060 8823
rect 22008 8780 22060 8789
rect 22192 8780 22244 8832
rect 23020 8780 23072 8832
rect 25596 8848 25648 8900
rect 25136 8823 25188 8832
rect 25136 8789 25145 8823
rect 25145 8789 25179 8823
rect 25179 8789 25188 8823
rect 25136 8780 25188 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 5080 8619 5132 8628
rect 5080 8585 5089 8619
rect 5089 8585 5123 8619
rect 5123 8585 5132 8619
rect 5080 8576 5132 8585
rect 6460 8576 6512 8628
rect 7656 8576 7708 8628
rect 7932 8619 7984 8628
rect 7932 8585 7941 8619
rect 7941 8585 7975 8619
rect 7975 8585 7984 8619
rect 7932 8576 7984 8585
rect 8392 8576 8444 8628
rect 9404 8576 9456 8628
rect 10140 8576 10192 8628
rect 13544 8619 13596 8628
rect 13544 8585 13553 8619
rect 13553 8585 13587 8619
rect 13587 8585 13596 8619
rect 13544 8576 13596 8585
rect 14740 8576 14792 8628
rect 15844 8576 15896 8628
rect 17500 8576 17552 8628
rect 17684 8576 17736 8628
rect 18420 8576 18472 8628
rect 19432 8619 19484 8628
rect 19432 8585 19441 8619
rect 19441 8585 19475 8619
rect 19475 8585 19484 8619
rect 19432 8576 19484 8585
rect 1216 8440 1268 8492
rect 1768 8440 1820 8492
rect 4344 8440 4396 8492
rect 14372 8551 14424 8560
rect 1676 8372 1728 8424
rect 2412 8372 2464 8424
rect 4896 8415 4948 8424
rect 1768 8347 1820 8356
rect 1768 8313 1777 8347
rect 1777 8313 1811 8347
rect 1811 8313 1820 8347
rect 1768 8304 1820 8313
rect 2964 8304 3016 8356
rect 4896 8381 4905 8415
rect 4905 8381 4939 8415
rect 4939 8381 4948 8415
rect 4896 8372 4948 8381
rect 5448 8415 5500 8424
rect 5448 8381 5457 8415
rect 5457 8381 5491 8415
rect 5491 8381 5500 8415
rect 5448 8372 5500 8381
rect 3516 8304 3568 8356
rect 1308 8236 1360 8288
rect 2688 8236 2740 8288
rect 2780 8236 2832 8288
rect 6276 8440 6328 8492
rect 11244 8483 11296 8492
rect 6828 8372 6880 8424
rect 8392 8372 8444 8424
rect 8852 8372 8904 8424
rect 11244 8449 11253 8483
rect 11253 8449 11287 8483
rect 11287 8449 11296 8483
rect 11244 8440 11296 8449
rect 11428 8483 11480 8492
rect 11428 8449 11437 8483
rect 11437 8449 11471 8483
rect 11471 8449 11480 8483
rect 11428 8440 11480 8449
rect 11152 8372 11204 8424
rect 6920 8304 6972 8356
rect 7564 8304 7616 8356
rect 8668 8304 8720 8356
rect 8392 8279 8444 8288
rect 8392 8245 8401 8279
rect 8401 8245 8435 8279
rect 8435 8245 8444 8279
rect 8392 8236 8444 8245
rect 9220 8304 9272 8356
rect 9772 8347 9824 8356
rect 9772 8313 9781 8347
rect 9781 8313 9815 8347
rect 9815 8313 9824 8347
rect 9772 8304 9824 8313
rect 12440 8372 12492 8424
rect 14372 8517 14381 8551
rect 14381 8517 14415 8551
rect 14415 8517 14424 8551
rect 14372 8508 14424 8517
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 14924 8415 14976 8424
rect 14924 8381 14933 8415
rect 14933 8381 14967 8415
rect 14967 8381 14976 8415
rect 14924 8372 14976 8381
rect 10784 8236 10836 8288
rect 16028 8372 16080 8424
rect 17408 8415 17460 8424
rect 17408 8381 17417 8415
rect 17417 8381 17451 8415
rect 17451 8381 17460 8415
rect 17408 8372 17460 8381
rect 19340 8508 19392 8560
rect 21180 8576 21232 8628
rect 22192 8619 22244 8628
rect 22192 8585 22201 8619
rect 22201 8585 22235 8619
rect 22235 8585 22244 8619
rect 22192 8576 22244 8585
rect 22928 8576 22980 8628
rect 23664 8619 23716 8628
rect 23664 8585 23673 8619
rect 23673 8585 23707 8619
rect 23707 8585 23716 8619
rect 23664 8576 23716 8585
rect 24952 8619 25004 8628
rect 24952 8585 24961 8619
rect 24961 8585 24995 8619
rect 24995 8585 25004 8619
rect 24952 8576 25004 8585
rect 26148 8619 26200 8628
rect 26148 8585 26157 8619
rect 26157 8585 26191 8619
rect 26191 8585 26200 8619
rect 26148 8576 26200 8585
rect 22008 8440 22060 8492
rect 22284 8440 22336 8492
rect 20260 8372 20312 8424
rect 11152 8279 11204 8288
rect 11152 8245 11161 8279
rect 11161 8245 11195 8279
rect 11195 8245 11204 8279
rect 11152 8236 11204 8245
rect 12440 8279 12492 8288
rect 12440 8245 12449 8279
rect 12449 8245 12483 8279
rect 12483 8245 12492 8279
rect 12440 8236 12492 8245
rect 13912 8236 13964 8288
rect 14096 8236 14148 8288
rect 14556 8236 14608 8288
rect 15384 8236 15436 8288
rect 15752 8236 15804 8288
rect 17316 8236 17368 8288
rect 18144 8304 18196 8356
rect 18512 8304 18564 8356
rect 18052 8236 18104 8288
rect 19524 8236 19576 8288
rect 21088 8372 21140 8424
rect 24124 8372 24176 8424
rect 25136 8372 25188 8424
rect 20720 8304 20772 8356
rect 23572 8304 23624 8356
rect 21732 8236 21784 8288
rect 21916 8279 21968 8288
rect 21916 8245 21925 8279
rect 21925 8245 21959 8279
rect 21959 8245 21968 8279
rect 21916 8236 21968 8245
rect 24768 8304 24820 8356
rect 25872 8236 25924 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 2504 8032 2556 8084
rect 5172 8032 5224 8084
rect 6276 8075 6328 8084
rect 6276 8041 6285 8075
rect 6285 8041 6319 8075
rect 6319 8041 6328 8075
rect 6276 8032 6328 8041
rect 7564 8075 7616 8084
rect 7564 8041 7573 8075
rect 7573 8041 7607 8075
rect 7607 8041 7616 8075
rect 7564 8032 7616 8041
rect 7656 8032 7708 8084
rect 9128 8032 9180 8084
rect 10140 8032 10192 8084
rect 10784 8075 10836 8084
rect 2780 8007 2832 8016
rect 2780 7973 2789 8007
rect 2789 7973 2823 8007
rect 2823 7973 2832 8007
rect 2780 7964 2832 7973
rect 5448 7964 5500 8016
rect 8300 7964 8352 8016
rect 9588 7964 9640 8016
rect 4988 7896 5040 7948
rect 6460 7896 6512 7948
rect 6920 7939 6972 7948
rect 6920 7905 6929 7939
rect 6929 7905 6963 7939
rect 6963 7905 6972 7939
rect 6920 7896 6972 7905
rect 7104 7896 7156 7948
rect 8760 7896 8812 7948
rect 9496 7896 9548 7948
rect 9864 7939 9916 7948
rect 9864 7905 9873 7939
rect 9873 7905 9907 7939
rect 9907 7905 9916 7939
rect 9864 7896 9916 7905
rect 10784 8041 10793 8075
rect 10793 8041 10827 8075
rect 10827 8041 10836 8075
rect 10784 8032 10836 8041
rect 12256 8032 12308 8084
rect 12992 8032 13044 8084
rect 13452 8032 13504 8084
rect 14096 8032 14148 8084
rect 14832 8032 14884 8084
rect 15292 8032 15344 8084
rect 15660 8032 15712 8084
rect 16212 8032 16264 8084
rect 17868 8032 17920 8084
rect 18144 8075 18196 8084
rect 18144 8041 18153 8075
rect 18153 8041 18187 8075
rect 18187 8041 18196 8075
rect 18144 8032 18196 8041
rect 19524 8032 19576 8084
rect 20628 8075 20680 8084
rect 20628 8041 20637 8075
rect 20637 8041 20671 8075
rect 20671 8041 20680 8075
rect 20628 8032 20680 8041
rect 21548 8075 21600 8084
rect 21548 8041 21557 8075
rect 21557 8041 21591 8075
rect 21591 8041 21600 8075
rect 21548 8032 21600 8041
rect 22928 8032 22980 8084
rect 24032 8075 24084 8084
rect 24032 8041 24041 8075
rect 24041 8041 24075 8075
rect 24075 8041 24084 8075
rect 24032 8032 24084 8041
rect 25228 8032 25280 8084
rect 26148 8075 26200 8084
rect 26148 8041 26157 8075
rect 26157 8041 26191 8075
rect 26191 8041 26200 8075
rect 26148 8032 26200 8041
rect 11428 7964 11480 8016
rect 12440 7964 12492 8016
rect 13820 7964 13872 8016
rect 17132 8007 17184 8016
rect 17132 7973 17141 8007
rect 17141 7973 17175 8007
rect 17175 7973 17184 8007
rect 17132 7964 17184 7973
rect 22100 8007 22152 8016
rect 22100 7973 22134 8007
rect 22134 7973 22152 8007
rect 22100 7964 22152 7973
rect 23756 7964 23808 8016
rect 10784 7896 10836 7948
rect 2136 7828 2188 7880
rect 2504 7828 2556 7880
rect 2964 7760 3016 7812
rect 3148 7828 3200 7880
rect 4896 7871 4948 7880
rect 4896 7837 4905 7871
rect 4905 7837 4939 7871
rect 4939 7837 4948 7871
rect 4896 7828 4948 7837
rect 8852 7828 8904 7880
rect 12348 7896 12400 7948
rect 12716 7896 12768 7948
rect 13452 7896 13504 7948
rect 13636 7871 13688 7880
rect 7012 7760 7064 7812
rect 9128 7760 9180 7812
rect 13636 7837 13645 7871
rect 13645 7837 13679 7871
rect 13679 7837 13688 7871
rect 13636 7828 13688 7837
rect 16028 7896 16080 7948
rect 17408 7896 17460 7948
rect 15476 7871 15528 7880
rect 15476 7837 15485 7871
rect 15485 7837 15519 7871
rect 15519 7837 15528 7871
rect 15476 7828 15528 7837
rect 17316 7871 17368 7880
rect 17316 7837 17325 7871
rect 17325 7837 17359 7871
rect 17359 7837 17368 7871
rect 23296 7896 23348 7948
rect 17316 7828 17368 7837
rect 14280 7760 14332 7812
rect 15292 7760 15344 7812
rect 1676 7735 1728 7744
rect 1676 7701 1685 7735
rect 1685 7701 1719 7735
rect 1719 7701 1728 7735
rect 1676 7692 1728 7701
rect 2136 7735 2188 7744
rect 2136 7701 2145 7735
rect 2145 7701 2179 7735
rect 2179 7701 2188 7735
rect 2136 7692 2188 7701
rect 3700 7735 3752 7744
rect 3700 7701 3709 7735
rect 3709 7701 3743 7735
rect 3743 7701 3752 7735
rect 3700 7692 3752 7701
rect 7748 7692 7800 7744
rect 8852 7692 8904 7744
rect 12256 7692 12308 7744
rect 12624 7735 12676 7744
rect 12624 7701 12633 7735
rect 12633 7701 12667 7735
rect 12667 7701 12676 7735
rect 12624 7692 12676 7701
rect 12808 7692 12860 7744
rect 21732 7828 21784 7880
rect 24124 7828 24176 7880
rect 24676 7896 24728 7948
rect 24768 7828 24820 7880
rect 18512 7692 18564 7744
rect 19432 7692 19484 7744
rect 20904 7692 20956 7744
rect 23940 7692 23992 7744
rect 26240 7692 26292 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 2044 7531 2096 7540
rect 2044 7497 2053 7531
rect 2053 7497 2087 7531
rect 2087 7497 2096 7531
rect 2044 7488 2096 7497
rect 7656 7488 7708 7540
rect 9588 7531 9640 7540
rect 9588 7497 9597 7531
rect 9597 7497 9631 7531
rect 9631 7497 9640 7531
rect 9588 7488 9640 7497
rect 9864 7531 9916 7540
rect 9864 7497 9873 7531
rect 9873 7497 9907 7531
rect 9907 7497 9916 7531
rect 9864 7488 9916 7497
rect 10784 7531 10836 7540
rect 10784 7497 10793 7531
rect 10793 7497 10827 7531
rect 10827 7497 10836 7531
rect 10784 7488 10836 7497
rect 11428 7488 11480 7540
rect 11888 7488 11940 7540
rect 12256 7531 12308 7540
rect 12256 7497 12265 7531
rect 12265 7497 12299 7531
rect 12299 7497 12308 7531
rect 12256 7488 12308 7497
rect 13636 7488 13688 7540
rect 16028 7531 16080 7540
rect 16028 7497 16037 7531
rect 16037 7497 16071 7531
rect 16071 7497 16080 7531
rect 16028 7488 16080 7497
rect 664 7420 716 7472
rect 1952 7420 2004 7472
rect 2136 7420 2188 7472
rect 4988 7420 5040 7472
rect 3700 7352 3752 7404
rect 4896 7352 4948 7404
rect 6920 7352 6972 7404
rect 8300 7420 8352 7472
rect 8852 7420 8904 7472
rect 7564 7352 7616 7404
rect 8944 7395 8996 7404
rect 8944 7361 8953 7395
rect 8953 7361 8987 7395
rect 8987 7361 8996 7395
rect 8944 7352 8996 7361
rect 10048 7420 10100 7472
rect 11060 7420 11112 7472
rect 13452 7463 13504 7472
rect 13452 7429 13461 7463
rect 13461 7429 13495 7463
rect 13495 7429 13504 7463
rect 13452 7420 13504 7429
rect 12624 7352 12676 7404
rect 12992 7395 13044 7404
rect 12992 7361 13001 7395
rect 13001 7361 13035 7395
rect 13035 7361 13044 7395
rect 12992 7352 13044 7361
rect 2504 7327 2556 7336
rect 2504 7293 2513 7327
rect 2513 7293 2547 7327
rect 2547 7293 2556 7327
rect 2504 7284 2556 7293
rect 4068 7327 4120 7336
rect 4068 7293 4077 7327
rect 4077 7293 4111 7327
rect 4111 7293 4120 7327
rect 4068 7284 4120 7293
rect 6368 7284 6420 7336
rect 8576 7284 8628 7336
rect 10692 7284 10744 7336
rect 11336 7284 11388 7336
rect 12808 7327 12860 7336
rect 12808 7293 12817 7327
rect 12817 7293 12851 7327
rect 12851 7293 12860 7327
rect 12808 7284 12860 7293
rect 14832 7284 14884 7336
rect 15016 7284 15068 7336
rect 16396 7284 16448 7336
rect 17040 7488 17092 7540
rect 20812 7531 20864 7540
rect 20812 7497 20821 7531
rect 20821 7497 20855 7531
rect 20855 7497 20864 7531
rect 20812 7488 20864 7497
rect 22100 7488 22152 7540
rect 23480 7488 23532 7540
rect 24768 7488 24820 7540
rect 26148 7531 26200 7540
rect 26148 7497 26157 7531
rect 26157 7497 26191 7531
rect 26191 7497 26200 7531
rect 26148 7488 26200 7497
rect 20720 7463 20772 7472
rect 20720 7429 20729 7463
rect 20729 7429 20763 7463
rect 20763 7429 20772 7463
rect 20720 7420 20772 7429
rect 18052 7352 18104 7404
rect 22468 7420 22520 7472
rect 26608 7420 26660 7472
rect 18604 7327 18656 7336
rect 18604 7293 18613 7327
rect 18613 7293 18647 7327
rect 18647 7293 18656 7327
rect 18604 7284 18656 7293
rect 21548 7352 21600 7404
rect 22100 7352 22152 7404
rect 22560 7352 22612 7404
rect 23296 7352 23348 7404
rect 23848 7352 23900 7404
rect 22008 7284 22060 7336
rect 23756 7284 23808 7336
rect 24768 7395 24820 7404
rect 24768 7361 24777 7395
rect 24777 7361 24811 7395
rect 24811 7361 24820 7395
rect 24768 7352 24820 7361
rect 1952 7148 2004 7200
rect 3148 7191 3200 7200
rect 3148 7157 3157 7191
rect 3157 7157 3191 7191
rect 3191 7157 3200 7191
rect 3148 7148 3200 7157
rect 4160 7216 4212 7268
rect 6000 7216 6052 7268
rect 7380 7216 7432 7268
rect 12072 7216 12124 7268
rect 14740 7216 14792 7268
rect 16764 7259 16816 7268
rect 16764 7225 16773 7259
rect 16773 7225 16807 7259
rect 16807 7225 16816 7259
rect 16764 7216 16816 7225
rect 17316 7259 17368 7268
rect 17316 7225 17325 7259
rect 17325 7225 17359 7259
rect 17359 7225 17368 7259
rect 17316 7216 17368 7225
rect 3976 7191 4028 7200
rect 3976 7157 3985 7191
rect 3985 7157 4019 7191
rect 4019 7157 4028 7191
rect 3976 7148 4028 7157
rect 5172 7191 5224 7200
rect 5172 7157 5181 7191
rect 5181 7157 5215 7191
rect 5215 7157 5224 7191
rect 5172 7148 5224 7157
rect 6644 7148 6696 7200
rect 8484 7191 8536 7200
rect 8484 7157 8493 7191
rect 8493 7157 8527 7191
rect 8527 7157 8536 7191
rect 8484 7148 8536 7157
rect 15200 7148 15252 7200
rect 15660 7191 15712 7200
rect 15660 7157 15669 7191
rect 15669 7157 15703 7191
rect 15703 7157 15712 7191
rect 15660 7148 15712 7157
rect 24124 7216 24176 7268
rect 20076 7148 20128 7200
rect 20352 7191 20404 7200
rect 20352 7157 20361 7191
rect 20361 7157 20395 7191
rect 20395 7157 20404 7191
rect 20352 7148 20404 7157
rect 22652 7191 22704 7200
rect 22652 7157 22661 7191
rect 22661 7157 22695 7191
rect 22695 7157 22704 7191
rect 22652 7148 22704 7157
rect 23480 7191 23532 7200
rect 23480 7157 23489 7191
rect 23489 7157 23523 7191
rect 23523 7157 23532 7191
rect 23480 7148 23532 7157
rect 25228 7148 25280 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 1768 6987 1820 6996
rect 1768 6953 1777 6987
rect 1777 6953 1811 6987
rect 1811 6953 1820 6987
rect 1768 6944 1820 6953
rect 2780 6944 2832 6996
rect 3976 6944 4028 6996
rect 4988 6987 5040 6996
rect 4988 6953 4997 6987
rect 4997 6953 5031 6987
rect 5031 6953 5040 6987
rect 4988 6944 5040 6953
rect 8576 6944 8628 6996
rect 9680 6944 9732 6996
rect 10048 6987 10100 6996
rect 10048 6953 10057 6987
rect 10057 6953 10091 6987
rect 10091 6953 10100 6987
rect 10048 6944 10100 6953
rect 10876 6944 10928 6996
rect 11336 6987 11388 6996
rect 11336 6953 11345 6987
rect 11345 6953 11379 6987
rect 11379 6953 11388 6987
rect 11336 6944 11388 6953
rect 11704 6987 11756 6996
rect 11704 6953 11713 6987
rect 11713 6953 11747 6987
rect 11747 6953 11756 6987
rect 11704 6944 11756 6953
rect 11796 6944 11848 6996
rect 12256 6944 12308 6996
rect 2596 6851 2648 6860
rect 2596 6817 2605 6851
rect 2605 6817 2639 6851
rect 2639 6817 2648 6851
rect 2596 6808 2648 6817
rect 5356 6808 5408 6860
rect 6644 6876 6696 6928
rect 5632 6851 5684 6860
rect 5632 6817 5641 6851
rect 5641 6817 5675 6851
rect 5675 6817 5684 6851
rect 8484 6876 8536 6928
rect 13728 6876 13780 6928
rect 15016 6944 15068 6996
rect 16212 6944 16264 6996
rect 17408 6944 17460 6996
rect 17776 6987 17828 6996
rect 17776 6953 17785 6987
rect 17785 6953 17819 6987
rect 17819 6953 17828 6987
rect 17776 6944 17828 6953
rect 20720 6944 20772 6996
rect 23848 6944 23900 6996
rect 26148 6987 26200 6996
rect 26148 6953 26157 6987
rect 26157 6953 26191 6987
rect 26191 6953 26200 6987
rect 26148 6944 26200 6953
rect 19432 6919 19484 6928
rect 5632 6808 5684 6817
rect 7012 6808 7064 6860
rect 10692 6808 10744 6860
rect 11520 6808 11572 6860
rect 12624 6808 12676 6860
rect 12900 6808 12952 6860
rect 13360 6851 13412 6860
rect 13360 6817 13369 6851
rect 13369 6817 13403 6851
rect 13403 6817 13412 6851
rect 13360 6808 13412 6817
rect 13820 6808 13872 6860
rect 19432 6885 19441 6919
rect 19441 6885 19475 6919
rect 19475 6885 19484 6919
rect 19432 6876 19484 6885
rect 21364 6876 21416 6928
rect 22652 6876 22704 6928
rect 24952 6876 25004 6928
rect 15936 6808 15988 6860
rect 16488 6808 16540 6860
rect 17224 6851 17276 6860
rect 17224 6817 17233 6851
rect 17233 6817 17267 6851
rect 17267 6817 17276 6851
rect 17224 6808 17276 6817
rect 17868 6851 17920 6860
rect 17868 6817 17877 6851
rect 17877 6817 17911 6851
rect 17911 6817 17920 6851
rect 17868 6808 17920 6817
rect 21824 6808 21876 6860
rect 22284 6808 22336 6860
rect 24124 6808 24176 6860
rect 2688 6783 2740 6792
rect 2688 6749 2697 6783
rect 2697 6749 2731 6783
rect 2731 6749 2740 6783
rect 2688 6740 2740 6749
rect 2780 6783 2832 6792
rect 2780 6749 2789 6783
rect 2789 6749 2823 6783
rect 2823 6749 2832 6783
rect 2780 6740 2832 6749
rect 5172 6740 5224 6792
rect 6000 6740 6052 6792
rect 7104 6740 7156 6792
rect 8484 6783 8536 6792
rect 8484 6749 8493 6783
rect 8493 6749 8527 6783
rect 8527 6749 8536 6783
rect 8484 6740 8536 6749
rect 8668 6783 8720 6792
rect 8668 6749 8677 6783
rect 8677 6749 8711 6783
rect 8711 6749 8720 6783
rect 8668 6740 8720 6749
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 7196 6672 7248 6724
rect 7564 6715 7616 6724
rect 7564 6681 7573 6715
rect 7573 6681 7607 6715
rect 7607 6681 7616 6715
rect 7564 6672 7616 6681
rect 8208 6672 8260 6724
rect 11888 6783 11940 6792
rect 11888 6749 11897 6783
rect 11897 6749 11931 6783
rect 11931 6749 11940 6783
rect 11888 6740 11940 6749
rect 13452 6783 13504 6792
rect 13452 6749 13461 6783
rect 13461 6749 13495 6783
rect 13495 6749 13504 6783
rect 13452 6740 13504 6749
rect 14648 6740 14700 6792
rect 10784 6672 10836 6724
rect 15108 6672 15160 6724
rect 15292 6715 15344 6724
rect 15292 6681 15301 6715
rect 15301 6681 15335 6715
rect 15335 6681 15344 6715
rect 15292 6672 15344 6681
rect 18052 6783 18104 6792
rect 18052 6749 18061 6783
rect 18061 6749 18095 6783
rect 18095 6749 18104 6783
rect 18052 6740 18104 6749
rect 18972 6740 19024 6792
rect 19524 6783 19576 6792
rect 19524 6749 19533 6783
rect 19533 6749 19567 6783
rect 19567 6749 19576 6783
rect 19524 6740 19576 6749
rect 20076 6740 20128 6792
rect 21364 6783 21416 6792
rect 21364 6749 21373 6783
rect 21373 6749 21407 6783
rect 21407 6749 21416 6783
rect 21364 6740 21416 6749
rect 21548 6783 21600 6792
rect 21548 6749 21557 6783
rect 21557 6749 21591 6783
rect 21591 6749 21600 6783
rect 21548 6740 21600 6749
rect 22100 6740 22152 6792
rect 22928 6783 22980 6792
rect 16488 6672 16540 6724
rect 19156 6672 19208 6724
rect 22284 6715 22336 6724
rect 22284 6681 22293 6715
rect 22293 6681 22327 6715
rect 22327 6681 22336 6715
rect 22284 6672 22336 6681
rect 22468 6715 22520 6724
rect 22468 6681 22477 6715
rect 22477 6681 22511 6715
rect 22511 6681 22520 6715
rect 22468 6672 22520 6681
rect 22928 6749 22937 6783
rect 22937 6749 22971 6783
rect 22971 6749 22980 6783
rect 22928 6740 22980 6749
rect 23204 6740 23256 6792
rect 24860 6808 24912 6860
rect 24032 6715 24084 6724
rect 24032 6681 24041 6715
rect 24041 6681 24075 6715
rect 24075 6681 24084 6715
rect 24032 6672 24084 6681
rect 1952 6604 2004 6656
rect 5264 6647 5316 6656
rect 5264 6613 5273 6647
rect 5273 6613 5307 6647
rect 5307 6613 5316 6647
rect 5264 6604 5316 6613
rect 7104 6647 7156 6656
rect 7104 6613 7113 6647
rect 7113 6613 7147 6647
rect 7147 6613 7156 6647
rect 7104 6604 7156 6613
rect 8024 6647 8076 6656
rect 8024 6613 8033 6647
rect 8033 6613 8067 6647
rect 8067 6613 8076 6647
rect 8024 6604 8076 6613
rect 8576 6604 8628 6656
rect 11888 6604 11940 6656
rect 12072 6604 12124 6656
rect 12716 6604 12768 6656
rect 13084 6604 13136 6656
rect 14188 6604 14240 6656
rect 14280 6604 14332 6656
rect 16304 6647 16356 6656
rect 16304 6613 16313 6647
rect 16313 6613 16347 6647
rect 16347 6613 16356 6647
rect 16304 6604 16356 6613
rect 17408 6647 17460 6656
rect 17408 6613 17417 6647
rect 17417 6613 17451 6647
rect 17451 6613 17460 6647
rect 17408 6604 17460 6613
rect 18512 6647 18564 6656
rect 18512 6613 18521 6647
rect 18521 6613 18555 6647
rect 18555 6613 18564 6647
rect 18512 6604 18564 6613
rect 18788 6647 18840 6656
rect 18788 6613 18797 6647
rect 18797 6613 18831 6647
rect 18831 6613 18840 6647
rect 18788 6604 18840 6613
rect 19984 6604 20036 6656
rect 20628 6604 20680 6656
rect 20996 6604 21048 6656
rect 21916 6647 21968 6656
rect 21916 6613 21925 6647
rect 21925 6613 21959 6647
rect 21959 6613 21968 6647
rect 21916 6604 21968 6613
rect 22192 6604 22244 6656
rect 25136 6672 25188 6724
rect 25412 6647 25464 6656
rect 25412 6613 25421 6647
rect 25421 6613 25455 6647
rect 25455 6613 25464 6647
rect 25412 6604 25464 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 2596 6400 2648 6452
rect 4160 6400 4212 6452
rect 2780 6332 2832 6384
rect 7012 6400 7064 6452
rect 9680 6443 9732 6452
rect 9680 6409 9689 6443
rect 9689 6409 9723 6443
rect 9723 6409 9732 6443
rect 9680 6400 9732 6409
rect 11520 6443 11572 6452
rect 11520 6409 11529 6443
rect 11529 6409 11563 6443
rect 11563 6409 11572 6443
rect 11520 6400 11572 6409
rect 11704 6400 11756 6452
rect 13360 6443 13412 6452
rect 13360 6409 13369 6443
rect 13369 6409 13403 6443
rect 13403 6409 13412 6443
rect 13360 6400 13412 6409
rect 13728 6400 13780 6452
rect 14280 6400 14332 6452
rect 15568 6400 15620 6452
rect 17868 6400 17920 6452
rect 19156 6443 19208 6452
rect 19156 6409 19165 6443
rect 19165 6409 19199 6443
rect 19199 6409 19208 6443
rect 19156 6400 19208 6409
rect 21640 6400 21692 6452
rect 22008 6400 22060 6452
rect 11336 6332 11388 6384
rect 11796 6332 11848 6384
rect 15016 6332 15068 6384
rect 15936 6332 15988 6384
rect 17132 6332 17184 6384
rect 19248 6332 19300 6384
rect 6000 6264 6052 6316
rect 8576 6307 8628 6316
rect 8576 6273 8585 6307
rect 8585 6273 8619 6307
rect 8619 6273 8628 6307
rect 8576 6264 8628 6273
rect 8668 6307 8720 6316
rect 8668 6273 8677 6307
rect 8677 6273 8711 6307
rect 8711 6273 8720 6307
rect 8668 6264 8720 6273
rect 1768 6196 1820 6248
rect 3608 6196 3660 6248
rect 2964 6128 3016 6180
rect 4988 6196 5040 6248
rect 5356 6239 5408 6248
rect 5356 6205 5365 6239
rect 5365 6205 5399 6239
rect 5399 6205 5408 6239
rect 5356 6196 5408 6205
rect 7564 6196 7616 6248
rect 8392 6196 8444 6248
rect 9680 6196 9732 6248
rect 10876 6196 10928 6248
rect 12716 6196 12768 6248
rect 14188 6239 14240 6248
rect 14188 6205 14222 6239
rect 14222 6205 14240 6239
rect 4804 6103 4856 6112
rect 4804 6069 4813 6103
rect 4813 6069 4847 6103
rect 4847 6069 4856 6103
rect 4804 6060 4856 6069
rect 4988 6103 5040 6112
rect 4988 6069 4997 6103
rect 4997 6069 5031 6103
rect 5031 6069 5040 6103
rect 4988 6060 5040 6069
rect 6000 6103 6052 6112
rect 6000 6069 6009 6103
rect 6009 6069 6043 6103
rect 6043 6069 6052 6103
rect 6000 6060 6052 6069
rect 7196 6103 7248 6112
rect 7196 6069 7205 6103
rect 7205 6069 7239 6103
rect 7239 6069 7248 6103
rect 7196 6060 7248 6069
rect 7656 6103 7708 6112
rect 7656 6069 7665 6103
rect 7665 6069 7699 6103
rect 7699 6069 7708 6103
rect 11060 6128 11112 6180
rect 12900 6171 12952 6180
rect 12900 6137 12909 6171
rect 12909 6137 12943 6171
rect 12943 6137 12952 6171
rect 12900 6128 12952 6137
rect 14188 6196 14240 6205
rect 16304 6264 16356 6316
rect 18512 6264 18564 6316
rect 19156 6264 19208 6316
rect 24676 6400 24728 6452
rect 25412 6400 25464 6452
rect 25596 6400 25648 6452
rect 24860 6332 24912 6384
rect 26240 6332 26292 6384
rect 20260 6196 20312 6248
rect 21916 6196 21968 6248
rect 14832 6128 14884 6180
rect 7656 6060 7708 6069
rect 8116 6103 8168 6112
rect 8116 6069 8125 6103
rect 8125 6069 8159 6103
rect 8159 6069 8168 6103
rect 8116 6060 8168 6069
rect 9864 6060 9916 6112
rect 13636 6060 13688 6112
rect 16028 6128 16080 6180
rect 15292 6103 15344 6112
rect 15292 6069 15301 6103
rect 15301 6069 15335 6103
rect 15335 6069 15344 6103
rect 15292 6060 15344 6069
rect 15936 6103 15988 6112
rect 15936 6069 15945 6103
rect 15945 6069 15979 6103
rect 15979 6069 15988 6103
rect 17960 6128 18012 6180
rect 18788 6128 18840 6180
rect 21640 6128 21692 6180
rect 22376 6128 22428 6180
rect 23756 6264 23808 6316
rect 23664 6196 23716 6248
rect 24860 6196 24912 6248
rect 23480 6171 23532 6180
rect 23480 6137 23489 6171
rect 23489 6137 23523 6171
rect 23523 6137 23532 6171
rect 23480 6128 23532 6137
rect 24768 6128 24820 6180
rect 15936 6060 15988 6069
rect 18972 6060 19024 6112
rect 19524 6103 19576 6112
rect 19524 6069 19533 6103
rect 19533 6069 19567 6103
rect 19567 6069 19576 6103
rect 19524 6060 19576 6069
rect 20720 6060 20772 6112
rect 21824 6103 21876 6112
rect 21824 6069 21833 6103
rect 21833 6069 21867 6103
rect 21867 6069 21876 6103
rect 21824 6060 21876 6069
rect 22928 6103 22980 6112
rect 22928 6069 22937 6103
rect 22937 6069 22971 6103
rect 22971 6069 22980 6103
rect 22928 6060 22980 6069
rect 25412 6103 25464 6112
rect 25412 6069 25421 6103
rect 25421 6069 25455 6103
rect 25455 6069 25464 6103
rect 25412 6060 25464 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 2688 5856 2740 5908
rect 2780 5856 2832 5908
rect 5172 5856 5224 5908
rect 6368 5899 6420 5908
rect 6368 5865 6377 5899
rect 6377 5865 6411 5899
rect 6411 5865 6420 5899
rect 6368 5856 6420 5865
rect 6828 5899 6880 5908
rect 6828 5865 6837 5899
rect 6837 5865 6871 5899
rect 6871 5865 6880 5899
rect 6828 5856 6880 5865
rect 8576 5856 8628 5908
rect 11060 5899 11112 5908
rect 11060 5865 11069 5899
rect 11069 5865 11103 5899
rect 11103 5865 11112 5899
rect 11060 5856 11112 5865
rect 11336 5899 11388 5908
rect 11336 5865 11345 5899
rect 11345 5865 11379 5899
rect 11379 5865 11388 5899
rect 11336 5856 11388 5865
rect 14648 5899 14700 5908
rect 14648 5865 14657 5899
rect 14657 5865 14691 5899
rect 14691 5865 14700 5899
rect 14648 5856 14700 5865
rect 15016 5899 15068 5908
rect 15016 5865 15025 5899
rect 15025 5865 15059 5899
rect 15059 5865 15068 5899
rect 15016 5856 15068 5865
rect 16672 5899 16724 5908
rect 1768 5763 1820 5772
rect 1768 5729 1777 5763
rect 1777 5729 1811 5763
rect 1811 5729 1820 5763
rect 1768 5720 1820 5729
rect 2044 5763 2096 5772
rect 2044 5729 2078 5763
rect 2078 5729 2096 5763
rect 2044 5720 2096 5729
rect 3608 5720 3660 5772
rect 5448 5788 5500 5840
rect 7564 5831 7616 5840
rect 7564 5797 7573 5831
rect 7573 5797 7607 5831
rect 7607 5797 7616 5831
rect 7564 5788 7616 5797
rect 8484 5788 8536 5840
rect 9772 5788 9824 5840
rect 10876 5788 10928 5840
rect 11428 5788 11480 5840
rect 4896 5763 4948 5772
rect 4896 5729 4930 5763
rect 4930 5729 4948 5763
rect 4896 5720 4948 5729
rect 6920 5763 6972 5772
rect 6920 5729 6929 5763
rect 6929 5729 6963 5763
rect 6963 5729 6972 5763
rect 6920 5720 6972 5729
rect 8300 5720 8352 5772
rect 9588 5720 9640 5772
rect 9680 5763 9732 5772
rect 9680 5729 9689 5763
rect 9689 5729 9723 5763
rect 9723 5729 9732 5763
rect 9680 5720 9732 5729
rect 7748 5652 7800 5704
rect 8116 5652 8168 5704
rect 8668 5695 8720 5704
rect 8668 5661 8677 5695
rect 8677 5661 8711 5695
rect 8711 5661 8720 5695
rect 8668 5652 8720 5661
rect 12440 5788 12492 5840
rect 14188 5788 14240 5840
rect 16672 5865 16681 5899
rect 16681 5865 16715 5899
rect 16715 5865 16724 5899
rect 16672 5856 16724 5865
rect 17132 5899 17184 5908
rect 17132 5865 17141 5899
rect 17141 5865 17175 5899
rect 17175 5865 17184 5899
rect 17132 5856 17184 5865
rect 17776 5856 17828 5908
rect 20076 5856 20128 5908
rect 20904 5899 20956 5908
rect 20904 5865 20913 5899
rect 20913 5865 20947 5899
rect 20947 5865 20956 5899
rect 20904 5856 20956 5865
rect 21364 5856 21416 5908
rect 22192 5856 22244 5908
rect 23664 5899 23716 5908
rect 23664 5865 23673 5899
rect 23673 5865 23707 5899
rect 23707 5865 23716 5899
rect 23664 5856 23716 5865
rect 24124 5899 24176 5908
rect 24124 5865 24133 5899
rect 24133 5865 24167 5899
rect 24167 5865 24176 5899
rect 24124 5856 24176 5865
rect 24676 5856 24728 5908
rect 25596 5856 25648 5908
rect 15752 5788 15804 5840
rect 17868 5788 17920 5840
rect 18052 5831 18104 5840
rect 18052 5797 18086 5831
rect 18086 5797 18104 5831
rect 18052 5788 18104 5797
rect 21824 5788 21876 5840
rect 26148 5831 26200 5840
rect 26148 5797 26157 5831
rect 26157 5797 26191 5831
rect 26191 5797 26200 5831
rect 26148 5788 26200 5797
rect 26332 5788 26384 5840
rect 11796 5720 11848 5772
rect 13176 5720 13228 5772
rect 14832 5720 14884 5772
rect 18328 5720 18380 5772
rect 18604 5720 18656 5772
rect 21548 5720 21600 5772
rect 22192 5763 22244 5772
rect 22192 5729 22226 5763
rect 22226 5729 22244 5763
rect 22192 5720 22244 5729
rect 22928 5720 22980 5772
rect 25044 5720 25096 5772
rect 13820 5652 13872 5704
rect 15016 5652 15068 5704
rect 20260 5652 20312 5704
rect 21732 5652 21784 5704
rect 23388 5652 23440 5704
rect 7564 5584 7616 5636
rect 8024 5627 8076 5636
rect 8024 5593 8033 5627
rect 8033 5593 8067 5627
rect 8067 5593 8076 5627
rect 8024 5584 8076 5593
rect 19340 5584 19392 5636
rect 6000 5559 6052 5568
rect 6000 5525 6009 5559
rect 6009 5525 6043 5559
rect 6043 5525 6052 5559
rect 6000 5516 6052 5525
rect 8208 5516 8260 5568
rect 10784 5516 10836 5568
rect 12532 5516 12584 5568
rect 19156 5559 19208 5568
rect 19156 5525 19165 5559
rect 19165 5525 19199 5559
rect 19199 5525 19208 5559
rect 19156 5516 19208 5525
rect 20996 5516 21048 5568
rect 21640 5516 21692 5568
rect 23572 5516 23624 5568
rect 24124 5516 24176 5568
rect 25136 5652 25188 5704
rect 25228 5516 25280 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 4620 5312 4672 5364
rect 5080 5312 5132 5364
rect 8116 5312 8168 5364
rect 11428 5355 11480 5364
rect 11428 5321 11437 5355
rect 11437 5321 11471 5355
rect 11471 5321 11480 5355
rect 11428 5312 11480 5321
rect 11796 5312 11848 5364
rect 2872 5244 2924 5296
rect 12072 5244 12124 5296
rect 12532 5244 12584 5296
rect 4896 5176 4948 5228
rect 3608 5108 3660 5160
rect 4804 5108 4856 5160
rect 6000 5176 6052 5228
rect 9680 5176 9732 5228
rect 9772 5176 9824 5228
rect 14096 5312 14148 5364
rect 15752 5312 15804 5364
rect 16488 5355 16540 5364
rect 16488 5321 16497 5355
rect 16497 5321 16531 5355
rect 16531 5321 16540 5355
rect 16488 5312 16540 5321
rect 16856 5355 16908 5364
rect 16856 5321 16865 5355
rect 16865 5321 16899 5355
rect 16899 5321 16908 5355
rect 16856 5312 16908 5321
rect 17868 5355 17920 5364
rect 17868 5321 17877 5355
rect 17877 5321 17911 5355
rect 17911 5321 17920 5355
rect 17868 5312 17920 5321
rect 20720 5355 20772 5364
rect 20720 5321 20729 5355
rect 20729 5321 20763 5355
rect 20763 5321 20772 5355
rect 20720 5312 20772 5321
rect 21088 5312 21140 5364
rect 22192 5355 22244 5364
rect 22192 5321 22201 5355
rect 22201 5321 22235 5355
rect 22235 5321 22244 5355
rect 22192 5312 22244 5321
rect 23480 5355 23532 5364
rect 23480 5321 23489 5355
rect 23489 5321 23523 5355
rect 23523 5321 23532 5355
rect 23480 5312 23532 5321
rect 25688 5312 25740 5364
rect 26148 5355 26200 5364
rect 26148 5321 26157 5355
rect 26157 5321 26191 5355
rect 26191 5321 26200 5355
rect 26148 5312 26200 5321
rect 14188 5219 14240 5228
rect 14188 5185 14197 5219
rect 14197 5185 14231 5219
rect 14231 5185 14240 5219
rect 14188 5176 14240 5185
rect 14832 5176 14884 5228
rect 20536 5176 20588 5228
rect 22100 5244 22152 5296
rect 23664 5244 23716 5296
rect 24308 5244 24360 5296
rect 25228 5244 25280 5296
rect 25596 5244 25648 5296
rect 25872 5244 25924 5296
rect 5448 5108 5500 5160
rect 8392 5108 8444 5160
rect 10048 5108 10100 5160
rect 7656 5083 7708 5092
rect 7656 5049 7665 5083
rect 7665 5049 7699 5083
rect 7699 5049 7708 5083
rect 7656 5040 7708 5049
rect 8852 5040 8904 5092
rect 9680 5040 9732 5092
rect 18328 5108 18380 5160
rect 20260 5108 20312 5160
rect 27160 5176 27212 5228
rect 24492 5108 24544 5160
rect 26056 5108 26108 5160
rect 1768 5015 1820 5024
rect 1768 4981 1777 5015
rect 1777 4981 1811 5015
rect 1811 4981 1820 5015
rect 1768 4972 1820 4981
rect 2044 4972 2096 5024
rect 2688 5015 2740 5024
rect 2688 4981 2697 5015
rect 2697 4981 2731 5015
rect 2731 4981 2740 5015
rect 2688 4972 2740 4981
rect 5080 5015 5132 5024
rect 5080 4981 5089 5015
rect 5089 4981 5123 5015
rect 5123 4981 5132 5015
rect 5080 4972 5132 4981
rect 5172 4972 5224 5024
rect 6460 4972 6512 5024
rect 6828 4972 6880 5024
rect 9128 5015 9180 5024
rect 9128 4981 9137 5015
rect 9137 4981 9171 5015
rect 9171 4981 9180 5015
rect 9128 4972 9180 4981
rect 9772 5015 9824 5024
rect 9772 4981 9781 5015
rect 9781 4981 9815 5015
rect 9815 4981 9824 5015
rect 9772 4972 9824 4981
rect 9956 5015 10008 5024
rect 9956 4981 9965 5015
rect 9965 4981 9999 5015
rect 9999 4981 10008 5015
rect 9956 4972 10008 4981
rect 11336 4972 11388 5024
rect 14832 5040 14884 5092
rect 19156 5040 19208 5092
rect 25044 5040 25096 5092
rect 25872 5040 25924 5092
rect 12624 5015 12676 5024
rect 12624 4981 12633 5015
rect 12633 4981 12667 5015
rect 12667 4981 12676 5015
rect 12624 4972 12676 4981
rect 12992 5015 13044 5024
rect 12992 4981 13001 5015
rect 13001 4981 13035 5015
rect 13035 4981 13044 5015
rect 12992 4972 13044 4981
rect 13544 5015 13596 5024
rect 13544 4981 13553 5015
rect 13553 4981 13587 5015
rect 13587 4981 13596 5015
rect 13544 4972 13596 4981
rect 19524 4972 19576 5024
rect 20076 4972 20128 5024
rect 20260 5015 20312 5024
rect 20260 4981 20269 5015
rect 20269 4981 20303 5015
rect 20303 4981 20312 5015
rect 20260 4972 20312 4981
rect 23020 5015 23072 5024
rect 23020 4981 23029 5015
rect 23029 4981 23063 5015
rect 23063 4981 23072 5015
rect 23020 4972 23072 4981
rect 23664 5015 23716 5024
rect 23664 4981 23673 5015
rect 23673 4981 23707 5015
rect 23707 4981 23716 5015
rect 23664 4972 23716 4981
rect 25688 4972 25740 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1216 4768 1268 4820
rect 1768 4768 1820 4820
rect 5080 4768 5132 4820
rect 7288 4811 7340 4820
rect 7288 4777 7297 4811
rect 7297 4777 7331 4811
rect 7331 4777 7340 4811
rect 7288 4768 7340 4777
rect 7748 4811 7800 4820
rect 7748 4777 7757 4811
rect 7757 4777 7791 4811
rect 7791 4777 7800 4811
rect 7748 4768 7800 4777
rect 8668 4768 8720 4820
rect 9128 4768 9180 4820
rect 9680 4811 9732 4820
rect 9680 4777 9689 4811
rect 9689 4777 9723 4811
rect 9723 4777 9732 4811
rect 9680 4768 9732 4777
rect 10048 4768 10100 4820
rect 13084 4811 13136 4820
rect 13084 4777 13093 4811
rect 13093 4777 13127 4811
rect 13127 4777 13136 4811
rect 13084 4768 13136 4777
rect 15016 4811 15068 4820
rect 15016 4777 15025 4811
rect 15025 4777 15059 4811
rect 15059 4777 15068 4811
rect 15016 4768 15068 4777
rect 15660 4811 15712 4820
rect 15660 4777 15669 4811
rect 15669 4777 15703 4811
rect 15703 4777 15712 4811
rect 15660 4768 15712 4777
rect 17960 4768 18012 4820
rect 19248 4768 19300 4820
rect 19432 4768 19484 4820
rect 20352 4811 20404 4820
rect 20352 4777 20361 4811
rect 20361 4777 20395 4811
rect 20395 4777 20404 4811
rect 20352 4768 20404 4777
rect 20720 4768 20772 4820
rect 20996 4768 21048 4820
rect 22192 4768 22244 4820
rect 22928 4811 22980 4820
rect 22928 4777 22937 4811
rect 22937 4777 22971 4811
rect 22971 4777 22980 4811
rect 22928 4768 22980 4777
rect 2228 4700 2280 4752
rect 4988 4700 5040 4752
rect 5540 4700 5592 4752
rect 2872 4632 2924 4684
rect 5264 4632 5316 4684
rect 6460 4700 6512 4752
rect 11520 4700 11572 4752
rect 12072 4700 12124 4752
rect 17316 4700 17368 4752
rect 23112 4700 23164 4752
rect 24124 4768 24176 4820
rect 24676 4768 24728 4820
rect 25136 4811 25188 4820
rect 25136 4777 25145 4811
rect 25145 4777 25179 4811
rect 25179 4777 25188 4811
rect 25136 4768 25188 4777
rect 26332 4768 26384 4820
rect 25504 4700 25556 4752
rect 6000 4632 6052 4684
rect 8484 4675 8536 4684
rect 8484 4641 8493 4675
rect 8493 4641 8527 4675
rect 8527 4641 8536 4675
rect 8484 4632 8536 4641
rect 10968 4632 11020 4684
rect 11428 4675 11480 4684
rect 11428 4641 11437 4675
rect 11437 4641 11471 4675
rect 11471 4641 11480 4675
rect 11428 4632 11480 4641
rect 2044 4564 2096 4616
rect 3792 4564 3844 4616
rect 2596 4496 2648 4548
rect 2780 4496 2832 4548
rect 8668 4539 8720 4548
rect 8668 4505 8677 4539
rect 8677 4505 8711 4539
rect 8711 4505 8720 4539
rect 8668 4496 8720 4505
rect 4804 4428 4856 4480
rect 5448 4471 5500 4480
rect 5448 4437 5457 4471
rect 5457 4437 5491 4471
rect 5491 4437 5500 4471
rect 5448 4428 5500 4437
rect 8300 4428 8352 4480
rect 10232 4607 10284 4616
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 12256 4632 12308 4684
rect 16212 4632 16264 4684
rect 16488 4632 16540 4684
rect 17776 4632 17828 4684
rect 19432 4675 19484 4684
rect 19432 4641 19441 4675
rect 19441 4641 19475 4675
rect 19475 4641 19484 4675
rect 19432 4632 19484 4641
rect 19984 4632 20036 4684
rect 20904 4632 20956 4684
rect 23296 4632 23348 4684
rect 10232 4564 10284 4573
rect 14096 4607 14148 4616
rect 14096 4573 14105 4607
rect 14105 4573 14139 4607
rect 14139 4573 14148 4607
rect 14096 4564 14148 4573
rect 14188 4607 14240 4616
rect 14188 4573 14197 4607
rect 14197 4573 14231 4607
rect 14231 4573 14240 4607
rect 15936 4607 15988 4616
rect 14188 4564 14240 4573
rect 15936 4573 15945 4607
rect 15945 4573 15979 4607
rect 15979 4573 15988 4607
rect 15936 4564 15988 4573
rect 17408 4564 17460 4616
rect 11428 4496 11480 4548
rect 13636 4539 13688 4548
rect 13636 4505 13645 4539
rect 13645 4505 13679 4539
rect 13679 4505 13688 4539
rect 13636 4496 13688 4505
rect 15292 4539 15344 4548
rect 15292 4505 15301 4539
rect 15301 4505 15335 4539
rect 15335 4505 15344 4539
rect 15292 4496 15344 4505
rect 17868 4496 17920 4548
rect 19524 4564 19576 4616
rect 22376 4564 22428 4616
rect 25136 4564 25188 4616
rect 24492 4496 24544 4548
rect 12348 4428 12400 4480
rect 12992 4428 13044 4480
rect 17040 4471 17092 4480
rect 17040 4437 17049 4471
rect 17049 4437 17083 4471
rect 17083 4437 17092 4471
rect 17040 4428 17092 4437
rect 18512 4471 18564 4480
rect 18512 4437 18521 4471
rect 18521 4437 18555 4471
rect 18555 4437 18564 4471
rect 18512 4428 18564 4437
rect 22100 4428 22152 4480
rect 23664 4471 23716 4480
rect 23664 4437 23673 4471
rect 23673 4437 23707 4471
rect 23707 4437 23716 4471
rect 23664 4428 23716 4437
rect 24860 4428 24912 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 2044 4267 2096 4276
rect 2044 4233 2053 4267
rect 2053 4233 2087 4267
rect 2087 4233 2096 4267
rect 2044 4224 2096 4233
rect 5448 4224 5500 4276
rect 9864 4267 9916 4276
rect 9864 4233 9873 4267
rect 9873 4233 9907 4267
rect 9907 4233 9916 4267
rect 9864 4224 9916 4233
rect 11520 4267 11572 4276
rect 11520 4233 11529 4267
rect 11529 4233 11563 4267
rect 11563 4233 11572 4267
rect 11520 4224 11572 4233
rect 2688 4156 2740 4208
rect 2044 4088 2096 4140
rect 2320 4088 2372 4140
rect 3332 4131 3384 4140
rect 3332 4097 3341 4131
rect 3341 4097 3375 4131
rect 3375 4097 3384 4131
rect 3332 4088 3384 4097
rect 4804 4156 4856 4208
rect 4988 4156 5040 4208
rect 8852 4156 8904 4208
rect 9404 4156 9456 4208
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 12716 4156 12768 4208
rect 11152 4088 11204 4140
rect 11612 4088 11664 4140
rect 2964 4020 3016 4072
rect 1860 3952 1912 4004
rect 7748 4020 7800 4072
rect 8392 4020 8444 4072
rect 9956 4020 10008 4072
rect 11980 4020 12032 4072
rect 3424 3952 3476 4004
rect 3884 3995 3936 4004
rect 3884 3961 3893 3995
rect 3893 3961 3927 3995
rect 3927 3961 3936 3995
rect 3884 3952 3936 3961
rect 5172 3952 5224 4004
rect 6000 3952 6052 4004
rect 9404 3952 9456 4004
rect 10232 3952 10284 4004
rect 10692 3952 10744 4004
rect 11336 3952 11388 4004
rect 1676 3927 1728 3936
rect 1676 3893 1685 3927
rect 1685 3893 1719 3927
rect 1719 3893 1728 3927
rect 1676 3884 1728 3893
rect 2872 3927 2924 3936
rect 2872 3893 2881 3927
rect 2881 3893 2915 3927
rect 2915 3893 2924 3927
rect 2872 3884 2924 3893
rect 4252 3927 4304 3936
rect 4252 3893 4261 3927
rect 4261 3893 4295 3927
rect 4295 3893 4304 3927
rect 4252 3884 4304 3893
rect 4712 3884 4764 3936
rect 6460 3884 6512 3936
rect 7380 3927 7432 3936
rect 7380 3893 7389 3927
rect 7389 3893 7423 3927
rect 7423 3893 7432 3927
rect 7380 3884 7432 3893
rect 7656 3927 7708 3936
rect 7656 3893 7665 3927
rect 7665 3893 7699 3927
rect 7699 3893 7708 3927
rect 7656 3884 7708 3893
rect 10048 3884 10100 3936
rect 10968 3884 11020 3936
rect 12072 3884 12124 3936
rect 14188 4224 14240 4276
rect 17408 4267 17460 4276
rect 17408 4233 17417 4267
rect 17417 4233 17451 4267
rect 17451 4233 17460 4267
rect 17408 4224 17460 4233
rect 15936 4199 15988 4208
rect 15936 4165 15945 4199
rect 15945 4165 15979 4199
rect 15979 4165 15988 4199
rect 15936 4156 15988 4165
rect 19248 4224 19300 4276
rect 22928 4224 22980 4276
rect 24676 4267 24728 4276
rect 24676 4233 24685 4267
rect 24685 4233 24719 4267
rect 24719 4233 24728 4267
rect 24676 4224 24728 4233
rect 25136 4267 25188 4276
rect 25136 4233 25145 4267
rect 25145 4233 25179 4267
rect 25179 4233 25188 4267
rect 25136 4224 25188 4233
rect 16856 4131 16908 4140
rect 16856 4097 16865 4131
rect 16865 4097 16899 4131
rect 16899 4097 16908 4131
rect 16856 4088 16908 4097
rect 12624 4020 12676 4072
rect 13728 4020 13780 4072
rect 14740 4020 14792 4072
rect 18788 4063 18840 4072
rect 12348 3952 12400 4004
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 14280 3952 14332 4004
rect 12440 3884 12492 3893
rect 17500 3952 17552 4004
rect 18788 4029 18797 4063
rect 18797 4029 18831 4063
rect 18831 4029 18840 4063
rect 18788 4020 18840 4029
rect 19432 4156 19484 4208
rect 20536 4131 20588 4140
rect 20536 4097 20545 4131
rect 20545 4097 20579 4131
rect 20579 4097 20588 4131
rect 20536 4088 20588 4097
rect 22284 4156 22336 4208
rect 25044 4156 25096 4208
rect 22376 4088 22428 4140
rect 23112 4088 23164 4140
rect 23480 4088 23532 4140
rect 19340 4020 19392 4072
rect 20628 4020 20680 4072
rect 24124 4063 24176 4072
rect 24124 4029 24133 4063
rect 24133 4029 24167 4063
rect 24167 4029 24176 4063
rect 24124 4020 24176 4029
rect 25228 4063 25280 4072
rect 25228 4029 25237 4063
rect 25237 4029 25271 4063
rect 25271 4029 25280 4063
rect 25228 4020 25280 4029
rect 26332 4063 26384 4072
rect 26332 4029 26341 4063
rect 26341 4029 26375 4063
rect 26375 4029 26384 4063
rect 26332 4020 26384 4029
rect 16304 3884 16356 3936
rect 16764 3927 16816 3936
rect 16764 3893 16773 3927
rect 16773 3893 16807 3927
rect 16807 3893 16816 3927
rect 16764 3884 16816 3893
rect 17776 3927 17828 3936
rect 17776 3893 17785 3927
rect 17785 3893 17819 3927
rect 17819 3893 17828 3927
rect 17776 3884 17828 3893
rect 18512 3884 18564 3936
rect 19340 3884 19392 3936
rect 20720 3952 20772 4004
rect 19984 3884 20036 3936
rect 21088 3884 21140 3936
rect 24032 3995 24084 4004
rect 24032 3961 24041 3995
rect 24041 3961 24075 3995
rect 24075 3961 24084 3995
rect 24032 3952 24084 3961
rect 24768 3952 24820 4004
rect 24952 3952 25004 4004
rect 21364 3884 21416 3936
rect 23480 3927 23532 3936
rect 23480 3893 23489 3927
rect 23489 3893 23523 3927
rect 23523 3893 23532 3927
rect 23480 3884 23532 3893
rect 23572 3884 23624 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1400 3723 1452 3732
rect 1400 3689 1409 3723
rect 1409 3689 1443 3723
rect 1443 3689 1452 3723
rect 1400 3680 1452 3689
rect 1676 3680 1728 3732
rect 2964 3723 3016 3732
rect 1584 3612 1636 3664
rect 2964 3689 2973 3723
rect 2973 3689 3007 3723
rect 3007 3689 3016 3723
rect 2964 3680 3016 3689
rect 3792 3723 3844 3732
rect 3792 3689 3801 3723
rect 3801 3689 3835 3723
rect 3835 3689 3844 3723
rect 3792 3680 3844 3689
rect 4068 3723 4120 3732
rect 4068 3689 4077 3723
rect 4077 3689 4111 3723
rect 4111 3689 4120 3723
rect 4068 3680 4120 3689
rect 5540 3723 5592 3732
rect 5540 3689 5549 3723
rect 5549 3689 5583 3723
rect 5583 3689 5592 3723
rect 5540 3680 5592 3689
rect 7380 3680 7432 3732
rect 8392 3680 8444 3732
rect 8484 3680 8536 3732
rect 9128 3680 9180 3732
rect 2872 3612 2924 3664
rect 6092 3612 6144 3664
rect 9588 3612 9640 3664
rect 9864 3612 9916 3664
rect 11336 3612 11388 3664
rect 11520 3612 11572 3664
rect 11796 3612 11848 3664
rect 12716 3612 12768 3664
rect 14372 3680 14424 3732
rect 14648 3723 14700 3732
rect 14648 3689 14657 3723
rect 14657 3689 14691 3723
rect 14691 3689 14700 3723
rect 14648 3680 14700 3689
rect 16764 3680 16816 3732
rect 19524 3723 19576 3732
rect 19524 3689 19533 3723
rect 19533 3689 19567 3723
rect 19567 3689 19576 3723
rect 19524 3680 19576 3689
rect 20168 3680 20220 3732
rect 20904 3723 20956 3732
rect 20904 3689 20913 3723
rect 20913 3689 20947 3723
rect 20947 3689 20956 3723
rect 20904 3680 20956 3689
rect 21916 3680 21968 3732
rect 22376 3723 22428 3732
rect 22376 3689 22385 3723
rect 22385 3689 22419 3723
rect 22419 3689 22428 3723
rect 22376 3680 22428 3689
rect 23020 3680 23072 3732
rect 24124 3680 24176 3732
rect 25780 3723 25832 3732
rect 25780 3689 25789 3723
rect 25789 3689 25823 3723
rect 25823 3689 25832 3723
rect 25780 3680 25832 3689
rect 26148 3723 26200 3732
rect 26148 3689 26157 3723
rect 26157 3689 26191 3723
rect 26191 3689 26200 3723
rect 26148 3680 26200 3689
rect 13452 3612 13504 3664
rect 15936 3612 15988 3664
rect 17316 3655 17368 3664
rect 17316 3621 17325 3655
rect 17325 3621 17359 3655
rect 17359 3621 17368 3655
rect 17316 3612 17368 3621
rect 18880 3612 18932 3664
rect 19340 3612 19392 3664
rect 21640 3612 21692 3664
rect 22928 3655 22980 3664
rect 22928 3621 22937 3655
rect 22937 3621 22971 3655
rect 22971 3621 22980 3655
rect 22928 3612 22980 3621
rect 24492 3655 24544 3664
rect 24492 3621 24501 3655
rect 24501 3621 24535 3655
rect 24535 3621 24544 3655
rect 24492 3612 24544 3621
rect 24768 3612 24820 3664
rect 3148 3544 3200 3596
rect 2228 3476 2280 3528
rect 1400 3340 1452 3392
rect 1952 3340 2004 3392
rect 5264 3544 5316 3596
rect 6000 3544 6052 3596
rect 6460 3544 6512 3596
rect 8024 3544 8076 3596
rect 9772 3544 9824 3596
rect 10968 3544 11020 3596
rect 11428 3544 11480 3596
rect 13084 3544 13136 3596
rect 14740 3544 14792 3596
rect 16396 3544 16448 3596
rect 16764 3544 16816 3596
rect 17592 3544 17644 3596
rect 19064 3544 19116 3596
rect 21272 3587 21324 3596
rect 21272 3553 21281 3587
rect 21281 3553 21315 3587
rect 21315 3553 21324 3587
rect 21272 3544 21324 3553
rect 22468 3544 22520 3596
rect 4712 3519 4764 3528
rect 4712 3485 4721 3519
rect 4721 3485 4755 3519
rect 4755 3485 4764 3519
rect 4712 3476 4764 3485
rect 5448 3476 5500 3528
rect 9404 3476 9456 3528
rect 11060 3476 11112 3528
rect 7288 3451 7340 3460
rect 7288 3417 7297 3451
rect 7297 3417 7331 3451
rect 7331 3417 7340 3451
rect 7288 3408 7340 3417
rect 9680 3451 9732 3460
rect 9680 3417 9689 3451
rect 9689 3417 9723 3451
rect 9723 3417 9732 3451
rect 9680 3408 9732 3417
rect 10048 3408 10100 3460
rect 10876 3408 10928 3460
rect 16856 3476 16908 3528
rect 6828 3340 6880 3392
rect 10784 3340 10836 3392
rect 11060 3383 11112 3392
rect 11060 3349 11069 3383
rect 11069 3349 11103 3383
rect 11103 3349 11112 3383
rect 12808 3408 12860 3460
rect 17500 3451 17552 3460
rect 17500 3417 17509 3451
rect 17509 3417 17543 3451
rect 17543 3417 17552 3451
rect 17500 3408 17552 3417
rect 17776 3476 17828 3528
rect 18328 3476 18380 3528
rect 20536 3476 20588 3528
rect 20720 3519 20772 3528
rect 20720 3485 20729 3519
rect 20729 3485 20763 3519
rect 20763 3485 20772 3519
rect 21548 3519 21600 3528
rect 20720 3476 20772 3485
rect 21548 3485 21557 3519
rect 21557 3485 21591 3519
rect 21591 3485 21600 3519
rect 21548 3476 21600 3485
rect 18604 3408 18656 3460
rect 22928 3476 22980 3528
rect 24676 3519 24728 3528
rect 24676 3485 24685 3519
rect 24685 3485 24719 3519
rect 24719 3485 24728 3519
rect 24676 3476 24728 3485
rect 14372 3383 14424 3392
rect 11060 3340 11112 3349
rect 14372 3349 14381 3383
rect 14381 3349 14415 3383
rect 14415 3349 14424 3383
rect 14372 3340 14424 3349
rect 15660 3340 15712 3392
rect 23756 3383 23808 3392
rect 23756 3349 23765 3383
rect 23765 3349 23799 3383
rect 23799 3349 23808 3383
rect 23756 3340 23808 3349
rect 24032 3383 24084 3392
rect 24032 3349 24041 3383
rect 24041 3349 24075 3383
rect 24075 3349 24084 3383
rect 24032 3340 24084 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1492 3136 1544 3188
rect 1676 3000 1728 3052
rect 2228 3000 2280 3052
rect 1768 2975 1820 2984
rect 1768 2941 1777 2975
rect 1777 2941 1811 2975
rect 1811 2941 1820 2975
rect 3332 3136 3384 3188
rect 4712 3136 4764 3188
rect 5264 3179 5316 3188
rect 5264 3145 5273 3179
rect 5273 3145 5307 3179
rect 5307 3145 5316 3179
rect 5264 3136 5316 3145
rect 6092 3136 6144 3188
rect 8208 3136 8260 3188
rect 9864 3179 9916 3188
rect 9864 3145 9873 3179
rect 9873 3145 9907 3179
rect 9907 3145 9916 3179
rect 12440 3179 12492 3188
rect 9864 3136 9916 3145
rect 7748 3068 7800 3120
rect 7656 3000 7708 3052
rect 9772 3068 9824 3120
rect 11336 3068 11388 3120
rect 11520 3068 11572 3120
rect 1768 2932 1820 2941
rect 3148 2932 3200 2984
rect 3608 2932 3660 2984
rect 3792 2975 3844 2984
rect 3792 2941 3826 2975
rect 3826 2941 3844 2975
rect 3792 2932 3844 2941
rect 7196 2932 7248 2984
rect 8024 2975 8076 2984
rect 8024 2941 8033 2975
rect 8033 2941 8067 2975
rect 8067 2941 8076 2975
rect 8024 2932 8076 2941
rect 8392 2932 8444 2984
rect 12440 3145 12449 3179
rect 12449 3145 12483 3179
rect 12483 3145 12492 3179
rect 12440 3136 12492 3145
rect 14832 3179 14884 3188
rect 14832 3145 14841 3179
rect 14841 3145 14875 3179
rect 14875 3145 14884 3179
rect 14832 3136 14884 3145
rect 8760 2975 8812 2984
rect 8760 2941 8783 2975
rect 8783 2941 8812 2975
rect 1584 2864 1636 2916
rect 2504 2864 2556 2916
rect 664 2796 716 2848
rect 5080 2796 5132 2848
rect 6276 2864 6328 2916
rect 6644 2907 6696 2916
rect 6644 2873 6653 2907
rect 6653 2873 6687 2907
rect 6687 2873 6696 2907
rect 6644 2864 6696 2873
rect 7932 2864 7984 2916
rect 8760 2932 8812 2941
rect 9956 2932 10008 2984
rect 11060 2932 11112 2984
rect 14372 3000 14424 3052
rect 15660 3136 15712 3188
rect 15936 3179 15988 3188
rect 15936 3145 15945 3179
rect 15945 3145 15979 3179
rect 15979 3145 15988 3179
rect 15936 3136 15988 3145
rect 18052 3179 18104 3188
rect 18052 3145 18061 3179
rect 18061 3145 18095 3179
rect 18095 3145 18104 3179
rect 18052 3136 18104 3145
rect 19524 3179 19576 3188
rect 19524 3145 19533 3179
rect 19533 3145 19567 3179
rect 19567 3145 19576 3179
rect 19524 3136 19576 3145
rect 20536 3136 20588 3188
rect 21180 3179 21232 3188
rect 21180 3145 21189 3179
rect 21189 3145 21223 3179
rect 21223 3145 21232 3179
rect 21180 3136 21232 3145
rect 25044 3179 25096 3188
rect 25044 3145 25053 3179
rect 25053 3145 25087 3179
rect 25087 3145 25096 3179
rect 25044 3136 25096 3145
rect 26332 3179 26384 3188
rect 26332 3145 26341 3179
rect 26341 3145 26375 3179
rect 26375 3145 26384 3179
rect 26332 3136 26384 3145
rect 16212 3068 16264 3120
rect 19064 3111 19116 3120
rect 19064 3077 19073 3111
rect 19073 3077 19107 3111
rect 19107 3077 19116 3111
rect 19064 3068 19116 3077
rect 19616 3111 19668 3120
rect 19616 3077 19625 3111
rect 19625 3077 19659 3111
rect 19659 3077 19668 3111
rect 19616 3068 19668 3077
rect 12808 2975 12860 2984
rect 12808 2941 12817 2975
rect 12817 2941 12851 2975
rect 12851 2941 12860 2975
rect 12808 2932 12860 2941
rect 13912 2932 13964 2984
rect 15292 2975 15344 2984
rect 15292 2941 15301 2975
rect 15301 2941 15335 2975
rect 15335 2941 15344 2975
rect 15292 2932 15344 2941
rect 16764 3000 16816 3052
rect 18604 3043 18656 3052
rect 18604 3009 18613 3043
rect 18613 3009 18647 3043
rect 18647 3009 18656 3043
rect 18604 3000 18656 3009
rect 20168 3043 20220 3052
rect 20168 3009 20177 3043
rect 20177 3009 20211 3043
rect 20211 3009 20220 3043
rect 20168 3000 20220 3009
rect 20812 3000 20864 3052
rect 21640 3043 21692 3052
rect 16304 2932 16356 2984
rect 16488 2975 16540 2984
rect 16488 2941 16497 2975
rect 16497 2941 16531 2975
rect 16531 2941 16540 2975
rect 16488 2932 16540 2941
rect 18880 2932 18932 2984
rect 20076 2975 20128 2984
rect 20076 2941 20085 2975
rect 20085 2941 20119 2975
rect 20119 2941 20128 2975
rect 20076 2932 20128 2941
rect 20720 2932 20772 2984
rect 9588 2864 9640 2916
rect 12716 2864 12768 2916
rect 13636 2864 13688 2916
rect 15568 2864 15620 2916
rect 18236 2864 18288 2916
rect 21640 3009 21649 3043
rect 21649 3009 21683 3043
rect 21683 3009 21692 3043
rect 21640 3000 21692 3009
rect 21456 2932 21508 2984
rect 22928 3000 22980 3052
rect 23020 3000 23072 3052
rect 23480 3000 23532 3052
rect 24676 3043 24728 3052
rect 24676 3009 24685 3043
rect 24685 3009 24719 3043
rect 24719 3009 24728 3043
rect 24676 3000 24728 3009
rect 23756 2932 23808 2984
rect 24032 2975 24084 2984
rect 24032 2941 24041 2975
rect 24041 2941 24075 2975
rect 24075 2941 24084 2975
rect 24032 2932 24084 2941
rect 25320 2932 25372 2984
rect 23940 2864 23992 2916
rect 25504 2907 25556 2916
rect 25504 2873 25513 2907
rect 25513 2873 25547 2907
rect 25547 2873 25556 2907
rect 25504 2864 25556 2873
rect 10968 2796 11020 2848
rect 12808 2796 12860 2848
rect 13452 2839 13504 2848
rect 13452 2805 13461 2839
rect 13461 2805 13495 2839
rect 13495 2805 13504 2839
rect 13452 2796 13504 2805
rect 14924 2839 14976 2848
rect 14924 2805 14933 2839
rect 14933 2805 14967 2839
rect 14967 2805 14976 2839
rect 14924 2796 14976 2805
rect 17500 2839 17552 2848
rect 17500 2805 17509 2839
rect 17509 2805 17543 2839
rect 17543 2805 17552 2839
rect 17500 2796 17552 2805
rect 17776 2796 17828 2848
rect 18144 2796 18196 2848
rect 18420 2839 18472 2848
rect 18420 2805 18429 2839
rect 18429 2805 18463 2839
rect 18463 2805 18472 2839
rect 18420 2796 18472 2805
rect 20076 2796 20128 2848
rect 20260 2796 20312 2848
rect 23020 2839 23072 2848
rect 23020 2805 23029 2839
rect 23029 2805 23063 2839
rect 23063 2805 23072 2839
rect 23020 2796 23072 2805
rect 23664 2839 23716 2848
rect 23664 2805 23673 2839
rect 23673 2805 23707 2839
rect 23707 2805 23716 2839
rect 23664 2796 23716 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 2136 2592 2188 2644
rect 3792 2592 3844 2644
rect 6000 2592 6052 2644
rect 7196 2635 7248 2644
rect 7196 2601 7205 2635
rect 7205 2601 7239 2635
rect 7239 2601 7248 2635
rect 7196 2592 7248 2601
rect 8852 2635 8904 2644
rect 8852 2601 8861 2635
rect 8861 2601 8895 2635
rect 8895 2601 8904 2635
rect 8852 2592 8904 2601
rect 9404 2592 9456 2644
rect 9588 2592 9640 2644
rect 1676 2524 1728 2576
rect 4620 2524 4672 2576
rect 5080 2524 5132 2576
rect 1400 2456 1452 2508
rect 3148 2456 3200 2508
rect 8392 2524 8444 2576
rect 9772 2524 9824 2576
rect 7748 2499 7800 2508
rect 2228 2388 2280 2440
rect 2964 2431 3016 2440
rect 2964 2397 2973 2431
rect 2973 2397 3007 2431
rect 3007 2397 3016 2431
rect 2964 2388 3016 2397
rect 7748 2465 7782 2499
rect 7782 2465 7800 2499
rect 7748 2456 7800 2465
rect 14004 2635 14056 2644
rect 11796 2524 11848 2576
rect 14004 2601 14013 2635
rect 14013 2601 14047 2635
rect 14047 2601 14056 2635
rect 14004 2592 14056 2601
rect 16396 2592 16448 2644
rect 18144 2635 18196 2644
rect 18144 2601 18153 2635
rect 18153 2601 18187 2635
rect 18187 2601 18196 2635
rect 18144 2592 18196 2601
rect 18696 2635 18748 2644
rect 18696 2601 18705 2635
rect 18705 2601 18739 2635
rect 18739 2601 18748 2635
rect 18696 2592 18748 2601
rect 14556 2567 14608 2576
rect 10600 2499 10652 2508
rect 10600 2465 10634 2499
rect 10634 2465 10652 2499
rect 10600 2456 10652 2465
rect 14556 2533 14565 2567
rect 14565 2533 14599 2567
rect 14599 2533 14608 2567
rect 14556 2524 14608 2533
rect 5448 2295 5500 2304
rect 5448 2261 5457 2295
rect 5457 2261 5491 2295
rect 5491 2261 5500 2295
rect 5448 2252 5500 2261
rect 14464 2388 14516 2440
rect 13728 2320 13780 2372
rect 15292 2295 15344 2304
rect 15292 2261 15301 2295
rect 15301 2261 15335 2295
rect 15335 2261 15344 2295
rect 16396 2388 16448 2440
rect 16764 2456 16816 2508
rect 18328 2456 18380 2508
rect 20168 2592 20220 2644
rect 20720 2592 20772 2644
rect 21640 2635 21692 2644
rect 21640 2601 21649 2635
rect 21649 2601 21683 2635
rect 21683 2601 21692 2635
rect 21640 2592 21692 2601
rect 22744 2635 22796 2644
rect 22744 2601 22753 2635
rect 22753 2601 22787 2635
rect 22787 2601 22796 2635
rect 22744 2592 22796 2601
rect 23940 2592 23992 2644
rect 20904 2567 20956 2576
rect 20904 2533 20913 2567
rect 20913 2533 20947 2567
rect 20947 2533 20956 2567
rect 20904 2524 20956 2533
rect 19984 2499 20036 2508
rect 19984 2465 19993 2499
rect 19993 2465 20027 2499
rect 20027 2465 20036 2499
rect 19984 2456 20036 2465
rect 24768 2592 24820 2644
rect 26424 2635 26476 2644
rect 26424 2601 26433 2635
rect 26433 2601 26467 2635
rect 26467 2601 26476 2635
rect 26424 2592 26476 2601
rect 23480 2456 23532 2508
rect 21732 2431 21784 2440
rect 21732 2397 21741 2431
rect 21741 2397 21775 2431
rect 21775 2397 21784 2431
rect 21732 2388 21784 2397
rect 23020 2388 23072 2440
rect 23664 2388 23716 2440
rect 24676 2431 24728 2440
rect 24676 2397 24685 2431
rect 24685 2397 24719 2431
rect 24719 2397 24728 2431
rect 24676 2388 24728 2397
rect 25596 2431 25648 2440
rect 25596 2397 25605 2431
rect 25605 2397 25639 2431
rect 25639 2397 25648 2431
rect 25596 2388 25648 2397
rect 15292 2252 15344 2261
rect 17132 2252 17184 2304
rect 17592 2295 17644 2304
rect 17592 2261 17601 2295
rect 17601 2261 17635 2295
rect 17635 2261 17644 2295
rect 17592 2252 17644 2261
rect 18328 2295 18380 2304
rect 18328 2261 18337 2295
rect 18337 2261 18371 2295
rect 18371 2261 18380 2295
rect 18328 2252 18380 2261
rect 20168 2295 20220 2304
rect 20168 2261 20177 2295
rect 20177 2261 20211 2295
rect 20211 2261 20220 2295
rect 20168 2252 20220 2261
rect 23020 2295 23072 2304
rect 23020 2261 23029 2295
rect 23029 2261 23063 2295
rect 23063 2261 23072 2295
rect 23020 2252 23072 2261
rect 23480 2295 23532 2304
rect 23480 2261 23489 2295
rect 23489 2261 23523 2295
rect 23523 2261 23532 2295
rect 23480 2252 23532 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 11520 2048 11572 2100
rect 13452 2048 13504 2100
rect 12532 1912 12584 1964
rect 18788 1912 18840 1964
rect 22652 552 22704 604
rect 22744 552 22796 604
rect 23756 552 23808 604
rect 25688 552 25740 604
<< metal2 >>
rect 294 27520 350 28000
rect 846 27520 902 28000
rect 1398 27520 1454 28000
rect 2042 27520 2098 28000
rect 2594 27520 2650 28000
rect 3146 27520 3202 28000
rect 3514 27704 3570 27713
rect 3514 27639 3570 27648
rect 3528 27606 3556 27639
rect 3516 27600 3568 27606
rect 3516 27542 3568 27548
rect 3790 27520 3846 28000
rect 4342 27520 4398 28000
rect 4894 27520 4950 28000
rect 5538 27520 5594 28000
rect 6090 27520 6146 28000
rect 6642 27520 6698 28000
rect 7286 27520 7342 28000
rect 7838 27520 7894 28000
rect 8390 27520 8446 28000
rect 9034 27520 9090 28000
rect 9128 27600 9180 27606
rect 9128 27542 9180 27548
rect 308 22273 336 27520
rect 860 23361 888 27520
rect 1412 27282 1440 27520
rect 1412 27254 1900 27282
rect 1674 27160 1730 27169
rect 1674 27095 1730 27104
rect 1490 26616 1546 26625
rect 1490 26551 1546 26560
rect 1504 24410 1532 26551
rect 1582 25392 1638 25401
rect 1582 25327 1638 25336
rect 1596 24954 1624 25327
rect 1584 24948 1636 24954
rect 1584 24890 1636 24896
rect 1582 24848 1638 24857
rect 1582 24783 1638 24792
rect 1492 24404 1544 24410
rect 1492 24346 1544 24352
rect 1398 24168 1454 24177
rect 1398 24103 1454 24112
rect 846 23352 902 23361
rect 846 23287 902 23296
rect 294 22264 350 22273
rect 294 22199 350 22208
rect 1412 21962 1440 24103
rect 1490 23080 1546 23089
rect 1490 23015 1546 23024
rect 1400 21956 1452 21962
rect 1400 21898 1452 21904
rect 1504 21690 1532 23015
rect 1596 22778 1624 24783
rect 1688 23866 1716 27095
rect 1676 23860 1728 23866
rect 1676 23802 1728 23808
rect 1676 23656 1728 23662
rect 1676 23598 1728 23604
rect 1688 23118 1716 23598
rect 1676 23112 1728 23118
rect 1674 23080 1676 23089
rect 1728 23080 1730 23089
rect 1674 23015 1730 23024
rect 1584 22772 1636 22778
rect 1584 22714 1636 22720
rect 1582 22536 1638 22545
rect 1582 22471 1638 22480
rect 1492 21684 1544 21690
rect 1492 21626 1544 21632
rect 1596 21146 1624 22471
rect 1584 21140 1636 21146
rect 1584 21082 1636 21088
rect 1872 20641 1900 27254
rect 2056 24426 2084 27520
rect 2608 27418 2636 27520
rect 2516 27390 2636 27418
rect 2228 25492 2280 25498
rect 2228 25434 2280 25440
rect 2240 24614 2268 25434
rect 2228 24608 2280 24614
rect 2228 24550 2280 24556
rect 2056 24398 2176 24426
rect 2044 24268 2096 24274
rect 2044 24210 2096 24216
rect 2056 23526 2084 24210
rect 2044 23520 2096 23526
rect 2044 23462 2096 23468
rect 2056 23225 2084 23462
rect 2042 23216 2098 23225
rect 2042 23151 2098 23160
rect 2148 22545 2176 24398
rect 2134 22536 2190 22545
rect 2134 22471 2190 22480
rect 2136 22432 2188 22438
rect 2136 22374 2188 22380
rect 2042 21584 2098 21593
rect 2042 21519 2044 21528
rect 2096 21519 2098 21528
rect 2044 21490 2096 21496
rect 2044 21004 2096 21010
rect 2044 20946 2096 20952
rect 1950 20768 2006 20777
rect 1950 20703 2006 20712
rect 1858 20632 1914 20641
rect 1858 20567 1914 20576
rect 1400 20256 1452 20262
rect 1400 20198 1452 20204
rect 1124 18692 1176 18698
rect 1124 18634 1176 18640
rect 848 18352 900 18358
rect 848 18294 900 18300
rect 860 13161 888 18294
rect 1030 17232 1086 17241
rect 1030 17167 1086 17176
rect 940 16244 992 16250
rect 940 16186 992 16192
rect 846 13152 902 13161
rect 846 13087 902 13096
rect 860 11257 888 13087
rect 952 11937 980 16186
rect 938 11928 994 11937
rect 938 11863 994 11872
rect 846 11248 902 11257
rect 846 11183 902 11192
rect 1044 10674 1072 17167
rect 1136 13705 1164 18634
rect 1412 16697 1440 20198
rect 1872 18970 1900 20567
rect 1860 18964 1912 18970
rect 1860 18906 1912 18912
rect 1964 18902 1992 20703
rect 2056 20534 2084 20946
rect 2044 20528 2096 20534
rect 2042 20496 2044 20505
rect 2096 20496 2098 20505
rect 2042 20431 2098 20440
rect 2044 19508 2096 19514
rect 2044 19450 2096 19456
rect 1952 18896 2004 18902
rect 1952 18838 2004 18844
rect 1952 18624 2004 18630
rect 1952 18566 2004 18572
rect 1964 18290 1992 18566
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 1584 18216 1636 18222
rect 2056 18170 2084 19450
rect 2148 19394 2176 22374
rect 2240 19514 2268 24550
rect 2320 23656 2372 23662
rect 2320 23598 2372 23604
rect 2332 23118 2360 23598
rect 2412 23180 2464 23186
rect 2412 23122 2464 23128
rect 2320 23112 2372 23118
rect 2320 23054 2372 23060
rect 2424 22438 2452 23122
rect 2412 22432 2464 22438
rect 2410 22400 2412 22409
rect 2464 22400 2466 22409
rect 2410 22335 2466 22344
rect 2320 22092 2372 22098
rect 2320 22034 2372 22040
rect 2332 21350 2360 22034
rect 2320 21344 2372 21350
rect 2320 21286 2372 21292
rect 2332 19825 2360 21286
rect 2516 21026 2544 27390
rect 2686 25936 2742 25945
rect 2686 25871 2742 25880
rect 2700 23866 2728 25871
rect 2688 23860 2740 23866
rect 2688 23802 2740 23808
rect 2686 22536 2742 22545
rect 2686 22471 2742 22480
rect 2700 22137 2728 22471
rect 2962 22264 3018 22273
rect 2962 22199 3018 22208
rect 2686 22128 2742 22137
rect 2686 22063 2742 22072
rect 2594 21856 2650 21865
rect 2594 21791 2650 21800
rect 2608 21146 2636 21791
rect 2780 21344 2832 21350
rect 2686 21312 2742 21321
rect 2780 21286 2832 21292
rect 2686 21247 2742 21256
rect 2596 21140 2648 21146
rect 2596 21082 2648 21088
rect 2516 20998 2636 21026
rect 2504 20392 2556 20398
rect 2504 20334 2556 20340
rect 2412 20256 2464 20262
rect 2410 20224 2412 20233
rect 2464 20224 2466 20233
rect 2410 20159 2466 20168
rect 2516 19990 2544 20334
rect 2608 19990 2636 20998
rect 2700 20602 2728 21247
rect 2688 20596 2740 20602
rect 2688 20538 2740 20544
rect 2504 19984 2556 19990
rect 2504 19926 2556 19932
rect 2596 19984 2648 19990
rect 2596 19926 2648 19932
rect 2318 19816 2374 19825
rect 2318 19751 2374 19760
rect 2320 19712 2372 19718
rect 2320 19654 2372 19660
rect 2228 19508 2280 19514
rect 2228 19450 2280 19456
rect 2148 19366 2268 19394
rect 1584 18158 1636 18164
rect 1492 18080 1544 18086
rect 1492 18022 1544 18028
rect 1398 16688 1454 16697
rect 1398 16623 1454 16632
rect 1400 15904 1452 15910
rect 1400 15846 1452 15852
rect 1216 15088 1268 15094
rect 1216 15030 1268 15036
rect 1122 13696 1178 13705
rect 1122 13631 1178 13640
rect 1124 12912 1176 12918
rect 1124 12854 1176 12860
rect 1136 12442 1164 12854
rect 1228 12782 1256 15030
rect 1412 14550 1440 15846
rect 1400 14544 1452 14550
rect 1400 14486 1452 14492
rect 1400 14272 1452 14278
rect 1400 14214 1452 14220
rect 1216 12776 1268 12782
rect 1216 12718 1268 12724
rect 1412 12646 1440 14214
rect 1400 12640 1452 12646
rect 1400 12582 1452 12588
rect 1504 12481 1532 18022
rect 1596 17338 1624 18158
rect 1964 18142 2084 18170
rect 1964 17814 1992 18142
rect 2240 18086 2268 19366
rect 2332 19174 2360 19654
rect 2792 19553 2820 21286
rect 2872 19712 2924 19718
rect 2872 19654 2924 19660
rect 2778 19544 2834 19553
rect 2778 19479 2834 19488
rect 2778 19408 2834 19417
rect 2778 19343 2834 19352
rect 2792 19242 2820 19343
rect 2780 19236 2832 19242
rect 2780 19178 2832 19184
rect 2884 19174 2912 19654
rect 2320 19168 2372 19174
rect 2320 19110 2372 19116
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 2044 18080 2096 18086
rect 2042 18048 2044 18057
rect 2228 18080 2280 18086
rect 2096 18048 2098 18057
rect 2228 18022 2280 18028
rect 2042 17983 2098 17992
rect 1952 17808 2004 17814
rect 1952 17750 2004 17756
rect 1676 17536 1728 17542
rect 1676 17478 1728 17484
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 1688 17066 1716 17478
rect 2228 17196 2280 17202
rect 2228 17138 2280 17144
rect 1676 17060 1728 17066
rect 1676 17002 1728 17008
rect 2240 16794 2268 17138
rect 2228 16788 2280 16794
rect 2228 16730 2280 16736
rect 1676 16720 1728 16726
rect 1676 16662 1728 16668
rect 1766 16688 1822 16697
rect 1688 15978 1716 16662
rect 1766 16623 1822 16632
rect 1780 16046 1808 16623
rect 1952 16584 2004 16590
rect 1952 16526 2004 16532
rect 2136 16584 2188 16590
rect 2332 16572 2360 19110
rect 2504 18624 2556 18630
rect 2504 18566 2556 18572
rect 2410 17912 2466 17921
rect 2410 17847 2412 17856
rect 2464 17847 2466 17856
rect 2412 17818 2464 17824
rect 2516 17105 2544 18566
rect 2884 18329 2912 19110
rect 2976 18970 3004 22199
rect 3160 21729 3188 27520
rect 3332 26240 3384 26246
rect 3332 26182 3384 26188
rect 3146 21720 3202 21729
rect 3146 21655 3202 21664
rect 3056 21480 3108 21486
rect 3056 21422 3108 21428
rect 3068 20913 3096 21422
rect 3148 21004 3200 21010
rect 3148 20946 3200 20952
rect 3054 20904 3110 20913
rect 3054 20839 3110 20848
rect 3160 20369 3188 20946
rect 3146 20360 3202 20369
rect 3146 20295 3148 20304
rect 3200 20295 3202 20304
rect 3148 20266 3200 20272
rect 3056 19168 3108 19174
rect 3056 19110 3108 19116
rect 2964 18964 3016 18970
rect 2964 18906 3016 18912
rect 2976 18426 3004 18906
rect 3068 18766 3096 19110
rect 3056 18760 3108 18766
rect 3056 18702 3108 18708
rect 2964 18420 3016 18426
rect 2964 18362 3016 18368
rect 2870 18320 2926 18329
rect 2596 18284 2648 18290
rect 2870 18255 2926 18264
rect 2596 18226 2648 18232
rect 2608 18057 2636 18226
rect 3068 18193 3096 18702
rect 3054 18184 3110 18193
rect 3054 18119 3110 18128
rect 2688 18080 2740 18086
rect 2594 18048 2650 18057
rect 2688 18022 2740 18028
rect 2594 17983 2650 17992
rect 2596 17808 2648 17814
rect 2596 17750 2648 17756
rect 2608 17338 2636 17750
rect 2700 17542 2728 18022
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2596 17332 2648 17338
rect 2596 17274 2648 17280
rect 2502 17096 2558 17105
rect 2502 17031 2558 17040
rect 2412 16992 2464 16998
rect 2412 16934 2464 16940
rect 2424 16726 2452 16934
rect 2412 16720 2464 16726
rect 2412 16662 2464 16668
rect 2332 16544 2452 16572
rect 2136 16526 2188 16532
rect 1860 16448 1912 16454
rect 1860 16390 1912 16396
rect 1768 16040 1820 16046
rect 1768 15982 1820 15988
rect 1676 15972 1728 15978
rect 1676 15914 1728 15920
rect 1872 15910 1900 16390
rect 1964 15910 1992 16526
rect 2044 16448 2096 16454
rect 2044 16390 2096 16396
rect 2056 16114 2084 16390
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 1860 15904 1912 15910
rect 1858 15872 1860 15881
rect 1952 15904 2004 15910
rect 1912 15872 1914 15881
rect 1952 15846 2004 15852
rect 1858 15807 1914 15816
rect 1676 15496 1728 15502
rect 2056 15484 2084 16050
rect 2148 15706 2176 16526
rect 2228 16040 2280 16046
rect 2228 15982 2280 15988
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 1676 15438 1728 15444
rect 1964 15456 2084 15484
rect 1688 14822 1716 15438
rect 1964 15366 1992 15456
rect 2148 15416 2176 15642
rect 2056 15388 2176 15416
rect 1768 15360 1820 15366
rect 1768 15302 1820 15308
rect 1952 15360 2004 15366
rect 1952 15302 2004 15308
rect 1676 14816 1728 14822
rect 1676 14758 1728 14764
rect 1688 14634 1716 14758
rect 1596 14606 1716 14634
rect 1490 12472 1546 12481
rect 1124 12436 1176 12442
rect 1490 12407 1546 12416
rect 1124 12378 1176 12384
rect 1400 12368 1452 12374
rect 1596 12356 1624 14606
rect 1780 14482 1808 15302
rect 1964 14822 1992 15302
rect 2056 14958 2084 15388
rect 2044 14952 2096 14958
rect 2044 14894 2096 14900
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1768 14476 1820 14482
rect 1768 14418 1820 14424
rect 1860 14408 1912 14414
rect 1860 14350 1912 14356
rect 1872 14278 1900 14350
rect 1860 14272 1912 14278
rect 1860 14214 1912 14220
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1400 12310 1452 12316
rect 1504 12328 1624 12356
rect 1032 10668 1084 10674
rect 1032 10610 1084 10616
rect 1216 8492 1268 8498
rect 1216 8434 1268 8440
rect 664 7472 716 7478
rect 664 7414 716 7420
rect 676 2854 704 7414
rect 1228 4826 1256 8434
rect 1308 8288 1360 8294
rect 1308 8230 1360 8236
rect 1216 4820 1268 4826
rect 1216 4762 1268 4768
rect 1214 3632 1270 3641
rect 1214 3567 1270 3576
rect 664 2848 716 2854
rect 664 2790 716 2796
rect 202 1728 258 1737
rect 202 1663 258 1672
rect 216 480 244 1663
rect 676 480 704 2790
rect 1228 480 1256 3567
rect 1320 3233 1348 8230
rect 1412 3738 1440 12310
rect 1400 3732 1452 3738
rect 1400 3674 1452 3680
rect 1400 3392 1452 3398
rect 1400 3334 1452 3340
rect 1306 3224 1362 3233
rect 1306 3159 1362 3168
rect 1412 2514 1440 3334
rect 1504 3194 1532 12328
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1596 9654 1624 10610
rect 1584 9648 1636 9654
rect 1584 9590 1636 9596
rect 1688 9518 1716 13874
rect 1768 13864 1820 13870
rect 1768 13806 1820 13812
rect 1780 13190 1808 13806
rect 1872 13734 1900 14214
rect 1860 13728 1912 13734
rect 1860 13670 1912 13676
rect 1768 13184 1820 13190
rect 1766 13152 1768 13161
rect 1820 13152 1822 13161
rect 1766 13087 1822 13096
rect 1872 12306 1900 13670
rect 1964 13002 1992 14758
rect 2056 13190 2084 14894
rect 2134 13832 2190 13841
rect 2134 13767 2136 13776
rect 2188 13767 2190 13776
rect 2136 13738 2188 13744
rect 2044 13184 2096 13190
rect 2044 13126 2096 13132
rect 1964 12974 2084 13002
rect 1950 12472 2006 12481
rect 1950 12407 2006 12416
rect 1860 12300 1912 12306
rect 1860 12242 1912 12248
rect 1872 11558 1900 12242
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1688 9178 1716 9454
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1596 3670 1624 8910
rect 1780 8498 1808 11290
rect 1860 11212 1912 11218
rect 1860 11154 1912 11160
rect 1872 10266 1900 11154
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 1860 9648 1912 9654
rect 1860 9590 1912 9596
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1766 8392 1822 8401
rect 1688 7750 1716 8366
rect 1766 8327 1768 8336
rect 1820 8327 1822 8336
rect 1768 8298 1820 8304
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1688 6236 1716 7686
rect 1780 7002 1808 8298
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 1768 6248 1820 6254
rect 1688 6208 1768 6236
rect 1768 6190 1820 6196
rect 1780 5778 1808 6190
rect 1768 5772 1820 5778
rect 1768 5714 1820 5720
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1780 4826 1808 4966
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 1674 4448 1730 4457
rect 1674 4383 1730 4392
rect 1688 3942 1716 4383
rect 1872 4010 1900 9590
rect 1964 7478 1992 12407
rect 2056 11200 2084 12974
rect 2148 12850 2176 13738
rect 2136 12844 2188 12850
rect 2136 12786 2188 12792
rect 2136 11620 2188 11626
rect 2136 11562 2188 11568
rect 2148 11354 2176 11562
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2136 11212 2188 11218
rect 2056 11172 2136 11200
rect 2136 11154 2188 11160
rect 2134 11112 2190 11121
rect 2134 11047 2190 11056
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 2056 7546 2084 8774
rect 2148 7886 2176 11047
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 2136 7744 2188 7750
rect 2136 7686 2188 7692
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 2148 7478 2176 7686
rect 1952 7472 2004 7478
rect 1952 7414 2004 7420
rect 2136 7472 2188 7478
rect 2136 7414 2188 7420
rect 1952 7200 2004 7206
rect 1952 7142 2004 7148
rect 1964 6662 1992 7142
rect 2240 6746 2268 15982
rect 2320 14000 2372 14006
rect 2320 13942 2372 13948
rect 2332 12374 2360 13942
rect 2320 12368 2372 12374
rect 2320 12310 2372 12316
rect 2332 11898 2360 12310
rect 2320 11892 2372 11898
rect 2320 11834 2372 11840
rect 2424 10112 2452 16544
rect 2504 15020 2556 15026
rect 2504 14962 2556 14968
rect 2516 14278 2544 14962
rect 2504 14272 2556 14278
rect 2504 14214 2556 14220
rect 2608 13462 2636 17274
rect 2700 17066 2728 17478
rect 2884 17134 2912 17614
rect 3056 17536 3108 17542
rect 3056 17478 3108 17484
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 2688 17060 2740 17066
rect 2688 17002 2740 17008
rect 2962 16960 3018 16969
rect 2962 16895 3018 16904
rect 2976 16794 3004 16895
rect 2964 16788 3016 16794
rect 2964 16730 3016 16736
rect 2964 16040 3016 16046
rect 2964 15982 3016 15988
rect 2688 15904 2740 15910
rect 2688 15846 2740 15852
rect 2596 13456 2648 13462
rect 2596 13398 2648 13404
rect 2700 13025 2728 15846
rect 2976 15366 3004 15982
rect 2964 15360 3016 15366
rect 2964 15302 3016 15308
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2792 14618 2820 14894
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 2780 14340 2832 14346
rect 2780 14282 2832 14288
rect 2792 14006 2820 14282
rect 2780 14000 2832 14006
rect 2780 13942 2832 13948
rect 2792 13870 2820 13942
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2870 13832 2926 13841
rect 2870 13767 2872 13776
rect 2924 13767 2926 13776
rect 2872 13738 2924 13744
rect 2780 13456 2832 13462
rect 2780 13398 2832 13404
rect 2686 13016 2742 13025
rect 2686 12951 2742 12960
rect 2792 12918 2820 13398
rect 2976 12986 3004 15302
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 2780 12912 2832 12918
rect 2778 12880 2780 12889
rect 2832 12880 2834 12889
rect 3068 12866 3096 17478
rect 3148 16992 3200 16998
rect 3148 16934 3200 16940
rect 3160 15586 3188 16934
rect 3344 16250 3372 26182
rect 3516 21684 3568 21690
rect 3516 21626 3568 21632
rect 3528 21146 3556 21626
rect 3804 21622 3832 27520
rect 4066 23624 4122 23633
rect 4066 23559 4122 23568
rect 4080 22778 4108 23559
rect 4068 22772 4120 22778
rect 4068 22714 4120 22720
rect 3792 21616 3844 21622
rect 3792 21558 3844 21564
rect 3516 21140 3568 21146
rect 3516 21082 3568 21088
rect 3884 20528 3936 20534
rect 3884 20470 3936 20476
rect 3608 20392 3660 20398
rect 3608 20334 3660 20340
rect 3620 19310 3648 20334
rect 3792 20256 3844 20262
rect 3792 20198 3844 20204
rect 3804 20097 3832 20198
rect 3790 20088 3846 20097
rect 3790 20023 3846 20032
rect 3608 19304 3660 19310
rect 3608 19246 3660 19252
rect 3698 19272 3754 19281
rect 3698 19207 3754 19216
rect 3712 18970 3740 19207
rect 3790 19136 3846 19145
rect 3790 19071 3846 19080
rect 3700 18964 3752 18970
rect 3700 18906 3752 18912
rect 3698 17776 3754 17785
rect 3698 17711 3754 17720
rect 3424 17196 3476 17202
rect 3424 17138 3476 17144
rect 3436 16590 3464 17138
rect 3608 17128 3660 17134
rect 3608 17070 3660 17076
rect 3516 16992 3568 16998
rect 3516 16934 3568 16940
rect 3424 16584 3476 16590
rect 3424 16526 3476 16532
rect 3436 16454 3464 16526
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 3436 16250 3464 16390
rect 3332 16244 3384 16250
rect 3332 16186 3384 16192
rect 3424 16244 3476 16250
rect 3424 16186 3476 16192
rect 3240 15972 3292 15978
rect 3240 15914 3292 15920
rect 3252 15745 3280 15914
rect 3238 15736 3294 15745
rect 3238 15671 3294 15680
rect 3160 15558 3280 15586
rect 3528 15570 3556 16934
rect 3148 15428 3200 15434
rect 3148 15370 3200 15376
rect 3160 13530 3188 15370
rect 3252 14822 3280 15558
rect 3516 15564 3568 15570
rect 3516 15506 3568 15512
rect 3424 15360 3476 15366
rect 3422 15328 3424 15337
rect 3476 15328 3478 15337
rect 3422 15263 3478 15272
rect 3516 14884 3568 14890
rect 3516 14826 3568 14832
rect 3240 14816 3292 14822
rect 3240 14758 3292 14764
rect 3252 13977 3280 14758
rect 3528 14618 3556 14826
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3238 13968 3294 13977
rect 3238 13903 3294 13912
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 3148 13388 3200 13394
rect 3148 13330 3200 13336
rect 2778 12815 2834 12824
rect 2884 12838 3096 12866
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 2516 11898 2544 12582
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2608 10810 2636 12718
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 2686 11656 2742 11665
rect 2686 11591 2688 11600
rect 2740 11591 2742 11600
rect 2688 11562 2740 11568
rect 2686 11520 2742 11529
rect 2686 11455 2742 11464
rect 2596 10804 2648 10810
rect 2596 10746 2648 10752
rect 2700 10606 2728 11455
rect 2792 11150 2820 12582
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2148 6718 2268 6746
rect 2332 10084 2452 10112
rect 2504 10124 2556 10130
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1860 4004 1912 4010
rect 1860 3946 1912 3952
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1858 3904 1914 3913
rect 1688 3738 1716 3878
rect 1858 3839 1914 3848
rect 1766 3768 1822 3777
rect 1676 3732 1728 3738
rect 1766 3703 1822 3712
rect 1676 3674 1728 3680
rect 1584 3664 1636 3670
rect 1584 3606 1636 3612
rect 1674 3224 1730 3233
rect 1492 3188 1544 3194
rect 1674 3159 1730 3168
rect 1492 3130 1544 3136
rect 1688 3058 1716 3159
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1780 2990 1808 3703
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 1584 2916 1636 2922
rect 1584 2858 1636 2864
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1412 2009 1440 2450
rect 1398 2000 1454 2009
rect 1398 1935 1454 1944
rect 1596 921 1624 2858
rect 1674 2680 1730 2689
rect 1674 2615 1730 2624
rect 1688 2582 1716 2615
rect 1676 2576 1728 2582
rect 1676 2518 1728 2524
rect 1582 912 1638 921
rect 1582 847 1638 856
rect 1872 626 1900 3839
rect 1964 3398 1992 6598
rect 2044 5772 2096 5778
rect 2044 5714 2096 5720
rect 2056 5030 2084 5714
rect 2044 5024 2096 5030
rect 2044 4966 2096 4972
rect 2056 4622 2084 4966
rect 2044 4616 2096 4622
rect 2044 4558 2096 4564
rect 2056 4282 2084 4558
rect 2044 4276 2096 4282
rect 2044 4218 2096 4224
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 2056 1601 2084 4082
rect 2148 2650 2176 6718
rect 2228 4752 2280 4758
rect 2228 4694 2280 4700
rect 2240 3534 2268 4694
rect 2332 4146 2360 10084
rect 2504 10066 2556 10072
rect 2410 10024 2466 10033
rect 2410 9959 2412 9968
rect 2464 9959 2466 9968
rect 2412 9930 2464 9936
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2424 8430 2452 9454
rect 2412 8424 2464 8430
rect 2412 8366 2464 8372
rect 2516 8090 2544 10066
rect 2608 9024 2636 10406
rect 2700 10266 2728 10542
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2792 10146 2820 10202
rect 2700 10130 2820 10146
rect 2688 10124 2820 10130
rect 2740 10118 2820 10124
rect 2688 10066 2740 10072
rect 2688 9920 2740 9926
rect 2688 9862 2740 9868
rect 2700 9178 2728 9862
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2688 9036 2740 9042
rect 2608 8996 2688 9024
rect 2688 8978 2740 8984
rect 2700 8294 2728 8978
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2792 8022 2820 8230
rect 2884 8129 2912 12838
rect 3160 12646 3188 13330
rect 3516 13320 3568 13326
rect 3514 13288 3516 13297
rect 3568 13288 3570 13297
rect 3436 13246 3514 13274
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2976 11354 3004 11494
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 2976 9450 3004 9998
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2976 8401 3004 8910
rect 2962 8392 3018 8401
rect 2962 8327 2964 8336
rect 3016 8327 3018 8336
rect 2964 8298 3016 8304
rect 2870 8120 2926 8129
rect 2870 8055 2926 8064
rect 2780 8016 2832 8022
rect 2780 7958 2832 7964
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2516 7342 2544 7822
rect 2504 7336 2556 7342
rect 2504 7278 2556 7284
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 2240 3058 2268 3470
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 2136 2644 2188 2650
rect 2136 2586 2188 2592
rect 2240 2446 2268 2994
rect 2318 2952 2374 2961
rect 2516 2922 2544 7278
rect 2792 7002 2820 7958
rect 2884 7857 2912 8055
rect 2870 7848 2926 7857
rect 2976 7818 3004 8298
rect 3160 7993 3188 12582
rect 3252 11665 3280 13126
rect 3436 12850 3464 13246
rect 3514 13223 3570 13232
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3528 12782 3556 13126
rect 3516 12776 3568 12782
rect 3516 12718 3568 12724
rect 3422 11792 3478 11801
rect 3422 11727 3478 11736
rect 3238 11656 3294 11665
rect 3238 11591 3294 11600
rect 3330 10568 3386 10577
rect 3330 10503 3386 10512
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 3252 10266 3280 10406
rect 3240 10260 3292 10266
rect 3240 10202 3292 10208
rect 3146 7984 3202 7993
rect 3146 7919 3202 7928
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 2870 7783 2926 7792
rect 2964 7812 3016 7818
rect 2964 7754 3016 7760
rect 3160 7206 3188 7822
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 2780 6996 2832 7002
rect 2780 6938 2832 6944
rect 2596 6860 2648 6866
rect 2596 6802 2648 6808
rect 2608 6458 2636 6802
rect 2688 6792 2740 6798
rect 2688 6734 2740 6740
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2608 4554 2636 6394
rect 2700 5914 2728 6734
rect 2792 6390 2820 6734
rect 2780 6384 2832 6390
rect 2780 6326 2832 6332
rect 2792 6168 2820 6326
rect 2964 6180 3016 6186
rect 2792 6140 2964 6168
rect 2792 5914 2820 6140
rect 2964 6122 3016 6128
rect 2688 5908 2740 5914
rect 2688 5850 2740 5856
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2700 5556 2728 5850
rect 2700 5528 2820 5556
rect 2688 5024 2740 5030
rect 2688 4966 2740 4972
rect 2596 4548 2648 4554
rect 2596 4490 2648 4496
rect 2700 4214 2728 4966
rect 2792 4554 2820 5528
rect 2872 5296 2924 5302
rect 2872 5238 2924 5244
rect 2884 4808 2912 5238
rect 2884 4780 3004 4808
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 2780 4548 2832 4554
rect 2780 4490 2832 4496
rect 2688 4208 2740 4214
rect 2688 4150 2740 4156
rect 2884 3942 2912 4626
rect 2976 4078 3004 4780
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2884 3670 2912 3878
rect 2976 3738 3004 4014
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2872 3664 2924 3670
rect 2872 3606 2924 3612
rect 3160 3602 3188 7142
rect 3344 4146 3372 10503
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3344 3194 3372 4082
rect 3436 4010 3464 11727
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3528 11218 3556 11494
rect 3516 11212 3568 11218
rect 3516 11154 3568 11160
rect 3620 11121 3648 17070
rect 3712 16153 3740 17711
rect 3698 16144 3754 16153
rect 3698 16079 3754 16088
rect 3700 15904 3752 15910
rect 3700 15846 3752 15852
rect 3712 11801 3740 15846
rect 3804 14929 3832 19071
rect 3896 18222 3924 20470
rect 4250 20224 4306 20233
rect 4250 20159 4306 20168
rect 4264 20058 4292 20159
rect 4252 20052 4304 20058
rect 4252 19994 4304 20000
rect 4252 19712 4304 19718
rect 4252 19654 4304 19660
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3988 19174 4016 19246
rect 3976 19168 4028 19174
rect 3976 19110 4028 19116
rect 3884 18216 3936 18222
rect 3884 18158 3936 18164
rect 3884 18080 3936 18086
rect 3884 18022 3936 18028
rect 3896 17678 3924 18022
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 3988 17490 4016 19110
rect 4068 18216 4120 18222
rect 4068 18158 4120 18164
rect 4080 17542 4108 18158
rect 3896 17462 4016 17490
rect 4068 17536 4120 17542
rect 4068 17478 4120 17484
rect 3790 14920 3846 14929
rect 3790 14855 3846 14864
rect 3896 13394 3924 17462
rect 3976 16992 4028 16998
rect 3976 16934 4028 16940
rect 3988 15337 4016 16934
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 3974 15328 4030 15337
rect 3974 15263 4030 15272
rect 4080 14958 4108 16390
rect 4172 15162 4200 16594
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 3988 13546 4016 14350
rect 3988 13530 4200 13546
rect 3988 13524 4212 13530
rect 3988 13518 4160 13524
rect 4160 13466 4212 13472
rect 4066 13424 4122 13433
rect 3884 13388 3936 13394
rect 3884 13330 3936 13336
rect 3976 13388 4028 13394
rect 4066 13359 4122 13368
rect 3976 13330 4028 13336
rect 3882 13152 3938 13161
rect 3882 13087 3938 13096
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3804 12442 3832 12786
rect 3792 12436 3844 12442
rect 3792 12378 3844 12384
rect 3698 11792 3754 11801
rect 3698 11727 3754 11736
rect 3606 11112 3662 11121
rect 3606 11047 3662 11056
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3804 10606 3832 10950
rect 3792 10600 3844 10606
rect 3792 10542 3844 10548
rect 3698 10296 3754 10305
rect 3698 10231 3754 10240
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3528 8362 3556 9318
rect 3712 8537 3740 10231
rect 3804 9926 3832 10542
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3804 9518 3832 9862
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3698 8528 3754 8537
rect 3698 8463 3754 8472
rect 3516 8356 3568 8362
rect 3516 8298 3568 8304
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 3712 7410 3740 7686
rect 3700 7404 3752 7410
rect 3700 7346 3752 7352
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3620 5778 3648 6190
rect 3896 6089 3924 13087
rect 3988 12442 4016 13330
rect 4080 13161 4108 13359
rect 4066 13152 4122 13161
rect 4066 13087 4122 13096
rect 4068 12912 4120 12918
rect 4068 12854 4120 12860
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 4080 12322 4108 12854
rect 4172 12442 4200 13466
rect 4160 12436 4212 12442
rect 4264 12424 4292 19654
rect 4356 19310 4384 27520
rect 4620 25968 4672 25974
rect 4620 25910 4672 25916
rect 4436 23520 4488 23526
rect 4436 23462 4488 23468
rect 4448 19496 4476 23462
rect 4448 19468 4568 19496
rect 4540 19360 4568 19468
rect 4448 19332 4568 19360
rect 4344 19304 4396 19310
rect 4342 19272 4344 19281
rect 4396 19272 4398 19281
rect 4342 19207 4398 19216
rect 4344 18284 4396 18290
rect 4344 18226 4396 18232
rect 4356 17882 4384 18226
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4356 16794 4384 17818
rect 4344 16788 4396 16794
rect 4344 16730 4396 16736
rect 4344 14476 4396 14482
rect 4344 14418 4396 14424
rect 4356 13870 4384 14418
rect 4344 13864 4396 13870
rect 4344 13806 4396 13812
rect 4344 12436 4396 12442
rect 4264 12396 4344 12424
rect 4160 12378 4212 12384
rect 4344 12378 4396 12384
rect 4080 12306 4200 12322
rect 4080 12300 4212 12306
rect 4080 12294 4160 12300
rect 4160 12242 4212 12248
rect 3974 11656 4030 11665
rect 3974 11591 4030 11600
rect 3988 11014 4016 11591
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 4068 10532 4120 10538
rect 4068 10474 4120 10480
rect 3974 10432 4030 10441
rect 3974 10367 4030 10376
rect 3988 9625 4016 10367
rect 3974 9616 4030 9625
rect 3974 9551 4030 9560
rect 4080 9382 4108 10474
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4080 8537 4108 9318
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4066 8528 4122 8537
rect 4356 8498 4384 8774
rect 4066 8463 4122 8472
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4448 7857 4476 19332
rect 4632 18952 4660 25910
rect 4908 23526 4936 27520
rect 5552 26178 5580 27520
rect 5540 26172 5592 26178
rect 5540 26114 5592 26120
rect 6104 26081 6132 27520
rect 6090 26072 6146 26081
rect 6090 26007 6146 26016
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 4896 23520 4948 23526
rect 4896 23462 4948 23468
rect 6656 23225 6684 27520
rect 6736 26104 6788 26110
rect 6736 26046 6788 26052
rect 6458 23216 6514 23225
rect 6458 23151 6514 23160
rect 6642 23216 6698 23225
rect 6642 23151 6698 23160
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5356 22568 5408 22574
rect 4710 22536 4766 22545
rect 5356 22510 5408 22516
rect 4710 22471 4766 22480
rect 4804 22500 4856 22506
rect 4724 22137 4752 22471
rect 4804 22442 4856 22448
rect 4816 22234 4844 22442
rect 5262 22400 5318 22409
rect 5262 22335 5318 22344
rect 4804 22228 4856 22234
rect 4804 22170 4856 22176
rect 4710 22128 4766 22137
rect 4710 22063 4766 22072
rect 4724 20058 4752 22063
rect 4816 21690 4844 22170
rect 4988 22092 5040 22098
rect 4988 22034 5040 22040
rect 4894 21720 4950 21729
rect 4804 21684 4856 21690
rect 4894 21655 4896 21664
rect 4804 21626 4856 21632
rect 4948 21655 4950 21664
rect 4896 21626 4948 21632
rect 4712 20052 4764 20058
rect 4712 19994 4764 20000
rect 4724 19514 4752 19994
rect 4816 19990 4844 21626
rect 4908 21418 4936 21626
rect 5000 21486 5028 22034
rect 4988 21480 5040 21486
rect 4988 21422 5040 21428
rect 4896 21412 4948 21418
rect 4896 21354 4948 21360
rect 4894 21176 4950 21185
rect 4894 21111 4896 21120
rect 4948 21111 4950 21120
rect 4896 21082 4948 21088
rect 5000 21026 5028 21422
rect 5172 21344 5224 21350
rect 5172 21286 5224 21292
rect 4908 20998 5028 21026
rect 4804 19984 4856 19990
rect 4804 19926 4856 19932
rect 4804 19848 4856 19854
rect 4804 19790 4856 19796
rect 4712 19508 4764 19514
rect 4712 19450 4764 19456
rect 4816 19446 4844 19790
rect 4804 19440 4856 19446
rect 4724 19388 4804 19394
rect 4724 19382 4856 19388
rect 4724 19366 4844 19382
rect 4724 18970 4752 19366
rect 4540 18924 4660 18952
rect 4712 18964 4764 18970
rect 4540 18222 4568 18924
rect 4712 18906 4764 18912
rect 4620 18828 4672 18834
rect 4620 18770 4672 18776
rect 4632 18426 4660 18770
rect 4620 18420 4672 18426
rect 4620 18362 4672 18368
rect 4528 18216 4580 18222
rect 4528 18158 4580 18164
rect 4632 16833 4660 18362
rect 4724 18290 4752 18906
rect 4712 18284 4764 18290
rect 4712 18226 4764 18232
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4618 16824 4674 16833
rect 4618 16759 4674 16768
rect 4724 16726 4752 16934
rect 4712 16720 4764 16726
rect 4712 16662 4764 16668
rect 4712 15632 4764 15638
rect 4712 15574 4764 15580
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4528 15360 4580 15366
rect 4528 15302 4580 15308
rect 4540 15026 4568 15302
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 4540 14550 4568 14962
rect 4632 14822 4660 15506
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4724 14550 4752 15574
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 4528 14544 4580 14550
rect 4528 14486 4580 14492
rect 4712 14544 4764 14550
rect 4712 14486 4764 14492
rect 4816 14074 4844 14894
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4908 13954 4936 20998
rect 4988 20936 5040 20942
rect 4988 20878 5040 20884
rect 5080 20936 5132 20942
rect 5080 20878 5132 20884
rect 5000 20641 5028 20878
rect 4986 20632 5042 20641
rect 4986 20567 5042 20576
rect 5000 20262 5028 20567
rect 5092 20330 5120 20878
rect 5184 20806 5212 21286
rect 5172 20800 5224 20806
rect 5172 20742 5224 20748
rect 5080 20324 5132 20330
rect 5080 20266 5132 20272
rect 4988 20256 5040 20262
rect 4988 20198 5040 20204
rect 4988 19916 5040 19922
rect 4988 19858 5040 19864
rect 5000 19174 5028 19858
rect 5092 19854 5120 20266
rect 5080 19848 5132 19854
rect 5080 19790 5132 19796
rect 5184 19310 5212 20742
rect 5276 20602 5304 22335
rect 5368 22166 5396 22510
rect 5356 22160 5408 22166
rect 5356 22102 5408 22108
rect 6276 21888 6328 21894
rect 6276 21830 6328 21836
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5540 21616 5592 21622
rect 5540 21558 5592 21564
rect 5552 21350 5580 21558
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 5540 21344 5592 21350
rect 5538 21312 5540 21321
rect 5592 21312 5594 21321
rect 5538 21247 5594 21256
rect 5368 21146 5580 21162
rect 5368 21140 5592 21146
rect 5368 21134 5540 21140
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 5264 20256 5316 20262
rect 5264 20198 5316 20204
rect 5276 19961 5304 20198
rect 5262 19952 5318 19961
rect 5262 19887 5318 19896
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 5368 19174 5396 21134
rect 5540 21082 5592 21088
rect 5448 21072 5500 21078
rect 5448 21014 5500 21020
rect 5538 21040 5594 21049
rect 5460 20346 5488 21014
rect 5538 20975 5540 20984
rect 5592 20975 5594 20984
rect 5540 20946 5592 20952
rect 5828 20942 5856 21490
rect 6090 21040 6146 21049
rect 6090 20975 6146 20984
rect 5816 20936 5868 20942
rect 5816 20878 5868 20884
rect 6000 20936 6052 20942
rect 6000 20878 6052 20884
rect 5540 20868 5592 20874
rect 5540 20810 5592 20816
rect 5552 20466 5580 20810
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 5724 20460 5776 20466
rect 5724 20402 5776 20408
rect 5460 20330 5580 20346
rect 5460 20324 5592 20330
rect 5460 20318 5540 20324
rect 4988 19168 5040 19174
rect 4988 19110 5040 19116
rect 5356 19168 5408 19174
rect 5356 19110 5408 19116
rect 5000 18737 5028 19110
rect 5460 18970 5488 20318
rect 5540 20266 5592 20272
rect 5736 19922 5764 20402
rect 6012 20262 6040 20878
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 5724 19916 5776 19922
rect 5724 19858 5776 19864
rect 5736 19825 5764 19858
rect 5538 19816 5594 19825
rect 5538 19751 5594 19760
rect 5722 19816 5778 19825
rect 5722 19751 5778 19760
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5264 18896 5316 18902
rect 5552 18873 5580 19751
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5264 18838 5316 18844
rect 5538 18864 5594 18873
rect 5080 18828 5132 18834
rect 5080 18770 5132 18776
rect 4986 18728 5042 18737
rect 4986 18663 5042 18672
rect 5092 18426 5120 18770
rect 5080 18420 5132 18426
rect 5080 18362 5132 18368
rect 5092 17678 5120 18362
rect 5276 17882 5304 18838
rect 5538 18799 5594 18808
rect 6012 18766 6040 20198
rect 6104 20058 6132 20975
rect 6184 20800 6236 20806
rect 6184 20742 6236 20748
rect 6092 20052 6144 20058
rect 6092 19994 6144 20000
rect 6092 19916 6144 19922
rect 6092 19858 6144 19864
rect 6104 19378 6132 19858
rect 6092 19372 6144 19378
rect 6092 19314 6144 19320
rect 6104 18902 6132 19314
rect 6196 18970 6224 20742
rect 6288 19242 6316 21830
rect 6472 19446 6500 23151
rect 6644 22636 6696 22642
rect 6644 22578 6696 22584
rect 6656 22438 6684 22578
rect 6644 22432 6696 22438
rect 6644 22374 6696 22380
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 6564 21146 6592 21830
rect 6656 21690 6684 22374
rect 6644 21684 6696 21690
rect 6644 21626 6696 21632
rect 6552 21140 6604 21146
rect 6552 21082 6604 21088
rect 6564 20602 6592 21082
rect 6552 20596 6604 20602
rect 6552 20538 6604 20544
rect 6644 20392 6696 20398
rect 6644 20334 6696 20340
rect 6656 19922 6684 20334
rect 6644 19916 6696 19922
rect 6644 19858 6696 19864
rect 6460 19440 6512 19446
rect 6460 19382 6512 19388
rect 6748 19258 6776 26046
rect 7300 23798 7328 27520
rect 7852 24970 7880 27520
rect 8114 25936 8170 25945
rect 8114 25871 8170 25880
rect 8024 25832 8076 25838
rect 7930 25800 7986 25809
rect 8024 25774 8076 25780
rect 7930 25735 7986 25744
rect 7760 24942 7880 24970
rect 7760 24721 7788 24942
rect 7746 24712 7802 24721
rect 7746 24647 7802 24656
rect 7564 24268 7616 24274
rect 7564 24210 7616 24216
rect 7288 23792 7340 23798
rect 7288 23734 7340 23740
rect 7576 23526 7604 24210
rect 7564 23520 7616 23526
rect 7564 23462 7616 23468
rect 7194 23352 7250 23361
rect 7194 23287 7196 23296
rect 7248 23287 7250 23296
rect 7196 23258 7248 23264
rect 7012 22976 7064 22982
rect 7012 22918 7064 22924
rect 7024 22506 7052 22918
rect 7208 22658 7236 23258
rect 7472 23180 7524 23186
rect 7472 23122 7524 23128
rect 7378 22944 7434 22953
rect 7378 22879 7434 22888
rect 7286 22672 7342 22681
rect 7208 22630 7286 22658
rect 7286 22607 7342 22616
rect 7104 22568 7156 22574
rect 7104 22510 7156 22516
rect 7012 22500 7064 22506
rect 7012 22442 7064 22448
rect 7024 22148 7052 22442
rect 7116 22273 7144 22510
rect 7300 22506 7328 22607
rect 7288 22500 7340 22506
rect 7288 22442 7340 22448
rect 7196 22432 7248 22438
rect 7196 22374 7248 22380
rect 7102 22264 7158 22273
rect 7102 22199 7158 22208
rect 7024 22120 7144 22148
rect 7116 22030 7144 22120
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 6920 21888 6972 21894
rect 6920 21830 6972 21836
rect 6828 21412 6880 21418
rect 6828 21354 6880 21360
rect 6840 20777 6868 21354
rect 6932 21185 6960 21830
rect 7116 21486 7144 21966
rect 7104 21480 7156 21486
rect 7104 21422 7156 21428
rect 6918 21176 6974 21185
rect 6918 21111 6974 21120
rect 6826 20768 6882 20777
rect 6826 20703 6882 20712
rect 6932 20466 6960 21111
rect 7208 21049 7236 22374
rect 7392 22216 7420 22879
rect 7484 22409 7512 23122
rect 7470 22400 7526 22409
rect 7470 22335 7526 22344
rect 7300 22188 7420 22216
rect 7194 21040 7250 21049
rect 7194 20975 7250 20984
rect 7300 20890 7328 22188
rect 7380 22092 7432 22098
rect 7380 22034 7432 22040
rect 7392 21690 7420 22034
rect 7380 21684 7432 21690
rect 7380 21626 7432 21632
rect 7024 20862 7328 20890
rect 6920 20460 6972 20466
rect 6920 20402 6972 20408
rect 6828 19984 6880 19990
rect 6828 19926 6880 19932
rect 6276 19236 6328 19242
rect 6276 19178 6328 19184
rect 6564 19230 6776 19258
rect 6368 19168 6420 19174
rect 6288 19116 6368 19122
rect 6288 19110 6420 19116
rect 6288 19094 6408 19110
rect 6184 18964 6236 18970
rect 6184 18906 6236 18912
rect 6092 18896 6144 18902
rect 6092 18838 6144 18844
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 6000 18760 6052 18766
rect 6000 18702 6052 18708
rect 5448 18080 5500 18086
rect 5552 18068 5580 18702
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 6012 18426 6040 18702
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 5500 18040 5580 18068
rect 5448 18022 5500 18028
rect 5552 17921 5580 18040
rect 5632 18080 5684 18086
rect 5632 18022 5684 18028
rect 5538 17912 5594 17921
rect 5264 17876 5316 17882
rect 5538 17847 5594 17856
rect 5264 17818 5316 17824
rect 5644 17785 5672 18022
rect 6000 17876 6052 17882
rect 6000 17818 6052 17824
rect 5630 17776 5686 17785
rect 5630 17711 5686 17720
rect 6012 17678 6040 17818
rect 6184 17740 6236 17746
rect 6184 17682 6236 17688
rect 4988 17672 5040 17678
rect 4988 17614 5040 17620
rect 5080 17672 5132 17678
rect 5080 17614 5132 17620
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 5000 17241 5028 17614
rect 5170 17368 5226 17377
rect 5170 17303 5226 17312
rect 5080 17264 5132 17270
rect 4986 17232 5042 17241
rect 5080 17206 5132 17212
rect 4986 17167 5042 17176
rect 5092 17134 5120 17206
rect 5184 17202 5212 17303
rect 5172 17196 5224 17202
rect 5172 17138 5224 17144
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 5080 17128 5132 17134
rect 5080 17070 5132 17076
rect 4988 17060 5040 17066
rect 4988 17002 5040 17008
rect 5000 16561 5028 17002
rect 4986 16552 5042 16561
rect 4986 16487 5042 16496
rect 4816 13926 4936 13954
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4540 12714 4568 13262
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4528 12708 4580 12714
rect 4528 12650 4580 12656
rect 4724 12374 4752 12718
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4528 9444 4580 9450
rect 4528 9386 4580 9392
rect 4066 7848 4122 7857
rect 4066 7783 4122 7792
rect 4434 7848 4490 7857
rect 4434 7783 4490 7792
rect 4080 7342 4108 7783
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 4160 7268 4212 7274
rect 4160 7210 4212 7216
rect 3976 7200 4028 7206
rect 3974 7168 3976 7177
rect 4028 7168 4030 7177
rect 3974 7103 4030 7112
rect 3988 7002 4016 7103
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 4172 6458 4200 7210
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 3882 6080 3938 6089
rect 3882 6015 3938 6024
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 3514 5536 3570 5545
rect 3514 5471 3570 5480
rect 3424 4004 3476 4010
rect 3424 3946 3476 3952
rect 3422 3224 3478 3233
rect 3332 3188 3384 3194
rect 3422 3159 3478 3168
rect 3332 3130 3384 3136
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 2318 2887 2374 2896
rect 2504 2916 2556 2922
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 2042 1592 2098 1601
rect 2042 1527 2098 1536
rect 1780 598 1900 626
rect 1780 480 1808 598
rect 2332 480 2360 2887
rect 2504 2858 2556 2864
rect 2870 2816 2926 2825
rect 2870 2751 2926 2760
rect 2884 480 2912 2751
rect 3160 2514 3188 2926
rect 3148 2508 3200 2514
rect 3148 2450 3200 2456
rect 2964 2440 3016 2446
rect 2962 2408 2964 2417
rect 3016 2408 3018 2417
rect 2962 2343 3018 2352
rect 3436 480 3464 3159
rect 3528 921 3556 5471
rect 3620 5166 3648 5714
rect 3608 5160 3660 5166
rect 3608 5102 3660 5108
rect 3620 2990 3648 5102
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3804 3738 3832 4558
rect 3884 4004 3936 4010
rect 3884 3946 3936 3952
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3790 3496 3846 3505
rect 3790 3431 3846 3440
rect 3804 2990 3832 3431
rect 3608 2984 3660 2990
rect 3608 2926 3660 2932
rect 3792 2984 3844 2990
rect 3792 2926 3844 2932
rect 3804 2650 3832 2926
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 3896 1465 3924 3946
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4066 3768 4122 3777
rect 4066 3703 4068 3712
rect 4120 3703 4122 3712
rect 4068 3674 4120 3680
rect 3974 3088 4030 3097
rect 3974 3023 4030 3032
rect 3882 1456 3938 1465
rect 3882 1391 3938 1400
rect 3514 912 3570 921
rect 3514 847 3570 856
rect 3988 480 4016 3023
rect 202 0 258 480
rect 662 0 718 480
rect 1214 0 1270 480
rect 1766 0 1822 480
rect 2318 0 2374 480
rect 2870 0 2926 480
rect 3422 0 3478 480
rect 3974 0 4030 480
rect 4264 377 4292 3878
rect 4540 480 4568 9386
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4632 2582 4660 5306
rect 4724 3942 4752 12310
rect 4816 10266 4844 13926
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4804 9988 4856 9994
rect 4804 9930 4856 9936
rect 4816 9722 4844 9930
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 5000 9654 5028 16487
rect 5092 12782 5120 17070
rect 5276 16640 5304 17138
rect 5184 16612 5304 16640
rect 5184 16454 5212 16612
rect 5172 16448 5224 16454
rect 5172 16390 5224 16396
rect 5184 15706 5212 16390
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 5368 14822 5396 16050
rect 5448 16040 5500 16046
rect 5552 16028 5580 17614
rect 6000 17536 6052 17542
rect 6000 17478 6052 17484
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5500 16000 5580 16028
rect 5448 15982 5500 15988
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5276 14278 5304 14758
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 5276 13394 5304 14214
rect 5460 14074 5488 15982
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5630 15872 5686 15881
rect 5552 15162 5580 15846
rect 5630 15807 5686 15816
rect 5644 15638 5672 15807
rect 5632 15632 5684 15638
rect 5632 15574 5684 15580
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6012 15162 6040 17478
rect 6196 17270 6224 17682
rect 6184 17264 6236 17270
rect 6184 17206 6236 17212
rect 6092 17196 6144 17202
rect 6092 17138 6144 17144
rect 6104 16794 6132 17138
rect 6288 16969 6316 19094
rect 6368 18896 6420 18902
rect 6368 18838 6420 18844
rect 6380 17542 6408 18838
rect 6368 17536 6420 17542
rect 6368 17478 6420 17484
rect 6458 17504 6514 17513
rect 6380 17338 6408 17478
rect 6458 17439 6514 17448
rect 6368 17332 6420 17338
rect 6368 17274 6420 17280
rect 6472 17218 6500 17439
rect 6380 17190 6500 17218
rect 6274 16960 6330 16969
rect 6274 16895 6330 16904
rect 6092 16788 6144 16794
rect 6092 16730 6144 16736
rect 6092 16584 6144 16590
rect 6092 16526 6144 16532
rect 6184 16584 6236 16590
rect 6184 16526 6236 16532
rect 6104 15978 6132 16526
rect 6092 15972 6144 15978
rect 6092 15914 6144 15920
rect 6196 15706 6224 16526
rect 6276 15904 6328 15910
rect 6276 15846 6328 15852
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6092 15428 6144 15434
rect 6092 15370 6144 15376
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 6000 15156 6052 15162
rect 6000 15098 6052 15104
rect 6104 15094 6132 15370
rect 6092 15088 6144 15094
rect 6092 15030 6144 15036
rect 6184 14816 6236 14822
rect 6184 14758 6236 14764
rect 6196 14550 6224 14758
rect 6184 14544 6236 14550
rect 6184 14486 6236 14492
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 6196 14074 6224 14486
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 6184 14068 6236 14074
rect 6184 14010 6236 14016
rect 5630 13968 5686 13977
rect 5630 13903 5686 13912
rect 5356 13728 5408 13734
rect 5356 13670 5408 13676
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5170 12880 5226 12889
rect 5276 12850 5304 13330
rect 5368 13258 5396 13670
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 5368 12866 5396 13194
rect 5552 13190 5580 13670
rect 5644 13530 5672 13903
rect 6000 13796 6052 13802
rect 6000 13738 6052 13744
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 6012 13258 6040 13738
rect 6000 13252 6052 13258
rect 6000 13194 6052 13200
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5552 12986 5580 13126
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6012 12986 6040 13194
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 5170 12815 5172 12824
rect 5224 12815 5226 12824
rect 5264 12844 5316 12850
rect 5172 12786 5224 12792
rect 5368 12838 5580 12866
rect 5264 12786 5316 12792
rect 5080 12776 5132 12782
rect 5080 12718 5132 12724
rect 5264 12708 5316 12714
rect 5264 12650 5316 12656
rect 5356 12708 5408 12714
rect 5356 12650 5408 12656
rect 5080 12164 5132 12170
rect 5080 12106 5132 12112
rect 5092 11830 5120 12106
rect 5080 11824 5132 11830
rect 5080 11766 5132 11772
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 5080 11280 5132 11286
rect 5080 11222 5132 11228
rect 5092 10742 5120 11222
rect 5080 10736 5132 10742
rect 5080 10678 5132 10684
rect 5184 10266 5212 11494
rect 5172 10260 5224 10266
rect 5172 10202 5224 10208
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 5184 8974 5212 9318
rect 5172 8968 5224 8974
rect 5078 8936 5134 8945
rect 5172 8910 5224 8916
rect 5078 8871 5134 8880
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4908 8430 4936 8774
rect 5092 8634 5120 8871
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 5184 8090 5212 8910
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 4896 7880 4948 7886
rect 4894 7848 4896 7857
rect 4948 7848 4950 7857
rect 4894 7783 4950 7792
rect 5000 7478 5028 7890
rect 4988 7472 5040 7478
rect 4988 7414 5040 7420
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4816 5166 4844 6054
rect 4908 5778 4936 7346
rect 5000 7002 5028 7414
rect 5276 7290 5304 12650
rect 5368 10810 5396 12650
rect 5446 12472 5502 12481
rect 5552 12442 5580 12838
rect 5446 12407 5502 12416
rect 5540 12436 5592 12442
rect 5460 12238 5488 12407
rect 5540 12378 5592 12384
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5460 11898 5488 12174
rect 6092 12096 6144 12102
rect 6090 12064 6092 12073
rect 6144 12064 6146 12073
rect 5622 11996 5918 12016
rect 6090 11999 6146 12008
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 6104 11694 6132 11999
rect 6196 11898 6224 12242
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 6092 11688 6144 11694
rect 5538 11656 5594 11665
rect 6092 11630 6144 11636
rect 5538 11591 5540 11600
rect 5592 11591 5594 11600
rect 5540 11562 5592 11568
rect 5552 11354 5580 11562
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 6092 11212 6144 11218
rect 6092 11154 6144 11160
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 6104 10130 6132 11154
rect 6196 10198 6224 11698
rect 6288 10742 6316 15846
rect 6380 13569 6408 17190
rect 6460 16992 6512 16998
rect 6460 16934 6512 16940
rect 6472 16182 6500 16934
rect 6564 16810 6592 19230
rect 6644 19168 6696 19174
rect 6644 19110 6696 19116
rect 6656 17814 6684 19110
rect 6734 19000 6790 19009
rect 6734 18935 6790 18944
rect 6644 17808 6696 17814
rect 6644 17750 6696 17756
rect 6656 17649 6684 17750
rect 6642 17640 6698 17649
rect 6642 17575 6698 17584
rect 6748 17338 6776 18935
rect 6840 18834 6868 19926
rect 7024 19310 7052 20862
rect 7196 20256 7248 20262
rect 7194 20224 7196 20233
rect 7248 20224 7250 20233
rect 7194 20159 7250 20168
rect 7208 19990 7236 20159
rect 7196 19984 7248 19990
rect 7196 19926 7248 19932
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7104 19440 7156 19446
rect 7104 19382 7156 19388
rect 7012 19304 7064 19310
rect 7012 19246 7064 19252
rect 7024 18970 7052 19246
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 7010 18864 7066 18873
rect 6828 18828 6880 18834
rect 6880 18788 6960 18816
rect 7010 18799 7066 18808
rect 6828 18770 6880 18776
rect 6828 18624 6880 18630
rect 6828 18566 6880 18572
rect 6840 18290 6868 18566
rect 6828 18284 6880 18290
rect 6828 18226 6880 18232
rect 6932 17882 6960 18788
rect 7024 18358 7052 18799
rect 7012 18352 7064 18358
rect 7012 18294 7064 18300
rect 6920 17876 6972 17882
rect 6840 17836 6920 17864
rect 6736 17332 6788 17338
rect 6736 17274 6788 17280
rect 6564 16782 6776 16810
rect 6642 16688 6698 16697
rect 6642 16623 6644 16632
rect 6696 16623 6698 16632
rect 6644 16594 6696 16600
rect 6552 16584 6604 16590
rect 6552 16526 6604 16532
rect 6460 16176 6512 16182
rect 6460 16118 6512 16124
rect 6564 15706 6592 16526
rect 6644 16516 6696 16522
rect 6644 16458 6696 16464
rect 6656 16250 6684 16458
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 6656 15881 6684 16186
rect 6642 15872 6698 15881
rect 6642 15807 6698 15816
rect 6552 15700 6604 15706
rect 6552 15642 6604 15648
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6564 14618 6592 15302
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6564 14414 6592 14554
rect 6644 14476 6696 14482
rect 6644 14418 6696 14424
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 6366 13560 6422 13569
rect 6366 13495 6422 13504
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6366 13152 6422 13161
rect 6366 13087 6422 13096
rect 6276 10736 6328 10742
rect 6276 10678 6328 10684
rect 6184 10192 6236 10198
rect 6184 10134 6236 10140
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 5460 9625 5488 10066
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 6012 9926 6040 9998
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5446 9616 5502 9625
rect 5446 9551 5502 9560
rect 5460 9178 5488 9551
rect 6012 9518 6040 9862
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 6012 9110 6040 9318
rect 6000 9104 6052 9110
rect 6000 9046 6052 9052
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 5460 8430 5488 8842
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5552 8276 5580 8978
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5460 8248 5580 8276
rect 6012 8265 6040 9046
rect 5998 8256 6054 8265
rect 5460 8022 5488 8248
rect 5998 8191 6054 8200
rect 5448 8016 5500 8022
rect 5448 7958 5500 7964
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5998 7576 6054 7585
rect 5998 7511 6054 7520
rect 5092 7262 5304 7290
rect 6012 7274 6040 7511
rect 6000 7268 6052 7274
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 5000 6254 5028 6938
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 4908 5234 4936 5714
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4804 5160 4856 5166
rect 4804 5102 4856 5108
rect 4816 4486 4844 5102
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4816 4214 4844 4422
rect 4908 4298 4936 5170
rect 5000 4758 5028 6054
rect 5092 5370 5120 7262
rect 6000 7210 6052 7216
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5184 6798 5212 7142
rect 5630 6896 5686 6905
rect 5356 6860 5408 6866
rect 5630 6831 5632 6840
rect 5356 6802 5408 6808
rect 5684 6831 5686 6840
rect 5632 6802 5684 6808
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5184 5914 5212 6734
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 5092 5114 5120 5306
rect 5092 5086 5212 5114
rect 5184 5030 5212 5086
rect 5080 5024 5132 5030
rect 5080 4966 5132 4972
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5092 4826 5120 4966
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 4988 4752 5040 4758
rect 4988 4694 5040 4700
rect 5276 4690 5304 6598
rect 5368 6254 5396 6802
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6012 6322 6040 6734
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 6012 6118 6040 6258
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 5448 5840 5500 5846
rect 5448 5782 5500 5788
rect 5460 5658 5488 5782
rect 5460 5630 5580 5658
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 5262 4584 5318 4593
rect 5262 4519 5318 4528
rect 4908 4270 5028 4298
rect 5000 4214 5028 4270
rect 4804 4208 4856 4214
rect 4804 4150 4856 4156
rect 4988 4208 5040 4214
rect 4988 4150 5040 4156
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 4724 3194 4752 3470
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 5092 2582 5120 2790
rect 4620 2576 4672 2582
rect 4620 2518 4672 2524
rect 5080 2576 5132 2582
rect 5080 2518 5132 2524
rect 5092 2009 5120 2518
rect 5078 2000 5134 2009
rect 5078 1935 5134 1944
rect 5184 1442 5212 3946
rect 5276 3602 5304 4519
rect 5460 4486 5488 5102
rect 5552 4758 5580 5630
rect 6012 5574 6040 6054
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6012 5234 6040 5510
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 5540 4752 5592 4758
rect 5540 4694 5592 4700
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5460 4282 5488 4422
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5538 4040 5594 4049
rect 6012 4010 6040 4626
rect 5538 3975 5594 3984
rect 6000 4004 6052 4010
rect 5552 3738 5580 3975
rect 6000 3946 6052 3952
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 6104 3670 6132 9862
rect 6196 9722 6224 10134
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6184 9716 6236 9722
rect 6184 9658 6236 9664
rect 6288 9586 6316 10066
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6288 8974 6316 9522
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6288 8498 6316 8774
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 6182 8256 6238 8265
rect 6182 8191 6238 8200
rect 6092 3664 6144 3670
rect 6092 3606 6144 3612
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 5276 3194 5304 3538
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5460 2310 5488 3470
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6012 2650 6040 3538
rect 6104 3194 6132 3606
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 5460 1714 5488 2246
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5460 1686 5672 1714
rect 5092 1414 5212 1442
rect 5092 480 5120 1414
rect 5644 480 5672 1686
rect 6196 480 6224 8191
rect 6288 8090 6316 8434
rect 6276 8084 6328 8090
rect 6276 8026 6328 8032
rect 6380 7342 6408 13087
rect 6472 12918 6500 13262
rect 6460 12912 6512 12918
rect 6460 12854 6512 12860
rect 6564 12850 6592 14350
rect 6656 14249 6684 14418
rect 6642 14240 6698 14249
rect 6642 14175 6698 14184
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6564 12730 6592 12786
rect 6472 12702 6592 12730
rect 6472 12238 6500 12702
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6564 12374 6592 12582
rect 6552 12368 6604 12374
rect 6552 12310 6604 12316
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6472 11762 6500 12174
rect 6564 11898 6592 12310
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6472 9489 6500 10950
rect 6656 10810 6684 14175
rect 6748 13394 6776 16782
rect 6840 15366 6868 17836
rect 6920 17818 6972 17824
rect 7116 17218 7144 19382
rect 7208 18834 7236 19654
rect 7286 19000 7342 19009
rect 7286 18935 7342 18944
rect 7196 18828 7248 18834
rect 7196 18770 7248 18776
rect 7208 18426 7236 18770
rect 7196 18420 7248 18426
rect 7196 18362 7248 18368
rect 7208 17882 7236 18362
rect 7196 17876 7248 17882
rect 7196 17818 7248 17824
rect 7024 17190 7144 17218
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6932 15026 6960 15642
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6840 14074 6868 14894
rect 7024 14657 7052 17190
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 7116 16114 7144 17070
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 7208 16697 7236 16730
rect 7194 16688 7250 16697
rect 7194 16623 7250 16632
rect 7104 16108 7156 16114
rect 7104 16050 7156 16056
rect 7196 15972 7248 15978
rect 7196 15914 7248 15920
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 7116 14890 7144 15438
rect 7104 14884 7156 14890
rect 7104 14826 7156 14832
rect 7010 14648 7066 14657
rect 7010 14583 7066 14592
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6840 13530 6868 13806
rect 7024 13530 7052 14583
rect 7116 13938 7144 14826
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 6748 13025 6776 13330
rect 6734 13016 6790 13025
rect 6734 12951 6736 12960
rect 6788 12951 6790 12960
rect 6736 12922 6788 12928
rect 6748 12891 6776 12922
rect 7208 12481 7236 15914
rect 7194 12472 7250 12481
rect 7194 12407 7250 12416
rect 6734 12336 6790 12345
rect 6734 12271 6790 12280
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6550 9888 6606 9897
rect 6550 9823 6606 9832
rect 6458 9480 6514 9489
rect 6564 9450 6592 9823
rect 6458 9415 6514 9424
rect 6552 9444 6604 9450
rect 6552 9386 6604 9392
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6472 8634 6500 8910
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6472 7954 6500 8570
rect 6642 7984 6698 7993
rect 6460 7948 6512 7954
rect 6642 7919 6698 7928
rect 6460 7890 6512 7896
rect 6656 7721 6684 7919
rect 6642 7712 6698 7721
rect 6642 7647 6698 7656
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6656 6934 6684 7142
rect 6644 6928 6696 6934
rect 6366 6896 6422 6905
rect 6644 6870 6696 6876
rect 6366 6831 6422 6840
rect 6380 5914 6408 6831
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6472 4758 6500 4966
rect 6460 4752 6512 4758
rect 6460 4694 6512 4700
rect 6472 3942 6500 4694
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6472 3602 6500 3878
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6642 2952 6698 2961
rect 6276 2916 6328 2922
rect 6642 2887 6644 2896
rect 6276 2858 6328 2864
rect 6696 2887 6698 2896
rect 6644 2858 6696 2864
rect 6288 1193 6316 2858
rect 6274 1184 6330 1193
rect 6274 1119 6330 1128
rect 6748 480 6776 12271
rect 6828 11552 6880 11558
rect 6826 11520 6828 11529
rect 6880 11520 6882 11529
rect 6826 11455 6882 11464
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6840 10606 6868 11290
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6840 9178 6868 10406
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6840 8430 6868 9114
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6932 8362 6960 11018
rect 7196 10600 7248 10606
rect 7300 10588 7328 18935
rect 7576 18737 7604 23462
rect 7654 22808 7710 22817
rect 7654 22743 7710 22752
rect 7668 22574 7696 22743
rect 7656 22568 7708 22574
rect 7656 22510 7708 22516
rect 7656 21344 7708 21350
rect 7656 21286 7708 21292
rect 7668 20058 7696 21286
rect 7656 20052 7708 20058
rect 7656 19994 7708 20000
rect 7668 19378 7696 19994
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7562 18728 7618 18737
rect 7562 18663 7618 18672
rect 7564 18624 7616 18630
rect 7564 18566 7616 18572
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 7484 17338 7512 18226
rect 7576 18086 7604 18566
rect 7564 18080 7616 18086
rect 7564 18022 7616 18028
rect 7564 17740 7616 17746
rect 7564 17682 7616 17688
rect 7472 17332 7524 17338
rect 7472 17274 7524 17280
rect 7576 17066 7604 17682
rect 7564 17060 7616 17066
rect 7564 17002 7616 17008
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7484 15910 7512 16526
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7484 13326 7512 14962
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7484 12714 7512 13126
rect 7472 12708 7524 12714
rect 7472 12650 7524 12656
rect 7576 12458 7604 17002
rect 7760 16794 7788 24647
rect 7944 24410 7972 25735
rect 7932 24404 7984 24410
rect 7932 24346 7984 24352
rect 8036 23866 8064 25774
rect 8024 23860 8076 23866
rect 8024 23802 8076 23808
rect 7840 23792 7892 23798
rect 8128 23746 8156 25871
rect 8404 24834 8432 27520
rect 8944 25764 8996 25770
rect 8944 25706 8996 25712
rect 8852 25152 8904 25158
rect 8852 25094 8904 25100
rect 8404 24806 8800 24834
rect 8668 24404 8720 24410
rect 8668 24346 8720 24352
rect 8680 24313 8708 24346
rect 8666 24304 8722 24313
rect 8300 24268 8352 24274
rect 8666 24239 8722 24248
rect 8300 24210 8352 24216
rect 7840 23734 7892 23740
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 7656 16652 7708 16658
rect 7656 16594 7708 16600
rect 7668 15910 7696 16594
rect 7760 16250 7788 16730
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 7668 15609 7696 15846
rect 7654 15600 7710 15609
rect 7654 15535 7710 15544
rect 7656 15360 7708 15366
rect 7654 15328 7656 15337
rect 7708 15328 7710 15337
rect 7654 15263 7710 15272
rect 7748 14340 7800 14346
rect 7748 14282 7800 14288
rect 7484 12430 7604 12458
rect 7378 11384 7434 11393
rect 7378 11319 7380 11328
rect 7432 11319 7434 11328
rect 7380 11290 7432 11296
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 7392 10849 7420 11154
rect 7378 10840 7434 10849
rect 7378 10775 7434 10784
rect 7380 10736 7432 10742
rect 7380 10678 7432 10684
rect 7248 10560 7328 10588
rect 7196 10542 7248 10548
rect 7392 8548 7420 10678
rect 7484 10554 7512 12430
rect 7562 12200 7618 12209
rect 7562 12135 7618 12144
rect 7576 11898 7604 12135
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 7576 10674 7604 11086
rect 7654 10976 7710 10985
rect 7654 10911 7710 10920
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7484 10526 7604 10554
rect 7208 8520 7420 8548
rect 7102 8392 7158 8401
rect 6920 8356 6972 8362
rect 7102 8327 7158 8336
rect 6920 8298 6972 8304
rect 6918 7984 6974 7993
rect 7116 7954 7144 8327
rect 6918 7919 6920 7928
rect 6972 7919 6974 7928
rect 7104 7948 7156 7954
rect 6920 7890 6972 7896
rect 7104 7890 7156 7896
rect 6932 7410 6960 7890
rect 7010 7848 7066 7857
rect 7010 7783 7012 7792
rect 7064 7783 7066 7792
rect 7012 7754 7064 7760
rect 7010 7440 7066 7449
rect 6920 7404 6972 7410
rect 7010 7375 7066 7384
rect 6920 7346 6972 7352
rect 7024 6866 7052 7375
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 6826 6624 6882 6633
rect 6826 6559 6882 6568
rect 6840 5914 6868 6559
rect 7024 6458 7052 6802
rect 7116 6798 7144 7890
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7208 6730 7236 8520
rect 7576 8480 7604 10526
rect 7668 10169 7696 10911
rect 7760 10742 7788 14282
rect 7852 11218 7880 23734
rect 7944 23718 8156 23746
rect 7944 19938 7972 23718
rect 8312 23594 8340 24210
rect 8300 23588 8352 23594
rect 8300 23530 8352 23536
rect 8312 23474 8340 23530
rect 8220 23446 8340 23474
rect 8220 23254 8248 23446
rect 8208 23248 8260 23254
rect 8208 23190 8260 23196
rect 8666 23216 8722 23225
rect 8666 23151 8722 23160
rect 8116 22636 8168 22642
rect 8116 22578 8168 22584
rect 8128 21962 8156 22578
rect 8208 22432 8260 22438
rect 8206 22400 8208 22409
rect 8260 22400 8262 22409
rect 8206 22335 8262 22344
rect 8390 21992 8446 22001
rect 8116 21956 8168 21962
rect 8390 21927 8446 21936
rect 8116 21898 8168 21904
rect 8208 21480 8260 21486
rect 8208 21422 8260 21428
rect 8024 21004 8076 21010
rect 8024 20946 8076 20952
rect 8036 20058 8064 20946
rect 8114 20632 8170 20641
rect 8114 20567 8170 20576
rect 8024 20052 8076 20058
rect 8024 19994 8076 20000
rect 7944 19910 8064 19938
rect 8036 19854 8064 19910
rect 8024 19848 8076 19854
rect 8024 19790 8076 19796
rect 8036 19174 8064 19790
rect 8024 19168 8076 19174
rect 8024 19110 8076 19116
rect 7932 18352 7984 18358
rect 7932 18294 7984 18300
rect 7944 18193 7972 18294
rect 7930 18184 7986 18193
rect 7930 18119 7986 18128
rect 7944 18086 7972 18119
rect 7932 18080 7984 18086
rect 7932 18022 7984 18028
rect 8036 16017 8064 19110
rect 8128 19009 8156 20567
rect 8220 19310 8248 21422
rect 8300 20868 8352 20874
rect 8300 20810 8352 20816
rect 8312 20602 8340 20810
rect 8300 20596 8352 20602
rect 8300 20538 8352 20544
rect 8404 20534 8432 21927
rect 8482 21312 8538 21321
rect 8482 21247 8538 21256
rect 8392 20528 8444 20534
rect 8392 20470 8444 20476
rect 8392 19916 8444 19922
rect 8392 19858 8444 19864
rect 8298 19816 8354 19825
rect 8298 19751 8354 19760
rect 8208 19304 8260 19310
rect 8208 19246 8260 19252
rect 8312 19242 8340 19751
rect 8404 19514 8432 19858
rect 8392 19508 8444 19514
rect 8392 19450 8444 19456
rect 8300 19236 8352 19242
rect 8300 19178 8352 19184
rect 8114 19000 8170 19009
rect 8312 18970 8340 19178
rect 8114 18935 8170 18944
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 8496 18902 8524 21247
rect 8680 21078 8708 23151
rect 8668 21072 8720 21078
rect 8668 21014 8720 21020
rect 8668 20460 8720 20466
rect 8668 20402 8720 20408
rect 8574 20088 8630 20097
rect 8574 20023 8630 20032
rect 8588 19700 8616 20023
rect 8680 19854 8708 20402
rect 8668 19848 8720 19854
rect 8668 19790 8720 19796
rect 8588 19672 8708 19700
rect 8484 18896 8536 18902
rect 8536 18856 8616 18884
rect 8484 18838 8536 18844
rect 8300 18352 8352 18358
rect 8300 18294 8352 18300
rect 8482 18320 8538 18329
rect 8208 18216 8260 18222
rect 8208 18158 8260 18164
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 8128 17105 8156 17478
rect 8220 17320 8248 18158
rect 8312 17490 8340 18294
rect 8482 18255 8538 18264
rect 8496 17882 8524 18255
rect 8588 18222 8616 18856
rect 8576 18216 8628 18222
rect 8576 18158 8628 18164
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8484 17876 8536 17882
rect 8484 17818 8536 17824
rect 8390 17776 8446 17785
rect 8390 17711 8392 17720
rect 8444 17711 8446 17720
rect 8392 17682 8444 17688
rect 8312 17462 8432 17490
rect 8300 17332 8352 17338
rect 8220 17292 8300 17320
rect 8300 17274 8352 17280
rect 8114 17096 8170 17105
rect 8114 17031 8170 17040
rect 8128 16998 8156 17031
rect 8116 16992 8168 16998
rect 8116 16934 8168 16940
rect 8404 16794 8432 17462
rect 8588 17134 8616 18022
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8482 16824 8538 16833
rect 8392 16788 8444 16794
rect 8588 16794 8616 17070
rect 8482 16759 8538 16768
rect 8576 16788 8628 16794
rect 8392 16730 8444 16736
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 8312 16114 8340 16390
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 8404 16046 8432 16730
rect 8392 16040 8444 16046
rect 8022 16008 8078 16017
rect 8022 15943 8078 15952
rect 8390 16008 8392 16017
rect 8444 16008 8446 16017
rect 8390 15943 8446 15952
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 8128 14414 8156 15506
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8220 15178 8248 15438
rect 8392 15360 8444 15366
rect 8392 15302 8444 15308
rect 8220 15162 8340 15178
rect 8220 15156 8352 15162
rect 8220 15150 8300 15156
rect 8300 15098 8352 15104
rect 8404 15042 8432 15302
rect 8220 15014 8432 15042
rect 8220 14958 8248 15014
rect 8496 14958 8524 16759
rect 8576 16730 8628 16736
rect 8576 16448 8628 16454
rect 8576 16390 8628 16396
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 8036 13938 8064 14214
rect 8024 13932 8076 13938
rect 8024 13874 8076 13880
rect 8588 13870 8616 16390
rect 8680 15638 8708 19672
rect 8772 17320 8800 24806
rect 8864 24614 8892 25094
rect 8852 24608 8904 24614
rect 8852 24550 8904 24556
rect 8864 24070 8892 24550
rect 8852 24064 8904 24070
rect 8852 24006 8904 24012
rect 8956 24018 8984 25706
rect 9048 24857 9076 27520
rect 9034 24848 9090 24857
rect 9034 24783 9090 24792
rect 8864 23882 8892 24006
rect 8956 23990 9076 24018
rect 8864 23854 8984 23882
rect 8956 23526 8984 23854
rect 8944 23520 8996 23526
rect 8850 23488 8906 23497
rect 8944 23462 8996 23468
rect 8850 23423 8906 23432
rect 8864 21434 8892 23423
rect 8956 22982 8984 23462
rect 8944 22976 8996 22982
rect 8944 22918 8996 22924
rect 8956 22030 8984 22918
rect 9048 22778 9076 23990
rect 9140 23866 9168 27542
rect 9586 27520 9642 28000
rect 10138 27520 10194 28000
rect 10782 27520 10838 28000
rect 11334 27520 11390 28000
rect 11886 27520 11942 28000
rect 12530 27520 12586 28000
rect 13082 27520 13138 28000
rect 13634 27520 13690 28000
rect 14278 27520 14334 28000
rect 14830 27520 14886 28000
rect 15382 27520 15438 28000
rect 16026 27520 16082 28000
rect 16578 27520 16634 28000
rect 17130 27520 17186 28000
rect 17774 27520 17830 28000
rect 18326 27520 18382 28000
rect 18878 27520 18934 28000
rect 19522 27520 19578 28000
rect 20074 27520 20130 28000
rect 20626 27520 20682 28000
rect 21270 27520 21326 28000
rect 21822 27520 21878 28000
rect 22374 27520 22430 28000
rect 23018 27520 23074 28000
rect 23570 27520 23626 28000
rect 24122 27520 24178 28000
rect 24766 27520 24822 28000
rect 25318 27520 25374 28000
rect 25870 27520 25926 28000
rect 26054 27704 26110 27713
rect 26054 27639 26110 27648
rect 9220 26036 9272 26042
rect 9220 25978 9272 25984
rect 9232 24954 9260 25978
rect 9494 24984 9550 24993
rect 9220 24948 9272 24954
rect 9220 24890 9272 24896
rect 9312 24948 9364 24954
rect 9494 24919 9550 24928
rect 9312 24890 9364 24896
rect 9128 23860 9180 23866
rect 9128 23802 9180 23808
rect 9324 23798 9352 24890
rect 9508 23866 9536 24919
rect 9496 23860 9548 23866
rect 9496 23802 9548 23808
rect 9312 23792 9364 23798
rect 9312 23734 9364 23740
rect 9508 23662 9536 23802
rect 9496 23656 9548 23662
rect 9496 23598 9548 23604
rect 9312 23180 9364 23186
rect 9312 23122 9364 23128
rect 9036 22772 9088 22778
rect 9036 22714 9088 22720
rect 9036 22568 9088 22574
rect 9036 22510 9088 22516
rect 8944 22024 8996 22030
rect 8944 21966 8996 21972
rect 8956 21554 8984 21966
rect 9048 21894 9076 22510
rect 9218 22128 9274 22137
rect 9218 22063 9274 22072
rect 9036 21888 9088 21894
rect 9036 21830 9088 21836
rect 9128 21888 9180 21894
rect 9128 21830 9180 21836
rect 8944 21548 8996 21554
rect 8944 21490 8996 21496
rect 8864 21406 8984 21434
rect 8852 21344 8904 21350
rect 8852 21286 8904 21292
rect 8864 20874 8892 21286
rect 8852 20868 8904 20874
rect 8852 20810 8904 20816
rect 8956 20584 8984 21406
rect 9048 21146 9076 21830
rect 9036 21140 9088 21146
rect 9036 21082 9088 21088
rect 8864 20556 8984 20584
rect 8864 18034 8892 20556
rect 8942 20360 8998 20369
rect 9140 20346 9168 21830
rect 8942 20295 8944 20304
rect 8996 20295 8998 20304
rect 9048 20318 9168 20346
rect 8944 20266 8996 20272
rect 9048 18714 9076 20318
rect 9128 20256 9180 20262
rect 9128 20198 9180 20204
rect 9140 19718 9168 20198
rect 9128 19712 9180 19718
rect 9126 19680 9128 19689
rect 9180 19680 9182 19689
rect 9126 19615 9182 19624
rect 9048 18686 9168 18714
rect 9034 18592 9090 18601
rect 9034 18527 9090 18536
rect 9048 18290 9076 18527
rect 9036 18284 9088 18290
rect 9036 18226 9088 18232
rect 8864 18006 8984 18034
rect 8850 17912 8906 17921
rect 8850 17847 8852 17856
rect 8904 17847 8906 17856
rect 8852 17818 8904 17824
rect 8772 17292 8892 17320
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8772 16658 8800 17138
rect 8760 16652 8812 16658
rect 8760 16594 8812 16600
rect 8668 15632 8720 15638
rect 8668 15574 8720 15580
rect 8864 15162 8892 17292
rect 8956 17270 8984 18006
rect 8944 17264 8996 17270
rect 8944 17206 8996 17212
rect 9034 17232 9090 17241
rect 9034 17167 9090 17176
rect 8942 17096 8998 17105
rect 8942 17031 8998 17040
rect 8852 15156 8904 15162
rect 8852 15098 8904 15104
rect 8956 15042 8984 17031
rect 9048 16794 9076 17167
rect 9036 16788 9088 16794
rect 9036 16730 9088 16736
rect 9034 15872 9090 15881
rect 9034 15807 9090 15816
rect 8772 15014 8984 15042
rect 8576 13864 8628 13870
rect 8022 13832 8078 13841
rect 8576 13806 8628 13812
rect 8022 13767 8078 13776
rect 8036 13530 8064 13767
rect 8588 13734 8616 13806
rect 8772 13802 8800 15014
rect 8850 14920 8906 14929
rect 8850 14855 8852 14864
rect 8904 14855 8906 14864
rect 8852 14826 8904 14832
rect 8864 14618 8892 14826
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8942 14512 8998 14521
rect 8942 14447 8998 14456
rect 8956 14278 8984 14447
rect 8944 14272 8996 14278
rect 8942 14240 8944 14249
rect 8996 14240 8998 14249
rect 8942 14175 8998 14184
rect 8852 14068 8904 14074
rect 8852 14010 8904 14016
rect 8760 13796 8812 13802
rect 8760 13738 8812 13744
rect 8576 13728 8628 13734
rect 8576 13670 8628 13676
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8300 13456 8352 13462
rect 8300 13398 8352 13404
rect 7932 13184 7984 13190
rect 7932 13126 7984 13132
rect 7944 12850 7972 13126
rect 8206 13016 8262 13025
rect 8206 12951 8262 12960
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 8024 12640 8076 12646
rect 8022 12608 8024 12617
rect 8076 12608 8078 12617
rect 8022 12543 8078 12552
rect 8114 12336 8170 12345
rect 8114 12271 8170 12280
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7944 11830 7972 12038
rect 7932 11824 7984 11830
rect 7932 11766 7984 11772
rect 7944 11694 7972 11766
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 8128 11354 8156 12271
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 7838 11112 7894 11121
rect 7838 11047 7894 11056
rect 8116 11076 8168 11082
rect 7748 10736 7800 10742
rect 7748 10678 7800 10684
rect 7654 10160 7710 10169
rect 7654 10095 7710 10104
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7668 8809 7696 8978
rect 7852 8838 7880 11047
rect 8116 11018 8168 11024
rect 7930 10568 7986 10577
rect 7930 10503 7932 10512
rect 7984 10503 7986 10512
rect 7932 10474 7984 10480
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 8036 9518 8064 9862
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 7932 9104 7984 9110
rect 7932 9046 7984 9052
rect 7840 8832 7892 8838
rect 7654 8800 7710 8809
rect 7840 8774 7892 8780
rect 7654 8735 7710 8744
rect 7668 8634 7696 8735
rect 7944 8673 7972 9046
rect 8036 8906 8064 9454
rect 8128 9450 8156 11018
rect 8116 9444 8168 9450
rect 8116 9386 8168 9392
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 7930 8664 7986 8673
rect 7656 8628 7708 8634
rect 7930 8599 7932 8608
rect 7656 8570 7708 8576
rect 7984 8599 7986 8608
rect 7932 8570 7984 8576
rect 7392 8452 7604 8480
rect 7286 7576 7342 7585
rect 7286 7511 7342 7520
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6828 5024 6880 5030
rect 6932 5012 6960 5714
rect 6880 4984 6960 5012
rect 6828 4966 6880 4972
rect 6826 4720 6882 4729
rect 6826 4655 6882 4664
rect 6840 4146 6868 4655
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6840 2145 6868 3334
rect 6826 2136 6882 2145
rect 6826 2071 6882 2080
rect 6932 1329 6960 4984
rect 6918 1320 6974 1329
rect 6918 1255 6974 1264
rect 4250 368 4306 377
rect 4250 303 4306 312
rect 4526 0 4582 480
rect 5078 0 5134 480
rect 5630 0 5686 480
rect 6182 0 6238 480
rect 6734 0 6790 480
rect 7116 377 7144 6598
rect 7194 6216 7250 6225
rect 7194 6151 7250 6160
rect 7208 6118 7236 6151
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 7300 5522 7328 7511
rect 7392 7274 7420 8452
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7576 8090 7604 8298
rect 7654 8120 7710 8129
rect 7564 8084 7616 8090
rect 7654 8055 7656 8064
rect 7564 8026 7616 8032
rect 7708 8055 7710 8064
rect 7656 8026 7708 8032
rect 7668 7546 7696 8026
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7380 7268 7432 7274
rect 7380 7210 7432 7216
rect 7576 6769 7604 7346
rect 7562 6760 7618 6769
rect 7562 6695 7564 6704
rect 7616 6695 7618 6704
rect 7564 6666 7616 6672
rect 7760 6633 7788 7686
rect 8220 7562 8248 12951
rect 8312 12442 8340 13398
rect 8390 12744 8446 12753
rect 8390 12679 8446 12688
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 8298 10840 8354 10849
rect 8298 10775 8300 10784
rect 8352 10775 8354 10784
rect 8300 10746 8352 10752
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8312 10266 8340 10542
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8298 9072 8354 9081
rect 8298 9007 8354 9016
rect 8312 8022 8340 9007
rect 8404 8634 8432 12679
rect 8680 12442 8708 13466
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 8482 11928 8538 11937
rect 8482 11863 8538 11872
rect 8496 11354 8524 11863
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8496 10606 8524 11154
rect 8484 10600 8536 10606
rect 8484 10542 8536 10548
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8404 8430 8432 8570
rect 8392 8424 8444 8430
rect 8496 8401 8524 10406
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8392 8366 8444 8372
rect 8482 8392 8538 8401
rect 8482 8327 8538 8336
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 7852 7534 8248 7562
rect 7746 6624 7802 6633
rect 7746 6559 7802 6568
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 7576 5846 7604 6190
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7564 5840 7616 5846
rect 7562 5808 7564 5817
rect 7616 5808 7618 5817
rect 7562 5743 7618 5752
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 7208 5494 7328 5522
rect 7208 3346 7236 5494
rect 7286 5400 7342 5409
rect 7286 5335 7342 5344
rect 7300 4826 7328 5335
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7392 3738 7420 3878
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7286 3496 7342 3505
rect 7286 3431 7288 3440
rect 7340 3431 7342 3440
rect 7288 3402 7340 3408
rect 7208 3318 7328 3346
rect 7194 3224 7250 3233
rect 7194 3159 7250 3168
rect 7208 2990 7236 3159
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 7208 2825 7236 2926
rect 7194 2816 7250 2825
rect 7194 2751 7250 2760
rect 7208 2650 7236 2751
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7300 480 7328 3318
rect 7102 368 7158 377
rect 7102 303 7158 312
rect 7286 0 7342 480
rect 7576 241 7604 5578
rect 7668 5098 7696 6054
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7656 5092 7708 5098
rect 7656 5034 7708 5040
rect 7760 4826 7788 5646
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7668 3058 7696 3878
rect 7760 3126 7788 4014
rect 7748 3120 7800 3126
rect 7748 3062 7800 3068
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 7668 2825 7696 2994
rect 7654 2816 7710 2825
rect 7654 2751 7710 2760
rect 7746 2680 7802 2689
rect 7746 2615 7802 2624
rect 7760 2514 7788 2615
rect 7748 2508 7800 2514
rect 7748 2450 7800 2456
rect 7852 480 7880 7534
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 8312 6882 8340 7414
rect 8220 6854 8340 6882
rect 8220 6730 8248 6854
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 8036 5953 8064 6598
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8022 5944 8078 5953
rect 8022 5879 8078 5888
rect 8128 5710 8156 6054
rect 8116 5704 8168 5710
rect 8022 5672 8078 5681
rect 8116 5646 8168 5652
rect 8022 5607 8024 5616
rect 8076 5607 8078 5616
rect 8024 5578 8076 5584
rect 8220 5574 8248 6666
rect 8404 6254 8432 8230
rect 8588 7342 8616 8910
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8680 8362 8708 8774
rect 8668 8356 8720 8362
rect 8668 8298 8720 8304
rect 8772 7954 8800 13738
rect 8864 13190 8892 14010
rect 9048 13546 9076 15807
rect 9140 14618 9168 18686
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 8956 13518 9076 13546
rect 8852 13184 8904 13190
rect 8852 13126 8904 13132
rect 8956 12866 8984 13518
rect 9034 13424 9090 13433
rect 9140 13394 9168 14554
rect 9034 13359 9090 13368
rect 9128 13388 9180 13394
rect 9048 12986 9076 13359
rect 9128 13330 9180 13336
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 9140 12918 9168 13126
rect 9128 12912 9180 12918
rect 8956 12838 9076 12866
rect 9128 12854 9180 12860
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8864 10674 8892 12582
rect 8942 11248 8998 11257
rect 8942 11183 8998 11192
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8864 9110 8892 10610
rect 8852 9104 8904 9110
rect 8852 9046 8904 9052
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8864 7886 8892 8366
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8864 7750 8892 7822
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8864 7478 8892 7686
rect 8852 7472 8904 7478
rect 8852 7414 8904 7420
rect 8956 7410 8984 11183
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 8496 6934 8524 7142
rect 8588 7002 8616 7278
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8484 6928 8536 6934
rect 8484 6870 8536 6876
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8496 6633 8524 6734
rect 8576 6656 8628 6662
rect 8482 6624 8538 6633
rect 8576 6598 8628 6604
rect 8482 6559 8538 6568
rect 8588 6322 8616 6598
rect 8680 6322 8708 6734
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8404 5828 8432 6190
rect 8588 5914 8616 6258
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8484 5840 8536 5846
rect 8404 5800 8484 5828
rect 8484 5782 8536 5788
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8208 5568 8260 5574
rect 7930 5536 7986 5545
rect 8208 5510 8260 5516
rect 7930 5471 7986 5480
rect 7944 2922 7972 5471
rect 8312 5386 8340 5714
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8128 5370 8340 5386
rect 8116 5364 8340 5370
rect 8168 5358 8340 5364
rect 8116 5306 8168 5312
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8300 4480 8352 4486
rect 8220 4428 8300 4434
rect 8220 4422 8352 4428
rect 8220 4406 8340 4422
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 8036 2990 8064 3538
rect 8220 3194 8248 4406
rect 8404 4078 8432 5102
rect 8680 4826 8708 5646
rect 8852 5092 8904 5098
rect 8852 5034 8904 5040
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8404 3738 8432 4014
rect 8496 3738 8524 4626
rect 8666 4584 8722 4593
rect 8666 4519 8668 4528
rect 8720 4519 8722 4528
rect 8668 4490 8720 4496
rect 8864 4214 8892 5034
rect 9048 4842 9076 12838
rect 9128 12776 9180 12782
rect 9128 12718 9180 12724
rect 9140 11830 9168 12718
rect 9128 11824 9180 11830
rect 9128 11766 9180 11772
rect 9232 11354 9260 22063
rect 9324 20602 9352 23122
rect 9496 23044 9548 23050
rect 9496 22986 9548 22992
rect 9404 22704 9456 22710
rect 9404 22646 9456 22652
rect 9416 22166 9444 22646
rect 9508 22642 9536 22986
rect 9496 22636 9548 22642
rect 9496 22578 9548 22584
rect 9404 22160 9456 22166
rect 9404 22102 9456 22108
rect 9416 21978 9444 22102
rect 9494 21992 9550 22001
rect 9416 21950 9494 21978
rect 9494 21927 9550 21936
rect 9600 21894 9628 27520
rect 9956 25900 10008 25906
rect 9956 25842 10008 25848
rect 9864 25288 9916 25294
rect 9864 25230 9916 25236
rect 9678 25120 9734 25129
rect 9678 25055 9734 25064
rect 9588 21888 9640 21894
rect 9588 21830 9640 21836
rect 9496 21412 9548 21418
rect 9496 21354 9548 21360
rect 9404 21344 9456 21350
rect 9404 21286 9456 21292
rect 9312 20596 9364 20602
rect 9312 20538 9364 20544
rect 9310 20496 9366 20505
rect 9416 20466 9444 21286
rect 9508 20942 9536 21354
rect 9692 21146 9720 25055
rect 9876 24886 9904 25230
rect 9864 24880 9916 24886
rect 9770 24848 9826 24857
rect 9864 24822 9916 24828
rect 9770 24783 9826 24792
rect 9680 21140 9732 21146
rect 9680 21082 9732 21088
rect 9588 21004 9640 21010
rect 9588 20946 9640 20952
rect 9496 20936 9548 20942
rect 9496 20878 9548 20884
rect 9600 20890 9628 20946
rect 9600 20862 9720 20890
rect 9496 20800 9548 20806
rect 9496 20742 9548 20748
rect 9310 20431 9366 20440
rect 9404 20460 9456 20466
rect 9324 18426 9352 20431
rect 9404 20402 9456 20408
rect 9508 20369 9536 20742
rect 9692 20602 9720 20862
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9678 20496 9734 20505
rect 9678 20431 9734 20440
rect 9494 20360 9550 20369
rect 9494 20295 9550 20304
rect 9588 20256 9640 20262
rect 9586 20224 9588 20233
rect 9640 20224 9642 20233
rect 9586 20159 9642 20168
rect 9588 19780 9640 19786
rect 9588 19722 9640 19728
rect 9494 19544 9550 19553
rect 9494 19479 9550 19488
rect 9404 19304 9456 19310
rect 9404 19246 9456 19252
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 9416 18222 9444 19246
rect 9404 18216 9456 18222
rect 9324 18176 9404 18204
rect 9324 17202 9352 18176
rect 9404 18158 9456 18164
rect 9402 17640 9458 17649
rect 9402 17575 9458 17584
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 9312 17060 9364 17066
rect 9312 17002 9364 17008
rect 9324 16561 9352 17002
rect 9416 16794 9444 17575
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 9310 16552 9366 16561
rect 9310 16487 9366 16496
rect 9402 15736 9458 15745
rect 9402 15671 9404 15680
rect 9456 15671 9458 15680
rect 9404 15642 9456 15648
rect 9402 15192 9458 15201
rect 9402 15127 9458 15136
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 9324 12345 9352 14418
rect 9416 13802 9444 15127
rect 9404 13796 9456 13802
rect 9404 13738 9456 13744
rect 9508 13394 9536 19479
rect 9600 18873 9628 19722
rect 9586 18864 9642 18873
rect 9586 18799 9642 18808
rect 9692 17898 9720 20431
rect 9784 18714 9812 24783
rect 9968 23746 9996 25842
rect 10048 24608 10100 24614
rect 10048 24550 10100 24556
rect 9876 23718 9996 23746
rect 9876 21010 9904 23718
rect 10060 23633 10088 24550
rect 10046 23624 10102 23633
rect 10046 23559 10102 23568
rect 10048 22772 10100 22778
rect 10048 22714 10100 22720
rect 9956 22432 10008 22438
rect 9956 22374 10008 22380
rect 9968 22098 9996 22374
rect 9956 22092 10008 22098
rect 9956 22034 10008 22040
rect 9968 21350 9996 22034
rect 10060 21894 10088 22714
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 10060 21418 10088 21830
rect 10048 21412 10100 21418
rect 10048 21354 10100 21360
rect 9956 21344 10008 21350
rect 10152 21298 10180 27520
rect 10796 26246 10824 27520
rect 11152 26308 11204 26314
rect 11152 26250 11204 26256
rect 10784 26240 10836 26246
rect 10784 26182 10836 26188
rect 10874 26208 10930 26217
rect 10874 26143 10930 26152
rect 10692 25696 10744 25702
rect 10692 25638 10744 25644
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10704 25498 10732 25638
rect 10888 25514 10916 26143
rect 10692 25492 10744 25498
rect 10692 25434 10744 25440
rect 10796 25486 10916 25514
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10232 24268 10284 24274
rect 10232 24210 10284 24216
rect 10244 23866 10272 24210
rect 10414 24168 10470 24177
rect 10796 24154 10824 25486
rect 10876 25356 10928 25362
rect 10876 25298 10928 25304
rect 10888 24614 10916 25298
rect 10876 24608 10928 24614
rect 10876 24550 10928 24556
rect 10414 24103 10416 24112
rect 10468 24103 10470 24112
rect 10704 24126 10824 24154
rect 10416 24074 10468 24080
rect 10704 23866 10732 24126
rect 10784 24064 10836 24070
rect 10784 24006 10836 24012
rect 10232 23860 10284 23866
rect 10232 23802 10284 23808
rect 10692 23860 10744 23866
rect 10692 23802 10744 23808
rect 10244 23769 10272 23802
rect 10230 23760 10286 23769
rect 10230 23695 10286 23704
rect 10796 23662 10824 24006
rect 10784 23656 10836 23662
rect 10784 23598 10836 23604
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10692 23180 10744 23186
rect 10692 23122 10744 23128
rect 10600 23112 10652 23118
rect 10600 23054 10652 23060
rect 10612 22778 10640 23054
rect 10600 22772 10652 22778
rect 10600 22714 10652 22720
rect 10704 22438 10732 23122
rect 10692 22432 10744 22438
rect 10692 22374 10744 22380
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10704 22166 10732 22374
rect 10692 22160 10744 22166
rect 10692 22102 10744 22108
rect 10690 21992 10746 22001
rect 10690 21927 10746 21936
rect 10704 21690 10732 21927
rect 10692 21684 10744 21690
rect 10692 21626 10744 21632
rect 10692 21480 10744 21486
rect 10692 21422 10744 21428
rect 9956 21286 10008 21292
rect 10060 21270 10180 21298
rect 9864 21004 9916 21010
rect 9864 20946 9916 20952
rect 9876 20058 9904 20946
rect 9956 20868 10008 20874
rect 9956 20810 10008 20816
rect 9864 20052 9916 20058
rect 9864 19994 9916 20000
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 9876 19145 9904 19790
rect 9862 19136 9918 19145
rect 9862 19071 9918 19080
rect 9862 19000 9918 19009
rect 9862 18935 9918 18944
rect 9876 18902 9904 18935
rect 9864 18896 9916 18902
rect 9864 18838 9916 18844
rect 9968 18834 9996 20810
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 9784 18686 9996 18714
rect 9864 18624 9916 18630
rect 9864 18566 9916 18572
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9600 17870 9720 17898
rect 9600 17626 9628 17870
rect 9680 17808 9732 17814
rect 9678 17776 9680 17785
rect 9732 17776 9734 17785
rect 9678 17711 9734 17720
rect 9784 17649 9812 18022
rect 9770 17640 9826 17649
rect 9600 17598 9720 17626
rect 9588 17128 9640 17134
rect 9588 17070 9640 17076
rect 9600 16590 9628 17070
rect 9588 16584 9640 16590
rect 9588 16526 9640 16532
rect 9692 16266 9720 17598
rect 9770 17575 9826 17584
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9600 16238 9720 16266
rect 9600 15586 9628 16238
rect 9678 16144 9734 16153
rect 9678 16079 9734 16088
rect 9692 15706 9720 16079
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9600 15558 9720 15586
rect 9588 14272 9640 14278
rect 9588 14214 9640 14220
rect 9600 13462 9628 14214
rect 9692 14090 9720 15558
rect 9784 14521 9812 17478
rect 9770 14512 9826 14521
rect 9770 14447 9826 14456
rect 9692 14062 9812 14090
rect 9680 13796 9732 13802
rect 9680 13738 9732 13744
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9692 13394 9720 13738
rect 9784 13705 9812 14062
rect 9770 13696 9826 13705
rect 9770 13631 9826 13640
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9496 13184 9548 13190
rect 9784 13138 9812 13466
rect 9496 13126 9548 13132
rect 9402 13016 9458 13025
rect 9402 12951 9458 12960
rect 9416 12782 9444 12951
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9310 12336 9366 12345
rect 9310 12271 9366 12280
rect 9508 12186 9536 13126
rect 9600 13110 9812 13138
rect 9600 12374 9628 13110
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9692 12442 9720 12718
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9588 12368 9640 12374
rect 9588 12310 9640 12316
rect 9324 12158 9536 12186
rect 9680 12164 9732 12170
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 9128 8832 9180 8838
rect 9324 8809 9352 12158
rect 9680 12106 9732 12112
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9416 11354 9444 12038
rect 9692 11744 9720 12106
rect 9600 11716 9720 11744
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9508 11121 9536 11494
rect 9494 11112 9550 11121
rect 9494 11047 9550 11056
rect 9508 10606 9536 11047
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9508 10130 9536 10542
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9600 9602 9628 11716
rect 9678 11656 9734 11665
rect 9678 11591 9734 11600
rect 9692 11354 9720 11591
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9692 10266 9720 11154
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9692 9761 9720 9862
rect 9678 9752 9734 9761
rect 9678 9687 9734 9696
rect 9600 9574 9720 9602
rect 9404 9104 9456 9110
rect 9404 9046 9456 9052
rect 9416 8974 9444 9046
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9128 8774 9180 8780
rect 9310 8800 9366 8809
rect 9140 8090 9168 8774
rect 9310 8735 9366 8744
rect 9220 8356 9272 8362
rect 9220 8298 9272 8304
rect 9232 8129 9260 8298
rect 9218 8120 9274 8129
rect 9128 8084 9180 8090
rect 9218 8055 9274 8064
rect 9128 8026 9180 8032
rect 9140 7818 9168 8026
rect 9218 7848 9274 7857
rect 9128 7812 9180 7818
rect 9218 7783 9274 7792
rect 9128 7754 9180 7760
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 8956 4814 9076 4842
rect 9140 4826 9168 4966
rect 9128 4820 9180 4826
rect 8852 4208 8904 4214
rect 8852 4150 8904 4156
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8404 2990 8432 3674
rect 8024 2984 8076 2990
rect 8022 2952 8024 2961
rect 8392 2984 8444 2990
rect 8076 2952 8078 2961
rect 7932 2916 7984 2922
rect 8392 2926 8444 2932
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 8022 2887 8078 2896
rect 7932 2858 7984 2864
rect 8404 2582 8432 2926
rect 8392 2576 8444 2582
rect 8772 2553 8800 2926
rect 8850 2816 8906 2825
rect 8850 2751 8906 2760
rect 8864 2650 8892 2751
rect 8852 2644 8904 2650
rect 8852 2586 8904 2592
rect 8392 2518 8444 2524
rect 8758 2544 8814 2553
rect 8758 2479 8814 2488
rect 8404 598 8524 626
rect 8404 480 8432 598
rect 7562 232 7618 241
rect 7562 167 7618 176
rect 7838 0 7894 480
rect 8390 0 8446 480
rect 8496 105 8524 598
rect 8956 480 8984 4814
rect 9128 4762 9180 4768
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9140 1057 9168 3674
rect 9232 3233 9260 7783
rect 9218 3224 9274 3233
rect 9218 3159 9274 3168
rect 9126 1048 9182 1057
rect 9126 983 9182 992
rect 8482 96 8538 105
rect 8482 31 8538 40
rect 8942 0 8998 480
rect 9324 105 9352 8735
rect 9416 8634 9444 8910
rect 9586 8664 9642 8673
rect 9404 8628 9456 8634
rect 9586 8599 9642 8608
rect 9404 8570 9456 8576
rect 9600 8022 9628 8599
rect 9588 8016 9640 8022
rect 9588 7958 9640 7964
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9404 4208 9456 4214
rect 9404 4150 9456 4156
rect 9416 4010 9444 4150
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 9416 3534 9444 3946
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9416 2650 9444 3470
rect 9404 2644 9456 2650
rect 9404 2586 9456 2592
rect 9508 480 9536 7890
rect 9600 7546 9628 7958
rect 9692 7857 9720 9574
rect 9784 9178 9812 12922
rect 9876 12714 9904 18566
rect 9968 16794 9996 18686
rect 10060 17338 10088 21270
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10140 21140 10192 21146
rect 10140 21082 10192 21088
rect 10048 17332 10100 17338
rect 10048 17274 10100 17280
rect 10152 17218 10180 21082
rect 10600 21072 10652 21078
rect 10600 21014 10652 21020
rect 10612 20913 10640 21014
rect 10704 21010 10732 21422
rect 10692 21004 10744 21010
rect 10692 20946 10744 20952
rect 10598 20904 10654 20913
rect 10598 20839 10654 20848
rect 10324 20800 10376 20806
rect 10324 20742 10376 20748
rect 10336 20398 10364 20742
rect 10324 20392 10376 20398
rect 10324 20334 10376 20340
rect 10612 20346 10640 20839
rect 10692 20800 10744 20806
rect 10692 20742 10744 20748
rect 10704 20466 10732 20742
rect 10796 20505 10824 23598
rect 10782 20496 10838 20505
rect 10692 20460 10744 20466
rect 10782 20431 10838 20440
rect 10692 20402 10744 20408
rect 10784 20392 10836 20398
rect 10612 20318 10732 20346
rect 10784 20334 10836 20340
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10232 19304 10284 19310
rect 10230 19272 10232 19281
rect 10284 19272 10286 19281
rect 10230 19207 10286 19216
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 10336 18630 10364 18770
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10336 18465 10364 18566
rect 10322 18456 10378 18465
rect 10322 18391 10378 18400
rect 10704 18154 10732 20318
rect 10796 19514 10824 20334
rect 10784 19508 10836 19514
rect 10784 19450 10836 19456
rect 10784 19304 10836 19310
rect 10784 19246 10836 19252
rect 10796 18714 10824 19246
rect 10888 18834 10916 24550
rect 11164 23254 11192 26250
rect 11244 24608 11296 24614
rect 11244 24550 11296 24556
rect 11256 24290 11284 24550
rect 11348 24426 11376 27520
rect 11794 26344 11850 26353
rect 11794 26279 11850 26288
rect 11808 25974 11836 26279
rect 11900 26110 11928 27520
rect 12348 26240 12400 26246
rect 12348 26182 12400 26188
rect 11888 26104 11940 26110
rect 11888 26046 11940 26052
rect 11796 25968 11848 25974
rect 11796 25910 11848 25916
rect 11888 25968 11940 25974
rect 11888 25910 11940 25916
rect 11518 25664 11574 25673
rect 11518 25599 11574 25608
rect 11426 24712 11482 24721
rect 11426 24647 11482 24656
rect 11440 24614 11468 24647
rect 11428 24608 11480 24614
rect 11428 24550 11480 24556
rect 11348 24398 11468 24426
rect 11532 24410 11560 25599
rect 11612 25356 11664 25362
rect 11612 25298 11664 25304
rect 11624 24614 11652 25298
rect 11612 24608 11664 24614
rect 11612 24550 11664 24556
rect 11256 24262 11376 24290
rect 11152 23248 11204 23254
rect 11152 23190 11204 23196
rect 10968 22976 11020 22982
rect 10968 22918 11020 22924
rect 10980 22574 11008 22918
rect 10968 22568 11020 22574
rect 11020 22516 11192 22522
rect 10968 22510 11192 22516
rect 10980 22494 11192 22510
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 11072 21350 11100 22374
rect 11164 21962 11192 22494
rect 11242 22400 11298 22409
rect 11242 22335 11298 22344
rect 11152 21956 11204 21962
rect 11152 21898 11204 21904
rect 11256 21434 11284 22335
rect 11164 21406 11284 21434
rect 11060 21344 11112 21350
rect 11060 21286 11112 21292
rect 11072 20058 11100 21286
rect 11164 21146 11192 21406
rect 11244 21344 11296 21350
rect 11244 21286 11296 21292
rect 11152 21140 11204 21146
rect 11152 21082 11204 21088
rect 11256 21078 11284 21286
rect 11244 21072 11296 21078
rect 11244 21014 11296 21020
rect 11256 20262 11284 21014
rect 11244 20256 11296 20262
rect 11244 20198 11296 20204
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 11152 19984 11204 19990
rect 11152 19926 11204 19932
rect 10966 19816 11022 19825
rect 10966 19751 11022 19760
rect 10980 19310 11008 19751
rect 11058 19680 11114 19689
rect 11058 19615 11114 19624
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 10968 19168 11020 19174
rect 10968 19110 11020 19116
rect 10980 19009 11008 19110
rect 10966 19000 11022 19009
rect 11072 18970 11100 19615
rect 11164 19378 11192 19926
rect 11256 19854 11284 20198
rect 11348 20097 11376 24262
rect 11334 20088 11390 20097
rect 11334 20023 11390 20032
rect 11334 19952 11390 19961
rect 11334 19887 11390 19896
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11256 19718 11284 19790
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 11256 19378 11284 19654
rect 11152 19372 11204 19378
rect 11152 19314 11204 19320
rect 11244 19372 11296 19378
rect 11244 19314 11296 19320
rect 11242 19272 11298 19281
rect 11242 19207 11244 19216
rect 11296 19207 11298 19216
rect 11244 19178 11296 19184
rect 11242 19136 11298 19145
rect 11242 19071 11298 19080
rect 10966 18935 11022 18944
rect 11060 18964 11112 18970
rect 11060 18906 11112 18912
rect 10876 18828 10928 18834
rect 10876 18770 10928 18776
rect 11152 18760 11204 18766
rect 10966 18728 11022 18737
rect 10796 18686 10916 18714
rect 10692 18148 10744 18154
rect 10692 18090 10744 18096
rect 10784 18148 10836 18154
rect 10784 18090 10836 18096
rect 10796 18034 10824 18090
rect 10704 18006 10824 18034
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10060 17190 10180 17218
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 9968 15978 9996 16594
rect 9956 15972 10008 15978
rect 9956 15914 10008 15920
rect 9954 15328 10010 15337
rect 9954 15263 10010 15272
rect 9968 15162 9996 15263
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9956 14340 10008 14346
rect 9956 14282 10008 14288
rect 9968 13870 9996 14282
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 9968 13258 9996 13806
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 9864 12708 9916 12714
rect 9864 12650 9916 12656
rect 9862 12608 9918 12617
rect 9862 12543 9918 12552
rect 9876 12442 9904 12543
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9876 11898 9904 12378
rect 9968 12238 9996 13194
rect 10060 13002 10088 17190
rect 10140 17060 10192 17066
rect 10140 17002 10192 17008
rect 10152 16794 10180 17002
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 10152 16250 10180 16730
rect 10232 16720 10284 16726
rect 10232 16662 10284 16668
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10244 15994 10272 16662
rect 10506 16280 10562 16289
rect 10506 16215 10508 16224
rect 10560 16215 10562 16224
rect 10508 16186 10560 16192
rect 10152 15966 10272 15994
rect 10152 14618 10180 15966
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10416 15632 10468 15638
rect 10416 15574 10468 15580
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 10336 15026 10364 15302
rect 10428 15065 10456 15574
rect 10704 15450 10732 18006
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 10796 15586 10824 17274
rect 10888 16096 10916 18686
rect 11152 18702 11204 18708
rect 10966 18663 11022 18672
rect 10980 18630 11008 18663
rect 10968 18624 11020 18630
rect 10968 18566 11020 18572
rect 11060 18148 11112 18154
rect 11060 18090 11112 18096
rect 10968 18080 11020 18086
rect 11072 18057 11100 18090
rect 10968 18022 11020 18028
rect 11058 18048 11114 18057
rect 10980 17814 11008 18022
rect 11058 17983 11114 17992
rect 11058 17912 11114 17921
rect 11058 17847 11114 17856
rect 10968 17808 11020 17814
rect 10968 17750 11020 17756
rect 11072 17746 11100 17847
rect 11060 17740 11112 17746
rect 11060 17682 11112 17688
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 10980 17270 11008 17614
rect 10968 17264 11020 17270
rect 10968 17206 11020 17212
rect 11072 17202 11100 17682
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 10888 16068 11100 16096
rect 10966 16008 11022 16017
rect 10966 15943 11022 15952
rect 10876 15904 10928 15910
rect 10874 15872 10876 15881
rect 10928 15872 10930 15881
rect 10874 15807 10930 15816
rect 10796 15558 10916 15586
rect 10704 15422 10824 15450
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10414 15056 10470 15065
rect 10324 15020 10376 15026
rect 10414 14991 10470 15000
rect 10324 14962 10376 14968
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 10152 14074 10180 14554
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 10138 13696 10194 13705
rect 10138 13631 10194 13640
rect 10152 13138 10180 13631
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 10152 13110 10272 13138
rect 10060 12986 10180 13002
rect 10060 12980 10192 12986
rect 10060 12974 10140 12980
rect 10140 12922 10192 12928
rect 10048 12912 10100 12918
rect 10244 12866 10272 13110
rect 10048 12854 10100 12860
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9968 12102 9996 12174
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9956 11824 10008 11830
rect 9956 11766 10008 11772
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9770 8392 9826 8401
rect 9770 8327 9772 8336
rect 9824 8327 9826 8336
rect 9772 8298 9824 8304
rect 9876 8072 9904 11698
rect 9784 8044 9904 8072
rect 9678 7848 9734 7857
rect 9678 7783 9734 7792
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9692 6458 9720 6938
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 9784 6202 9812 8044
rect 9864 7948 9916 7954
rect 9864 7890 9916 7896
rect 9876 7857 9904 7890
rect 9862 7848 9918 7857
rect 9862 7783 9918 7792
rect 9876 7546 9904 7783
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9876 7177 9904 7482
rect 9862 7168 9918 7177
rect 9862 7103 9918 7112
rect 9968 6644 9996 11766
rect 10060 10266 10088 12854
rect 10152 12838 10272 12866
rect 10336 12850 10364 13330
rect 10704 12850 10732 15302
rect 10796 13870 10824 15422
rect 10888 15337 10916 15558
rect 10874 15328 10930 15337
rect 10874 15263 10930 15272
rect 10980 14890 11008 15943
rect 11072 15638 11100 16068
rect 11060 15632 11112 15638
rect 11060 15574 11112 15580
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 11072 14958 11100 15438
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 10968 14884 11020 14890
rect 10968 14826 11020 14832
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 10968 14544 11020 14550
rect 10968 14486 11020 14492
rect 11072 14498 11100 14758
rect 11164 14618 11192 18702
rect 11256 18222 11284 19071
rect 11244 18216 11296 18222
rect 11244 18158 11296 18164
rect 11256 17338 11284 18158
rect 11348 17814 11376 19887
rect 11336 17808 11388 17814
rect 11336 17750 11388 17756
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 11244 17332 11296 17338
rect 11244 17274 11296 17280
rect 11348 16794 11376 17614
rect 11336 16788 11388 16794
rect 11336 16730 11388 16736
rect 11242 16552 11298 16561
rect 11242 16487 11298 16496
rect 11336 16516 11388 16522
rect 11256 15570 11284 16487
rect 11336 16458 11388 16464
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11348 15416 11376 16458
rect 11440 16017 11468 24398
rect 11520 24404 11572 24410
rect 11520 24346 11572 24352
rect 11612 24268 11664 24274
rect 11612 24210 11664 24216
rect 11624 23526 11652 24210
rect 11704 24132 11756 24138
rect 11704 24074 11756 24080
rect 11796 24132 11848 24138
rect 11796 24074 11848 24080
rect 11716 23730 11744 24074
rect 11704 23724 11756 23730
rect 11704 23666 11756 23672
rect 11612 23520 11664 23526
rect 11612 23462 11664 23468
rect 11624 22953 11652 23462
rect 11610 22944 11666 22953
rect 11610 22879 11666 22888
rect 11612 22772 11664 22778
rect 11612 22714 11664 22720
rect 11518 22536 11574 22545
rect 11518 22471 11574 22480
rect 11532 22166 11560 22471
rect 11520 22160 11572 22166
rect 11520 22102 11572 22108
rect 11518 20768 11574 20777
rect 11518 20703 11574 20712
rect 11532 20058 11560 20703
rect 11520 20052 11572 20058
rect 11520 19994 11572 20000
rect 11532 19961 11560 19994
rect 11518 19952 11574 19961
rect 11518 19887 11574 19896
rect 11624 19904 11652 22714
rect 11716 20505 11744 23666
rect 11808 23050 11836 24074
rect 11900 23322 11928 25910
rect 12164 25900 12216 25906
rect 12164 25842 12216 25848
rect 12176 25242 12204 25842
rect 12360 25650 12388 26182
rect 12268 25622 12388 25650
rect 12268 25498 12296 25622
rect 12256 25492 12308 25498
rect 12256 25434 12308 25440
rect 12348 25492 12400 25498
rect 12348 25434 12400 25440
rect 12360 25242 12388 25434
rect 12176 25214 12388 25242
rect 12256 24608 12308 24614
rect 12256 24550 12308 24556
rect 11980 23588 12032 23594
rect 11980 23530 12032 23536
rect 11888 23316 11940 23322
rect 11888 23258 11940 23264
rect 11888 23180 11940 23186
rect 11888 23122 11940 23128
rect 11796 23044 11848 23050
rect 11796 22986 11848 22992
rect 11808 22098 11836 22986
rect 11900 22438 11928 23122
rect 11888 22432 11940 22438
rect 11888 22374 11940 22380
rect 11900 22137 11928 22374
rect 11886 22128 11942 22137
rect 11796 22092 11848 22098
rect 11886 22063 11942 22072
rect 11796 22034 11848 22040
rect 11702 20496 11758 20505
rect 11702 20431 11758 20440
rect 11704 19916 11756 19922
rect 11532 19514 11560 19887
rect 11624 19876 11704 19904
rect 11704 19858 11756 19864
rect 11610 19816 11666 19825
rect 11610 19751 11666 19760
rect 11520 19508 11572 19514
rect 11520 19450 11572 19456
rect 11624 19394 11652 19751
rect 11532 19366 11652 19394
rect 11532 18902 11560 19366
rect 11808 19281 11836 22034
rect 11886 20224 11942 20233
rect 11886 20159 11942 20168
rect 11900 19825 11928 20159
rect 11886 19816 11942 19825
rect 11886 19751 11942 19760
rect 11992 19292 12020 23530
rect 12072 23112 12124 23118
rect 12072 23054 12124 23060
rect 12084 22778 12112 23054
rect 12072 22772 12124 22778
rect 12072 22714 12124 22720
rect 12072 21956 12124 21962
rect 12072 21898 12124 21904
rect 12084 19378 12112 21898
rect 12268 20097 12296 24550
rect 12348 24268 12400 24274
rect 12348 24210 12400 24216
rect 12360 23526 12388 24210
rect 12348 23520 12400 23526
rect 12346 23488 12348 23497
rect 12400 23488 12402 23497
rect 12346 23423 12402 23432
rect 12440 22568 12492 22574
rect 12346 22536 12402 22545
rect 12544 22545 12572 27520
rect 12716 25356 12768 25362
rect 12716 25298 12768 25304
rect 12440 22510 12492 22516
rect 12530 22536 12586 22545
rect 12346 22471 12402 22480
rect 12360 22030 12388 22471
rect 12348 22024 12400 22030
rect 12348 21966 12400 21972
rect 12360 21554 12388 21966
rect 12348 21548 12400 21554
rect 12348 21490 12400 21496
rect 12360 20641 12388 21490
rect 12346 20632 12402 20641
rect 12346 20567 12402 20576
rect 12452 20448 12480 22510
rect 12530 22471 12586 22480
rect 12728 22420 12756 25298
rect 12898 24984 12954 24993
rect 12898 24919 12954 24928
rect 12912 24449 12940 24919
rect 12992 24608 13044 24614
rect 12992 24550 13044 24556
rect 12898 24440 12954 24449
rect 12898 24375 12954 24384
rect 12808 24064 12860 24070
rect 12808 24006 12860 24012
rect 12820 23526 12848 24006
rect 12808 23520 12860 23526
rect 13004 23497 13032 24550
rect 12808 23462 12860 23468
rect 12990 23488 13046 23497
rect 12990 23423 13046 23432
rect 12900 22976 12952 22982
rect 12900 22918 12952 22924
rect 12912 22642 12940 22918
rect 12900 22636 12952 22642
rect 12900 22578 12952 22584
rect 12360 20420 12480 20448
rect 12544 22392 12756 22420
rect 12254 20088 12310 20097
rect 12360 20074 12388 20420
rect 12438 20360 12494 20369
rect 12438 20295 12494 20304
rect 12452 20262 12480 20295
rect 12440 20256 12492 20262
rect 12440 20198 12492 20204
rect 12360 20046 12480 20074
rect 12254 20023 12310 20032
rect 12348 19984 12400 19990
rect 12348 19926 12400 19932
rect 12256 19780 12308 19786
rect 12256 19722 12308 19728
rect 12268 19446 12296 19722
rect 12256 19440 12308 19446
rect 12256 19382 12308 19388
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 11794 19272 11850 19281
rect 11704 19236 11756 19242
rect 11794 19207 11850 19216
rect 11900 19264 12020 19292
rect 11704 19178 11756 19184
rect 11520 18896 11572 18902
rect 11520 18838 11572 18844
rect 11716 18766 11744 19178
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 11808 18902 11836 19110
rect 11900 18986 11928 19264
rect 12072 19236 12124 19242
rect 12072 19178 12124 19184
rect 11980 19168 12032 19174
rect 11978 19136 11980 19145
rect 12032 19136 12034 19145
rect 11978 19071 12034 19080
rect 11900 18958 12020 18986
rect 11796 18896 11848 18902
rect 11796 18838 11848 18844
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 11704 18760 11756 18766
rect 11888 18760 11940 18766
rect 11704 18702 11756 18708
rect 11794 18728 11850 18737
rect 11532 18222 11560 18702
rect 11612 18624 11664 18630
rect 11612 18566 11664 18572
rect 11520 18216 11572 18222
rect 11520 18158 11572 18164
rect 11426 16008 11482 16017
rect 11426 15943 11482 15952
rect 11426 15736 11482 15745
rect 11426 15671 11482 15680
rect 11440 15502 11468 15671
rect 11428 15496 11480 15502
rect 11428 15438 11480 15444
rect 11256 15388 11376 15416
rect 11256 15094 11284 15388
rect 11428 15360 11480 15366
rect 11334 15328 11390 15337
rect 11428 15302 11480 15308
rect 11334 15263 11390 15272
rect 11244 15088 11296 15094
rect 11244 15030 11296 15036
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 11256 14521 11284 14894
rect 11242 14512 11298 14521
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10888 13938 10916 14214
rect 10980 14113 11008 14486
rect 11072 14470 11192 14498
rect 11058 14376 11114 14385
rect 11058 14311 11114 14320
rect 10966 14104 11022 14113
rect 10966 14039 11022 14048
rect 10968 14000 11020 14006
rect 10968 13942 11020 13948
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10876 13796 10928 13802
rect 10876 13738 10928 13744
rect 10888 13705 10916 13738
rect 10874 13696 10930 13705
rect 10874 13631 10930 13640
rect 10782 13560 10838 13569
rect 10782 13495 10784 13504
rect 10836 13495 10838 13504
rect 10784 13466 10836 13472
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 10888 13025 10916 13194
rect 10874 13016 10930 13025
rect 10874 12951 10930 12960
rect 10782 12880 10838 12889
rect 10152 12170 10180 12838
rect 10244 12714 10272 12838
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 10692 12844 10744 12850
rect 10782 12815 10838 12824
rect 10692 12786 10744 12792
rect 10232 12708 10284 12714
rect 10232 12650 10284 12656
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10704 12345 10732 12786
rect 10796 12442 10824 12815
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 10414 12336 10470 12345
rect 10324 12300 10376 12306
rect 10414 12271 10470 12280
rect 10690 12336 10746 12345
rect 10888 12322 10916 12582
rect 10690 12271 10746 12280
rect 10796 12294 10916 12322
rect 10324 12242 10376 12248
rect 10140 12164 10192 12170
rect 10140 12106 10192 12112
rect 10230 12064 10286 12073
rect 10230 11999 10286 12008
rect 10244 11898 10272 11999
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10138 11792 10194 11801
rect 10138 11727 10194 11736
rect 10152 11558 10180 11727
rect 10336 11626 10364 12242
rect 10428 12073 10456 12271
rect 10796 12238 10824 12294
rect 10980 12238 11008 13942
rect 11072 12458 11100 14311
rect 11164 14006 11192 14470
rect 11242 14447 11298 14456
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11152 14000 11204 14006
rect 11256 13977 11284 14214
rect 11152 13942 11204 13948
rect 11242 13968 11298 13977
rect 11164 13274 11192 13942
rect 11242 13903 11298 13912
rect 11348 13802 11376 15263
rect 11440 14414 11468 15302
rect 11428 14408 11480 14414
rect 11428 14350 11480 14356
rect 11440 13841 11468 14350
rect 11426 13832 11482 13841
rect 11336 13796 11388 13802
rect 11426 13767 11482 13776
rect 11336 13738 11388 13744
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 11256 13394 11284 13670
rect 11348 13530 11376 13738
rect 11532 13716 11560 18158
rect 11624 16114 11652 18566
rect 11716 18086 11744 18702
rect 11888 18702 11940 18708
rect 11794 18663 11850 18672
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11702 17912 11758 17921
rect 11702 17847 11758 17856
rect 11716 17513 11744 17847
rect 11702 17504 11758 17513
rect 11702 17439 11758 17448
rect 11808 16538 11836 18663
rect 11900 17814 11928 18702
rect 11888 17808 11940 17814
rect 11888 17750 11940 17756
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 11716 16510 11836 16538
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 11612 15564 11664 15570
rect 11612 15506 11664 15512
rect 11624 15201 11652 15506
rect 11610 15192 11666 15201
rect 11610 15127 11612 15136
rect 11664 15127 11666 15136
rect 11612 15098 11664 15104
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11440 13688 11560 13716
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 11244 13388 11296 13394
rect 11244 13330 11296 13336
rect 11164 13246 11376 13274
rect 11244 13184 11296 13190
rect 11244 13126 11296 13132
rect 11256 12850 11284 13126
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 11152 12708 11204 12714
rect 11152 12650 11204 12656
rect 11164 12617 11192 12650
rect 11150 12608 11206 12617
rect 11150 12543 11206 12552
rect 11072 12430 11192 12458
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10414 12064 10470 12073
rect 10414 11999 10470 12008
rect 10520 11762 10548 12174
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10612 11676 10640 11834
rect 10704 11830 10732 12038
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 10612 11648 10732 11676
rect 10324 11620 10376 11626
rect 10324 11562 10376 11568
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 10152 11354 10180 11494
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10600 11212 10652 11218
rect 10600 11154 10652 11160
rect 10324 11076 10376 11082
rect 10324 11018 10376 11024
rect 10336 10810 10364 11018
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10612 10713 10640 11154
rect 10598 10704 10654 10713
rect 10598 10639 10600 10648
rect 10652 10639 10654 10648
rect 10600 10610 10652 10616
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 10060 9722 10088 10202
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 10152 9654 10180 10202
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 10244 9518 10272 9998
rect 10232 9512 10284 9518
rect 10232 9454 10284 9460
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10152 8090 10180 8570
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10046 7712 10102 7721
rect 10046 7647 10102 7656
rect 10060 7478 10088 7647
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 10060 7002 10088 7414
rect 10704 7342 10732 11648
rect 10796 10266 10824 12038
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10796 9217 10824 9318
rect 10782 9208 10838 9217
rect 10782 9143 10838 9152
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10796 8090 10824 8230
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10888 8004 10916 11494
rect 10980 11082 11008 11698
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 10968 10260 11020 10266
rect 11072 10248 11100 11018
rect 11164 10606 11192 12430
rect 11348 12322 11376 13246
rect 11256 12294 11376 12322
rect 11256 11898 11284 12294
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11348 11937 11376 12174
rect 11334 11928 11390 11937
rect 11244 11892 11296 11898
rect 11334 11863 11390 11872
rect 11244 11834 11296 11840
rect 11242 11656 11298 11665
rect 11242 11591 11298 11600
rect 11256 11558 11284 11591
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11348 11370 11376 11494
rect 11256 11342 11376 11370
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 11020 10220 11100 10248
rect 10968 10202 11020 10208
rect 10966 9752 11022 9761
rect 10966 9687 11022 9696
rect 10980 8838 11008 9687
rect 11072 9586 11100 10220
rect 11164 9722 11192 10406
rect 11256 9897 11284 11342
rect 11440 11234 11468 13688
rect 11520 13456 11572 13462
rect 11624 13433 11652 14418
rect 11716 13462 11744 16510
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11808 16250 11836 16390
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 11796 16108 11848 16114
rect 11796 16050 11848 16056
rect 11704 13456 11756 13462
rect 11520 13398 11572 13404
rect 11610 13424 11666 13433
rect 11532 12646 11560 13398
rect 11704 13398 11756 13404
rect 11610 13359 11666 13368
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11532 12209 11560 12242
rect 11518 12200 11574 12209
rect 11518 12135 11574 12144
rect 11532 11354 11560 12135
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11440 11206 11560 11234
rect 11428 11008 11480 11014
rect 11428 10950 11480 10956
rect 11440 10674 11468 10950
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 11336 10464 11388 10470
rect 11334 10432 11336 10441
rect 11388 10432 11390 10441
rect 11334 10367 11390 10376
rect 11440 9926 11468 10610
rect 11428 9920 11480 9926
rect 11242 9888 11298 9897
rect 11428 9862 11480 9868
rect 11242 9823 11298 9832
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 11242 9616 11298 9625
rect 11060 9580 11112 9586
rect 11242 9551 11298 9560
rect 11060 9522 11112 9528
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 11058 9344 11114 9353
rect 11058 9279 11114 9288
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10888 7976 11008 8004
rect 10784 7948 10836 7954
rect 10836 7908 10916 7936
rect 10784 7890 10836 7896
rect 10782 7712 10838 7721
rect 10782 7647 10838 7656
rect 10796 7546 10824 7647
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 10704 6866 10732 7278
rect 10888 7002 10916 7908
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10140 6792 10192 6798
rect 10138 6760 10140 6769
rect 10192 6760 10194 6769
rect 10138 6695 10194 6704
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 9968 6616 10180 6644
rect 9692 5778 9720 6190
rect 9784 6174 9996 6202
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9772 5840 9824 5846
rect 9772 5782 9824 5788
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9600 4706 9628 5714
rect 9692 5234 9720 5714
rect 9784 5234 9812 5782
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9680 5092 9732 5098
rect 9680 5034 9732 5040
rect 9692 4826 9720 5034
rect 9784 5030 9812 5170
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9600 4678 9720 4706
rect 9586 4176 9642 4185
rect 9586 4111 9642 4120
rect 9600 3670 9628 4111
rect 9588 3664 9640 3670
rect 9588 3606 9640 3612
rect 9692 3466 9720 4678
rect 9876 4282 9904 6054
rect 9968 5137 9996 6174
rect 10046 5944 10102 5953
rect 10046 5879 10102 5888
rect 10060 5166 10088 5879
rect 10048 5160 10100 5166
rect 9954 5128 10010 5137
rect 10048 5102 10100 5108
rect 9954 5063 10010 5072
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 9968 4078 9996 4966
rect 10060 4826 10088 5102
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 10048 3936 10100 3942
rect 10046 3904 10048 3913
rect 10100 3904 10102 3913
rect 10046 3839 10102 3848
rect 9862 3768 9918 3777
rect 9862 3703 9918 3712
rect 9876 3670 9904 3703
rect 9864 3664 9916 3670
rect 9864 3606 9916 3612
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9784 3126 9812 3538
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 9588 2916 9640 2922
rect 9588 2858 9640 2864
rect 9600 2650 9628 2858
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9784 2582 9812 3062
rect 9876 2689 9904 3130
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 9968 2825 9996 2926
rect 9954 2816 10010 2825
rect 9954 2751 10010 2760
rect 9862 2680 9918 2689
rect 9862 2615 9918 2624
rect 9772 2576 9824 2582
rect 9772 2518 9824 2524
rect 10060 480 10088 3402
rect 10152 1442 10180 6616
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10690 5672 10746 5681
rect 10690 5607 10746 5616
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10244 4010 10272 4558
rect 10704 4010 10732 5607
rect 10796 5574 10824 6666
rect 10888 6254 10916 6938
rect 10876 6248 10928 6254
rect 10876 6190 10928 6196
rect 10888 5846 10916 6190
rect 10876 5840 10928 5846
rect 10876 5782 10928 5788
rect 10784 5568 10836 5574
rect 10980 5556 11008 7976
rect 11072 7585 11100 9279
rect 11164 9178 11192 9386
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 11150 8664 11206 8673
rect 11150 8599 11206 8608
rect 11164 8430 11192 8599
rect 11256 8498 11284 9551
rect 11440 9110 11468 9862
rect 11428 9104 11480 9110
rect 11334 9072 11390 9081
rect 11428 9046 11480 9052
rect 11334 9007 11390 9016
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11152 8424 11204 8430
rect 11348 8378 11376 9007
rect 11428 8492 11480 8498
rect 11428 8434 11480 8440
rect 11152 8366 11204 8372
rect 11164 8294 11192 8366
rect 11256 8350 11376 8378
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11058 7576 11114 7585
rect 11058 7511 11114 7520
rect 11060 7472 11112 7478
rect 11058 7440 11060 7449
rect 11112 7440 11114 7449
rect 11058 7375 11114 7384
rect 11060 6180 11112 6186
rect 11060 6122 11112 6128
rect 11072 5914 11100 6122
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 10784 5510 10836 5516
rect 10888 5528 11008 5556
rect 10232 4004 10284 4010
rect 10232 3946 10284 3952
rect 10692 4004 10744 4010
rect 10692 3946 10744 3952
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10796 3398 10824 5510
rect 10888 3466 10916 5528
rect 11164 5386 11192 8230
rect 11256 5545 11284 8350
rect 11440 8022 11468 8434
rect 11428 8016 11480 8022
rect 11428 7958 11480 7964
rect 11440 7546 11468 7958
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11348 7002 11376 7278
rect 11336 6996 11388 7002
rect 11336 6938 11388 6944
rect 11532 6866 11560 11206
rect 11624 10044 11652 12718
rect 11716 12238 11744 12786
rect 11808 12628 11836 16050
rect 11900 15881 11928 16594
rect 11886 15872 11942 15881
rect 11886 15807 11942 15816
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11900 15162 11928 15438
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11900 14550 11928 15098
rect 11888 14544 11940 14550
rect 11888 14486 11940 14492
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 11900 14074 11928 14350
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11900 12753 11928 14010
rect 11992 12782 12020 18958
rect 12084 17082 12112 19178
rect 12162 18864 12218 18873
rect 12162 18799 12218 18808
rect 12176 18601 12204 18799
rect 12162 18592 12218 18601
rect 12162 18527 12218 18536
rect 12256 18352 12308 18358
rect 12360 18329 12388 19926
rect 12256 18294 12308 18300
rect 12346 18320 12402 18329
rect 12164 18080 12216 18086
rect 12164 18022 12216 18028
rect 12176 17921 12204 18022
rect 12162 17912 12218 17921
rect 12162 17847 12218 17856
rect 12268 17270 12296 18294
rect 12346 18255 12402 18264
rect 12452 18170 12480 20046
rect 12544 19514 12572 22392
rect 12716 22024 12768 22030
rect 12716 21966 12768 21972
rect 12808 22024 12860 22030
rect 12808 21966 12860 21972
rect 12728 21078 12756 21966
rect 12820 21690 12848 21966
rect 12808 21684 12860 21690
rect 12808 21626 12860 21632
rect 12716 21072 12768 21078
rect 12716 21014 12768 21020
rect 12728 20466 12756 21014
rect 12820 20777 12848 21626
rect 12806 20768 12862 20777
rect 12806 20703 12862 20712
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12808 20256 12860 20262
rect 12808 20198 12860 20204
rect 12820 20097 12848 20198
rect 12806 20088 12862 20097
rect 12806 20023 12808 20032
rect 12860 20023 12862 20032
rect 12808 19994 12860 20000
rect 12716 19916 12768 19922
rect 12716 19858 12768 19864
rect 12622 19816 12678 19825
rect 12622 19751 12678 19760
rect 12532 19508 12584 19514
rect 12532 19450 12584 19456
rect 12636 19417 12664 19751
rect 12622 19408 12678 19417
rect 12622 19343 12678 19352
rect 12728 19224 12756 19858
rect 12820 19553 12848 19994
rect 12806 19544 12862 19553
rect 12912 19514 12940 22578
rect 12992 21480 13044 21486
rect 12992 21422 13044 21428
rect 13004 19990 13032 21422
rect 12992 19984 13044 19990
rect 12992 19926 13044 19932
rect 13004 19854 13032 19926
rect 12992 19848 13044 19854
rect 12992 19790 13044 19796
rect 12806 19479 12862 19488
rect 12900 19508 12952 19514
rect 12900 19450 12952 19456
rect 12728 19196 12848 19224
rect 12624 19168 12676 19174
rect 12624 19110 12676 19116
rect 12714 19136 12770 19145
rect 12532 18760 12584 18766
rect 12530 18728 12532 18737
rect 12584 18728 12586 18737
rect 12530 18663 12586 18672
rect 12532 18624 12584 18630
rect 12636 18612 12664 19110
rect 12820 19122 12848 19196
rect 13004 19122 13032 19790
rect 12770 19094 12848 19122
rect 12912 19094 13032 19122
rect 12714 19071 12770 19080
rect 12808 18828 12860 18834
rect 12912 18816 12940 19094
rect 12990 19000 13046 19009
rect 12990 18935 13046 18944
rect 13004 18902 13032 18935
rect 12992 18896 13044 18902
rect 12992 18838 13044 18844
rect 12860 18788 12940 18816
rect 12808 18770 12860 18776
rect 12584 18584 12664 18612
rect 12714 18592 12770 18601
rect 12532 18566 12584 18572
rect 12360 18142 12480 18170
rect 12256 17264 12308 17270
rect 12256 17206 12308 17212
rect 12084 17054 12296 17082
rect 12072 16720 12124 16726
rect 12072 16662 12124 16668
rect 12084 16250 12112 16662
rect 12072 16244 12124 16250
rect 12072 16186 12124 16192
rect 12162 14920 12218 14929
rect 12162 14855 12218 14864
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 12084 14074 12112 14554
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 12072 13932 12124 13938
rect 12072 13874 12124 13880
rect 11980 12776 12032 12782
rect 11886 12744 11942 12753
rect 11980 12718 12032 12724
rect 11886 12679 11942 12688
rect 11980 12640 12032 12646
rect 11808 12600 11928 12628
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11702 11928 11758 11937
rect 11702 11863 11758 11872
rect 11716 11694 11744 11863
rect 11794 11792 11850 11801
rect 11794 11727 11850 11736
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 11808 11286 11836 11727
rect 11900 11540 11928 12600
rect 11980 12582 12032 12588
rect 11992 11665 12020 12582
rect 11978 11656 12034 11665
rect 11978 11591 12034 11600
rect 11900 11512 12020 11540
rect 11796 11280 11848 11286
rect 11796 11222 11848 11228
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11716 10198 11744 11154
rect 11808 10742 11836 11222
rect 11796 10736 11848 10742
rect 11796 10678 11848 10684
rect 11704 10192 11756 10198
rect 11702 10160 11704 10169
rect 11756 10160 11758 10169
rect 11702 10095 11758 10104
rect 11888 10056 11940 10062
rect 11624 10016 11744 10044
rect 11610 9888 11666 9897
rect 11610 9823 11666 9832
rect 11520 6860 11572 6866
rect 11520 6802 11572 6808
rect 11532 6497 11560 6802
rect 11518 6488 11574 6497
rect 11518 6423 11520 6432
rect 11572 6423 11574 6432
rect 11520 6394 11572 6400
rect 11336 6384 11388 6390
rect 11532 6363 11560 6394
rect 11336 6326 11388 6332
rect 11348 5914 11376 6326
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11428 5840 11480 5846
rect 11428 5782 11480 5788
rect 11242 5536 11298 5545
rect 11242 5471 11298 5480
rect 11164 5358 11284 5386
rect 11440 5370 11468 5782
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 10980 4570 11008 4626
rect 10980 4542 11100 4570
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 10980 3602 11008 3878
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10876 3460 10928 3466
rect 10876 3402 10928 3408
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10980 2854 11008 3538
rect 11072 3534 11100 4542
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 11072 2990 11100 3334
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 10612 2281 10640 2450
rect 10598 2272 10654 2281
rect 10598 2207 10654 2216
rect 10152 1414 10640 1442
rect 10612 480 10640 1414
rect 11164 480 11192 4082
rect 11256 2972 11284 5358
rect 11428 5364 11480 5370
rect 11428 5306 11480 5312
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11348 4185 11376 4966
rect 11440 4690 11468 5306
rect 11520 4752 11572 4758
rect 11520 4694 11572 4700
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11428 4548 11480 4554
rect 11428 4490 11480 4496
rect 11334 4176 11390 4185
rect 11334 4111 11390 4120
rect 11336 4004 11388 4010
rect 11336 3946 11388 3952
rect 11348 3670 11376 3946
rect 11336 3664 11388 3670
rect 11336 3606 11388 3612
rect 11348 3126 11376 3606
rect 11440 3602 11468 4490
rect 11532 4282 11560 4694
rect 11520 4276 11572 4282
rect 11520 4218 11572 4224
rect 11532 4026 11560 4218
rect 11624 4146 11652 9823
rect 11716 7936 11744 10016
rect 11888 9998 11940 10004
rect 11900 9761 11928 9998
rect 11886 9752 11942 9761
rect 11886 9687 11942 9696
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11808 9178 11836 9522
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11900 8906 11928 9687
rect 11888 8900 11940 8906
rect 11888 8842 11940 8848
rect 11992 8809 12020 11512
rect 12084 11150 12112 13874
rect 12072 11144 12124 11150
rect 12070 11112 12072 11121
rect 12124 11112 12126 11121
rect 12070 11047 12126 11056
rect 12084 11021 12112 11047
rect 12176 10962 12204 14855
rect 12268 13716 12296 17054
rect 12360 16266 12388 18142
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12452 16454 12480 18022
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12544 16289 12572 18566
rect 12714 18527 12770 18536
rect 12622 17640 12678 17649
rect 12622 17575 12678 17584
rect 12530 16280 12586 16289
rect 12360 16238 12480 16266
rect 12348 14068 12400 14074
rect 12348 14010 12400 14016
rect 12360 13841 12388 14010
rect 12346 13832 12402 13841
rect 12346 13767 12402 13776
rect 12268 13688 12388 13716
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12268 12442 12296 13466
rect 12256 12436 12308 12442
rect 12256 12378 12308 12384
rect 12256 12164 12308 12170
rect 12256 12106 12308 12112
rect 12268 11558 12296 12106
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 12360 11370 12388 13688
rect 12452 13530 12480 16238
rect 12530 16215 12586 16224
rect 12636 14074 12664 17575
rect 12728 17066 12756 18527
rect 13004 18426 13032 18838
rect 12992 18420 13044 18426
rect 12992 18362 13044 18368
rect 12808 18284 12860 18290
rect 12808 18226 12860 18232
rect 12820 17814 12848 18226
rect 13096 18034 13124 27520
rect 13452 26104 13504 26110
rect 13452 26046 13504 26052
rect 13360 25152 13412 25158
rect 13360 25094 13412 25100
rect 13372 24698 13400 25094
rect 13464 24886 13492 26046
rect 13544 25900 13596 25906
rect 13544 25842 13596 25848
rect 13556 25129 13584 25842
rect 13542 25120 13598 25129
rect 13542 25055 13598 25064
rect 13452 24880 13504 24886
rect 13452 24822 13504 24828
rect 13176 24676 13228 24682
rect 13372 24670 13584 24698
rect 13176 24618 13228 24624
rect 13188 22114 13216 24618
rect 13360 24608 13412 24614
rect 13360 24550 13412 24556
rect 13372 24070 13400 24550
rect 13452 24404 13504 24410
rect 13452 24346 13504 24352
rect 13360 24064 13412 24070
rect 13360 24006 13412 24012
rect 13268 23180 13320 23186
rect 13268 23122 13320 23128
rect 13280 22778 13308 23122
rect 13372 23050 13400 24006
rect 13464 23225 13492 24346
rect 13556 23769 13584 24670
rect 13542 23760 13598 23769
rect 13542 23695 13598 23704
rect 13556 23662 13584 23695
rect 13544 23656 13596 23662
rect 13544 23598 13596 23604
rect 13450 23216 13506 23225
rect 13450 23151 13506 23160
rect 13452 23112 13504 23118
rect 13452 23054 13504 23060
rect 13360 23044 13412 23050
rect 13360 22986 13412 22992
rect 13268 22772 13320 22778
rect 13268 22714 13320 22720
rect 13464 22234 13492 23054
rect 13544 23044 13596 23050
rect 13544 22986 13596 22992
rect 13452 22228 13504 22234
rect 13452 22170 13504 22176
rect 13450 22128 13506 22137
rect 13188 22086 13308 22114
rect 13280 22080 13308 22086
rect 13280 22052 13400 22080
rect 13450 22063 13506 22072
rect 13268 21888 13320 21894
rect 13268 21830 13320 21836
rect 13280 21350 13308 21830
rect 13268 21344 13320 21350
rect 13268 21286 13320 21292
rect 13176 20324 13228 20330
rect 13176 20266 13228 20272
rect 13188 19802 13216 20266
rect 13280 19922 13308 21286
rect 13268 19916 13320 19922
rect 13268 19858 13320 19864
rect 13188 19774 13308 19802
rect 13174 19272 13230 19281
rect 13174 19207 13230 19216
rect 13188 18086 13216 19207
rect 13004 18006 13124 18034
rect 13176 18080 13228 18086
rect 13176 18022 13228 18028
rect 12808 17808 12860 17814
rect 12808 17750 12860 17756
rect 12716 17060 12768 17066
rect 12716 17002 12768 17008
rect 12820 15910 12848 17750
rect 12900 17740 12952 17746
rect 12900 17682 12952 17688
rect 12912 16998 12940 17682
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12912 16794 12940 16934
rect 12900 16788 12952 16794
rect 12900 16730 12952 16736
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12820 15745 12848 15846
rect 12806 15736 12862 15745
rect 12806 15671 12862 15680
rect 12900 15700 12952 15706
rect 12714 15600 12770 15609
rect 12714 15535 12770 15544
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12452 12850 12480 13330
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12452 11762 12480 12786
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12440 11756 12492 11762
rect 12440 11698 12492 11704
rect 12544 11626 12572 12038
rect 12532 11620 12584 11626
rect 12532 11562 12584 11568
rect 12084 10934 12204 10962
rect 12268 11342 12388 11370
rect 11978 8800 12034 8809
rect 11978 8735 12034 8744
rect 11716 7908 11836 7936
rect 11702 7848 11758 7857
rect 11702 7783 11758 7792
rect 11716 7002 11744 7783
rect 11808 7002 11836 7908
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11796 6996 11848 7002
rect 11796 6938 11848 6944
rect 11716 6458 11744 6938
rect 11900 6798 11928 7482
rect 11888 6792 11940 6798
rect 11808 6752 11888 6780
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11808 6390 11836 6752
rect 11888 6734 11940 6740
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11796 6384 11848 6390
rect 11796 6326 11848 6332
rect 11796 5772 11848 5778
rect 11796 5714 11848 5720
rect 11702 5536 11758 5545
rect 11702 5471 11758 5480
rect 11612 4140 11664 4146
rect 11612 4082 11664 4088
rect 11532 3998 11652 4026
rect 11518 3768 11574 3777
rect 11518 3703 11574 3712
rect 11532 3670 11560 3703
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 11428 3596 11480 3602
rect 11428 3538 11480 3544
rect 11532 3126 11560 3606
rect 11336 3120 11388 3126
rect 11520 3120 11572 3126
rect 11336 3062 11388 3068
rect 11518 3088 11520 3097
rect 11572 3088 11574 3097
rect 11518 3023 11574 3032
rect 11256 2944 11468 2972
rect 11440 2666 11468 2944
rect 11440 2638 11560 2666
rect 11532 2106 11560 2638
rect 11520 2100 11572 2106
rect 11520 2042 11572 2048
rect 11532 1737 11560 2042
rect 11518 1728 11574 1737
rect 11518 1663 11574 1672
rect 11624 1465 11652 3998
rect 11610 1456 11666 1465
rect 11610 1391 11666 1400
rect 11716 480 11744 5471
rect 11808 5370 11836 5714
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11794 4856 11850 4865
rect 11794 4791 11850 4800
rect 11808 4321 11836 4791
rect 11794 4312 11850 4321
rect 11794 4247 11850 4256
rect 11796 3664 11848 3670
rect 11796 3606 11848 3612
rect 11808 2689 11836 3606
rect 11794 2680 11850 2689
rect 11794 2615 11850 2624
rect 11808 2582 11836 2615
rect 11796 2576 11848 2582
rect 11796 2518 11848 2524
rect 11900 1737 11928 6598
rect 11992 5001 12020 8735
rect 12084 7274 12112 10934
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12176 9382 12204 10066
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12268 8242 12296 11342
rect 12728 11268 12756 15535
rect 12820 14618 12848 15671
rect 12900 15642 12952 15648
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12820 13734 12848 14214
rect 12912 13938 12940 15642
rect 13004 15609 13032 18006
rect 13084 17876 13136 17882
rect 13084 17818 13136 17824
rect 13096 17678 13124 17818
rect 13084 17672 13136 17678
rect 13084 17614 13136 17620
rect 13096 16250 13124 17614
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 12990 15600 13046 15609
rect 12990 15535 13046 15544
rect 12992 14612 13044 14618
rect 12992 14554 13044 14560
rect 13004 13938 13032 14554
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 12808 13728 12860 13734
rect 12808 13670 12860 13676
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12820 13530 12848 13670
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12806 13288 12862 13297
rect 12806 13223 12808 13232
rect 12860 13223 12862 13232
rect 12808 13194 12860 13200
rect 12820 12714 12848 13194
rect 12808 12708 12860 12714
rect 12808 12650 12860 12656
rect 12912 12594 12940 13670
rect 13096 13462 13124 14350
rect 13084 13456 13136 13462
rect 12346 11248 12402 11257
rect 12346 11183 12348 11192
rect 12400 11183 12402 11192
rect 12636 11240 12756 11268
rect 12820 12566 12940 12594
rect 13004 13416 13084 13444
rect 12348 11154 12400 11160
rect 12346 11112 12402 11121
rect 12346 11047 12348 11056
rect 12400 11047 12402 11056
rect 12348 11018 12400 11024
rect 12348 10464 12400 10470
rect 12348 10406 12400 10412
rect 12360 9450 12388 10406
rect 12438 9752 12494 9761
rect 12438 9687 12440 9696
rect 12492 9687 12494 9696
rect 12440 9658 12492 9664
rect 12348 9444 12400 9450
rect 12348 9386 12400 9392
rect 12438 9072 12494 9081
rect 12438 9007 12494 9016
rect 12452 8430 12480 9007
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12176 8214 12296 8242
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12072 7268 12124 7274
rect 12072 7210 12124 7216
rect 12084 6662 12112 7210
rect 12072 6656 12124 6662
rect 12072 6598 12124 6604
rect 12070 6080 12126 6089
rect 12070 6015 12126 6024
rect 12084 5302 12112 6015
rect 12072 5296 12124 5302
rect 12072 5238 12124 5244
rect 11978 4992 12034 5001
rect 11978 4927 12034 4936
rect 12084 4758 12112 5238
rect 12072 4752 12124 4758
rect 12072 4694 12124 4700
rect 12176 4570 12204 8214
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12268 7750 12296 8026
rect 12452 8022 12480 8230
rect 12440 8016 12492 8022
rect 12440 7958 12492 7964
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12268 7546 12296 7686
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12268 4690 12296 6938
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 11992 4542 12204 4570
rect 12360 4570 12388 7890
rect 12636 7834 12664 11240
rect 12820 10985 12848 12566
rect 12806 10976 12862 10985
rect 12806 10911 12862 10920
rect 13004 10588 13032 13416
rect 13084 13398 13136 13404
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 12820 10560 13032 10588
rect 12716 9444 12768 9450
rect 12716 9386 12768 9392
rect 12728 9178 12756 9386
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 12728 7954 12756 9114
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 12820 7834 12848 10560
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 13004 8498 13032 8910
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13004 8090 13032 8434
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 12636 7806 12756 7834
rect 12820 7806 12940 7834
rect 12624 7744 12676 7750
rect 12622 7712 12624 7721
rect 12676 7712 12678 7721
rect 12622 7647 12678 7656
rect 12636 7410 12664 7647
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 12440 5840 12492 5846
rect 12440 5782 12492 5788
rect 12452 4842 12480 5782
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 12544 5302 12572 5510
rect 12636 5409 12664 6802
rect 12728 6746 12756 7806
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12820 7342 12848 7686
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12912 6866 12940 7806
rect 13004 7410 13032 8026
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 13096 6746 13124 11834
rect 13188 11218 13216 17070
rect 13280 16833 13308 19774
rect 13266 16824 13322 16833
rect 13266 16759 13322 16768
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 13280 11694 13308 16594
rect 13372 13308 13400 22052
rect 13464 19310 13492 22063
rect 13452 19304 13504 19310
rect 13452 19246 13504 19252
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 13464 18873 13492 19110
rect 13450 18864 13506 18873
rect 13450 18799 13506 18808
rect 13452 18420 13504 18426
rect 13452 18362 13504 18368
rect 13464 17882 13492 18362
rect 13452 17876 13504 17882
rect 13452 17818 13504 17824
rect 13452 17604 13504 17610
rect 13452 17546 13504 17552
rect 13464 16522 13492 17546
rect 13452 16516 13504 16522
rect 13452 16458 13504 16464
rect 13464 15638 13492 16458
rect 13452 15632 13504 15638
rect 13452 15574 13504 15580
rect 13464 15162 13492 15574
rect 13452 15156 13504 15162
rect 13452 15098 13504 15104
rect 13452 14952 13504 14958
rect 13450 14920 13452 14929
rect 13504 14920 13506 14929
rect 13450 14855 13506 14864
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13464 14657 13492 14758
rect 13450 14648 13506 14657
rect 13450 14583 13506 14592
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13464 14006 13492 14418
rect 13452 14000 13504 14006
rect 13450 13968 13452 13977
rect 13504 13968 13506 13977
rect 13450 13903 13506 13912
rect 13452 13456 13504 13462
rect 13450 13424 13452 13433
rect 13504 13424 13506 13433
rect 13450 13359 13506 13368
rect 13372 13280 13492 13308
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 13188 10742 13216 11154
rect 13176 10736 13228 10742
rect 13176 10678 13228 10684
rect 13174 9208 13230 9217
rect 13174 9143 13230 9152
rect 13268 9172 13320 9178
rect 13188 9110 13216 9143
rect 13268 9114 13320 9120
rect 13176 9104 13228 9110
rect 13176 9046 13228 9052
rect 12728 6718 12848 6746
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12728 6254 12756 6598
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 12622 5400 12678 5409
rect 12622 5335 12678 5344
rect 12532 5296 12584 5302
rect 12532 5238 12584 5244
rect 12622 5128 12678 5137
rect 12622 5063 12678 5072
rect 12636 5030 12664 5063
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12452 4814 12664 4842
rect 12360 4542 12572 4570
rect 11992 4078 12020 4542
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 12254 4312 12310 4321
rect 12254 4247 12310 4256
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 12084 2009 12112 3878
rect 12070 2000 12126 2009
rect 12070 1935 12126 1944
rect 11886 1728 11942 1737
rect 11886 1663 11942 1672
rect 12268 480 12296 4247
rect 12360 4010 12388 4422
rect 12438 4040 12494 4049
rect 12348 4004 12400 4010
rect 12438 3975 12494 3984
rect 12348 3946 12400 3952
rect 12452 3942 12480 3975
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12438 3360 12494 3369
rect 12438 3295 12494 3304
rect 12452 3194 12480 3295
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12544 1970 12572 4542
rect 12636 4078 12664 4814
rect 12728 4214 12756 6190
rect 12820 5681 12848 6718
rect 13004 6718 13124 6746
rect 12900 6180 12952 6186
rect 12900 6122 12952 6128
rect 12912 5817 12940 6122
rect 13004 6089 13032 6718
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 12990 6080 13046 6089
rect 12990 6015 13046 6024
rect 12898 5808 12954 5817
rect 12898 5743 12954 5752
rect 12806 5672 12862 5681
rect 12806 5607 12862 5616
rect 12716 4208 12768 4214
rect 12716 4150 12768 4156
rect 12624 4072 12676 4078
rect 12624 4014 12676 4020
rect 12716 3664 12768 3670
rect 12716 3606 12768 3612
rect 12728 2922 12756 3606
rect 12820 3466 12848 5607
rect 13004 5273 13032 6015
rect 12990 5264 13046 5273
rect 12990 5199 13046 5208
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 13004 4729 13032 4966
rect 13096 4826 13124 6598
rect 13174 5808 13230 5817
rect 13174 5743 13176 5752
rect 13228 5743 13230 5752
rect 13176 5714 13228 5720
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 12990 4720 13046 4729
rect 12990 4655 13046 4664
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 12808 3460 12860 3466
rect 12808 3402 12860 3408
rect 12820 2990 12848 3402
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 12716 2916 12768 2922
rect 12716 2858 12768 2864
rect 12808 2848 12860 2854
rect 12808 2790 12860 2796
rect 12532 1964 12584 1970
rect 12532 1906 12584 1912
rect 12820 480 12848 2790
rect 13004 2281 13032 4422
rect 13280 3618 13308 9114
rect 13372 6866 13400 12922
rect 13464 9178 13492 13280
rect 13556 11898 13584 22986
rect 13648 17241 13676 27520
rect 13820 25764 13872 25770
rect 13820 25706 13872 25712
rect 13832 25498 13860 25706
rect 13728 25492 13780 25498
rect 13728 25434 13780 25440
rect 13820 25492 13872 25498
rect 13820 25434 13872 25440
rect 14096 25492 14148 25498
rect 14096 25434 14148 25440
rect 13740 24886 13768 25434
rect 13728 24880 13780 24886
rect 13728 24822 13780 24828
rect 14004 24812 14056 24818
rect 14004 24754 14056 24760
rect 13820 24404 13872 24410
rect 13820 24346 13872 24352
rect 13832 23866 13860 24346
rect 13912 24200 13964 24206
rect 13912 24142 13964 24148
rect 13820 23860 13872 23866
rect 13820 23802 13872 23808
rect 13728 23724 13780 23730
rect 13728 23666 13780 23672
rect 13740 23118 13768 23666
rect 13728 23112 13780 23118
rect 13728 23054 13780 23060
rect 13740 22506 13768 23054
rect 13924 22982 13952 24142
rect 14016 23050 14044 24754
rect 14108 24410 14136 25434
rect 14292 24993 14320 27520
rect 14464 26308 14516 26314
rect 14464 26250 14516 26256
rect 14476 25945 14504 26250
rect 14462 25936 14518 25945
rect 14462 25871 14518 25880
rect 14372 25288 14424 25294
rect 14372 25230 14424 25236
rect 14648 25288 14700 25294
rect 14648 25230 14700 25236
rect 14278 24984 14334 24993
rect 14384 24954 14412 25230
rect 14556 25220 14608 25226
rect 14556 25162 14608 25168
rect 14278 24919 14334 24928
rect 14372 24948 14424 24954
rect 14372 24890 14424 24896
rect 14280 24812 14332 24818
rect 14280 24754 14332 24760
rect 14096 24404 14148 24410
rect 14096 24346 14148 24352
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 14108 23594 14136 24142
rect 14096 23588 14148 23594
rect 14096 23530 14148 23536
rect 14004 23044 14056 23050
rect 14004 22986 14056 22992
rect 13912 22976 13964 22982
rect 13912 22918 13964 22924
rect 13818 22672 13874 22681
rect 13818 22607 13874 22616
rect 13832 22574 13860 22607
rect 13820 22568 13872 22574
rect 13820 22510 13872 22516
rect 13728 22500 13780 22506
rect 13728 22442 13780 22448
rect 13740 21418 13768 22442
rect 13924 22234 13952 22918
rect 13912 22228 13964 22234
rect 13912 22170 13964 22176
rect 14004 22160 14056 22166
rect 14004 22102 14056 22108
rect 13912 22024 13964 22030
rect 13912 21966 13964 21972
rect 13924 21418 13952 21966
rect 13728 21412 13780 21418
rect 13728 21354 13780 21360
rect 13912 21412 13964 21418
rect 13912 21354 13964 21360
rect 13740 20874 13768 21354
rect 13820 21004 13872 21010
rect 13820 20946 13872 20952
rect 13728 20868 13780 20874
rect 13728 20810 13780 20816
rect 13740 20058 13768 20810
rect 13832 20602 13860 20946
rect 13820 20596 13872 20602
rect 13820 20538 13872 20544
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 13728 19916 13780 19922
rect 13728 19858 13780 19864
rect 13740 18970 13768 19858
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 13728 18964 13780 18970
rect 13728 18906 13780 18912
rect 13832 18850 13860 19246
rect 13924 19174 13952 21354
rect 13912 19168 13964 19174
rect 13912 19110 13964 19116
rect 13740 18822 13860 18850
rect 13740 18601 13768 18822
rect 13820 18692 13872 18698
rect 13820 18634 13872 18640
rect 13726 18592 13782 18601
rect 13726 18527 13782 18536
rect 13728 18352 13780 18358
rect 13728 18294 13780 18300
rect 13740 17921 13768 18294
rect 13726 17912 13782 17921
rect 13726 17847 13782 17856
rect 13832 17626 13860 18634
rect 14016 18426 14044 22102
rect 14108 21690 14136 23530
rect 14186 22808 14242 22817
rect 14186 22743 14242 22752
rect 14096 21684 14148 21690
rect 14096 21626 14148 21632
rect 14094 21176 14150 21185
rect 14094 21111 14150 21120
rect 14108 21078 14136 21111
rect 14096 21072 14148 21078
rect 14096 21014 14148 21020
rect 14200 20754 14228 22743
rect 14292 21350 14320 24754
rect 14464 24744 14516 24750
rect 14464 24686 14516 24692
rect 14476 24585 14504 24686
rect 14462 24576 14518 24585
rect 14462 24511 14518 24520
rect 14372 22636 14424 22642
rect 14372 22578 14424 22584
rect 14280 21344 14332 21350
rect 14280 21286 14332 21292
rect 14280 21072 14332 21078
rect 14280 21014 14332 21020
rect 14108 20726 14228 20754
rect 14108 19310 14136 20726
rect 14186 20632 14242 20641
rect 14186 20567 14188 20576
rect 14240 20567 14242 20576
rect 14188 20538 14240 20544
rect 14188 19508 14240 19514
rect 14188 19450 14240 19456
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 14200 19156 14228 19450
rect 14108 19128 14228 19156
rect 14004 18420 14056 18426
rect 14004 18362 14056 18368
rect 13912 18216 13964 18222
rect 13912 18158 13964 18164
rect 13740 17598 13860 17626
rect 13634 17232 13690 17241
rect 13634 17167 13690 17176
rect 13636 16992 13688 16998
rect 13636 16934 13688 16940
rect 13648 16658 13676 16934
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 13636 16516 13688 16522
rect 13636 16458 13688 16464
rect 13648 16289 13676 16458
rect 13634 16280 13690 16289
rect 13634 16215 13690 16224
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13648 15570 13676 16050
rect 13636 15564 13688 15570
rect 13636 15506 13688 15512
rect 13634 15464 13690 15473
rect 13634 15399 13690 15408
rect 13648 14550 13676 15399
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13648 14074 13676 14214
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 13634 13832 13690 13841
rect 13634 13767 13690 13776
rect 13648 12986 13676 13767
rect 13740 13258 13768 17598
rect 13924 17542 13952 18158
rect 13820 17536 13872 17542
rect 13820 17478 13872 17484
rect 13912 17536 13964 17542
rect 14108 17513 14136 19128
rect 14186 18320 14242 18329
rect 14186 18255 14242 18264
rect 14200 17882 14228 18255
rect 14188 17876 14240 17882
rect 14188 17818 14240 17824
rect 13912 17478 13964 17484
rect 14094 17504 14150 17513
rect 13832 13569 13860 17478
rect 13924 16697 13952 17478
rect 14094 17439 14150 17448
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 13910 16688 13966 16697
rect 13910 16623 13966 16632
rect 13924 16590 13952 16623
rect 13912 16584 13964 16590
rect 13912 16526 13964 16532
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13924 14958 13952 15438
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 13912 14544 13964 14550
rect 13912 14486 13964 14492
rect 13924 14006 13952 14486
rect 13912 14000 13964 14006
rect 13912 13942 13964 13948
rect 13818 13560 13874 13569
rect 13818 13495 13874 13504
rect 13832 13326 13860 13495
rect 13910 13424 13966 13433
rect 13910 13359 13912 13368
rect 13964 13359 13966 13368
rect 13912 13330 13964 13336
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13728 13252 13780 13258
rect 13728 13194 13780 13200
rect 13726 13152 13782 13161
rect 13726 13087 13782 13096
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13634 12336 13690 12345
rect 13634 12271 13690 12280
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13544 11620 13596 11626
rect 13544 11562 13596 11568
rect 13556 10577 13584 11562
rect 13648 11354 13676 12271
rect 13740 11898 13768 13087
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 13832 11762 13860 12718
rect 14016 12374 14044 17274
rect 14186 17232 14242 17241
rect 14186 17167 14242 17176
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 14108 16726 14136 16934
rect 14096 16720 14148 16726
rect 14096 16662 14148 16668
rect 14108 15162 14136 16662
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 14108 13462 14136 14758
rect 14096 13456 14148 13462
rect 14094 13424 14096 13433
rect 14148 13424 14150 13433
rect 14094 13359 14150 13368
rect 14096 12436 14148 12442
rect 14096 12378 14148 12384
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13912 11688 13964 11694
rect 13818 11656 13874 11665
rect 13912 11630 13964 11636
rect 13818 11591 13874 11600
rect 13832 11558 13860 11591
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13924 11354 13952 11630
rect 13636 11348 13688 11354
rect 13912 11348 13964 11354
rect 13636 11290 13688 11296
rect 13740 11308 13912 11336
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13542 10568 13598 10577
rect 13542 10503 13598 10512
rect 13556 9994 13584 10503
rect 13648 10266 13676 11154
rect 13740 10810 13768 11308
rect 13912 11290 13964 11296
rect 14016 11234 14044 12310
rect 13832 11206 14044 11234
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13544 9988 13596 9994
rect 13544 9930 13596 9936
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 13464 8090 13492 8978
rect 13556 8974 13584 9318
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13556 8634 13584 8910
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13648 7970 13676 8774
rect 13832 8106 13860 11206
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 13924 10266 13952 11086
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 13912 9104 13964 9110
rect 13912 9046 13964 9052
rect 13924 8294 13952 9046
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13832 8078 13952 8106
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13556 7942 13676 7970
rect 13820 8016 13872 8022
rect 13820 7958 13872 7964
rect 13464 7478 13492 7890
rect 13452 7472 13504 7478
rect 13452 7414 13504 7420
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 13372 6458 13400 6802
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13358 4992 13414 5001
rect 13358 4927 13414 4936
rect 13372 4185 13400 4927
rect 13358 4176 13414 4185
rect 13358 4111 13414 4120
rect 13096 3602 13308 3618
rect 13084 3596 13308 3602
rect 13136 3590 13308 3596
rect 13084 3538 13136 3544
rect 12990 2272 13046 2281
rect 12990 2207 13046 2216
rect 13372 480 13400 4111
rect 13464 3754 13492 6734
rect 13556 5250 13584 7942
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13648 7546 13676 7822
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13634 7032 13690 7041
rect 13634 6967 13690 6976
rect 13648 6118 13676 6967
rect 13728 6928 13780 6934
rect 13728 6870 13780 6876
rect 13740 6458 13768 6870
rect 13832 6866 13860 7958
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13740 5545 13768 6394
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13726 5536 13782 5545
rect 13726 5471 13782 5480
rect 13832 5386 13860 5646
rect 13740 5358 13860 5386
rect 13556 5222 13676 5250
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13556 4865 13584 4966
rect 13542 4856 13598 4865
rect 13542 4791 13598 4800
rect 13648 4706 13676 5222
rect 13556 4678 13676 4706
rect 13556 4049 13584 4678
rect 13634 4584 13690 4593
rect 13634 4519 13636 4528
rect 13688 4519 13690 4528
rect 13636 4490 13688 4496
rect 13740 4162 13768 5358
rect 13648 4134 13768 4162
rect 13542 4040 13598 4049
rect 13542 3975 13598 3984
rect 13464 3726 13584 3754
rect 13452 3664 13504 3670
rect 13452 3606 13504 3612
rect 13464 2854 13492 3606
rect 13556 3505 13584 3726
rect 13542 3496 13598 3505
rect 13542 3431 13598 3440
rect 13648 2922 13676 4134
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13636 2916 13688 2922
rect 13636 2858 13688 2864
rect 13452 2848 13504 2854
rect 13452 2790 13504 2796
rect 13464 2106 13492 2790
rect 13740 2378 13768 4014
rect 13924 2990 13952 8078
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 14016 2836 14044 10950
rect 14108 8786 14136 12378
rect 14200 9654 14228 17167
rect 14292 16969 14320 21014
rect 14384 20602 14412 22578
rect 14372 20596 14424 20602
rect 14372 20538 14424 20544
rect 14370 19000 14426 19009
rect 14370 18935 14426 18944
rect 14384 18086 14412 18935
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14372 17672 14424 17678
rect 14372 17614 14424 17620
rect 14384 16980 14412 17614
rect 14476 17338 14504 24511
rect 14568 24392 14596 25162
rect 14660 24954 14688 25230
rect 14740 25152 14792 25158
rect 14740 25094 14792 25100
rect 14752 24954 14780 25094
rect 14648 24948 14700 24954
rect 14648 24890 14700 24896
rect 14740 24948 14792 24954
rect 14740 24890 14792 24896
rect 14844 24818 14872 27520
rect 15292 25356 15344 25362
rect 15292 25298 15344 25304
rect 15304 25226 15332 25298
rect 15292 25220 15344 25226
rect 15292 25162 15344 25168
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15292 24948 15344 24954
rect 15292 24890 15344 24896
rect 15108 24880 15160 24886
rect 14922 24848 14978 24857
rect 14832 24812 14884 24818
rect 15108 24822 15160 24828
rect 14922 24783 14978 24792
rect 14832 24754 14884 24760
rect 14832 24676 14884 24682
rect 14832 24618 14884 24624
rect 14568 24364 14780 24392
rect 14648 24268 14700 24274
rect 14648 24210 14700 24216
rect 14660 23526 14688 24210
rect 14648 23520 14700 23526
rect 14648 23462 14700 23468
rect 14556 22568 14608 22574
rect 14556 22510 14608 22516
rect 14568 22030 14596 22510
rect 14556 22024 14608 22030
rect 14556 21966 14608 21972
rect 14660 21962 14688 23462
rect 14752 22522 14780 24364
rect 14844 23361 14872 24618
rect 14936 24614 14964 24783
rect 15120 24614 15148 24822
rect 14924 24608 14976 24614
rect 15108 24608 15160 24614
rect 14924 24550 14976 24556
rect 15106 24576 15108 24585
rect 15160 24576 15162 24585
rect 15106 24511 15162 24520
rect 15304 24342 15332 24890
rect 15292 24336 15344 24342
rect 15292 24278 15344 24284
rect 15292 24200 15344 24206
rect 15292 24142 15344 24148
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15200 23724 15252 23730
rect 15200 23666 15252 23672
rect 15212 23474 15240 23666
rect 15028 23446 15240 23474
rect 14830 23352 14886 23361
rect 14830 23287 14886 23296
rect 15028 23254 15056 23446
rect 15304 23338 15332 24142
rect 15120 23322 15332 23338
rect 15108 23316 15332 23322
rect 15160 23310 15332 23316
rect 15108 23258 15160 23264
rect 15016 23248 15068 23254
rect 15016 23190 15068 23196
rect 15290 23216 15346 23225
rect 15290 23151 15346 23160
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14752 22494 14872 22522
rect 14740 22432 14792 22438
rect 14740 22374 14792 22380
rect 14648 21956 14700 21962
rect 14648 21898 14700 21904
rect 14556 21344 14608 21350
rect 14556 21286 14608 21292
rect 14568 19514 14596 21286
rect 14648 20256 14700 20262
rect 14648 20198 14700 20204
rect 14660 19990 14688 20198
rect 14648 19984 14700 19990
rect 14646 19952 14648 19961
rect 14700 19952 14702 19961
rect 14646 19887 14702 19896
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 14568 18902 14596 19314
rect 14556 18896 14608 18902
rect 14556 18838 14608 18844
rect 14568 18290 14596 18838
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14568 17814 14596 18226
rect 14556 17808 14608 17814
rect 14556 17750 14608 17756
rect 14464 17332 14516 17338
rect 14464 17274 14516 17280
rect 14464 17128 14516 17134
rect 14462 17096 14464 17105
rect 14516 17096 14518 17105
rect 14462 17031 14518 17040
rect 14278 16960 14334 16969
rect 14384 16952 14504 16980
rect 14278 16895 14334 16904
rect 14370 16824 14426 16833
rect 14370 16759 14372 16768
rect 14424 16759 14426 16768
rect 14372 16730 14424 16736
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14292 13920 14320 16526
rect 14384 16250 14412 16526
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 14370 16144 14426 16153
rect 14370 16079 14426 16088
rect 14384 15978 14412 16079
rect 14372 15972 14424 15978
rect 14372 15914 14424 15920
rect 14384 15706 14412 15914
rect 14476 15706 14504 16952
rect 14568 16726 14596 17750
rect 14648 17740 14700 17746
rect 14648 17682 14700 17688
rect 14660 17270 14688 17682
rect 14752 17678 14780 22374
rect 14844 22098 14872 22494
rect 15108 22432 15160 22438
rect 15108 22374 15160 22380
rect 15120 22273 15148 22374
rect 15106 22264 15162 22273
rect 15106 22199 15162 22208
rect 14832 22092 14884 22098
rect 14832 22034 14884 22040
rect 14844 21486 14872 22034
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14832 21480 14884 21486
rect 14832 21422 14884 21428
rect 15304 21010 15332 23151
rect 15292 21004 15344 21010
rect 15292 20946 15344 20952
rect 14832 20868 14884 20874
rect 14832 20810 14884 20816
rect 14844 20482 14872 20810
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15106 20496 15162 20505
rect 14844 20466 14964 20482
rect 14844 20460 14976 20466
rect 14844 20454 14924 20460
rect 15106 20431 15162 20440
rect 14924 20402 14976 20408
rect 14830 20360 14886 20369
rect 14830 20295 14886 20304
rect 14844 19961 14872 20295
rect 15120 20058 15148 20431
rect 15108 20052 15160 20058
rect 15108 19994 15160 20000
rect 14830 19952 14886 19961
rect 14830 19887 14886 19896
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15200 19440 15252 19446
rect 15200 19382 15252 19388
rect 15212 19156 15240 19382
rect 15304 19310 15332 20946
rect 15396 20890 15424 27520
rect 15934 26072 15990 26081
rect 15934 26007 15990 26016
rect 15948 24993 15976 26007
rect 15934 24984 15990 24993
rect 15934 24919 15990 24928
rect 15476 24812 15528 24818
rect 15476 24754 15528 24760
rect 15488 24410 15516 24754
rect 15566 24440 15622 24449
rect 15476 24404 15528 24410
rect 15566 24375 15568 24384
rect 15476 24346 15528 24352
rect 15620 24375 15622 24384
rect 15844 24404 15896 24410
rect 15568 24346 15620 24352
rect 15844 24346 15896 24352
rect 15660 24064 15712 24070
rect 15660 24006 15712 24012
rect 15752 24064 15804 24070
rect 15752 24006 15804 24012
rect 15474 23896 15530 23905
rect 15474 23831 15476 23840
rect 15528 23831 15530 23840
rect 15476 23802 15528 23808
rect 15474 23624 15530 23633
rect 15474 23559 15530 23568
rect 15488 21078 15516 23559
rect 15672 23497 15700 24006
rect 15658 23488 15714 23497
rect 15658 23423 15714 23432
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 15672 22953 15700 23054
rect 15658 22944 15714 22953
rect 15658 22879 15714 22888
rect 15672 22778 15700 22879
rect 15660 22772 15712 22778
rect 15660 22714 15712 22720
rect 15672 22080 15700 22714
rect 15580 22052 15700 22080
rect 15580 21298 15608 22052
rect 15580 21270 15700 21298
rect 15476 21072 15528 21078
rect 15476 21014 15528 21020
rect 15396 20862 15516 20890
rect 15384 20800 15436 20806
rect 15384 20742 15436 20748
rect 15396 20602 15424 20742
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15384 19916 15436 19922
rect 15384 19858 15436 19864
rect 15396 19378 15424 19858
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15212 19128 15332 19156
rect 14832 18624 14884 18630
rect 14832 18566 14884 18572
rect 14844 17728 14872 18566
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15108 18080 15160 18086
rect 15160 18028 15240 18034
rect 15108 18022 15240 18028
rect 15120 18006 15240 18022
rect 15106 17912 15162 17921
rect 15106 17847 15108 17856
rect 15160 17847 15162 17856
rect 15108 17818 15160 17824
rect 15212 17762 15240 18006
rect 15304 17882 15332 19128
rect 15384 18828 15436 18834
rect 15384 18770 15436 18776
rect 15396 18426 15424 18770
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15384 18148 15436 18154
rect 15384 18090 15436 18096
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15212 17734 15332 17762
rect 14844 17700 14964 17728
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 14830 17640 14886 17649
rect 14936 17610 14964 17700
rect 14830 17575 14886 17584
rect 14924 17604 14976 17610
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14648 17264 14700 17270
rect 14648 17206 14700 17212
rect 14648 17128 14700 17134
rect 14646 17096 14648 17105
rect 14700 17096 14702 17105
rect 14646 17031 14702 17040
rect 14660 16794 14688 17031
rect 14752 16969 14780 17478
rect 14844 17338 14872 17575
rect 14924 17546 14976 17552
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14832 17332 14884 17338
rect 14832 17274 14884 17280
rect 15200 17128 15252 17134
rect 15200 17070 15252 17076
rect 15108 16992 15160 16998
rect 14738 16960 14794 16969
rect 15108 16934 15160 16940
rect 14738 16895 14794 16904
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 14556 16720 14608 16726
rect 14556 16662 14608 16668
rect 15120 16522 15148 16934
rect 15212 16697 15240 17070
rect 15198 16688 15254 16697
rect 15198 16623 15200 16632
rect 15252 16623 15254 16632
rect 15200 16594 15252 16600
rect 15212 16563 15240 16594
rect 15108 16516 15160 16522
rect 15108 16458 15160 16464
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14738 16280 14794 16289
rect 14956 16272 15252 16292
rect 14738 16215 14794 16224
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 14384 15586 14412 15642
rect 14384 15558 14596 15586
rect 14372 15428 14424 15434
rect 14372 15370 14424 15376
rect 14384 15026 14412 15370
rect 14372 15020 14424 15026
rect 14372 14962 14424 14968
rect 14464 15020 14516 15026
rect 14464 14962 14516 14968
rect 14476 14618 14504 14962
rect 14464 14612 14516 14618
rect 14464 14554 14516 14560
rect 14476 14414 14504 14554
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14476 13977 14504 14350
rect 14462 13968 14518 13977
rect 14292 13892 14412 13920
rect 14462 13903 14518 13912
rect 14280 13456 14332 13462
rect 14280 13398 14332 13404
rect 14292 11286 14320 13398
rect 14384 12481 14412 13892
rect 14464 13864 14516 13870
rect 14462 13832 14464 13841
rect 14516 13832 14518 13841
rect 14462 13767 14518 13776
rect 14568 13326 14596 15558
rect 14646 15192 14702 15201
rect 14646 15127 14702 15136
rect 14660 14074 14688 15127
rect 14752 14634 14780 16215
rect 15304 15570 15332 17734
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 14832 15360 14884 15366
rect 14832 15302 14884 15308
rect 14844 14793 14872 15302
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15106 15056 15162 15065
rect 15106 14991 15162 15000
rect 14830 14784 14886 14793
rect 14830 14719 14886 14728
rect 14752 14606 14872 14634
rect 15120 14618 15148 14991
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 14738 14240 14794 14249
rect 14738 14175 14794 14184
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14646 13968 14702 13977
rect 14646 13903 14648 13912
rect 14700 13903 14702 13912
rect 14648 13874 14700 13880
rect 14660 13326 14688 13874
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14568 12986 14596 13262
rect 14646 13016 14702 13025
rect 14556 12980 14608 12986
rect 14646 12951 14702 12960
rect 14556 12922 14608 12928
rect 14464 12640 14516 12646
rect 14464 12582 14516 12588
rect 14370 12472 14426 12481
rect 14370 12407 14426 12416
rect 14476 12356 14504 12582
rect 14384 12328 14504 12356
rect 14280 11280 14332 11286
rect 14280 11222 14332 11228
rect 14384 11218 14412 12328
rect 14464 12232 14516 12238
rect 14660 12220 14688 12951
rect 14464 12174 14516 12180
rect 14568 12192 14688 12220
rect 14476 12073 14504 12174
rect 14462 12064 14518 12073
rect 14462 11999 14518 12008
rect 14568 11830 14596 12192
rect 14646 11928 14702 11937
rect 14646 11863 14702 11872
rect 14556 11824 14608 11830
rect 14556 11766 14608 11772
rect 14568 11694 14596 11766
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 14372 11212 14424 11218
rect 14372 11154 14424 11160
rect 14280 11076 14332 11082
rect 14280 11018 14332 11024
rect 14292 10606 14320 11018
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14384 10470 14412 11154
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14292 9722 14320 10066
rect 14384 9897 14412 10406
rect 14464 9920 14516 9926
rect 14370 9888 14426 9897
rect 14464 9862 14516 9868
rect 14370 9823 14426 9832
rect 14280 9716 14332 9722
rect 14280 9658 14332 9664
rect 14188 9648 14240 9654
rect 14188 9590 14240 9596
rect 14372 8900 14424 8906
rect 14372 8842 14424 8848
rect 14108 8758 14320 8786
rect 14186 8664 14242 8673
rect 14186 8599 14242 8608
rect 14096 8288 14148 8294
rect 14096 8230 14148 8236
rect 14108 8090 14136 8230
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 14200 6746 14228 8599
rect 14292 8242 14320 8758
rect 14384 8566 14412 8842
rect 14372 8560 14424 8566
rect 14370 8528 14372 8537
rect 14424 8528 14426 8537
rect 14370 8463 14426 8472
rect 14292 8214 14412 8242
rect 14278 8120 14334 8129
rect 14278 8055 14334 8064
rect 14292 7818 14320 8055
rect 14280 7812 14332 7818
rect 14280 7754 14332 7760
rect 14384 7154 14412 8214
rect 14476 7698 14504 9862
rect 14568 8294 14596 11630
rect 14660 11558 14688 11863
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14660 11354 14688 11494
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 14646 10840 14702 10849
rect 14646 10775 14702 10784
rect 14660 10130 14688 10775
rect 14648 10124 14700 10130
rect 14648 10066 14700 10072
rect 14752 9654 14780 14175
rect 14844 11014 14872 14606
rect 15108 14612 15160 14618
rect 15108 14554 15160 14560
rect 15304 14550 15332 14758
rect 15292 14544 15344 14550
rect 15106 14512 15162 14521
rect 15292 14486 15344 14492
rect 15106 14447 15162 14456
rect 15120 14346 15148 14447
rect 15290 14376 15346 14385
rect 15108 14340 15160 14346
rect 15290 14311 15292 14320
rect 15108 14282 15160 14288
rect 15344 14311 15346 14320
rect 15292 14282 15344 14288
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15290 13968 15346 13977
rect 15290 13903 15346 13912
rect 15304 13326 15332 13903
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15304 12782 15332 13262
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 14924 12708 14976 12714
rect 14924 12650 14976 12656
rect 14936 12481 14964 12650
rect 14922 12472 14978 12481
rect 14922 12407 14978 12416
rect 15304 12306 15332 12718
rect 15396 12617 15424 18090
rect 15488 15706 15516 20862
rect 15566 20632 15622 20641
rect 15566 20567 15622 20576
rect 15476 15700 15528 15706
rect 15476 15642 15528 15648
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 15382 12608 15438 12617
rect 15382 12543 15438 12552
rect 15382 12336 15438 12345
rect 15292 12300 15344 12306
rect 15382 12271 15438 12280
rect 15292 12242 15344 12248
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15200 11620 15252 11626
rect 15200 11562 15252 11568
rect 15212 11150 15240 11562
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 14832 11008 14884 11014
rect 14832 10950 14884 10956
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14832 10736 14884 10742
rect 14830 10704 14832 10713
rect 15200 10736 15252 10742
rect 14884 10704 14886 10713
rect 15200 10678 15252 10684
rect 14830 10639 14886 10648
rect 15212 10554 15240 10678
rect 15304 10674 15332 12038
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15212 10526 15332 10554
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15212 10266 15240 10406
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 15106 9616 15162 9625
rect 15106 9551 15162 9560
rect 14660 9518 14688 9549
rect 15120 9518 15148 9551
rect 14648 9512 14700 9518
rect 14646 9480 14648 9489
rect 15108 9512 15160 9518
rect 14700 9480 14702 9489
rect 14646 9415 14702 9424
rect 14830 9480 14886 9489
rect 15108 9454 15160 9460
rect 14830 9415 14886 9424
rect 15016 9444 15068 9450
rect 14660 9178 14688 9415
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14844 9058 14872 9415
rect 15016 9386 15068 9392
rect 15028 9217 15056 9386
rect 15014 9208 15070 9217
rect 15120 9178 15148 9454
rect 15014 9143 15070 9152
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 14660 9030 14872 9058
rect 14660 8673 14688 9030
rect 14830 8936 14886 8945
rect 14830 8871 14886 8880
rect 14646 8664 14702 8673
rect 14646 8599 14702 8608
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14476 7670 14596 7698
rect 14384 7126 14504 7154
rect 14370 7032 14426 7041
rect 14370 6967 14426 6976
rect 14108 6718 14228 6746
rect 14108 5370 14136 6718
rect 14188 6656 14240 6662
rect 14188 6598 14240 6604
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14200 6254 14228 6598
rect 14292 6458 14320 6598
rect 14280 6452 14332 6458
rect 14280 6394 14332 6400
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 14188 5840 14240 5846
rect 14188 5782 14240 5788
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 14200 5234 14228 5782
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 14200 4706 14228 5170
rect 14200 4678 14320 4706
rect 14096 4616 14148 4622
rect 14094 4584 14096 4593
rect 14188 4616 14240 4622
rect 14148 4584 14150 4593
rect 14188 4558 14240 4564
rect 14094 4519 14150 4528
rect 14200 4282 14228 4558
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 14292 4010 14320 4678
rect 14280 4004 14332 4010
rect 14280 3946 14332 3952
rect 14384 3738 14412 6967
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 14384 3058 14412 3334
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 13924 2808 14044 2836
rect 14370 2816 14426 2825
rect 13728 2372 13780 2378
rect 13728 2314 13780 2320
rect 13452 2100 13504 2106
rect 13452 2042 13504 2048
rect 13924 480 13952 2808
rect 14370 2751 14426 2760
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 14016 2553 14044 2586
rect 14002 2544 14058 2553
rect 14002 2479 14058 2488
rect 14384 480 14412 2751
rect 14476 2666 14504 7126
rect 14568 3777 14596 7670
rect 14752 7274 14780 8570
rect 14844 8090 14872 8871
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15106 8528 15162 8537
rect 15106 8463 15162 8472
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14936 7834 14964 8366
rect 15120 7857 15148 8463
rect 15304 8090 15332 10526
rect 15396 9178 15424 12271
rect 15384 9172 15436 9178
rect 15384 9114 15436 9120
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 14844 7806 14964 7834
rect 15106 7848 15162 7857
rect 14844 7342 14872 7806
rect 15106 7783 15162 7792
rect 15290 7848 15346 7857
rect 15290 7783 15292 7792
rect 15344 7783 15346 7792
rect 15292 7754 15344 7760
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 14740 7268 14792 7274
rect 14740 7210 14792 7216
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 14660 6633 14688 6734
rect 14646 6624 14702 6633
rect 14646 6559 14702 6568
rect 14660 5914 14688 6559
rect 14844 6186 14872 7278
rect 15028 7002 15056 7278
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15016 6996 15068 7002
rect 15016 6938 15068 6944
rect 15108 6724 15160 6730
rect 15212 6712 15240 7142
rect 15290 6896 15346 6905
rect 15290 6831 15346 6840
rect 15304 6730 15332 6831
rect 15160 6684 15240 6712
rect 15292 6724 15344 6730
rect 15108 6666 15160 6672
rect 15292 6666 15344 6672
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15016 6384 15068 6390
rect 15016 6326 15068 6332
rect 14832 6180 14884 6186
rect 14832 6122 14884 6128
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14844 5778 14872 6122
rect 15028 5914 15056 6326
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15016 5908 15068 5914
rect 15016 5850 15068 5856
rect 14832 5772 14884 5778
rect 14832 5714 14884 5720
rect 14844 5250 14872 5714
rect 15028 5710 15056 5850
rect 15304 5817 15332 6054
rect 15290 5808 15346 5817
rect 15290 5743 15346 5752
rect 15016 5704 15068 5710
rect 15016 5646 15068 5652
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14752 5234 14872 5250
rect 14752 5228 14884 5234
rect 14752 5222 14832 5228
rect 14646 4856 14702 4865
rect 14646 4791 14702 4800
rect 14554 3768 14610 3777
rect 14660 3738 14688 4791
rect 14752 4078 14780 5222
rect 14832 5170 14884 5176
rect 14832 5092 14884 5098
rect 14832 5034 14884 5040
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 14554 3703 14610 3712
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14752 3602 14780 4014
rect 14740 3596 14792 3602
rect 14740 3538 14792 3544
rect 14844 3194 14872 5034
rect 15014 4992 15070 5001
rect 15014 4927 15070 4936
rect 15028 4826 15056 4927
rect 15016 4820 15068 4826
rect 15016 4762 15068 4768
rect 15292 4548 15344 4554
rect 15292 4490 15344 4496
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14832 3188 14884 3194
rect 14832 3130 14884 3136
rect 15304 2990 15332 4490
rect 15292 2984 15344 2990
rect 14922 2952 14978 2961
rect 15396 2972 15424 8230
rect 15488 8106 15516 15506
rect 15580 10538 15608 20567
rect 15672 16250 15700 21270
rect 15660 16244 15712 16250
rect 15660 16186 15712 16192
rect 15660 15972 15712 15978
rect 15660 15914 15712 15920
rect 15672 15745 15700 15914
rect 15658 15736 15714 15745
rect 15658 15671 15714 15680
rect 15660 15428 15712 15434
rect 15660 15370 15712 15376
rect 15672 15162 15700 15370
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 15658 14648 15714 14657
rect 15658 14583 15660 14592
rect 15712 14583 15714 14592
rect 15660 14554 15712 14560
rect 15672 14074 15700 14554
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 15764 12986 15792 24006
rect 15856 23866 15884 24346
rect 15844 23860 15896 23866
rect 15844 23802 15896 23808
rect 15948 23769 15976 24919
rect 16040 24857 16068 27520
rect 16120 26308 16172 26314
rect 16120 26250 16172 26256
rect 16132 26081 16160 26250
rect 16118 26072 16174 26081
rect 16592 26042 16620 27520
rect 16118 26007 16174 26016
rect 16580 26036 16632 26042
rect 16580 25978 16632 25984
rect 17144 25838 17172 27520
rect 17132 25832 17184 25838
rect 17132 25774 17184 25780
rect 17224 25764 17276 25770
rect 17224 25706 17276 25712
rect 17038 25528 17094 25537
rect 16212 25492 16264 25498
rect 17094 25486 17172 25514
rect 17038 25463 17094 25472
rect 16212 25434 16264 25440
rect 16120 25356 16172 25362
rect 16120 25298 16172 25304
rect 16026 24848 16082 24857
rect 16026 24783 16082 24792
rect 16132 24614 16160 25298
rect 16224 24682 16252 25434
rect 16580 25424 16632 25430
rect 16580 25366 16632 25372
rect 16304 25356 16356 25362
rect 16304 25298 16356 25304
rect 16316 24750 16344 25298
rect 16488 25288 16540 25294
rect 16488 25230 16540 25236
rect 16396 24812 16448 24818
rect 16396 24754 16448 24760
rect 16304 24744 16356 24750
rect 16304 24686 16356 24692
rect 16212 24676 16264 24682
rect 16212 24618 16264 24624
rect 16120 24608 16172 24614
rect 16120 24550 16172 24556
rect 16028 24064 16080 24070
rect 16028 24006 16080 24012
rect 15934 23760 15990 23769
rect 15934 23695 15990 23704
rect 15936 23656 15988 23662
rect 15934 23624 15936 23633
rect 15988 23624 15990 23633
rect 15934 23559 15990 23568
rect 15844 23248 15896 23254
rect 15844 23190 15896 23196
rect 15856 22438 15884 23190
rect 15936 23112 15988 23118
rect 15934 23080 15936 23089
rect 15988 23080 15990 23089
rect 16040 23066 16068 24006
rect 15990 23038 16068 23066
rect 15934 23015 15990 23024
rect 15936 22636 15988 22642
rect 15936 22578 15988 22584
rect 15844 22432 15896 22438
rect 15842 22400 15844 22409
rect 15896 22400 15898 22409
rect 15842 22335 15898 22344
rect 15844 22160 15896 22166
rect 15844 22102 15896 22108
rect 15856 22030 15884 22102
rect 15844 22024 15896 22030
rect 15844 21966 15896 21972
rect 15856 20641 15884 21966
rect 15948 21894 15976 22578
rect 16040 22166 16068 23038
rect 16132 22166 16160 24550
rect 16224 23662 16252 24618
rect 16304 24608 16356 24614
rect 16304 24550 16356 24556
rect 16316 23769 16344 24550
rect 16408 24070 16436 24754
rect 16500 24206 16528 25230
rect 16592 24750 16620 25366
rect 16764 25152 16816 25158
rect 16764 25094 16816 25100
rect 16580 24744 16632 24750
rect 16580 24686 16632 24692
rect 16672 24676 16724 24682
rect 16672 24618 16724 24624
rect 16488 24200 16540 24206
rect 16540 24160 16620 24188
rect 16488 24142 16540 24148
rect 16396 24064 16448 24070
rect 16396 24006 16448 24012
rect 16302 23760 16358 23769
rect 16302 23695 16358 23704
rect 16488 23724 16540 23730
rect 16488 23666 16540 23672
rect 16212 23656 16264 23662
rect 16212 23598 16264 23604
rect 16396 23656 16448 23662
rect 16396 23598 16448 23604
rect 16304 23588 16356 23594
rect 16304 23530 16356 23536
rect 16212 22976 16264 22982
rect 16212 22918 16264 22924
rect 16028 22160 16080 22166
rect 16028 22102 16080 22108
rect 16120 22160 16172 22166
rect 16120 22102 16172 22108
rect 16026 21992 16082 22001
rect 16026 21927 16082 21936
rect 15936 21888 15988 21894
rect 15936 21830 15988 21836
rect 15948 20942 15976 21830
rect 15936 20936 15988 20942
rect 15936 20878 15988 20884
rect 15842 20632 15898 20641
rect 15842 20567 15898 20576
rect 15948 20534 15976 20878
rect 15936 20528 15988 20534
rect 15936 20470 15988 20476
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 15856 19718 15884 20402
rect 15948 20398 15976 20470
rect 15936 20392 15988 20398
rect 15936 20334 15988 20340
rect 15936 20256 15988 20262
rect 15936 20198 15988 20204
rect 15844 19712 15896 19718
rect 15844 19654 15896 19660
rect 15856 19310 15884 19654
rect 15844 19304 15896 19310
rect 15844 19246 15896 19252
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15856 18834 15884 19110
rect 15844 18828 15896 18834
rect 15844 18770 15896 18776
rect 15948 18426 15976 20198
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 15856 17649 15884 18022
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 15842 17640 15898 17649
rect 15842 17575 15898 17584
rect 15948 16998 15976 17818
rect 15936 16992 15988 16998
rect 15936 16934 15988 16940
rect 15948 16289 15976 16934
rect 15934 16280 15990 16289
rect 15934 16215 15990 16224
rect 15936 15904 15988 15910
rect 15934 15872 15936 15881
rect 15988 15872 15990 15881
rect 15934 15807 15990 15816
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 15844 15632 15896 15638
rect 15844 15574 15896 15580
rect 15856 15094 15884 15574
rect 15844 15088 15896 15094
rect 15844 15030 15896 15036
rect 15844 14952 15896 14958
rect 15844 14894 15896 14900
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15658 12744 15714 12753
rect 15658 12679 15714 12688
rect 15672 11529 15700 12679
rect 15764 12374 15792 12922
rect 15856 12442 15884 14894
rect 15948 13530 15976 15642
rect 15936 13524 15988 13530
rect 15936 13466 15988 13472
rect 16040 13297 16068 21927
rect 16026 13288 16082 13297
rect 16026 13223 16082 13232
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 15752 12368 15804 12374
rect 15752 12310 15804 12316
rect 15934 12336 15990 12345
rect 15764 11937 15792 12310
rect 15934 12271 15990 12280
rect 15750 11928 15806 11937
rect 15750 11863 15806 11872
rect 15658 11520 15714 11529
rect 15658 11455 15714 11464
rect 15764 11354 15792 11863
rect 15948 11558 15976 12271
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 15660 11280 15712 11286
rect 15660 11222 15712 11228
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15566 10296 15622 10305
rect 15566 10231 15622 10240
rect 15580 8378 15608 10231
rect 15672 10198 15700 11222
rect 15750 11112 15806 11121
rect 15750 11047 15806 11056
rect 15764 10742 15792 11047
rect 15752 10736 15804 10742
rect 15752 10678 15804 10684
rect 15752 10532 15804 10538
rect 15752 10474 15804 10480
rect 15660 10192 15712 10198
rect 15660 10134 15712 10140
rect 15658 10024 15714 10033
rect 15658 9959 15714 9968
rect 15672 9178 15700 9959
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 15764 9058 15792 10474
rect 15844 10464 15896 10470
rect 15842 10432 15844 10441
rect 15896 10432 15898 10441
rect 15842 10367 15898 10376
rect 15764 9030 15884 9058
rect 15752 8968 15804 8974
rect 15750 8936 15752 8945
rect 15804 8936 15806 8945
rect 15750 8871 15806 8880
rect 15856 8634 15884 9030
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15580 8350 15884 8378
rect 15752 8288 15804 8294
rect 15752 8230 15804 8236
rect 15488 8078 15608 8106
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15488 7313 15516 7822
rect 15474 7304 15530 7313
rect 15474 7239 15530 7248
rect 15580 6458 15608 8078
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15672 7313 15700 8026
rect 15658 7304 15714 7313
rect 15658 7239 15714 7248
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 15672 6361 15700 7142
rect 15658 6352 15714 6361
rect 15658 6287 15714 6296
rect 15566 6216 15622 6225
rect 15566 6151 15622 6160
rect 15396 2944 15516 2972
rect 15292 2926 15344 2932
rect 14922 2887 14978 2896
rect 14936 2854 14964 2887
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 14476 2638 14872 2666
rect 14556 2576 14608 2582
rect 14554 2544 14556 2553
rect 14608 2544 14610 2553
rect 14554 2479 14610 2488
rect 14464 2440 14516 2446
rect 14462 2408 14464 2417
rect 14516 2408 14518 2417
rect 14462 2343 14518 2352
rect 14844 1986 14872 2638
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15304 2009 15332 2246
rect 15290 2000 15346 2009
rect 14844 1958 14964 1986
rect 14936 480 14964 1958
rect 15290 1935 15346 1944
rect 15488 480 15516 2944
rect 15580 2922 15608 6151
rect 15764 5846 15792 8230
rect 15752 5840 15804 5846
rect 15752 5782 15804 5788
rect 15764 5370 15792 5782
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15658 4856 15714 4865
rect 15856 4842 15884 8350
rect 15948 7993 15976 11494
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 16040 10033 16068 10746
rect 16026 10024 16082 10033
rect 16026 9959 16082 9968
rect 16026 9072 16082 9081
rect 16026 9007 16082 9016
rect 16040 8430 16068 9007
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 15934 7984 15990 7993
rect 15934 7919 15990 7928
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 16040 7585 16068 7890
rect 16026 7576 16082 7585
rect 16026 7511 16028 7520
rect 16080 7511 16082 7520
rect 16028 7482 16080 7488
rect 16026 7304 16082 7313
rect 16026 7239 16082 7248
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15948 6390 15976 6802
rect 15936 6384 15988 6390
rect 15936 6326 15988 6332
rect 16040 6186 16068 7239
rect 16028 6180 16080 6186
rect 16028 6122 16080 6128
rect 15936 6112 15988 6118
rect 15934 6080 15936 6089
rect 15988 6080 15990 6089
rect 15934 6015 15990 6024
rect 15856 4814 16068 4842
rect 15658 4791 15660 4800
rect 15712 4791 15714 4800
rect 15660 4762 15712 4768
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 15948 4214 15976 4558
rect 15936 4208 15988 4214
rect 15936 4150 15988 4156
rect 15948 3670 15976 4150
rect 15936 3664 15988 3670
rect 15936 3606 15988 3612
rect 15660 3392 15712 3398
rect 15660 3334 15712 3340
rect 15672 3194 15700 3334
rect 15948 3194 15976 3606
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 15568 2916 15620 2922
rect 15568 2858 15620 2864
rect 16040 480 16068 4814
rect 16132 921 16160 22102
rect 16224 17218 16252 22918
rect 16316 21865 16344 23530
rect 16408 22545 16436 23598
rect 16500 23202 16528 23666
rect 16592 23322 16620 24160
rect 16684 24070 16712 24618
rect 16776 24614 16804 25094
rect 17038 24848 17094 24857
rect 17038 24783 17094 24792
rect 16764 24608 16816 24614
rect 16764 24550 16816 24556
rect 16854 24576 16910 24585
rect 16672 24064 16724 24070
rect 16672 24006 16724 24012
rect 16776 23866 16804 24550
rect 16854 24511 16910 24520
rect 16868 24410 16896 24511
rect 16856 24404 16908 24410
rect 16856 24346 16908 24352
rect 16948 24268 17000 24274
rect 16948 24210 17000 24216
rect 16856 24064 16908 24070
rect 16856 24006 16908 24012
rect 16764 23860 16816 23866
rect 16764 23802 16816 23808
rect 16580 23316 16632 23322
rect 16580 23258 16632 23264
rect 16868 23225 16896 24006
rect 16960 23526 16988 24210
rect 17052 23798 17080 24783
rect 17144 24041 17172 25486
rect 17130 24032 17186 24041
rect 17130 23967 17186 23976
rect 17040 23792 17092 23798
rect 17040 23734 17092 23740
rect 17144 23662 17172 23967
rect 17132 23656 17184 23662
rect 17132 23598 17184 23604
rect 16948 23520 17000 23526
rect 16948 23462 17000 23468
rect 16854 23216 16910 23225
rect 16500 23174 16712 23202
rect 16394 22536 16450 22545
rect 16394 22471 16450 22480
rect 16580 22500 16632 22506
rect 16580 22442 16632 22448
rect 16396 22432 16448 22438
rect 16396 22374 16448 22380
rect 16408 22234 16436 22374
rect 16396 22228 16448 22234
rect 16396 22170 16448 22176
rect 16302 21856 16358 21865
rect 16302 21791 16358 21800
rect 16302 21720 16358 21729
rect 16302 21655 16358 21664
rect 16316 20482 16344 21655
rect 16408 21321 16436 22170
rect 16592 21457 16620 22442
rect 16578 21448 16634 21457
rect 16578 21383 16634 21392
rect 16684 21350 16712 23174
rect 16854 23151 16910 23160
rect 16764 22092 16816 22098
rect 16764 22034 16816 22040
rect 16856 22092 16908 22098
rect 16856 22034 16908 22040
rect 16776 21622 16804 22034
rect 16764 21616 16816 21622
rect 16764 21558 16816 21564
rect 16764 21412 16816 21418
rect 16764 21354 16816 21360
rect 16672 21344 16724 21350
rect 16394 21312 16450 21321
rect 16672 21286 16724 21292
rect 16394 21247 16450 21256
rect 16396 21140 16448 21146
rect 16396 21082 16448 21088
rect 16408 20777 16436 21082
rect 16580 21004 16632 21010
rect 16580 20946 16632 20952
rect 16592 20890 16620 20946
rect 16500 20862 16620 20890
rect 16394 20768 16450 20777
rect 16394 20703 16450 20712
rect 16500 20602 16528 20862
rect 16488 20596 16540 20602
rect 16488 20538 16540 20544
rect 16316 20454 16528 20482
rect 16396 20392 16448 20398
rect 16396 20334 16448 20340
rect 16408 19922 16436 20334
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 16408 19514 16436 19858
rect 16396 19508 16448 19514
rect 16396 19450 16448 19456
rect 16302 19272 16358 19281
rect 16302 19207 16358 19216
rect 16316 18970 16344 19207
rect 16408 18970 16436 19450
rect 16304 18964 16356 18970
rect 16304 18906 16356 18912
rect 16396 18964 16448 18970
rect 16500 18952 16528 20454
rect 16776 20346 16804 21354
rect 16684 20318 16804 20346
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 16592 19310 16620 19994
rect 16684 19417 16712 20318
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16776 19990 16804 20198
rect 16764 19984 16816 19990
rect 16764 19926 16816 19932
rect 16776 19514 16804 19926
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16670 19408 16726 19417
rect 16670 19343 16726 19352
rect 16580 19304 16632 19310
rect 16868 19258 16896 22034
rect 16580 19246 16632 19252
rect 16684 19230 16896 19258
rect 16500 18924 16620 18952
rect 16396 18906 16448 18912
rect 16304 18624 16356 18630
rect 16304 18566 16356 18572
rect 16316 18193 16344 18566
rect 16302 18184 16358 18193
rect 16302 18119 16358 18128
rect 16408 17882 16436 18906
rect 16486 18864 16542 18873
rect 16486 18799 16542 18808
rect 16500 18766 16528 18799
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16592 18612 16620 18924
rect 16500 18584 16620 18612
rect 16396 17876 16448 17882
rect 16396 17818 16448 17824
rect 16500 17610 16528 18584
rect 16580 18352 16632 18358
rect 16580 18294 16632 18300
rect 16592 18193 16620 18294
rect 16578 18184 16634 18193
rect 16578 18119 16634 18128
rect 16592 18086 16620 18119
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16224 17190 16528 17218
rect 16394 16688 16450 16697
rect 16304 16652 16356 16658
rect 16224 16612 16304 16640
rect 16224 16182 16252 16612
rect 16394 16623 16450 16632
rect 16304 16594 16356 16600
rect 16304 16244 16356 16250
rect 16304 16186 16356 16192
rect 16212 16176 16264 16182
rect 16212 16118 16264 16124
rect 16212 15972 16264 15978
rect 16212 15914 16264 15920
rect 16224 15706 16252 15914
rect 16212 15700 16264 15706
rect 16212 15642 16264 15648
rect 16210 15600 16266 15609
rect 16210 15535 16212 15544
rect 16264 15535 16266 15544
rect 16212 15506 16264 15512
rect 16224 15026 16252 15506
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 16212 14884 16264 14890
rect 16212 14826 16264 14832
rect 16224 12918 16252 14826
rect 16212 12912 16264 12918
rect 16212 12854 16264 12860
rect 16224 12646 16252 12854
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 16224 9518 16252 12378
rect 16316 10810 16344 16186
rect 16408 15502 16436 16623
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16396 15088 16448 15094
rect 16396 15030 16448 15036
rect 16408 14929 16436 15030
rect 16394 14920 16450 14929
rect 16394 14855 16450 14864
rect 16394 14512 16450 14521
rect 16394 14447 16450 14456
rect 16408 14074 16436 14447
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16396 13796 16448 13802
rect 16396 13738 16448 13744
rect 16408 13394 16436 13738
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16408 12782 16436 13330
rect 16396 12776 16448 12782
rect 16396 12718 16448 12724
rect 16396 12640 16448 12646
rect 16396 12582 16448 12588
rect 16408 12209 16436 12582
rect 16394 12200 16450 12209
rect 16394 12135 16450 12144
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16408 11898 16436 12038
rect 16396 11892 16448 11898
rect 16396 11834 16448 11840
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16408 10305 16436 10406
rect 16394 10296 16450 10305
rect 16394 10231 16450 10240
rect 16500 9704 16528 17190
rect 16580 17060 16632 17066
rect 16580 17002 16632 17008
rect 16592 16794 16620 17002
rect 16580 16788 16632 16794
rect 16580 16730 16632 16736
rect 16580 15564 16632 15570
rect 16580 15506 16632 15512
rect 16592 15162 16620 15506
rect 16580 15156 16632 15162
rect 16580 15098 16632 15104
rect 16592 12850 16620 15098
rect 16684 14634 16712 19230
rect 16856 19168 16908 19174
rect 16856 19110 16908 19116
rect 16764 18964 16816 18970
rect 16764 18906 16816 18912
rect 16776 18290 16804 18906
rect 16868 18834 16896 19110
rect 16856 18828 16908 18834
rect 16856 18770 16908 18776
rect 16764 18284 16816 18290
rect 16764 18226 16816 18232
rect 16868 17882 16896 18770
rect 16856 17876 16908 17882
rect 16856 17818 16908 17824
rect 16764 17536 16816 17542
rect 16764 17478 16816 17484
rect 16776 16454 16804 17478
rect 16960 17241 16988 23462
rect 17236 23322 17264 25706
rect 17316 25356 17368 25362
rect 17316 25298 17368 25304
rect 17328 24614 17356 25298
rect 17592 24744 17644 24750
rect 17788 24698 17816 27520
rect 17866 26344 17922 26353
rect 17866 26279 17922 26288
rect 17880 25158 17908 26279
rect 18144 26172 18196 26178
rect 18144 26114 18196 26120
rect 17868 25152 17920 25158
rect 17868 25094 17920 25100
rect 18050 24984 18106 24993
rect 18050 24919 18106 24928
rect 17592 24686 17644 24692
rect 17316 24608 17368 24614
rect 17316 24550 17368 24556
rect 17224 23316 17276 23322
rect 17224 23258 17276 23264
rect 17132 23180 17184 23186
rect 17132 23122 17184 23128
rect 17144 22438 17172 23122
rect 17236 22778 17264 23258
rect 17224 22772 17276 22778
rect 17224 22714 17276 22720
rect 17224 22636 17276 22642
rect 17224 22578 17276 22584
rect 17132 22432 17184 22438
rect 17130 22400 17132 22409
rect 17184 22400 17186 22409
rect 17130 22335 17186 22344
rect 17132 21616 17184 21622
rect 17130 21584 17132 21593
rect 17184 21584 17186 21593
rect 17130 21519 17186 21528
rect 17132 21344 17184 21350
rect 17132 21286 17184 21292
rect 17040 20936 17092 20942
rect 17040 20878 17092 20884
rect 17052 20505 17080 20878
rect 17038 20496 17094 20505
rect 17038 20431 17094 20440
rect 17144 20346 17172 21286
rect 17052 20318 17172 20346
rect 16946 17232 17002 17241
rect 16946 17167 17002 17176
rect 17052 17116 17080 20318
rect 17132 18080 17184 18086
rect 17132 18022 17184 18028
rect 16868 17088 17080 17116
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16776 16289 16804 16390
rect 16762 16280 16818 16289
rect 16762 16215 16818 16224
rect 16762 15056 16818 15065
rect 16762 14991 16764 15000
rect 16816 14991 16818 15000
rect 16764 14962 16816 14968
rect 16764 14884 16816 14890
rect 16764 14826 16816 14832
rect 16776 14793 16804 14826
rect 16762 14784 16818 14793
rect 16762 14719 16818 14728
rect 16684 14606 16804 14634
rect 16672 14476 16724 14482
rect 16672 14418 16724 14424
rect 16684 13802 16712 14418
rect 16672 13796 16724 13802
rect 16672 13738 16724 13744
rect 16670 13560 16726 13569
rect 16670 13495 16726 13504
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16684 12714 16712 13495
rect 16580 12708 16632 12714
rect 16580 12650 16632 12656
rect 16672 12708 16724 12714
rect 16672 12650 16724 12656
rect 16592 12442 16620 12650
rect 16776 12594 16804 14606
rect 16868 14482 16896 17088
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 17052 16250 17080 16594
rect 17040 16244 17092 16250
rect 17040 16186 17092 16192
rect 17144 16130 17172 18022
rect 17052 16102 17172 16130
rect 16948 15360 17000 15366
rect 16948 15302 17000 15308
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16868 13530 16896 13806
rect 16960 13802 16988 15302
rect 17052 15162 17080 16102
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 17144 15745 17172 15846
rect 17130 15736 17186 15745
rect 17130 15671 17186 15680
rect 17040 15156 17092 15162
rect 17040 15098 17092 15104
rect 17132 15020 17184 15026
rect 17132 14962 17184 14968
rect 17144 14550 17172 14962
rect 17132 14544 17184 14550
rect 17132 14486 17184 14492
rect 17040 14476 17092 14482
rect 17040 14418 17092 14424
rect 16948 13796 17000 13802
rect 16948 13738 17000 13744
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 16856 13252 16908 13258
rect 16856 13194 16908 13200
rect 16684 12566 16804 12594
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16592 10282 16620 12174
rect 16684 10470 16712 12566
rect 16762 12336 16818 12345
rect 16762 12271 16818 12280
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16592 10254 16712 10282
rect 16580 10192 16632 10198
rect 16580 10134 16632 10140
rect 16316 9676 16528 9704
rect 16212 9512 16264 9518
rect 16212 9454 16264 9460
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16224 8090 16252 9114
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 16210 7576 16266 7585
rect 16210 7511 16266 7520
rect 16224 7002 16252 7511
rect 16212 6996 16264 7002
rect 16212 6938 16264 6944
rect 16224 4842 16252 6938
rect 16316 6769 16344 9676
rect 16592 9602 16620 10134
rect 16684 10044 16712 10254
rect 16776 10198 16804 12271
rect 16868 11286 16896 13194
rect 16960 12986 16988 13738
rect 17052 13530 17080 14418
rect 17144 13938 17172 14486
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17130 13832 17186 13841
rect 17130 13767 17132 13776
rect 17184 13767 17186 13776
rect 17132 13738 17184 13744
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 17038 13424 17094 13433
rect 17144 13394 17172 13738
rect 17038 13359 17094 13368
rect 17132 13388 17184 13394
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 16948 12708 17000 12714
rect 16948 12650 17000 12656
rect 16960 12442 16988 12650
rect 17052 12481 17080 13359
rect 17132 13330 17184 13336
rect 17144 12986 17172 13330
rect 17236 13297 17264 22578
rect 17328 21593 17356 24550
rect 17408 24336 17460 24342
rect 17408 24278 17460 24284
rect 17420 23798 17448 24278
rect 17604 23798 17632 24686
rect 17696 24670 17816 24698
rect 17696 24313 17724 24670
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17682 24304 17738 24313
rect 17682 24239 17738 24248
rect 17408 23792 17460 23798
rect 17408 23734 17460 23740
rect 17592 23792 17644 23798
rect 17592 23734 17644 23740
rect 17408 23112 17460 23118
rect 17408 23054 17460 23060
rect 17314 21584 17370 21593
rect 17314 21519 17370 21528
rect 17420 21026 17448 23054
rect 17592 22976 17644 22982
rect 17592 22918 17644 22924
rect 17500 22432 17552 22438
rect 17500 22374 17552 22380
rect 17512 21418 17540 22374
rect 17500 21412 17552 21418
rect 17500 21354 17552 21360
rect 17420 20998 17540 21026
rect 17408 20936 17460 20942
rect 17408 20878 17460 20884
rect 17316 20800 17368 20806
rect 17316 20742 17368 20748
rect 17328 20466 17356 20742
rect 17316 20460 17368 20466
rect 17316 20402 17368 20408
rect 17420 20262 17448 20878
rect 17408 20256 17460 20262
rect 17408 20198 17460 20204
rect 17420 19174 17448 20198
rect 17408 19168 17460 19174
rect 17408 19110 17460 19116
rect 17408 18624 17460 18630
rect 17408 18566 17460 18572
rect 17316 18148 17368 18154
rect 17316 18090 17368 18096
rect 17222 13288 17278 13297
rect 17222 13223 17278 13232
rect 17224 13184 17276 13190
rect 17224 13126 17276 13132
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 17038 12472 17094 12481
rect 16948 12436 17000 12442
rect 17038 12407 17094 12416
rect 16948 12378 17000 12384
rect 17040 12368 17092 12374
rect 17040 12310 17092 12316
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 16856 11280 16908 11286
rect 16856 11222 16908 11228
rect 16856 11076 16908 11082
rect 16960 11064 16988 11698
rect 17052 11354 17080 12310
rect 17130 11928 17186 11937
rect 17130 11863 17186 11872
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 16908 11036 16988 11064
rect 16856 11018 16908 11024
rect 16764 10192 16816 10198
rect 16764 10134 16816 10140
rect 16684 10016 16804 10044
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 16684 9722 16712 9862
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 16500 9586 16620 9602
rect 16488 9580 16620 9586
rect 16540 9574 16620 9580
rect 16488 9522 16540 9528
rect 16488 9444 16540 9450
rect 16488 9386 16540 9392
rect 16500 9178 16528 9386
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16408 8838 16436 8869
rect 16396 8832 16448 8838
rect 16394 8800 16396 8809
rect 16448 8800 16450 8809
rect 16394 8735 16450 8744
rect 16408 7342 16436 8735
rect 16396 7336 16448 7342
rect 16396 7278 16448 7284
rect 16500 6866 16528 9114
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 16302 6760 16358 6769
rect 16302 6695 16358 6704
rect 16488 6724 16540 6730
rect 16488 6666 16540 6672
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 16316 6322 16344 6598
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16500 5370 16528 6666
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 16224 4814 16436 4842
rect 16212 4684 16264 4690
rect 16212 4626 16264 4632
rect 16224 3126 16252 4626
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16212 3120 16264 3126
rect 16212 3062 16264 3068
rect 16316 2990 16344 3878
rect 16408 3602 16436 4814
rect 16488 4684 16540 4690
rect 16488 4626 16540 4632
rect 16396 3596 16448 3602
rect 16396 3538 16448 3544
rect 16394 3496 16450 3505
rect 16394 3431 16450 3440
rect 16304 2984 16356 2990
rect 16304 2926 16356 2932
rect 16408 2650 16436 3431
rect 16500 2990 16528 4626
rect 16488 2984 16540 2990
rect 16488 2926 16540 2932
rect 16592 2825 16620 9318
rect 16776 7392 16804 10016
rect 16868 9586 16896 11018
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16856 9580 16908 9586
rect 16856 9522 16908 9528
rect 16868 9178 16896 9522
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 16960 9042 16988 10406
rect 17052 10062 17080 10610
rect 17040 10056 17092 10062
rect 17040 9998 17092 10004
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 17144 8106 17172 11863
rect 17236 8974 17264 13126
rect 17328 12646 17356 18090
rect 17420 17882 17448 18566
rect 17408 17876 17460 17882
rect 17408 17818 17460 17824
rect 17408 17740 17460 17746
rect 17408 17682 17460 17688
rect 17420 17202 17448 17682
rect 17408 17196 17460 17202
rect 17408 17138 17460 17144
rect 17420 16794 17448 17138
rect 17408 16788 17460 16794
rect 17408 16730 17460 16736
rect 17408 15020 17460 15026
rect 17408 14962 17460 14968
rect 17420 14550 17448 14962
rect 17408 14544 17460 14550
rect 17408 14486 17460 14492
rect 17420 14074 17448 14486
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17314 12472 17370 12481
rect 17314 12407 17316 12416
rect 17368 12407 17370 12416
rect 17316 12378 17368 12384
rect 17420 11801 17448 13466
rect 17512 12424 17540 20998
rect 17604 17241 17632 22918
rect 17684 22772 17736 22778
rect 17684 22714 17736 22720
rect 17696 22098 17724 22714
rect 17684 22092 17736 22098
rect 17684 22034 17736 22040
rect 17684 21956 17736 21962
rect 17684 21898 17736 21904
rect 17696 21026 17724 21898
rect 17788 21146 17816 24550
rect 18064 24410 18092 24919
rect 18052 24404 18104 24410
rect 18052 24346 18104 24352
rect 18050 24304 18106 24313
rect 18050 24239 18106 24248
rect 17960 23724 18012 23730
rect 17960 23666 18012 23672
rect 17868 23248 17920 23254
rect 17868 23190 17920 23196
rect 17880 22166 17908 23190
rect 17868 22160 17920 22166
rect 17868 22102 17920 22108
rect 17868 22024 17920 22030
rect 17868 21966 17920 21972
rect 17880 21350 17908 21966
rect 17868 21344 17920 21350
rect 17868 21286 17920 21292
rect 17776 21140 17828 21146
rect 17776 21082 17828 21088
rect 17696 20998 17816 21026
rect 17684 19168 17736 19174
rect 17682 19136 17684 19145
rect 17736 19136 17738 19145
rect 17682 19071 17738 19080
rect 17684 18964 17736 18970
rect 17684 18906 17736 18912
rect 17696 18426 17724 18906
rect 17684 18420 17736 18426
rect 17684 18362 17736 18368
rect 17682 17776 17738 17785
rect 17682 17711 17738 17720
rect 17590 17232 17646 17241
rect 17590 17167 17646 17176
rect 17696 17066 17724 17711
rect 17684 17060 17736 17066
rect 17684 17002 17736 17008
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17604 14618 17632 15982
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17696 15026 17724 15438
rect 17684 15020 17736 15026
rect 17684 14962 17736 14968
rect 17684 14884 17736 14890
rect 17684 14826 17736 14832
rect 17592 14612 17644 14618
rect 17592 14554 17644 14560
rect 17604 13530 17632 14554
rect 17592 13524 17644 13530
rect 17592 13466 17644 13472
rect 17590 13424 17646 13433
rect 17590 13359 17646 13368
rect 17604 13258 17632 13359
rect 17592 13252 17644 13258
rect 17592 13194 17644 13200
rect 17696 12986 17724 14826
rect 17684 12980 17736 12986
rect 17684 12922 17736 12928
rect 17788 12764 17816 20998
rect 17880 20641 17908 21286
rect 17866 20632 17922 20641
rect 17866 20567 17922 20576
rect 17868 20528 17920 20534
rect 17866 20496 17868 20505
rect 17920 20496 17922 20505
rect 17866 20431 17922 20440
rect 17868 20256 17920 20262
rect 17868 20198 17920 20204
rect 17880 19825 17908 20198
rect 17866 19816 17922 19825
rect 17866 19751 17922 19760
rect 17972 18426 18000 23666
rect 18064 21894 18092 24239
rect 18156 23662 18184 26114
rect 18340 25702 18368 27520
rect 18892 26110 18920 27520
rect 19536 26246 19564 27520
rect 19524 26240 19576 26246
rect 19524 26182 19576 26188
rect 18880 26104 18932 26110
rect 18880 26046 18932 26052
rect 19524 25832 19576 25838
rect 19524 25774 19576 25780
rect 19156 25764 19208 25770
rect 19156 25706 19208 25712
rect 18328 25696 18380 25702
rect 18328 25638 18380 25644
rect 19064 25356 19116 25362
rect 19064 25298 19116 25304
rect 18420 25220 18472 25226
rect 18420 25162 18472 25168
rect 18328 23792 18380 23798
rect 18328 23734 18380 23740
rect 18144 23656 18196 23662
rect 18144 23598 18196 23604
rect 18156 23322 18184 23598
rect 18144 23316 18196 23322
rect 18144 23258 18196 23264
rect 18156 23202 18184 23258
rect 18156 23174 18276 23202
rect 18142 23080 18198 23089
rect 18142 23015 18198 23024
rect 18156 22710 18184 23015
rect 18144 22704 18196 22710
rect 18144 22646 18196 22652
rect 18248 22642 18276 23174
rect 18340 22642 18368 23734
rect 18432 23508 18460 25162
rect 19076 24614 19104 25298
rect 19064 24608 19116 24614
rect 19064 24550 19116 24556
rect 19076 24449 19104 24550
rect 19062 24440 19118 24449
rect 18512 24404 18564 24410
rect 19168 24410 19196 25706
rect 19062 24375 19118 24384
rect 19156 24404 19208 24410
rect 18512 24346 18564 24352
rect 19156 24346 19208 24352
rect 19340 24404 19392 24410
rect 19340 24346 19392 24352
rect 18524 23662 18552 24346
rect 19156 24268 19208 24274
rect 19156 24210 19208 24216
rect 18604 24200 18656 24206
rect 18604 24142 18656 24148
rect 19064 24200 19116 24206
rect 19064 24142 19116 24148
rect 18616 23730 18644 24142
rect 18604 23724 18656 23730
rect 18656 23684 18736 23712
rect 18604 23666 18656 23672
rect 18512 23656 18564 23662
rect 18512 23598 18564 23604
rect 18432 23480 18552 23508
rect 18418 23352 18474 23361
rect 18418 23287 18420 23296
rect 18472 23287 18474 23296
rect 18420 23258 18472 23264
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 18328 22636 18380 22642
rect 18328 22578 18380 22584
rect 18144 22568 18196 22574
rect 18144 22510 18196 22516
rect 18234 22536 18290 22545
rect 18156 22137 18184 22510
rect 18234 22471 18290 22480
rect 18142 22128 18198 22137
rect 18142 22063 18198 22072
rect 18248 21962 18276 22471
rect 18328 22432 18380 22438
rect 18328 22374 18380 22380
rect 18418 22400 18474 22409
rect 18236 21956 18288 21962
rect 18236 21898 18288 21904
rect 18052 21888 18104 21894
rect 18052 21830 18104 21836
rect 18052 21344 18104 21350
rect 18052 21286 18104 21292
rect 18142 21312 18198 21321
rect 18064 21185 18092 21286
rect 18142 21247 18198 21256
rect 18050 21176 18106 21185
rect 18156 21146 18184 21247
rect 18050 21111 18106 21120
rect 18144 21140 18196 21146
rect 18144 21082 18196 21088
rect 18234 21040 18290 21049
rect 18234 20975 18290 20984
rect 18144 20936 18196 20942
rect 18064 20884 18144 20890
rect 18064 20878 18196 20884
rect 18064 20862 18184 20878
rect 18064 19700 18092 20862
rect 18144 20528 18196 20534
rect 18144 20470 18196 20476
rect 18156 20233 18184 20470
rect 18142 20224 18198 20233
rect 18142 20159 18198 20168
rect 18248 20058 18276 20975
rect 18236 20052 18288 20058
rect 18236 19994 18288 20000
rect 18236 19712 18288 19718
rect 18064 19680 18236 19700
rect 18288 19680 18290 19689
rect 18064 19672 18234 19680
rect 18234 19615 18290 19624
rect 18236 19236 18288 19242
rect 18236 19178 18288 19184
rect 18144 18624 18196 18630
rect 18144 18566 18196 18572
rect 17960 18420 18012 18426
rect 17960 18362 18012 18368
rect 17866 18184 17922 18193
rect 17866 18119 17922 18128
rect 17880 16794 17908 18119
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 17868 16788 17920 16794
rect 17868 16730 17920 16736
rect 17972 16504 18000 17818
rect 18050 17504 18106 17513
rect 18050 17439 18106 17448
rect 18064 17338 18092 17439
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 18050 17232 18106 17241
rect 18050 17167 18106 17176
rect 18064 17134 18092 17167
rect 18052 17128 18104 17134
rect 18052 17070 18104 17076
rect 18064 16658 18092 17070
rect 18156 16697 18184 18566
rect 18142 16688 18198 16697
rect 18052 16652 18104 16658
rect 18142 16623 18198 16632
rect 18052 16594 18104 16600
rect 17880 16476 18000 16504
rect 17880 16250 17908 16476
rect 17958 16416 18014 16425
rect 17958 16351 18014 16360
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 17868 15564 17920 15570
rect 17972 15552 18000 16351
rect 18064 16182 18092 16594
rect 18052 16176 18104 16182
rect 18052 16118 18104 16124
rect 18052 15904 18104 15910
rect 18052 15846 18104 15852
rect 17920 15524 18000 15552
rect 17868 15506 17920 15512
rect 17880 15094 17908 15506
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 17868 15088 17920 15094
rect 17868 15030 17920 15036
rect 17972 14890 18000 15370
rect 18064 15337 18092 15846
rect 18050 15328 18106 15337
rect 18248 15314 18276 19178
rect 18050 15263 18106 15272
rect 18156 15286 18276 15314
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 17960 14884 18012 14890
rect 17960 14826 18012 14832
rect 17868 14816 17920 14822
rect 17868 14758 17920 14764
rect 17880 13870 17908 14758
rect 18064 14657 18092 14894
rect 18050 14648 18106 14657
rect 18050 14583 18106 14592
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 18064 13870 18092 14214
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 17958 13560 18014 13569
rect 17958 13495 18014 13504
rect 17972 13462 18000 13495
rect 17960 13456 18012 13462
rect 17960 13398 18012 13404
rect 18064 13394 18092 13806
rect 18052 13388 18104 13394
rect 18052 13330 18104 13336
rect 17958 12880 18014 12889
rect 17958 12815 18014 12824
rect 17788 12736 17908 12764
rect 17684 12708 17736 12714
rect 17684 12650 17736 12656
rect 17512 12396 17632 12424
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17512 11898 17540 12242
rect 17604 12238 17632 12396
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 17592 12096 17644 12102
rect 17592 12038 17644 12044
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17406 11792 17462 11801
rect 17462 11750 17540 11778
rect 17406 11727 17462 11736
rect 17316 11552 17368 11558
rect 17314 11520 17316 11529
rect 17368 11520 17370 11529
rect 17314 11455 17370 11464
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 17052 8078 17172 8106
rect 17052 7546 17080 8078
rect 17132 8016 17184 8022
rect 17130 7984 17132 7993
rect 17184 7984 17186 7993
rect 17130 7919 17186 7928
rect 17040 7540 17092 7546
rect 17040 7482 17092 7488
rect 16684 7364 16804 7392
rect 16684 5914 16712 7364
rect 16762 7304 16818 7313
rect 16762 7239 16764 7248
rect 16816 7239 16818 7248
rect 16764 7210 16816 7216
rect 16854 7032 16910 7041
rect 16854 6967 16910 6976
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 16684 3369 16712 5850
rect 16868 5370 16896 6967
rect 17236 6866 17264 8774
rect 17328 8294 17356 11290
rect 17408 11076 17460 11082
rect 17408 11018 17460 11024
rect 17420 8673 17448 11018
rect 17512 10606 17540 11750
rect 17500 10600 17552 10606
rect 17500 10542 17552 10548
rect 17512 10169 17540 10542
rect 17498 10160 17554 10169
rect 17498 10095 17554 10104
rect 17498 9208 17554 9217
rect 17498 9143 17500 9152
rect 17552 9143 17554 9152
rect 17500 9114 17552 9120
rect 17406 8664 17462 8673
rect 17512 8634 17540 9114
rect 17406 8599 17462 8608
rect 17500 8628 17552 8634
rect 17420 8430 17448 8599
rect 17500 8570 17552 8576
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 17316 8288 17368 8294
rect 17316 8230 17368 8236
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 17316 7880 17368 7886
rect 17420 7857 17448 7890
rect 17316 7822 17368 7828
rect 17406 7848 17462 7857
rect 17328 7274 17356 7822
rect 17406 7783 17462 7792
rect 17316 7268 17368 7274
rect 17316 7210 17368 7216
rect 17420 7002 17448 7783
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 17236 6769 17264 6802
rect 17038 6760 17094 6769
rect 17038 6695 17094 6704
rect 17222 6760 17278 6769
rect 17222 6695 17278 6704
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 16868 4146 16896 5306
rect 17052 5273 17080 6695
rect 17408 6656 17460 6662
rect 17406 6624 17408 6633
rect 17460 6624 17462 6633
rect 17406 6559 17462 6568
rect 17132 6384 17184 6390
rect 17132 6326 17184 6332
rect 17144 5914 17172 6326
rect 17132 5908 17184 5914
rect 17132 5850 17184 5856
rect 17038 5264 17094 5273
rect 17038 5199 17094 5208
rect 17316 4752 17368 4758
rect 17316 4694 17368 4700
rect 17406 4720 17462 4729
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16776 3738 16804 3878
rect 16764 3732 16816 3738
rect 16764 3674 16816 3680
rect 16764 3596 16816 3602
rect 16764 3538 16816 3544
rect 16670 3360 16726 3369
rect 16670 3295 16726 3304
rect 16776 3176 16804 3538
rect 16856 3528 16908 3534
rect 16854 3496 16856 3505
rect 17052 3505 17080 4422
rect 17328 4185 17356 4694
rect 17406 4655 17462 4664
rect 17420 4622 17448 4655
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17420 4282 17448 4558
rect 17408 4276 17460 4282
rect 17408 4218 17460 4224
rect 17314 4176 17370 4185
rect 17314 4111 17370 4120
rect 17328 3670 17356 4111
rect 17604 4049 17632 12038
rect 17696 11257 17724 12650
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17682 11248 17738 11257
rect 17682 11183 17738 11192
rect 17788 11082 17816 12174
rect 17776 11076 17828 11082
rect 17776 11018 17828 11024
rect 17682 10976 17738 10985
rect 17682 10911 17738 10920
rect 17696 9466 17724 10911
rect 17788 10713 17816 11018
rect 17774 10704 17830 10713
rect 17774 10639 17830 10648
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17788 9654 17816 10066
rect 17776 9648 17828 9654
rect 17776 9590 17828 9596
rect 17696 9438 17816 9466
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17696 8634 17724 8910
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 17788 7002 17816 9438
rect 17880 9081 17908 12736
rect 17972 12481 18000 12815
rect 17958 12472 18014 12481
rect 17958 12407 18014 12416
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 17972 11762 18000 12038
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17960 11620 18012 11626
rect 17960 11562 18012 11568
rect 17972 11150 18000 11562
rect 18052 11212 18104 11218
rect 18052 11154 18104 11160
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 17972 9897 18000 11086
rect 18064 10985 18092 11154
rect 18156 11014 18184 15286
rect 18234 15192 18290 15201
rect 18234 15127 18290 15136
rect 18248 13977 18276 15127
rect 18234 13968 18290 13977
rect 18234 13903 18290 13912
rect 18248 13326 18276 13903
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 18236 11212 18288 11218
rect 18236 11154 18288 11160
rect 18144 11008 18196 11014
rect 18050 10976 18106 10985
rect 18144 10950 18196 10956
rect 18050 10911 18106 10920
rect 18050 10840 18106 10849
rect 18248 10810 18276 11154
rect 18050 10775 18106 10784
rect 18236 10804 18288 10810
rect 18064 10266 18092 10775
rect 18236 10746 18288 10752
rect 18142 10704 18198 10713
rect 18142 10639 18198 10648
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 17958 9888 18014 9897
rect 17958 9823 18014 9832
rect 18064 9722 18092 10202
rect 18052 9716 18104 9722
rect 18052 9658 18104 9664
rect 18156 9450 18184 10639
rect 18340 10282 18368 22374
rect 18418 22335 18474 22344
rect 18432 22166 18460 22335
rect 18420 22160 18472 22166
rect 18420 22102 18472 22108
rect 18420 21888 18472 21894
rect 18420 21830 18472 21836
rect 18432 21350 18460 21830
rect 18524 21570 18552 23480
rect 18602 23488 18658 23497
rect 18602 23423 18658 23432
rect 18616 22420 18644 23423
rect 18708 23322 18736 23684
rect 18788 23656 18840 23662
rect 18788 23598 18840 23604
rect 18696 23316 18748 23322
rect 18696 23258 18748 23264
rect 18696 23180 18748 23186
rect 18696 23122 18748 23128
rect 18708 22574 18736 23122
rect 18696 22568 18748 22574
rect 18696 22510 18748 22516
rect 18616 22392 18736 22420
rect 18604 22160 18656 22166
rect 18604 22102 18656 22108
rect 18616 21690 18644 22102
rect 18708 22030 18736 22392
rect 18696 22024 18748 22030
rect 18696 21966 18748 21972
rect 18604 21684 18656 21690
rect 18604 21626 18656 21632
rect 18708 21622 18736 21966
rect 18696 21616 18748 21622
rect 18524 21542 18644 21570
rect 18696 21558 18748 21564
rect 18510 21448 18566 21457
rect 18510 21383 18566 21392
rect 18420 21344 18472 21350
rect 18420 21286 18472 21292
rect 18432 21049 18460 21286
rect 18418 21040 18474 21049
rect 18418 20975 18474 20984
rect 18418 20768 18474 20777
rect 18418 20703 18474 20712
rect 18432 20398 18460 20703
rect 18524 20398 18552 21383
rect 18420 20392 18472 20398
rect 18420 20334 18472 20340
rect 18512 20392 18564 20398
rect 18512 20334 18564 20340
rect 18616 20244 18644 21542
rect 18696 21004 18748 21010
rect 18696 20946 18748 20952
rect 18432 20216 18644 20244
rect 18432 16810 18460 20216
rect 18512 19916 18564 19922
rect 18512 19858 18564 19864
rect 18524 18630 18552 19858
rect 18708 19825 18736 20946
rect 18694 19816 18750 19825
rect 18694 19751 18750 19760
rect 18604 19168 18656 19174
rect 18604 19110 18656 19116
rect 18512 18624 18564 18630
rect 18616 18601 18644 19110
rect 18512 18566 18564 18572
rect 18602 18592 18658 18601
rect 18524 18329 18552 18566
rect 18602 18527 18658 18536
rect 18510 18320 18566 18329
rect 18694 18320 18750 18329
rect 18510 18255 18566 18264
rect 18616 18278 18694 18306
rect 18512 17808 18564 17814
rect 18512 17750 18564 17756
rect 18524 17241 18552 17750
rect 18510 17232 18566 17241
rect 18510 17167 18566 17176
rect 18512 17128 18564 17134
rect 18512 17070 18564 17076
rect 18524 16969 18552 17070
rect 18616 17066 18644 18278
rect 18694 18255 18750 18264
rect 18694 17640 18750 17649
rect 18694 17575 18750 17584
rect 18708 17202 18736 17575
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 18604 17060 18656 17066
rect 18604 17002 18656 17008
rect 18510 16960 18566 16969
rect 18510 16895 18566 16904
rect 18616 16833 18644 17002
rect 18602 16824 18658 16833
rect 18432 16782 18552 16810
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18432 16046 18460 16390
rect 18420 16040 18472 16046
rect 18418 16008 18420 16017
rect 18472 16008 18474 16017
rect 18418 15943 18474 15952
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18432 12714 18460 15098
rect 18524 13297 18552 16782
rect 18602 16759 18658 16768
rect 18604 16176 18656 16182
rect 18604 16118 18656 16124
rect 18616 15502 18644 16118
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 18708 15570 18736 16050
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 18604 15496 18656 15502
rect 18604 15438 18656 15444
rect 18696 14476 18748 14482
rect 18696 14418 18748 14424
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 18616 13870 18644 14214
rect 18604 13864 18656 13870
rect 18604 13806 18656 13812
rect 18708 13734 18736 14418
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 18510 13288 18566 13297
rect 18510 13223 18566 13232
rect 18420 12708 18472 12714
rect 18420 12650 18472 12656
rect 18708 10810 18736 13670
rect 18696 10804 18748 10810
rect 18696 10746 18748 10752
rect 18708 10606 18736 10746
rect 18696 10600 18748 10606
rect 18696 10542 18748 10548
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18248 10254 18368 10282
rect 18144 9444 18196 9450
rect 18144 9386 18196 9392
rect 17866 9072 17922 9081
rect 17866 9007 17922 9016
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 17972 8922 18000 8978
rect 17880 8894 18000 8922
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 17880 8090 17908 8894
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 17868 8084 17920 8090
rect 17868 8026 17920 8032
rect 17972 7290 18000 8774
rect 18064 8294 18092 8910
rect 18144 8356 18196 8362
rect 18144 8298 18196 8304
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 18064 7410 18092 8230
rect 18156 8090 18184 8298
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18052 7404 18104 7410
rect 18052 7346 18104 7352
rect 17972 7262 18184 7290
rect 17866 7168 17922 7177
rect 17866 7103 17922 7112
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 17788 5914 17816 6938
rect 17880 6866 17908 7103
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 17880 6458 17908 6802
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 17960 6180 18012 6186
rect 17960 6122 18012 6128
rect 17776 5908 17828 5914
rect 17776 5850 17828 5856
rect 17868 5840 17920 5846
rect 17868 5782 17920 5788
rect 17880 5370 17908 5782
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 17774 4720 17830 4729
rect 17774 4655 17776 4664
rect 17828 4655 17830 4664
rect 17776 4626 17828 4632
rect 17880 4554 17908 5306
rect 17972 4826 18000 6122
rect 18064 5846 18092 6734
rect 18052 5840 18104 5846
rect 18052 5782 18104 5788
rect 17960 4820 18012 4826
rect 17960 4762 18012 4768
rect 18050 4584 18106 4593
rect 17868 4548 17920 4554
rect 18050 4519 18106 4528
rect 17868 4490 17920 4496
rect 17406 4040 17462 4049
rect 17590 4040 17646 4049
rect 17406 3975 17462 3984
rect 17500 4004 17552 4010
rect 17316 3664 17368 3670
rect 17316 3606 17368 3612
rect 16908 3496 16910 3505
rect 16854 3431 16910 3440
rect 17038 3496 17094 3505
rect 17038 3431 17094 3440
rect 16684 3148 16804 3176
rect 16578 2816 16634 2825
rect 16578 2751 16634 2760
rect 16684 2666 16712 3148
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 16396 2644 16448 2650
rect 16396 2586 16448 2592
rect 16592 2638 16712 2666
rect 16408 2446 16436 2586
rect 16396 2440 16448 2446
rect 16396 2382 16448 2388
rect 16118 912 16174 921
rect 16118 847 16174 856
rect 16592 480 16620 2638
rect 16776 2514 16804 2994
rect 17420 2961 17448 3975
rect 17590 3975 17646 3984
rect 17500 3946 17552 3952
rect 17512 3466 17540 3946
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17788 3641 17816 3878
rect 17774 3632 17830 3641
rect 17592 3596 17644 3602
rect 17774 3567 17830 3576
rect 17592 3538 17644 3544
rect 17500 3460 17552 3466
rect 17500 3402 17552 3408
rect 17406 2952 17462 2961
rect 17406 2887 17462 2896
rect 17500 2848 17552 2854
rect 17498 2816 17500 2825
rect 17552 2816 17554 2825
rect 17498 2751 17554 2760
rect 16764 2508 16816 2514
rect 16764 2450 16816 2456
rect 17604 2310 17632 3538
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 17788 2854 17816 3470
rect 18064 3194 18092 4519
rect 18156 4185 18184 7262
rect 18142 4176 18198 4185
rect 18142 4111 18198 4120
rect 18248 3777 18276 10254
rect 18328 10192 18380 10198
rect 18328 10134 18380 10140
rect 18340 9761 18368 10134
rect 18510 9888 18566 9897
rect 18510 9823 18566 9832
rect 18326 9752 18382 9761
rect 18326 9687 18328 9696
rect 18380 9687 18382 9696
rect 18328 9658 18380 9664
rect 18328 9512 18380 9518
rect 18328 9454 18380 9460
rect 18340 6225 18368 9454
rect 18418 9344 18474 9353
rect 18418 9279 18474 9288
rect 18432 8634 18460 9279
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18326 6216 18382 6225
rect 18326 6151 18382 6160
rect 18328 5772 18380 5778
rect 18328 5714 18380 5720
rect 18340 5166 18368 5714
rect 18328 5160 18380 5166
rect 18328 5102 18380 5108
rect 18234 3768 18290 3777
rect 18234 3703 18290 3712
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18340 3369 18368 3470
rect 18326 3360 18382 3369
rect 18326 3295 18382 3304
rect 18052 3188 18104 3194
rect 18052 3130 18104 3136
rect 18236 2916 18288 2922
rect 18236 2858 18288 2864
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 18156 2650 18184 2790
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 17132 2304 17184 2310
rect 17132 2246 17184 2252
rect 17592 2304 17644 2310
rect 17592 2246 17644 2252
rect 17144 480 17172 2246
rect 17604 1873 17632 2246
rect 17590 1864 17646 1873
rect 17590 1799 17646 1808
rect 17604 598 17724 626
rect 9310 96 9366 105
rect 9310 31 9366 40
rect 9494 0 9550 480
rect 10046 0 10102 480
rect 10598 0 10654 480
rect 11150 0 11206 480
rect 11702 0 11758 480
rect 12254 0 12310 480
rect 12806 0 12862 480
rect 13358 0 13414 480
rect 13910 0 13966 480
rect 14370 0 14426 480
rect 14922 0 14978 480
rect 15474 0 15530 480
rect 16026 0 16082 480
rect 16578 0 16634 480
rect 17130 0 17186 480
rect 17604 377 17632 598
rect 17696 480 17724 598
rect 18248 480 18276 2858
rect 18432 2854 18460 8570
rect 18524 8362 18552 9823
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 18616 9178 18644 9454
rect 18604 9172 18656 9178
rect 18604 9114 18656 9120
rect 18512 8356 18564 8362
rect 18512 8298 18564 8304
rect 18524 7750 18552 8298
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18524 7324 18552 7686
rect 18604 7336 18656 7342
rect 18524 7296 18604 7324
rect 18604 7278 18656 7284
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18524 6322 18552 6598
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18616 5778 18644 7278
rect 18604 5772 18656 5778
rect 18604 5714 18656 5720
rect 18512 4480 18564 4486
rect 18512 4422 18564 4428
rect 18524 3942 18552 4422
rect 18512 3936 18564 3942
rect 18512 3878 18564 3884
rect 18420 2848 18472 2854
rect 18420 2790 18472 2796
rect 18326 2544 18382 2553
rect 18326 2479 18328 2488
rect 18380 2479 18382 2488
rect 18328 2450 18380 2456
rect 18328 2304 18380 2310
rect 18328 2246 18380 2252
rect 18340 1737 18368 2246
rect 18524 2009 18552 3878
rect 18708 3641 18736 10406
rect 18800 9178 18828 23598
rect 18880 23112 18932 23118
rect 18880 23054 18932 23060
rect 18892 21894 18920 23054
rect 19076 22817 19104 24142
rect 19168 23526 19196 24210
rect 19156 23520 19208 23526
rect 19156 23462 19208 23468
rect 19062 22808 19118 22817
rect 19062 22743 19118 22752
rect 19352 22522 19380 24346
rect 19168 22494 19380 22522
rect 18972 21956 19024 21962
rect 18972 21898 19024 21904
rect 18880 21888 18932 21894
rect 18880 21830 18932 21836
rect 18880 21548 18932 21554
rect 18880 21490 18932 21496
rect 18892 20942 18920 21490
rect 18880 20936 18932 20942
rect 18880 20878 18932 20884
rect 18878 20496 18934 20505
rect 18878 20431 18934 20440
rect 18892 17626 18920 20431
rect 18984 20058 19012 21898
rect 19062 21856 19118 21865
rect 19062 21791 19118 21800
rect 19076 21486 19104 21791
rect 19064 21480 19116 21486
rect 19064 21422 19116 21428
rect 19064 20800 19116 20806
rect 19064 20742 19116 20748
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 18984 19310 19012 19994
rect 19076 19854 19104 20742
rect 19064 19848 19116 19854
rect 19064 19790 19116 19796
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 19076 18902 19104 19790
rect 19064 18896 19116 18902
rect 19064 18838 19116 18844
rect 18972 18624 19024 18630
rect 18972 18566 19024 18572
rect 18984 18465 19012 18566
rect 18970 18456 19026 18465
rect 18970 18391 19026 18400
rect 19076 18290 19104 18838
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 19064 18080 19116 18086
rect 19062 18048 19064 18057
rect 19116 18048 19118 18057
rect 19062 17983 19118 17992
rect 18892 17598 19104 17626
rect 18880 17536 18932 17542
rect 18880 17478 18932 17484
rect 18892 16726 18920 17478
rect 18880 16720 18932 16726
rect 18878 16688 18880 16697
rect 18972 16720 19024 16726
rect 18932 16688 18934 16697
rect 18972 16662 19024 16668
rect 18878 16623 18934 16632
rect 18892 16250 18920 16623
rect 18880 16244 18932 16250
rect 18880 16186 18932 16192
rect 18880 14952 18932 14958
rect 18880 14894 18932 14900
rect 18892 14618 18920 14894
rect 18880 14612 18932 14618
rect 18880 14554 18932 14560
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 18892 12889 18920 13126
rect 18878 12880 18934 12889
rect 18878 12815 18880 12824
rect 18932 12815 18934 12824
rect 18880 12786 18932 12792
rect 18984 12730 19012 16662
rect 19076 16096 19104 17598
rect 19168 16726 19196 22494
rect 19432 22432 19484 22438
rect 19430 22400 19432 22409
rect 19484 22400 19486 22409
rect 19430 22335 19486 22344
rect 19536 22098 19564 25774
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19984 25356 20036 25362
rect 19984 25298 20036 25304
rect 19996 24614 20024 25298
rect 19984 24608 20036 24614
rect 19984 24550 20036 24556
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19616 24064 19668 24070
rect 19616 24006 19668 24012
rect 19628 23662 19656 24006
rect 19616 23656 19668 23662
rect 19616 23598 19668 23604
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19614 23216 19670 23225
rect 19614 23151 19670 23160
rect 19628 22778 19656 23151
rect 19616 22772 19668 22778
rect 19616 22714 19668 22720
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19524 22092 19576 22098
rect 19524 22034 19576 22040
rect 19248 21888 19300 21894
rect 19248 21830 19300 21836
rect 19260 21010 19288 21830
rect 19338 21584 19394 21593
rect 19338 21519 19394 21528
rect 19248 21004 19300 21010
rect 19248 20946 19300 20952
rect 19248 20256 19300 20262
rect 19248 20198 19300 20204
rect 19260 18222 19288 20198
rect 19352 19310 19380 21519
rect 19522 21448 19578 21457
rect 19522 21383 19578 21392
rect 19536 21146 19564 21383
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19524 21140 19576 21146
rect 19524 21082 19576 21088
rect 19706 21040 19762 21049
rect 19706 20975 19708 20984
rect 19760 20975 19762 20984
rect 19708 20946 19760 20952
rect 19432 20392 19484 20398
rect 19432 20334 19484 20340
rect 19444 19718 19472 20334
rect 19720 20330 19748 20946
rect 19890 20904 19946 20913
rect 19890 20839 19892 20848
rect 19944 20839 19946 20848
rect 19892 20810 19944 20816
rect 19708 20324 19760 20330
rect 19708 20266 19760 20272
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19536 19417 19564 20198
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19614 19952 19670 19961
rect 19614 19887 19670 19896
rect 19522 19408 19578 19417
rect 19522 19343 19578 19352
rect 19340 19304 19392 19310
rect 19628 19258 19656 19887
rect 19708 19712 19760 19718
rect 19708 19654 19760 19660
rect 19720 19281 19748 19654
rect 19340 19246 19392 19252
rect 19536 19230 19656 19258
rect 19706 19272 19762 19281
rect 19340 19168 19392 19174
rect 19340 19110 19392 19116
rect 19248 18216 19300 18222
rect 19248 18158 19300 18164
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 19260 17338 19288 18022
rect 19248 17332 19300 17338
rect 19248 17274 19300 17280
rect 19248 17128 19300 17134
rect 19352 17116 19380 19110
rect 19430 18864 19486 18873
rect 19536 18850 19564 19230
rect 19706 19207 19762 19216
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19536 18822 19656 18850
rect 19430 18799 19432 18808
rect 19484 18799 19486 18808
rect 19432 18770 19484 18776
rect 19524 18760 19576 18766
rect 19524 18702 19576 18708
rect 19432 18692 19484 18698
rect 19432 18634 19484 18640
rect 19444 17921 19472 18634
rect 19430 17912 19486 17921
rect 19536 17882 19564 18702
rect 19628 18290 19656 18822
rect 19616 18284 19668 18290
rect 19616 18226 19668 18232
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19996 17882 20024 24550
rect 20088 24177 20116 27520
rect 20350 25256 20406 25265
rect 20350 25191 20406 25200
rect 20168 24744 20220 24750
rect 20168 24686 20220 24692
rect 20074 24168 20130 24177
rect 20074 24103 20130 24112
rect 20180 23730 20208 24686
rect 20364 23866 20392 25191
rect 20640 24721 20668 27520
rect 21284 25906 21312 27520
rect 21272 25900 21324 25906
rect 21272 25842 21324 25848
rect 21364 25492 21416 25498
rect 21364 25434 21416 25440
rect 20720 24880 20772 24886
rect 20720 24822 20772 24828
rect 20626 24712 20682 24721
rect 20626 24647 20682 24656
rect 20732 23866 20760 24822
rect 21088 24608 21140 24614
rect 21088 24550 21140 24556
rect 21100 24313 21128 24550
rect 21376 24410 21404 25434
rect 21732 24608 21784 24614
rect 21836 24596 21864 27520
rect 21916 25696 21968 25702
rect 21916 25638 21968 25644
rect 21928 25498 21956 25638
rect 21916 25492 21968 25498
rect 21916 25434 21968 25440
rect 22008 25356 22060 25362
rect 22008 25298 22060 25304
rect 22020 24614 22048 25298
rect 21784 24568 21864 24596
rect 22008 24608 22060 24614
rect 21732 24550 21784 24556
rect 22008 24550 22060 24556
rect 21364 24404 21416 24410
rect 21364 24346 21416 24352
rect 21180 24336 21232 24342
rect 21086 24304 21142 24313
rect 21180 24278 21232 24284
rect 21086 24239 21142 24248
rect 20352 23860 20404 23866
rect 20352 23802 20404 23808
rect 20720 23860 20772 23866
rect 20720 23802 20772 23808
rect 20168 23724 20220 23730
rect 20168 23666 20220 23672
rect 20364 23662 20392 23802
rect 20352 23656 20404 23662
rect 20352 23598 20404 23604
rect 20168 23520 20220 23526
rect 20168 23462 20220 23468
rect 20076 23180 20128 23186
rect 20076 23122 20128 23128
rect 20088 22642 20116 23122
rect 20076 22636 20128 22642
rect 20076 22578 20128 22584
rect 20076 22432 20128 22438
rect 20076 22374 20128 22380
rect 20088 22030 20116 22374
rect 20076 22024 20128 22030
rect 20076 21966 20128 21972
rect 20074 21720 20130 21729
rect 20074 21655 20076 21664
rect 20128 21655 20130 21664
rect 20076 21626 20128 21632
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 20088 20369 20116 20402
rect 20074 20360 20130 20369
rect 20074 20295 20130 20304
rect 20088 20058 20116 20295
rect 20076 20052 20128 20058
rect 20076 19994 20128 20000
rect 20088 19446 20116 19994
rect 20076 19440 20128 19446
rect 20076 19382 20128 19388
rect 19430 17847 19486 17856
rect 19524 17876 19576 17882
rect 19444 17338 19472 17847
rect 19524 17818 19576 17824
rect 19984 17876 20036 17882
rect 19984 17818 20036 17824
rect 20076 17808 20128 17814
rect 20074 17776 20076 17785
rect 20128 17776 20130 17785
rect 19984 17740 20036 17746
rect 20074 17711 20130 17720
rect 19984 17682 20036 17688
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19300 17088 19380 17116
rect 19248 17070 19300 17076
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19156 16720 19208 16726
rect 19156 16662 19208 16668
rect 19076 16068 19288 16096
rect 19064 15972 19116 15978
rect 19064 15914 19116 15920
rect 19076 14770 19104 15914
rect 19156 15564 19208 15570
rect 19156 15506 19208 15512
rect 19168 15473 19196 15506
rect 19154 15464 19210 15473
rect 19154 15399 19210 15408
rect 19168 15162 19196 15399
rect 19156 15156 19208 15162
rect 19156 15098 19208 15104
rect 19076 14742 19196 14770
rect 19064 14612 19116 14618
rect 19064 14554 19116 14560
rect 19076 12850 19104 14554
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 18892 12702 19012 12730
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 18788 6656 18840 6662
rect 18788 6598 18840 6604
rect 18800 6186 18828 6598
rect 18788 6180 18840 6186
rect 18788 6122 18840 6128
rect 18788 4072 18840 4078
rect 18788 4014 18840 4020
rect 18694 3632 18750 3641
rect 18694 3567 18750 3576
rect 18694 3496 18750 3505
rect 18604 3460 18656 3466
rect 18694 3431 18750 3440
rect 18604 3402 18656 3408
rect 18616 3058 18644 3402
rect 18708 3233 18736 3431
rect 18800 3369 18828 4014
rect 18892 3670 18920 12702
rect 19076 12442 19104 12786
rect 19168 12442 19196 14742
rect 19260 14482 19288 16068
rect 19248 14476 19300 14482
rect 19248 14418 19300 14424
rect 19352 14414 19380 16934
rect 19444 16153 19472 17138
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19524 16788 19576 16794
rect 19524 16730 19576 16736
rect 19430 16144 19486 16153
rect 19430 16079 19486 16088
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19340 14408 19392 14414
rect 19338 14376 19340 14385
rect 19392 14376 19394 14385
rect 19338 14311 19394 14320
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19260 13394 19288 14214
rect 19444 14074 19472 14962
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19338 13560 19394 13569
rect 19338 13495 19394 13504
rect 19352 13394 19380 13495
rect 19444 13462 19472 14010
rect 19432 13456 19484 13462
rect 19432 13398 19484 13404
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19444 12986 19472 13398
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19064 12436 19116 12442
rect 19064 12378 19116 12384
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 19340 12232 19392 12238
rect 19340 12174 19392 12180
rect 19352 11626 19380 12174
rect 19536 11694 19564 16730
rect 19616 16652 19668 16658
rect 19616 16594 19668 16600
rect 19628 16153 19656 16594
rect 19614 16144 19670 16153
rect 19614 16079 19670 16088
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19996 15586 20024 17682
rect 20076 16992 20128 16998
rect 20076 16934 20128 16940
rect 20088 15609 20116 16934
rect 19904 15558 20024 15586
rect 20074 15600 20130 15609
rect 19904 15094 19932 15558
rect 20074 15535 20130 15544
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 19892 15088 19944 15094
rect 19892 15030 19944 15036
rect 19996 14822 20024 15438
rect 20076 15428 20128 15434
rect 20076 15370 20128 15376
rect 20088 15042 20116 15370
rect 20180 15162 20208 23462
rect 21192 23322 21220 24278
rect 21376 23882 21404 24346
rect 21548 24200 21600 24206
rect 21548 24142 21600 24148
rect 21376 23866 21496 23882
rect 21376 23860 21508 23866
rect 21376 23854 21456 23860
rect 21456 23802 21508 23808
rect 21364 23520 21416 23526
rect 21364 23462 21416 23468
rect 21180 23316 21232 23322
rect 21180 23258 21232 23264
rect 21180 23180 21232 23186
rect 21180 23122 21232 23128
rect 20352 22976 20404 22982
rect 20352 22918 20404 22924
rect 20720 22976 20772 22982
rect 20720 22918 20772 22924
rect 20364 22506 20392 22918
rect 20352 22500 20404 22506
rect 20352 22442 20404 22448
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 20272 19310 20300 22170
rect 20364 21690 20392 22442
rect 20732 22234 20760 22918
rect 21192 22438 21220 23122
rect 21180 22432 21232 22438
rect 21180 22374 21232 22380
rect 21086 22264 21142 22273
rect 20720 22228 20772 22234
rect 21086 22199 21142 22208
rect 20720 22170 20772 22176
rect 20628 22092 20680 22098
rect 20628 22034 20680 22040
rect 20444 22024 20496 22030
rect 20444 21966 20496 21972
rect 20352 21684 20404 21690
rect 20352 21626 20404 21632
rect 20456 19961 20484 21966
rect 20442 19952 20498 19961
rect 20442 19887 20498 19896
rect 20534 19816 20590 19825
rect 20534 19751 20590 19760
rect 20352 19712 20404 19718
rect 20352 19654 20404 19660
rect 20364 19378 20392 19654
rect 20352 19372 20404 19378
rect 20352 19314 20404 19320
rect 20260 19304 20312 19310
rect 20260 19246 20312 19252
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 20272 18630 20300 19110
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 20272 16674 20300 18566
rect 20364 18290 20392 19314
rect 20442 18864 20498 18873
rect 20442 18799 20498 18808
rect 20352 18284 20404 18290
rect 20352 18226 20404 18232
rect 20364 17882 20392 18226
rect 20352 17876 20404 17882
rect 20352 17818 20404 17824
rect 20350 17776 20406 17785
rect 20350 17711 20352 17720
rect 20404 17711 20406 17720
rect 20352 17682 20404 17688
rect 20352 17060 20404 17066
rect 20352 17002 20404 17008
rect 20364 16794 20392 17002
rect 20352 16788 20404 16794
rect 20352 16730 20404 16736
rect 20272 16646 20392 16674
rect 20258 16008 20314 16017
rect 20258 15943 20314 15952
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20088 15014 20208 15042
rect 20074 14920 20130 14929
rect 20180 14890 20208 15014
rect 20074 14855 20076 14864
rect 20128 14855 20130 14864
rect 20168 14884 20220 14890
rect 20076 14826 20128 14832
rect 20168 14826 20220 14832
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19996 14521 20024 14758
rect 20088 14618 20116 14826
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 19982 14512 20038 14521
rect 19714 14476 19766 14482
rect 20272 14498 20300 15943
rect 20364 15502 20392 16646
rect 20352 15496 20404 15502
rect 20352 15438 20404 15444
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 20364 14958 20392 15302
rect 20352 14952 20404 14958
rect 20352 14894 20404 14900
rect 20352 14816 20404 14822
rect 20352 14758 20404 14764
rect 19982 14447 20038 14456
rect 20088 14470 20300 14498
rect 19714 14418 19766 14424
rect 19720 14113 19748 14418
rect 19984 14408 20036 14414
rect 19984 14350 20036 14356
rect 19706 14104 19762 14113
rect 19706 14039 19708 14048
rect 19760 14039 19762 14048
rect 19708 14010 19760 14016
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19996 13530 20024 14350
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 20088 12764 20116 14470
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 20180 12918 20208 14350
rect 20364 14226 20392 14758
rect 20456 14346 20484 18799
rect 20548 16697 20576 19751
rect 20640 19514 20668 22034
rect 20996 22024 21048 22030
rect 20996 21966 21048 21972
rect 20904 21888 20956 21894
rect 20904 21830 20956 21836
rect 20916 21554 20944 21830
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 21008 21146 21036 21966
rect 21100 21962 21128 22199
rect 21088 21956 21140 21962
rect 21088 21898 21140 21904
rect 21192 21842 21220 22374
rect 21192 21814 21312 21842
rect 20996 21140 21048 21146
rect 20996 21082 21048 21088
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 20732 20505 20760 20946
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 21008 20777 21036 20878
rect 20994 20768 21050 20777
rect 20994 20703 21050 20712
rect 21008 20602 21036 20703
rect 20996 20596 21048 20602
rect 20996 20538 21048 20544
rect 20718 20496 20774 20505
rect 20718 20431 20720 20440
rect 20772 20431 20774 20440
rect 20720 20402 20772 20408
rect 20812 20256 20864 20262
rect 20718 20224 20774 20233
rect 20812 20198 20864 20204
rect 21180 20256 21232 20262
rect 21180 20198 21232 20204
rect 20718 20159 20774 20168
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20732 19258 20760 20159
rect 20824 19961 20852 20198
rect 20810 19952 20866 19961
rect 20810 19887 20866 19896
rect 20904 19712 20956 19718
rect 20904 19654 20956 19660
rect 21088 19712 21140 19718
rect 21192 19689 21220 20198
rect 21088 19654 21140 19660
rect 21178 19680 21234 19689
rect 20916 19417 20944 19654
rect 21100 19530 21128 19654
rect 21178 19615 21234 19624
rect 21100 19502 21220 19530
rect 20902 19408 20958 19417
rect 20902 19343 20958 19352
rect 21192 19258 21220 19502
rect 20640 18970 20668 19246
rect 20732 19230 20944 19258
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20628 18964 20680 18970
rect 20628 18906 20680 18912
rect 20534 16688 20590 16697
rect 20534 16623 20590 16632
rect 20536 16584 20588 16590
rect 20536 16526 20588 16532
rect 20548 16250 20576 16526
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20548 15502 20576 16186
rect 20640 15745 20668 18906
rect 20732 18737 20760 19110
rect 20718 18728 20774 18737
rect 20718 18663 20774 18672
rect 20812 18624 20864 18630
rect 20812 18566 20864 18572
rect 20718 18184 20774 18193
rect 20718 18119 20720 18128
rect 20772 18119 20774 18128
rect 20720 18090 20772 18096
rect 20718 18048 20774 18057
rect 20718 17983 20774 17992
rect 20626 15736 20682 15745
rect 20626 15671 20682 15680
rect 20626 15600 20682 15609
rect 20626 15535 20628 15544
rect 20680 15535 20682 15544
rect 20628 15506 20680 15512
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 20548 14414 20576 15438
rect 20628 15088 20680 15094
rect 20628 15030 20680 15036
rect 20640 14618 20668 15030
rect 20628 14612 20680 14618
rect 20628 14554 20680 14560
rect 20626 14512 20682 14521
rect 20626 14447 20682 14456
rect 20536 14408 20588 14414
rect 20536 14350 20588 14356
rect 20444 14340 20496 14346
rect 20444 14282 20496 14288
rect 20364 14198 20576 14226
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20258 13016 20314 13025
rect 20258 12951 20260 12960
rect 20312 12951 20314 12960
rect 20260 12922 20312 12928
rect 20168 12912 20220 12918
rect 20168 12854 20220 12860
rect 20088 12736 20208 12764
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19984 12096 20036 12102
rect 19984 12038 20036 12044
rect 19524 11688 19576 11694
rect 19524 11630 19576 11636
rect 19340 11620 19392 11626
rect 19340 11562 19392 11568
rect 19352 11014 19380 11562
rect 19524 11552 19576 11558
rect 19524 11494 19576 11500
rect 19536 11150 19564 11494
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19996 11354 20024 12038
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 20076 11212 20128 11218
rect 20076 11154 20128 11160
rect 19524 11144 19576 11150
rect 19524 11086 19576 11092
rect 19432 11076 19484 11082
rect 19432 11018 19484 11024
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 19352 10470 19380 10950
rect 19340 10464 19392 10470
rect 19260 10424 19340 10452
rect 19154 10296 19210 10305
rect 19154 10231 19156 10240
rect 19208 10231 19210 10240
rect 19156 10202 19208 10208
rect 18972 9988 19024 9994
rect 18972 9930 19024 9936
rect 18984 9586 19012 9930
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 19168 9450 19196 10202
rect 19260 9586 19288 10424
rect 19340 10406 19392 10412
rect 19444 9654 19472 11018
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19522 10160 19578 10169
rect 19522 10095 19524 10104
rect 19576 10095 19578 10104
rect 19616 10124 19668 10130
rect 19524 10066 19576 10072
rect 19616 10066 19668 10072
rect 19432 9648 19484 9654
rect 19338 9616 19394 9625
rect 19248 9580 19300 9586
rect 19432 9590 19484 9596
rect 19338 9551 19394 9560
rect 19248 9522 19300 9528
rect 19156 9444 19208 9450
rect 19156 9386 19208 9392
rect 19156 8968 19208 8974
rect 19156 8910 19208 8916
rect 18972 6792 19024 6798
rect 18972 6734 19024 6740
rect 18984 6474 19012 6734
rect 19168 6730 19196 8910
rect 19352 8566 19380 9551
rect 19432 9376 19484 9382
rect 19430 9344 19432 9353
rect 19628 9364 19656 10066
rect 19984 9920 20036 9926
rect 19984 9862 20036 9868
rect 19892 9512 19944 9518
rect 19890 9480 19892 9489
rect 19944 9480 19946 9489
rect 19890 9415 19946 9424
rect 19484 9344 19656 9364
rect 19486 9336 19656 9344
rect 19430 9279 19486 9288
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19430 9072 19486 9081
rect 19996 9042 20024 9862
rect 20088 9654 20116 11154
rect 20076 9648 20128 9654
rect 20076 9590 20128 9596
rect 19430 9007 19486 9016
rect 19984 9036 20036 9042
rect 19444 8634 19472 9007
rect 19984 8978 20036 8984
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19340 8560 19392 8566
rect 19340 8502 19392 8508
rect 19536 8294 19564 8910
rect 19524 8288 19576 8294
rect 19524 8230 19576 8236
rect 19536 8090 19564 8230
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 19432 7744 19484 7750
rect 19432 7686 19484 7692
rect 19444 6934 19472 7686
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19432 6928 19484 6934
rect 19430 6896 19432 6905
rect 19484 6896 19486 6905
rect 19430 6831 19486 6840
rect 20088 6798 20116 7142
rect 19524 6792 19576 6798
rect 19522 6760 19524 6769
rect 20076 6792 20128 6798
rect 19576 6760 19578 6769
rect 19156 6724 19208 6730
rect 20076 6734 20128 6740
rect 19522 6695 19578 6704
rect 19156 6666 19208 6672
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19154 6488 19210 6497
rect 18984 6446 19154 6474
rect 19154 6423 19156 6432
rect 19208 6423 19210 6432
rect 19156 6394 19208 6400
rect 19248 6384 19300 6390
rect 19248 6326 19300 6332
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 18972 6112 19024 6118
rect 18972 6054 19024 6060
rect 18984 5681 19012 6054
rect 18970 5672 19026 5681
rect 18970 5607 19026 5616
rect 19168 5574 19196 6258
rect 19260 6066 19288 6326
rect 19524 6112 19576 6118
rect 19260 6038 19472 6066
rect 19524 6054 19576 6060
rect 19340 5636 19392 5642
rect 19340 5578 19392 5584
rect 19156 5568 19208 5574
rect 19156 5510 19208 5516
rect 19168 5098 19196 5510
rect 19156 5092 19208 5098
rect 19156 5034 19208 5040
rect 19168 4706 19196 5034
rect 19248 4820 19300 4826
rect 19352 4808 19380 5578
rect 19444 4826 19472 6038
rect 19536 5030 19564 6054
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19524 5024 19576 5030
rect 19524 4966 19576 4972
rect 19300 4780 19380 4808
rect 19248 4762 19300 4768
rect 19168 4678 19288 4706
rect 19260 4282 19288 4678
rect 19248 4276 19300 4282
rect 19248 4218 19300 4224
rect 19260 3924 19288 4218
rect 19352 4078 19380 4780
rect 19432 4820 19484 4826
rect 19432 4762 19484 4768
rect 19432 4684 19484 4690
rect 19432 4626 19484 4632
rect 19444 4214 19472 4626
rect 19536 4622 19564 4966
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19996 4690 20024 6598
rect 20088 5914 20116 6734
rect 20076 5908 20128 5914
rect 20076 5850 20128 5856
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 19984 4684 20036 4690
rect 19984 4626 20036 4632
rect 19524 4616 19576 4622
rect 19524 4558 19576 4564
rect 19982 4584 20038 4593
rect 19982 4519 20038 4528
rect 19432 4208 19484 4214
rect 19432 4150 19484 4156
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 19996 3942 20024 4519
rect 19340 3936 19392 3942
rect 19260 3896 19340 3924
rect 19984 3936 20036 3942
rect 19340 3878 19392 3884
rect 19430 3904 19486 3913
rect 19984 3878 20036 3884
rect 19430 3839 19486 3848
rect 19338 3768 19394 3777
rect 19338 3703 19394 3712
rect 19352 3670 19380 3703
rect 18880 3664 18932 3670
rect 18880 3606 18932 3612
rect 19340 3664 19392 3670
rect 19340 3606 19392 3612
rect 18786 3360 18842 3369
rect 18786 3295 18842 3304
rect 18694 3224 18750 3233
rect 18694 3159 18750 3168
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18708 2650 18736 3159
rect 18892 2990 18920 3606
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 19076 3126 19104 3538
rect 19064 3120 19116 3126
rect 19064 3062 19116 3068
rect 18880 2984 18932 2990
rect 18880 2926 18932 2932
rect 18696 2644 18748 2650
rect 18696 2586 18748 2592
rect 18510 2000 18566 2009
rect 18510 1935 18566 1944
rect 18788 1964 18840 1970
rect 18788 1906 18840 1912
rect 18326 1728 18382 1737
rect 18326 1663 18382 1672
rect 18800 480 18828 1906
rect 19444 1306 19472 3839
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19536 3194 19564 3674
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 19616 3120 19668 3126
rect 19614 3088 19616 3097
rect 19668 3088 19670 3097
rect 19614 3023 19670 3032
rect 20088 2990 20116 4966
rect 20180 3738 20208 12736
rect 20260 12164 20312 12170
rect 20260 12106 20312 12112
rect 20272 11762 20300 12106
rect 20260 11756 20312 11762
rect 20260 11698 20312 11704
rect 20260 11552 20312 11558
rect 20260 11494 20312 11500
rect 20272 11082 20300 11494
rect 20260 11076 20312 11082
rect 20260 11018 20312 11024
rect 20260 10600 20312 10606
rect 20260 10542 20312 10548
rect 20272 8838 20300 10542
rect 20260 8832 20312 8838
rect 20260 8774 20312 8780
rect 20272 8430 20300 8774
rect 20260 8424 20312 8430
rect 20260 8366 20312 8372
rect 20364 8129 20392 14010
rect 20444 13184 20496 13190
rect 20444 13126 20496 13132
rect 20456 10180 20484 13126
rect 20548 10282 20576 14198
rect 20640 14113 20668 14447
rect 20626 14104 20682 14113
rect 20732 14074 20760 17983
rect 20626 14039 20682 14048
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20626 13968 20682 13977
rect 20626 13903 20682 13912
rect 20640 11898 20668 13903
rect 20720 13864 20772 13870
rect 20718 13832 20720 13841
rect 20772 13832 20774 13841
rect 20718 13767 20774 13776
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20628 11688 20680 11694
rect 20628 11630 20680 11636
rect 20640 10826 20668 11630
rect 20732 11257 20760 13126
rect 20824 12374 20852 18566
rect 20916 18222 20944 19230
rect 21100 19230 21220 19258
rect 20904 18216 20956 18222
rect 20904 18158 20956 18164
rect 20916 18086 20944 18158
rect 20904 18080 20956 18086
rect 20904 18022 20956 18028
rect 20916 17762 20944 18022
rect 20916 17734 21036 17762
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 20916 16998 20944 17614
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20916 14074 20944 16934
rect 21008 16017 21036 17734
rect 20994 16008 21050 16017
rect 20994 15943 21050 15952
rect 20996 15904 21048 15910
rect 20996 15846 21048 15852
rect 21008 15473 21036 15846
rect 20994 15464 21050 15473
rect 20994 15399 21050 15408
rect 21008 15201 21036 15399
rect 20994 15192 21050 15201
rect 20994 15127 21050 15136
rect 20994 14648 21050 14657
rect 20994 14583 21050 14592
rect 20904 14068 20956 14074
rect 20904 14010 20956 14016
rect 21008 13462 21036 14583
rect 20996 13456 21048 13462
rect 20996 13398 21048 13404
rect 20994 12744 21050 12753
rect 20994 12679 20996 12688
rect 21048 12679 21050 12688
rect 20996 12650 21048 12656
rect 20996 12436 21048 12442
rect 20996 12378 21048 12384
rect 20812 12368 20864 12374
rect 20812 12310 20864 12316
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20810 12200 20866 12209
rect 20810 12135 20866 12144
rect 20718 11248 20774 11257
rect 20718 11183 20774 11192
rect 20640 10810 20760 10826
rect 20640 10804 20772 10810
rect 20640 10798 20720 10804
rect 20720 10746 20772 10752
rect 20824 10742 20852 12135
rect 20916 11529 20944 12242
rect 20902 11520 20958 11529
rect 20902 11455 20958 11464
rect 20902 10976 20958 10985
rect 20902 10911 20958 10920
rect 20812 10736 20864 10742
rect 20812 10678 20864 10684
rect 20812 10600 20864 10606
rect 20812 10542 20864 10548
rect 20548 10254 20760 10282
rect 20456 10152 20576 10180
rect 20444 9988 20496 9994
rect 20444 9930 20496 9936
rect 20350 8120 20406 8129
rect 20350 8055 20406 8064
rect 20350 7576 20406 7585
rect 20350 7511 20406 7520
rect 20364 7206 20392 7511
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 20260 6248 20312 6254
rect 20260 6190 20312 6196
rect 20272 5710 20300 6190
rect 20456 5953 20484 9930
rect 20548 9466 20576 10152
rect 20628 10124 20680 10130
rect 20628 10066 20680 10072
rect 20640 9586 20668 10066
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20548 9438 20668 9466
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20548 9217 20576 9318
rect 20534 9208 20590 9217
rect 20534 9143 20536 9152
rect 20588 9143 20590 9152
rect 20536 9114 20588 9120
rect 20548 9083 20576 9114
rect 20536 9036 20588 9042
rect 20536 8978 20588 8984
rect 20548 8673 20576 8978
rect 20640 8906 20668 9438
rect 20628 8900 20680 8906
rect 20628 8842 20680 8848
rect 20732 8786 20760 10254
rect 20824 9194 20852 10542
rect 20916 9926 20944 10911
rect 20904 9920 20956 9926
rect 20904 9862 20956 9868
rect 20916 9450 20944 9862
rect 20904 9444 20956 9450
rect 20904 9386 20956 9392
rect 21008 9382 21036 12378
rect 21100 12288 21128 19230
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 21192 18057 21220 19110
rect 21178 18048 21234 18057
rect 21178 17983 21234 17992
rect 21180 17604 21232 17610
rect 21180 17546 21232 17552
rect 21192 16998 21220 17546
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 21192 15570 21220 16934
rect 21180 15564 21232 15570
rect 21180 15506 21232 15512
rect 21180 15088 21232 15094
rect 21178 15056 21180 15065
rect 21232 15056 21234 15065
rect 21178 14991 21234 15000
rect 21180 14476 21232 14482
rect 21180 14418 21232 14424
rect 21192 14278 21220 14418
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 21192 14006 21220 14214
rect 21180 14000 21232 14006
rect 21180 13942 21232 13948
rect 21178 13288 21234 13297
rect 21178 13223 21234 13232
rect 21192 12986 21220 13223
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21100 12260 21220 12288
rect 21086 12200 21142 12209
rect 21086 12135 21088 12144
rect 21140 12135 21142 12144
rect 21088 12106 21140 12112
rect 21086 11656 21142 11665
rect 21086 11591 21142 11600
rect 21100 10810 21128 11591
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 20824 9166 21036 9194
rect 20904 9036 20956 9042
rect 20904 8978 20956 8984
rect 20640 8758 20760 8786
rect 20812 8832 20864 8838
rect 20812 8774 20864 8780
rect 20534 8664 20590 8673
rect 20534 8599 20590 8608
rect 20640 8514 20668 8758
rect 20548 8486 20668 8514
rect 20548 7562 20576 8486
rect 20640 8362 20760 8378
rect 20640 8356 20772 8362
rect 20640 8350 20720 8356
rect 20640 8090 20668 8350
rect 20720 8298 20772 8304
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20824 7993 20852 8774
rect 20810 7984 20866 7993
rect 20810 7919 20866 7928
rect 20810 7848 20866 7857
rect 20810 7783 20866 7792
rect 20548 7534 20760 7562
rect 20824 7546 20852 7783
rect 20916 7750 20944 8978
rect 20904 7744 20956 7750
rect 20904 7686 20956 7692
rect 20732 7478 20760 7534
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20720 7472 20772 7478
rect 20720 7414 20772 7420
rect 20732 7002 20760 7414
rect 20720 6996 20772 7002
rect 20720 6938 20772 6944
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20442 5944 20498 5953
rect 20442 5879 20498 5888
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 20272 5166 20300 5646
rect 20350 5264 20406 5273
rect 20350 5199 20406 5208
rect 20536 5228 20588 5234
rect 20260 5160 20312 5166
rect 20260 5102 20312 5108
rect 20260 5024 20312 5030
rect 20260 4966 20312 4972
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 20168 3052 20220 3058
rect 20168 2994 20220 3000
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 20076 2848 20128 2854
rect 20074 2816 20076 2825
rect 20128 2816 20130 2825
rect 19622 2748 19918 2768
rect 20074 2751 20130 2760
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 20180 2650 20208 2994
rect 20272 2854 20300 4966
rect 20364 4826 20392 5199
rect 20536 5170 20588 5176
rect 20352 4820 20404 4826
rect 20352 4762 20404 4768
rect 20548 4146 20576 5170
rect 20640 4808 20668 6598
rect 20810 6352 20866 6361
rect 20810 6287 20866 6296
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20732 5370 20760 6054
rect 20824 5794 20852 6287
rect 20916 5914 20944 7686
rect 21008 6746 21036 9166
rect 21100 8430 21128 10610
rect 21192 9722 21220 12260
rect 21180 9716 21232 9722
rect 21180 9658 21232 9664
rect 21284 9586 21312 21814
rect 21376 20330 21404 23462
rect 21560 23202 21588 24142
rect 21822 23488 21878 23497
rect 21822 23423 21878 23432
rect 21468 23174 21588 23202
rect 21468 22982 21496 23174
rect 21548 23112 21600 23118
rect 21548 23054 21600 23060
rect 21456 22976 21508 22982
rect 21456 22918 21508 22924
rect 21364 20324 21416 20330
rect 21364 20266 21416 20272
rect 21364 18760 21416 18766
rect 21362 18728 21364 18737
rect 21416 18728 21418 18737
rect 21362 18663 21418 18672
rect 21376 18426 21404 18663
rect 21364 18420 21416 18426
rect 21364 18362 21416 18368
rect 21362 18320 21418 18329
rect 21362 18255 21418 18264
rect 21376 18086 21404 18255
rect 21364 18080 21416 18086
rect 21364 18022 21416 18028
rect 21364 17740 21416 17746
rect 21364 17682 21416 17688
rect 21376 16794 21404 17682
rect 21364 16788 21416 16794
rect 21364 16730 21416 16736
rect 21376 13258 21404 16730
rect 21364 13252 21416 13258
rect 21364 13194 21416 13200
rect 21362 11656 21418 11665
rect 21362 11591 21418 11600
rect 21376 11257 21404 11591
rect 21362 11248 21418 11257
rect 21362 11183 21418 11192
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 21376 10266 21404 11086
rect 21468 10606 21496 22918
rect 21560 22438 21588 23054
rect 21836 22778 21864 23423
rect 22020 23338 22048 24550
rect 22190 23896 22246 23905
rect 22190 23831 22246 23840
rect 22020 23310 22140 23338
rect 21916 22976 21968 22982
rect 21916 22918 21968 22924
rect 21824 22772 21876 22778
rect 21824 22714 21876 22720
rect 21822 22672 21878 22681
rect 21822 22607 21878 22616
rect 21548 22432 21600 22438
rect 21548 22374 21600 22380
rect 21560 22166 21588 22374
rect 21836 22166 21864 22607
rect 21548 22160 21600 22166
rect 21548 22102 21600 22108
rect 21732 22160 21784 22166
rect 21732 22102 21784 22108
rect 21824 22160 21876 22166
rect 21824 22102 21876 22108
rect 21640 21684 21692 21690
rect 21640 21626 21692 21632
rect 21652 21457 21680 21626
rect 21638 21448 21694 21457
rect 21638 21383 21694 21392
rect 21638 20632 21694 20641
rect 21638 20567 21694 20576
rect 21652 20466 21680 20567
rect 21640 20460 21692 20466
rect 21640 20402 21692 20408
rect 21640 20256 21692 20262
rect 21640 20198 21692 20204
rect 21548 19848 21600 19854
rect 21548 19790 21600 19796
rect 21560 18630 21588 19790
rect 21652 19718 21680 20198
rect 21640 19712 21692 19718
rect 21640 19654 21692 19660
rect 21640 18760 21692 18766
rect 21640 18702 21692 18708
rect 21548 18624 21600 18630
rect 21548 18566 21600 18572
rect 21652 17898 21680 18702
rect 21560 17870 21680 17898
rect 21560 17814 21588 17870
rect 21548 17808 21600 17814
rect 21548 17750 21600 17756
rect 21560 17649 21588 17750
rect 21546 17640 21602 17649
rect 21546 17575 21602 17584
rect 21640 17536 21692 17542
rect 21640 17478 21692 17484
rect 21548 17196 21600 17202
rect 21548 17138 21600 17144
rect 21560 16998 21588 17138
rect 21548 16992 21600 16998
rect 21548 16934 21600 16940
rect 21560 16726 21588 16934
rect 21548 16720 21600 16726
rect 21548 16662 21600 16668
rect 21560 16182 21588 16662
rect 21548 16176 21600 16182
rect 21548 16118 21600 16124
rect 21652 15745 21680 17478
rect 21638 15736 21694 15745
rect 21638 15671 21694 15680
rect 21546 15328 21602 15337
rect 21546 15263 21602 15272
rect 21560 15162 21588 15263
rect 21548 15156 21600 15162
rect 21548 15098 21600 15104
rect 21548 14816 21600 14822
rect 21548 14758 21600 14764
rect 21560 14278 21588 14758
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 21548 14272 21600 14278
rect 21546 14240 21548 14249
rect 21600 14240 21602 14249
rect 21546 14175 21602 14184
rect 21652 14113 21680 14350
rect 21638 14104 21694 14113
rect 21638 14039 21694 14048
rect 21640 13456 21692 13462
rect 21640 13398 21692 13404
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 21560 12628 21588 13330
rect 21652 12782 21680 13398
rect 21640 12776 21692 12782
rect 21640 12718 21692 12724
rect 21560 12600 21680 12628
rect 21652 12102 21680 12600
rect 21640 12096 21692 12102
rect 21546 12064 21602 12073
rect 21640 12038 21692 12044
rect 21546 11999 21602 12008
rect 21456 10600 21508 10606
rect 21456 10542 21508 10548
rect 21364 10260 21416 10266
rect 21364 10202 21416 10208
rect 21272 9580 21324 9586
rect 21272 9522 21324 9528
rect 21560 9500 21588 11999
rect 21468 9472 21588 9500
rect 21180 9376 21232 9382
rect 21180 9318 21232 9324
rect 21364 9376 21416 9382
rect 21364 9318 21416 9324
rect 21192 9178 21220 9318
rect 21180 9172 21232 9178
rect 21180 9114 21232 9120
rect 21180 8968 21232 8974
rect 21180 8910 21232 8916
rect 21192 8634 21220 8910
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 21088 8424 21140 8430
rect 21088 8366 21140 8372
rect 21376 6934 21404 9318
rect 21468 8838 21496 9472
rect 21548 8900 21600 8906
rect 21548 8842 21600 8848
rect 21456 8832 21508 8838
rect 21456 8774 21508 8780
rect 21560 8090 21588 8842
rect 21548 8084 21600 8090
rect 21548 8026 21600 8032
rect 21560 7410 21588 8026
rect 21548 7404 21600 7410
rect 21548 7346 21600 7352
rect 21364 6928 21416 6934
rect 21364 6870 21416 6876
rect 21364 6792 21416 6798
rect 21008 6718 21128 6746
rect 21364 6734 21416 6740
rect 21548 6792 21600 6798
rect 21548 6734 21600 6740
rect 20996 6656 21048 6662
rect 20996 6598 21048 6604
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 20824 5766 20944 5794
rect 20720 5364 20772 5370
rect 20720 5306 20772 5312
rect 20720 4820 20772 4826
rect 20640 4780 20720 4808
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 20640 4078 20668 4780
rect 20916 4808 20944 5766
rect 21008 5574 21036 6598
rect 20996 5568 21048 5574
rect 20996 5510 21048 5516
rect 21008 4826 21036 5510
rect 21100 5370 21128 6718
rect 21376 6633 21404 6734
rect 21362 6624 21418 6633
rect 21362 6559 21418 6568
rect 21376 5914 21404 6559
rect 21364 5908 21416 5914
rect 21364 5850 21416 5856
rect 21560 5778 21588 6734
rect 21652 6458 21680 12038
rect 21744 11626 21772 22102
rect 21822 21992 21878 22001
rect 21822 21927 21878 21936
rect 21836 20602 21864 21927
rect 21824 20596 21876 20602
rect 21824 20538 21876 20544
rect 21824 19372 21876 19378
rect 21824 19314 21876 19320
rect 21836 18970 21864 19314
rect 21928 19009 21956 22918
rect 22112 22166 22140 23310
rect 22100 22160 22152 22166
rect 22100 22102 22152 22108
rect 22008 22092 22060 22098
rect 22008 22034 22060 22040
rect 22020 21690 22048 22034
rect 22112 21690 22140 22102
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 22100 21684 22152 21690
rect 22100 21626 22152 21632
rect 22008 21480 22060 21486
rect 22100 21480 22152 21486
rect 22008 21422 22060 21428
rect 22098 21448 22100 21457
rect 22152 21448 22154 21457
rect 22020 21332 22048 21422
rect 22098 21383 22154 21392
rect 22020 21304 22140 21332
rect 22112 20058 22140 21304
rect 22100 20052 22152 20058
rect 22100 19994 22152 20000
rect 22008 19916 22060 19922
rect 22008 19858 22060 19864
rect 21914 19000 21970 19009
rect 21824 18964 21876 18970
rect 21914 18935 21970 18944
rect 21824 18906 21876 18912
rect 21824 18828 21876 18834
rect 21824 18770 21876 18776
rect 21836 18057 21864 18770
rect 21916 18692 21968 18698
rect 21916 18634 21968 18640
rect 21928 18329 21956 18634
rect 22020 18578 22048 19858
rect 22204 18970 22232 23831
rect 22284 22432 22336 22438
rect 22284 22374 22336 22380
rect 22296 22234 22324 22374
rect 22284 22228 22336 22234
rect 22284 22170 22336 22176
rect 22388 22137 22416 27520
rect 22928 25492 22980 25498
rect 22928 25434 22980 25440
rect 22744 25356 22796 25362
rect 22744 25298 22796 25304
rect 22650 25120 22706 25129
rect 22650 25055 22706 25064
rect 22560 24064 22612 24070
rect 22560 24006 22612 24012
rect 22468 23520 22520 23526
rect 22468 23462 22520 23468
rect 22480 23118 22508 23462
rect 22468 23112 22520 23118
rect 22468 23054 22520 23060
rect 22374 22128 22430 22137
rect 22374 22063 22430 22072
rect 22284 22024 22336 22030
rect 22282 21992 22284 22001
rect 22336 21992 22338 22001
rect 22282 21927 22338 21936
rect 22296 21622 22324 21927
rect 22480 21894 22508 23054
rect 22468 21888 22520 21894
rect 22468 21830 22520 21836
rect 22284 21616 22336 21622
rect 22284 21558 22336 21564
rect 22376 21548 22428 21554
rect 22376 21490 22428 21496
rect 22282 21448 22338 21457
rect 22282 21383 22338 21392
rect 22296 21078 22324 21383
rect 22284 21072 22336 21078
rect 22284 21014 22336 21020
rect 22388 20942 22416 21490
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22284 20800 22336 20806
rect 22282 20768 22284 20777
rect 22336 20768 22338 20777
rect 22282 20703 22338 20712
rect 22388 20466 22416 20878
rect 22376 20460 22428 20466
rect 22376 20402 22428 20408
rect 22284 20324 22336 20330
rect 22284 20266 22336 20272
rect 22376 20324 22428 20330
rect 22376 20266 22428 20272
rect 22296 19378 22324 20266
rect 22284 19372 22336 19378
rect 22284 19314 22336 19320
rect 22192 18964 22244 18970
rect 22192 18906 22244 18912
rect 22100 18828 22152 18834
rect 22100 18770 22152 18776
rect 22112 18578 22140 18770
rect 22020 18550 22140 18578
rect 21914 18320 21970 18329
rect 21914 18255 21970 18264
rect 21914 18184 21970 18193
rect 21914 18119 21970 18128
rect 21822 18048 21878 18057
rect 21822 17983 21878 17992
rect 21822 17912 21878 17921
rect 21822 17847 21878 17856
rect 21836 17814 21864 17847
rect 21824 17808 21876 17814
rect 21824 17750 21876 17756
rect 21824 17128 21876 17134
rect 21824 17070 21876 17076
rect 21836 13870 21864 17070
rect 21928 16250 21956 18119
rect 22020 17882 22048 18550
rect 22100 18352 22152 18358
rect 22100 18294 22152 18300
rect 22008 17876 22060 17882
rect 22008 17818 22060 17824
rect 22006 17776 22062 17785
rect 22006 17711 22062 17720
rect 22020 17610 22048 17711
rect 22008 17604 22060 17610
rect 22008 17546 22060 17552
rect 22008 16992 22060 16998
rect 22008 16934 22060 16940
rect 21916 16244 21968 16250
rect 21916 16186 21968 16192
rect 22020 15910 22048 16934
rect 22112 16250 22140 18294
rect 22204 17882 22232 18906
rect 22284 18624 22336 18630
rect 22388 18601 22416 20266
rect 22284 18566 22336 18572
rect 22374 18592 22430 18601
rect 22296 18358 22324 18566
rect 22374 18527 22430 18536
rect 22284 18352 22336 18358
rect 22284 18294 22336 18300
rect 22192 17876 22244 17882
rect 22192 17818 22244 17824
rect 22376 17740 22428 17746
rect 22376 17682 22428 17688
rect 22388 17513 22416 17682
rect 22374 17504 22430 17513
rect 22374 17439 22430 17448
rect 22376 17332 22428 17338
rect 22376 17274 22428 17280
rect 22388 16794 22416 17274
rect 22376 16788 22428 16794
rect 22376 16730 22428 16736
rect 22480 16674 22508 21830
rect 22296 16646 22508 16674
rect 22100 16244 22152 16250
rect 22100 16186 22152 16192
rect 22100 15972 22152 15978
rect 22100 15914 22152 15920
rect 22008 15904 22060 15910
rect 22008 15846 22060 15852
rect 22112 15706 22140 15914
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 22204 15706 22232 15846
rect 22100 15700 22152 15706
rect 22100 15642 22152 15648
rect 22192 15700 22244 15706
rect 22192 15642 22244 15648
rect 22296 15586 22324 16646
rect 22376 16584 22428 16590
rect 22376 16526 22428 16532
rect 22008 15564 22060 15570
rect 22008 15506 22060 15512
rect 22112 15558 22324 15586
rect 22020 15162 22048 15506
rect 22008 15156 22060 15162
rect 22008 15098 22060 15104
rect 22008 14272 22060 14278
rect 22008 14214 22060 14220
rect 21824 13864 21876 13870
rect 21824 13806 21876 13812
rect 22020 13530 22048 14214
rect 22008 13524 22060 13530
rect 21928 13484 22008 13512
rect 21928 12986 21956 13484
rect 22008 13466 22060 13472
rect 21916 12980 21968 12986
rect 21916 12922 21968 12928
rect 21822 12880 21878 12889
rect 21822 12815 21878 12824
rect 21836 11898 21864 12815
rect 21928 12374 21956 12922
rect 21916 12368 21968 12374
rect 21916 12310 21968 12316
rect 22006 12336 22062 12345
rect 22006 12271 22062 12280
rect 21916 12232 21968 12238
rect 21916 12174 21968 12180
rect 21824 11892 21876 11898
rect 21824 11834 21876 11840
rect 21732 11620 21784 11626
rect 21732 11562 21784 11568
rect 21824 11552 21876 11558
rect 21824 11494 21876 11500
rect 21836 10690 21864 11494
rect 21744 10662 21864 10690
rect 21744 8401 21772 10662
rect 21928 9654 21956 12174
rect 22020 12102 22048 12271
rect 22008 12096 22060 12102
rect 22008 12038 22060 12044
rect 22008 11756 22060 11762
rect 22008 11698 22060 11704
rect 22020 11354 22048 11698
rect 22008 11348 22060 11354
rect 22008 11290 22060 11296
rect 22006 10976 22062 10985
rect 22006 10911 22062 10920
rect 22020 10742 22048 10911
rect 22008 10736 22060 10742
rect 22008 10678 22060 10684
rect 21824 9648 21876 9654
rect 21824 9590 21876 9596
rect 21916 9648 21968 9654
rect 21916 9590 21968 9596
rect 21836 8974 21864 9590
rect 21824 8968 21876 8974
rect 21824 8910 21876 8916
rect 21730 8392 21786 8401
rect 21730 8327 21786 8336
rect 21732 8288 21784 8294
rect 21836 8276 21864 8910
rect 22008 8832 22060 8838
rect 22008 8774 22060 8780
rect 22020 8498 22048 8774
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 21784 8248 21864 8276
rect 21916 8288 21968 8294
rect 21732 8230 21784 8236
rect 21916 8230 21968 8236
rect 21744 7886 21772 8230
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 21640 6452 21692 6458
rect 21640 6394 21692 6400
rect 21652 6186 21680 6394
rect 21640 6180 21692 6186
rect 21640 6122 21692 6128
rect 21548 5772 21600 5778
rect 21548 5714 21600 5720
rect 21178 5672 21234 5681
rect 21178 5607 21234 5616
rect 21088 5364 21140 5370
rect 21088 5306 21140 5312
rect 20720 4762 20772 4768
rect 20824 4780 20944 4808
rect 20996 4820 21048 4826
rect 20628 4072 20680 4078
rect 20442 4040 20498 4049
rect 20628 4014 20680 4020
rect 20442 3975 20498 3984
rect 20720 4004 20772 4010
rect 20260 2848 20312 2854
rect 20260 2790 20312 2796
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 19996 1873 20024 2450
rect 20168 2304 20220 2310
rect 20168 2246 20220 2252
rect 19982 1864 20038 1873
rect 19982 1799 20038 1808
rect 20180 1737 20208 2246
rect 20166 1728 20222 1737
rect 20166 1663 20222 1672
rect 19444 1278 19932 1306
rect 19352 598 19472 626
rect 19352 480 19380 598
rect 17590 368 17646 377
rect 17590 303 17646 312
rect 17682 0 17738 480
rect 18234 0 18290 480
rect 18786 0 18842 480
rect 19338 0 19394 480
rect 19444 241 19472 598
rect 19904 480 19932 1278
rect 20456 480 20484 3975
rect 20720 3946 20772 3952
rect 20732 3534 20760 3946
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20548 3194 20576 3470
rect 20536 3188 20588 3194
rect 20536 3130 20588 3136
rect 20824 3058 20852 4780
rect 20996 4762 21048 4768
rect 21192 4706 21220 5607
rect 21454 5264 21510 5273
rect 21454 5199 21510 5208
rect 20904 4684 20956 4690
rect 20904 4626 20956 4632
rect 21008 4678 21220 4706
rect 20916 4049 20944 4626
rect 20902 4040 20958 4049
rect 20902 3975 20958 3984
rect 20916 3738 20944 3975
rect 20904 3732 20956 3738
rect 20904 3674 20956 3680
rect 21008 3618 21036 4678
rect 21178 4448 21234 4457
rect 21178 4383 21234 4392
rect 21088 3936 21140 3942
rect 21088 3878 21140 3884
rect 20916 3590 21036 3618
rect 20812 3052 20864 3058
rect 20812 2994 20864 3000
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 20732 2650 20760 2926
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 20916 2582 20944 3590
rect 20994 3496 21050 3505
rect 20994 3431 21050 3440
rect 20904 2576 20956 2582
rect 20904 2518 20956 2524
rect 21008 480 21036 3431
rect 19430 232 19486 241
rect 19430 167 19486 176
rect 19890 0 19946 480
rect 20442 0 20498 480
rect 20994 0 21050 480
rect 21100 105 21128 3878
rect 21192 3194 21220 4383
rect 21364 3936 21416 3942
rect 21284 3896 21364 3924
rect 21284 3602 21312 3896
rect 21364 3878 21416 3884
rect 21272 3596 21324 3602
rect 21272 3538 21324 3544
rect 21284 3505 21312 3538
rect 21270 3496 21326 3505
rect 21270 3431 21326 3440
rect 21180 3188 21232 3194
rect 21180 3130 21232 3136
rect 21468 2990 21496 5199
rect 21560 3534 21588 5714
rect 21652 5574 21680 6122
rect 21744 5710 21772 7822
rect 21824 6860 21876 6866
rect 21824 6802 21876 6808
rect 21836 6118 21864 6802
rect 21928 6662 21956 8230
rect 22112 8022 22140 15558
rect 22284 15088 22336 15094
rect 22284 15030 22336 15036
rect 22192 13728 22244 13734
rect 22192 13670 22244 13676
rect 22204 13326 22232 13670
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 22296 12442 22324 15030
rect 22284 12436 22336 12442
rect 22284 12378 22336 12384
rect 22282 12336 22338 12345
rect 22282 12271 22338 12280
rect 22192 10464 22244 10470
rect 22192 10406 22244 10412
rect 22204 9994 22232 10406
rect 22192 9988 22244 9994
rect 22192 9930 22244 9936
rect 22296 9761 22324 12271
rect 22282 9752 22338 9761
rect 22282 9687 22338 9696
rect 22284 9648 22336 9654
rect 22284 9590 22336 9596
rect 22192 9376 22244 9382
rect 22192 9318 22244 9324
rect 22204 9178 22232 9318
rect 22192 9172 22244 9178
rect 22192 9114 22244 9120
rect 22192 8832 22244 8838
rect 22190 8800 22192 8809
rect 22244 8800 22246 8809
rect 22190 8735 22246 8744
rect 22190 8664 22246 8673
rect 22190 8599 22192 8608
rect 22244 8599 22246 8608
rect 22192 8570 22244 8576
rect 22296 8498 22324 9590
rect 22284 8492 22336 8498
rect 22284 8434 22336 8440
rect 22100 8016 22152 8022
rect 22100 7958 22152 7964
rect 22006 7576 22062 7585
rect 22112 7546 22140 7958
rect 22006 7511 22062 7520
rect 22100 7540 22152 7546
rect 22020 7342 22048 7511
rect 22152 7500 22232 7528
rect 22100 7482 22152 7488
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 22008 7336 22060 7342
rect 22008 7278 22060 7284
rect 21916 6656 21968 6662
rect 21916 6598 21968 6604
rect 21928 6497 21956 6598
rect 21914 6488 21970 6497
rect 22020 6458 22048 7278
rect 22112 6798 22140 7346
rect 22100 6792 22152 6798
rect 22100 6734 22152 6740
rect 21914 6423 21970 6432
rect 22008 6452 22060 6458
rect 21928 6254 21956 6423
rect 22008 6394 22060 6400
rect 21916 6248 21968 6254
rect 21916 6190 21968 6196
rect 21824 6112 21876 6118
rect 21824 6054 21876 6060
rect 21836 5846 21864 6054
rect 21824 5840 21876 5846
rect 21824 5782 21876 5788
rect 21732 5704 21784 5710
rect 21732 5646 21784 5652
rect 21640 5568 21692 5574
rect 21640 5510 21692 5516
rect 22112 5302 22140 6734
rect 22204 6662 22232 7500
rect 22284 6860 22336 6866
rect 22284 6802 22336 6808
rect 22296 6730 22324 6802
rect 22284 6724 22336 6730
rect 22284 6666 22336 6672
rect 22192 6656 22244 6662
rect 22192 6598 22244 6604
rect 22204 5914 22232 6598
rect 22192 5908 22244 5914
rect 22192 5850 22244 5856
rect 22192 5772 22244 5778
rect 22192 5714 22244 5720
rect 22204 5370 22232 5714
rect 22192 5364 22244 5370
rect 22192 5306 22244 5312
rect 22100 5296 22152 5302
rect 22100 5238 22152 5244
rect 22204 4826 22232 5306
rect 22192 4820 22244 4826
rect 22192 4762 22244 4768
rect 22100 4480 22152 4486
rect 21928 4440 22100 4468
rect 21928 3738 21956 4440
rect 22100 4422 22152 4428
rect 22296 4214 22324 6666
rect 22388 6304 22416 16526
rect 22468 16448 22520 16454
rect 22468 16390 22520 16396
rect 22480 16114 22508 16390
rect 22468 16108 22520 16114
rect 22468 16050 22520 16056
rect 22466 15192 22522 15201
rect 22466 15127 22522 15136
rect 22480 13462 22508 15127
rect 22468 13456 22520 13462
rect 22468 13398 22520 13404
rect 22480 12646 22508 13398
rect 22468 12640 22520 12646
rect 22468 12582 22520 12588
rect 22468 12436 22520 12442
rect 22468 12378 22520 12384
rect 22480 10130 22508 12378
rect 22468 10124 22520 10130
rect 22468 10066 22520 10072
rect 22480 7478 22508 10066
rect 22468 7472 22520 7478
rect 22468 7414 22520 7420
rect 22572 7410 22600 24006
rect 22664 17338 22692 25055
rect 22756 24070 22784 25298
rect 22940 25226 22968 25434
rect 23032 25430 23060 27520
rect 23386 27160 23442 27169
rect 23386 27095 23442 27104
rect 23202 26616 23258 26625
rect 23202 26551 23258 26560
rect 23020 25424 23072 25430
rect 23020 25366 23072 25372
rect 22928 25220 22980 25226
rect 22928 25162 22980 25168
rect 22836 24608 22888 24614
rect 22836 24550 22888 24556
rect 22744 24064 22796 24070
rect 22744 24006 22796 24012
rect 22756 21457 22784 24006
rect 22742 21448 22798 21457
rect 22742 21383 22798 21392
rect 22744 21344 22796 21350
rect 22744 21286 22796 21292
rect 22756 20874 22784 21286
rect 22744 20868 22796 20874
rect 22744 20810 22796 20816
rect 22756 19394 22784 20810
rect 22848 20330 22876 24550
rect 23112 24200 23164 24206
rect 23112 24142 23164 24148
rect 22928 23792 22980 23798
rect 22928 23734 22980 23740
rect 22836 20324 22888 20330
rect 22836 20266 22888 20272
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 22848 19514 22876 19858
rect 22940 19854 22968 23734
rect 23020 23520 23072 23526
rect 23020 23462 23072 23468
rect 23032 22273 23060 23462
rect 23018 22264 23074 22273
rect 23018 22199 23074 22208
rect 23018 21992 23074 22001
rect 23018 21927 23074 21936
rect 22928 19848 22980 19854
rect 22928 19790 22980 19796
rect 22836 19508 22888 19514
rect 22836 19450 22888 19456
rect 22756 19366 22876 19394
rect 22744 19304 22796 19310
rect 22744 19246 22796 19252
rect 22652 17332 22704 17338
rect 22652 17274 22704 17280
rect 22756 17048 22784 19246
rect 22664 17020 22784 17048
rect 22664 15094 22692 17020
rect 22742 16960 22798 16969
rect 22742 16895 22798 16904
rect 22756 16658 22784 16895
rect 22744 16652 22796 16658
rect 22744 16594 22796 16600
rect 22744 16176 22796 16182
rect 22744 16118 22796 16124
rect 22756 15434 22784 16118
rect 22744 15428 22796 15434
rect 22744 15370 22796 15376
rect 22756 15162 22784 15370
rect 22744 15156 22796 15162
rect 22744 15098 22796 15104
rect 22652 15088 22704 15094
rect 22652 15030 22704 15036
rect 22742 15056 22798 15065
rect 22742 14991 22798 15000
rect 22652 14952 22704 14958
rect 22652 14894 22704 14900
rect 22664 13025 22692 14894
rect 22756 14074 22784 14991
rect 22744 14068 22796 14074
rect 22744 14010 22796 14016
rect 22744 13728 22796 13734
rect 22744 13670 22796 13676
rect 22650 13016 22706 13025
rect 22650 12951 22706 12960
rect 22650 12880 22706 12889
rect 22650 12815 22706 12824
rect 22664 12714 22692 12815
rect 22652 12708 22704 12714
rect 22652 12650 22704 12656
rect 22652 12368 22704 12374
rect 22652 12310 22704 12316
rect 22560 7404 22612 7410
rect 22560 7346 22612 7352
rect 22664 7324 22692 12310
rect 22756 11354 22784 13670
rect 22848 12753 22876 19366
rect 22940 19310 22968 19790
rect 22928 19304 22980 19310
rect 22928 19246 22980 19252
rect 22926 18592 22982 18601
rect 22926 18527 22982 18536
rect 22940 16425 22968 18527
rect 22926 16416 22982 16425
rect 22926 16351 22982 16360
rect 22926 16280 22982 16289
rect 22926 16215 22982 16224
rect 22940 15366 22968 16215
rect 22928 15360 22980 15366
rect 22928 15302 22980 15308
rect 22940 14006 22968 15302
rect 23032 14074 23060 21927
rect 23124 21593 23152 24142
rect 23216 23866 23244 26551
rect 23296 25152 23348 25158
rect 23296 25094 23348 25100
rect 23308 24596 23336 25094
rect 23400 24818 23428 27095
rect 23584 25945 23612 27520
rect 23570 25936 23626 25945
rect 23570 25871 23626 25880
rect 24032 25356 24084 25362
rect 24032 25298 24084 25304
rect 23848 25288 23900 25294
rect 23848 25230 23900 25236
rect 23860 25158 23888 25230
rect 23848 25152 23900 25158
rect 23848 25094 23900 25100
rect 23860 24886 23888 25094
rect 23848 24880 23900 24886
rect 23848 24822 23900 24828
rect 23388 24812 23440 24818
rect 23388 24754 23440 24760
rect 23480 24608 23532 24614
rect 23308 24568 23480 24596
rect 23296 24064 23348 24070
rect 23296 24006 23348 24012
rect 23204 23860 23256 23866
rect 23204 23802 23256 23808
rect 23204 22636 23256 22642
rect 23204 22578 23256 22584
rect 23216 22098 23244 22578
rect 23204 22092 23256 22098
rect 23204 22034 23256 22040
rect 23204 21956 23256 21962
rect 23204 21898 23256 21904
rect 23216 21690 23244 21898
rect 23204 21684 23256 21690
rect 23204 21626 23256 21632
rect 23110 21584 23166 21593
rect 23110 21519 23166 21528
rect 23204 20460 23256 20466
rect 23204 20402 23256 20408
rect 23112 20256 23164 20262
rect 23112 20198 23164 20204
rect 23124 20097 23152 20198
rect 23110 20088 23166 20097
rect 23110 20023 23166 20032
rect 23216 19854 23244 20402
rect 23308 19854 23336 24006
rect 23400 23633 23428 24568
rect 23480 24550 23532 24556
rect 23756 24608 23808 24614
rect 23756 24550 23808 24556
rect 23480 24132 23532 24138
rect 23480 24074 23532 24080
rect 23386 23624 23442 23633
rect 23386 23559 23442 23568
rect 23388 22976 23440 22982
rect 23492 22964 23520 24074
rect 23572 24064 23624 24070
rect 23572 24006 23624 24012
rect 23440 22936 23520 22964
rect 23388 22918 23440 22924
rect 23400 21554 23428 22918
rect 23480 22432 23532 22438
rect 23480 22374 23532 22380
rect 23492 22273 23520 22374
rect 23478 22264 23534 22273
rect 23478 22199 23534 22208
rect 23480 22024 23532 22030
rect 23480 21966 23532 21972
rect 23388 21548 23440 21554
rect 23388 21490 23440 21496
rect 23492 21350 23520 21966
rect 23480 21344 23532 21350
rect 23480 21286 23532 21292
rect 23388 21140 23440 21146
rect 23388 21082 23440 21088
rect 23400 20369 23428 21082
rect 23492 21049 23520 21286
rect 23478 21040 23534 21049
rect 23478 20975 23534 20984
rect 23386 20360 23442 20369
rect 23386 20295 23442 20304
rect 23480 20256 23532 20262
rect 23480 20198 23532 20204
rect 23492 19922 23520 20198
rect 23480 19916 23532 19922
rect 23480 19858 23532 19864
rect 23204 19848 23256 19854
rect 23204 19790 23256 19796
rect 23296 19848 23348 19854
rect 23296 19790 23348 19796
rect 23216 19145 23244 19790
rect 23388 19780 23440 19786
rect 23388 19722 23440 19728
rect 23296 19168 23348 19174
rect 23202 19136 23258 19145
rect 23296 19110 23348 19116
rect 23202 19071 23258 19080
rect 23216 18902 23244 19071
rect 23204 18896 23256 18902
rect 23204 18838 23256 18844
rect 23308 18766 23336 19110
rect 23112 18760 23164 18766
rect 23112 18702 23164 18708
rect 23296 18760 23348 18766
rect 23296 18702 23348 18708
rect 23124 18358 23152 18702
rect 23308 18601 23336 18702
rect 23294 18592 23350 18601
rect 23294 18527 23350 18536
rect 23400 18426 23428 19722
rect 23478 19680 23534 19689
rect 23478 19615 23534 19624
rect 23492 18970 23520 19615
rect 23480 18964 23532 18970
rect 23480 18906 23532 18912
rect 23480 18828 23532 18834
rect 23480 18770 23532 18776
rect 23388 18420 23440 18426
rect 23388 18362 23440 18368
rect 23112 18352 23164 18358
rect 23112 18294 23164 18300
rect 23294 18320 23350 18329
rect 23124 18086 23152 18294
rect 23294 18255 23350 18264
rect 23112 18080 23164 18086
rect 23112 18022 23164 18028
rect 23124 17524 23152 18022
rect 23308 17882 23336 18255
rect 23296 17876 23348 17882
rect 23296 17818 23348 17824
rect 23204 17740 23256 17746
rect 23204 17682 23256 17688
rect 23216 17649 23244 17682
rect 23202 17640 23258 17649
rect 23202 17575 23258 17584
rect 23124 17496 23244 17524
rect 23110 17232 23166 17241
rect 23110 17167 23112 17176
rect 23164 17167 23166 17176
rect 23112 17138 23164 17144
rect 23110 16960 23166 16969
rect 23110 16895 23166 16904
rect 23124 14958 23152 16895
rect 23112 14952 23164 14958
rect 23112 14894 23164 14900
rect 23112 14816 23164 14822
rect 23112 14758 23164 14764
rect 23124 14414 23152 14758
rect 23112 14408 23164 14414
rect 23112 14350 23164 14356
rect 23110 14104 23166 14113
rect 23020 14068 23072 14074
rect 23110 14039 23166 14048
rect 23020 14010 23072 14016
rect 22928 14000 22980 14006
rect 22928 13942 22980 13948
rect 22940 13530 22968 13942
rect 23032 13870 23060 14010
rect 23020 13864 23072 13870
rect 23020 13806 23072 13812
rect 22928 13524 22980 13530
rect 22928 13466 22980 13472
rect 23124 13394 23152 14039
rect 23216 13569 23244 17496
rect 23308 17241 23336 17818
rect 23388 17672 23440 17678
rect 23388 17614 23440 17620
rect 23294 17232 23350 17241
rect 23294 17167 23350 17176
rect 23296 16992 23348 16998
rect 23296 16934 23348 16940
rect 23308 16522 23336 16934
rect 23400 16833 23428 17614
rect 23492 17610 23520 18770
rect 23480 17604 23532 17610
rect 23480 17546 23532 17552
rect 23480 17060 23532 17066
rect 23480 17002 23532 17008
rect 23386 16824 23442 16833
rect 23386 16759 23388 16768
rect 23440 16759 23442 16768
rect 23388 16730 23440 16736
rect 23400 16699 23428 16730
rect 23296 16516 23348 16522
rect 23296 16458 23348 16464
rect 23308 15162 23336 16458
rect 23386 16416 23442 16425
rect 23386 16351 23442 16360
rect 23400 16250 23428 16351
rect 23492 16250 23520 17002
rect 23584 16561 23612 24006
rect 23664 23520 23716 23526
rect 23664 23462 23716 23468
rect 23676 21078 23704 23462
rect 23768 21690 23796 24550
rect 23848 24268 23900 24274
rect 23848 24210 23900 24216
rect 23860 24177 23888 24210
rect 23846 24168 23902 24177
rect 24044 24138 24072 25298
rect 24136 24857 24164 27520
rect 24674 25936 24730 25945
rect 24674 25871 24730 25880
rect 24216 25152 24268 25158
rect 24216 25094 24268 25100
rect 24122 24848 24178 24857
rect 24122 24783 24178 24792
rect 24124 24676 24176 24682
rect 24124 24618 24176 24624
rect 23846 24103 23902 24112
rect 24032 24132 24084 24138
rect 24032 24074 24084 24080
rect 24136 24070 24164 24618
rect 24124 24064 24176 24070
rect 24122 24032 24124 24041
rect 24176 24032 24178 24041
rect 24122 23967 24178 23976
rect 24228 23866 24256 25094
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24688 24954 24716 25871
rect 24780 25430 24808 27520
rect 25136 25968 25188 25974
rect 25136 25910 25188 25916
rect 24768 25424 24820 25430
rect 24768 25366 24820 25372
rect 24768 25288 24820 25294
rect 24768 25230 24820 25236
rect 24676 24948 24728 24954
rect 24676 24890 24728 24896
rect 24780 24596 24808 25230
rect 24860 24608 24912 24614
rect 24780 24576 24860 24596
rect 24912 24576 24914 24585
rect 24780 24568 24858 24576
rect 24858 24511 24914 24520
rect 25044 24268 25096 24274
rect 25044 24210 25096 24216
rect 24952 24200 25004 24206
rect 24952 24142 25004 24148
rect 24860 24132 24912 24138
rect 24860 24074 24912 24080
rect 24676 24064 24728 24070
rect 24872 24018 24900 24074
rect 24676 24006 24728 24012
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24216 23860 24268 23866
rect 24216 23802 24268 23808
rect 24308 23724 24360 23730
rect 24308 23666 24360 23672
rect 24320 23633 24348 23666
rect 24306 23624 24362 23633
rect 24124 23588 24176 23594
rect 24306 23559 24362 23568
rect 24124 23530 24176 23536
rect 24136 23497 24164 23530
rect 24308 23520 24360 23526
rect 24122 23488 24178 23497
rect 24308 23462 24360 23468
rect 24122 23423 24178 23432
rect 24320 23254 24348 23462
rect 24308 23248 24360 23254
rect 24308 23190 24360 23196
rect 23848 23180 23900 23186
rect 23848 23122 23900 23128
rect 23860 22710 23888 23122
rect 23940 23112 23992 23118
rect 23940 23054 23992 23060
rect 24124 23112 24176 23118
rect 24124 23054 24176 23060
rect 23848 22704 23900 22710
rect 23848 22646 23900 22652
rect 23846 22536 23902 22545
rect 23846 22471 23902 22480
rect 23756 21684 23808 21690
rect 23756 21626 23808 21632
rect 23664 21072 23716 21078
rect 23664 21014 23716 21020
rect 23756 21004 23808 21010
rect 23756 20946 23808 20952
rect 23664 20936 23716 20942
rect 23664 20878 23716 20884
rect 23676 20398 23704 20878
rect 23664 20392 23716 20398
rect 23664 20334 23716 20340
rect 23676 19514 23704 20334
rect 23768 20262 23796 20946
rect 23756 20256 23808 20262
rect 23756 20198 23808 20204
rect 23664 19508 23716 19514
rect 23664 19450 23716 19456
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 23676 18290 23704 18906
rect 23754 18456 23810 18465
rect 23754 18391 23756 18400
rect 23808 18391 23810 18400
rect 23756 18362 23808 18368
rect 23664 18284 23716 18290
rect 23664 18226 23716 18232
rect 23860 18222 23888 22471
rect 23952 22234 23980 23054
rect 24136 22642 24164 23054
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24124 22636 24176 22642
rect 24124 22578 24176 22584
rect 24492 22636 24544 22642
rect 24492 22578 24544 22584
rect 24400 22500 24452 22506
rect 24400 22442 24452 22448
rect 24412 22409 24440 22442
rect 24398 22400 24454 22409
rect 24398 22335 24454 22344
rect 23940 22228 23992 22234
rect 23940 22170 23992 22176
rect 24124 22160 24176 22166
rect 24122 22128 24124 22137
rect 24176 22128 24178 22137
rect 23940 22092 23992 22098
rect 24122 22063 24178 22072
rect 24398 22128 24454 22137
rect 24504 22114 24532 22578
rect 24454 22086 24532 22114
rect 24398 22063 24454 22072
rect 23940 22034 23992 22040
rect 23952 21457 23980 22034
rect 24412 22030 24440 22063
rect 24400 22024 24452 22030
rect 24400 21966 24452 21972
rect 24688 21894 24716 24006
rect 24780 23990 24900 24018
rect 24780 23050 24808 23990
rect 24860 23860 24912 23866
rect 24860 23802 24912 23808
rect 24768 23044 24820 23050
rect 24768 22986 24820 22992
rect 24872 22760 24900 23802
rect 24964 23798 24992 24142
rect 24952 23792 25004 23798
rect 24952 23734 25004 23740
rect 25056 23730 25084 24210
rect 25044 23724 25096 23730
rect 25044 23666 25096 23672
rect 25148 23202 25176 25910
rect 25332 24721 25360 27520
rect 25778 26208 25834 26217
rect 25778 26143 25834 26152
rect 25410 25392 25466 25401
rect 25594 25392 25650 25401
rect 25466 25350 25544 25378
rect 25410 25327 25466 25336
rect 25410 24848 25466 24857
rect 25410 24783 25466 24792
rect 25318 24712 25374 24721
rect 25318 24647 25374 24656
rect 25320 24608 25372 24614
rect 25320 24550 25372 24556
rect 25332 24206 25360 24550
rect 25320 24200 25372 24206
rect 25226 24168 25282 24177
rect 25320 24142 25372 24148
rect 25226 24103 25282 24112
rect 25240 23322 25268 24103
rect 25424 23866 25452 24783
rect 25412 23860 25464 23866
rect 25412 23802 25464 23808
rect 25228 23316 25280 23322
rect 25228 23258 25280 23264
rect 25044 23180 25096 23186
rect 25148 23174 25360 23202
rect 25044 23122 25096 23128
rect 25056 23089 25084 23122
rect 25042 23080 25098 23089
rect 25042 23015 25098 23024
rect 25056 22778 25084 23015
rect 25044 22772 25096 22778
rect 24872 22732 24992 22760
rect 24768 22704 24820 22710
rect 24820 22652 24900 22658
rect 24768 22646 24900 22652
rect 24780 22630 24900 22646
rect 24766 22536 24822 22545
rect 24766 22471 24822 22480
rect 24216 21888 24268 21894
rect 24216 21830 24268 21836
rect 24676 21888 24728 21894
rect 24676 21830 24728 21836
rect 24228 21486 24256 21830
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24676 21684 24728 21690
rect 24676 21626 24728 21632
rect 24216 21480 24268 21486
rect 23938 21448 23994 21457
rect 24216 21422 24268 21428
rect 23938 21383 23994 21392
rect 23940 21344 23992 21350
rect 23940 21286 23992 21292
rect 23952 19990 23980 21286
rect 24032 21004 24084 21010
rect 24032 20946 24084 20952
rect 24044 20058 24072 20946
rect 24124 20868 24176 20874
rect 24124 20810 24176 20816
rect 24136 20466 24164 20810
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24216 20528 24268 20534
rect 24584 20528 24636 20534
rect 24268 20488 24348 20516
rect 24216 20470 24268 20476
rect 24124 20460 24176 20466
rect 24124 20402 24176 20408
rect 24032 20052 24084 20058
rect 24032 19994 24084 20000
rect 23940 19984 23992 19990
rect 23940 19926 23992 19932
rect 24032 19916 24084 19922
rect 24032 19858 24084 19864
rect 23940 19372 23992 19378
rect 23940 19314 23992 19320
rect 23952 18902 23980 19314
rect 23940 18896 23992 18902
rect 23940 18838 23992 18844
rect 23848 18216 23900 18222
rect 23848 18158 23900 18164
rect 23756 18148 23808 18154
rect 23756 18090 23808 18096
rect 23768 17762 23796 18090
rect 23860 17882 23888 18158
rect 23938 18048 23994 18057
rect 23938 17983 23994 17992
rect 23848 17876 23900 17882
rect 23848 17818 23900 17824
rect 23768 17734 23888 17762
rect 23754 17368 23810 17377
rect 23754 17303 23756 17312
rect 23808 17303 23810 17312
rect 23756 17274 23808 17280
rect 23664 17196 23716 17202
rect 23664 17138 23716 17144
rect 23676 16794 23704 17138
rect 23756 16992 23808 16998
rect 23756 16934 23808 16940
rect 23664 16788 23716 16794
rect 23664 16730 23716 16736
rect 23662 16688 23718 16697
rect 23662 16623 23718 16632
rect 23570 16552 23626 16561
rect 23570 16487 23626 16496
rect 23388 16244 23440 16250
rect 23388 16186 23440 16192
rect 23480 16244 23532 16250
rect 23480 16186 23532 16192
rect 23388 16108 23440 16114
rect 23388 16050 23440 16056
rect 23296 15156 23348 15162
rect 23296 15098 23348 15104
rect 23400 14278 23428 16050
rect 23480 16040 23532 16046
rect 23480 15982 23532 15988
rect 23492 15094 23520 15982
rect 23572 15972 23624 15978
rect 23572 15914 23624 15920
rect 23584 15706 23612 15914
rect 23572 15700 23624 15706
rect 23572 15642 23624 15648
rect 23676 15144 23704 16623
rect 23584 15116 23704 15144
rect 23480 15088 23532 15094
rect 23480 15030 23532 15036
rect 23478 14920 23534 14929
rect 23478 14855 23534 14864
rect 23388 14272 23440 14278
rect 23388 14214 23440 14220
rect 23492 13818 23520 14855
rect 23296 13796 23348 13802
rect 23296 13738 23348 13744
rect 23400 13790 23520 13818
rect 23202 13560 23258 13569
rect 23202 13495 23258 13504
rect 23308 13462 23336 13738
rect 23296 13456 23348 13462
rect 23296 13398 23348 13404
rect 23112 13388 23164 13394
rect 23032 13348 23112 13376
rect 22928 13184 22980 13190
rect 22928 13126 22980 13132
rect 22940 12986 22968 13126
rect 22928 12980 22980 12986
rect 22928 12922 22980 12928
rect 22926 12880 22982 12889
rect 23032 12850 23060 13348
rect 23112 13330 23164 13336
rect 23202 13152 23258 13161
rect 23202 13087 23258 13096
rect 22926 12815 22982 12824
rect 23020 12844 23072 12850
rect 22834 12744 22890 12753
rect 22834 12679 22890 12688
rect 22836 12640 22888 12646
rect 22836 12582 22888 12588
rect 22848 11762 22876 12582
rect 22836 11756 22888 11762
rect 22836 11698 22888 11704
rect 22836 11620 22888 11626
rect 22836 11562 22888 11568
rect 22744 11348 22796 11354
rect 22744 11290 22796 11296
rect 22744 11212 22796 11218
rect 22744 11154 22796 11160
rect 22756 10742 22784 11154
rect 22744 10736 22796 10742
rect 22742 10704 22744 10713
rect 22796 10704 22798 10713
rect 22742 10639 22798 10648
rect 22742 10296 22798 10305
rect 22742 10231 22744 10240
rect 22796 10231 22798 10240
rect 22744 10202 22796 10208
rect 22744 10124 22796 10130
rect 22744 10066 22796 10072
rect 22756 9722 22784 10066
rect 22744 9716 22796 9722
rect 22744 9658 22796 9664
rect 22756 9518 22784 9658
rect 22744 9512 22796 9518
rect 22744 9454 22796 9460
rect 22848 9217 22876 11562
rect 22834 9208 22890 9217
rect 22834 9143 22890 9152
rect 22940 9110 22968 12815
rect 23020 12786 23072 12792
rect 23112 12776 23164 12782
rect 23112 12718 23164 12724
rect 23020 12708 23072 12714
rect 23020 12650 23072 12656
rect 23032 12306 23060 12650
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 23032 11762 23060 12242
rect 23020 11756 23072 11762
rect 23020 11698 23072 11704
rect 23018 11656 23074 11665
rect 23018 11591 23074 11600
rect 23032 11354 23060 11591
rect 23020 11348 23072 11354
rect 23020 11290 23072 11296
rect 23020 11212 23072 11218
rect 23020 11154 23072 11160
rect 23032 10266 23060 11154
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 23020 10056 23072 10062
rect 23018 10024 23020 10033
rect 23072 10024 23074 10033
rect 23018 9959 23074 9968
rect 23020 9920 23072 9926
rect 23020 9862 23072 9868
rect 22928 9104 22980 9110
rect 22928 9046 22980 9052
rect 22940 8634 22968 9046
rect 23032 8838 23060 9862
rect 23020 8832 23072 8838
rect 23020 8774 23072 8780
rect 22928 8628 22980 8634
rect 22928 8570 22980 8576
rect 22834 8120 22890 8129
rect 22940 8090 22968 8570
rect 22834 8055 22890 8064
rect 22928 8084 22980 8090
rect 22664 7296 22784 7324
rect 22652 7200 22704 7206
rect 22652 7142 22704 7148
rect 22664 6934 22692 7142
rect 22652 6928 22704 6934
rect 22466 6896 22522 6905
rect 22652 6870 22704 6876
rect 22466 6831 22522 6840
rect 22480 6730 22508 6831
rect 22468 6724 22520 6730
rect 22468 6666 22520 6672
rect 22388 6276 22508 6304
rect 22376 6180 22428 6186
rect 22376 6122 22428 6128
rect 22388 4622 22416 6122
rect 22376 4616 22428 4622
rect 22376 4558 22428 4564
rect 22284 4208 22336 4214
rect 22098 4176 22154 4185
rect 22284 4150 22336 4156
rect 22388 4146 22416 4558
rect 22098 4111 22154 4120
rect 22376 4140 22428 4146
rect 21916 3732 21968 3738
rect 21916 3674 21968 3680
rect 21640 3664 21692 3670
rect 21640 3606 21692 3612
rect 21548 3528 21600 3534
rect 21548 3470 21600 3476
rect 21546 3088 21602 3097
rect 21652 3058 21680 3606
rect 21546 3023 21602 3032
rect 21640 3052 21692 3058
rect 21456 2984 21508 2990
rect 21456 2926 21508 2932
rect 21560 480 21588 3023
rect 21640 2994 21692 3000
rect 21638 2680 21694 2689
rect 21638 2615 21640 2624
rect 21692 2615 21694 2624
rect 21640 2586 21692 2592
rect 21732 2440 21784 2446
rect 21730 2408 21732 2417
rect 21784 2408 21786 2417
rect 21730 2343 21786 2352
rect 22112 480 22140 4111
rect 22376 4082 22428 4088
rect 22388 3738 22416 4082
rect 22376 3732 22428 3738
rect 22376 3674 22428 3680
rect 22480 3602 22508 6276
rect 22468 3596 22520 3602
rect 22468 3538 22520 3544
rect 22756 2650 22784 7296
rect 22848 3652 22876 8055
rect 22928 8026 22980 8032
rect 22928 6792 22980 6798
rect 22928 6734 22980 6740
rect 22940 6118 22968 6734
rect 22928 6112 22980 6118
rect 22928 6054 22980 6060
rect 22940 5778 22968 6054
rect 22928 5772 22980 5778
rect 22928 5714 22980 5720
rect 22940 4826 22968 5714
rect 23020 5024 23072 5030
rect 23020 4966 23072 4972
rect 22928 4820 22980 4826
rect 22928 4762 22980 4768
rect 22940 4282 22968 4762
rect 22928 4276 22980 4282
rect 22928 4218 22980 4224
rect 23032 3738 23060 4966
rect 23124 4758 23152 12718
rect 23216 11898 23244 13087
rect 23296 12708 23348 12714
rect 23296 12650 23348 12656
rect 23204 11892 23256 11898
rect 23204 11834 23256 11840
rect 23204 11688 23256 11694
rect 23202 11656 23204 11665
rect 23256 11656 23258 11665
rect 23202 11591 23258 11600
rect 23204 11348 23256 11354
rect 23204 11290 23256 11296
rect 23216 10130 23244 11290
rect 23308 11082 23336 12650
rect 23400 12306 23428 13790
rect 23480 13388 23532 13394
rect 23480 13330 23532 13336
rect 23492 12986 23520 13330
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23584 12714 23612 15116
rect 23664 15020 23716 15026
rect 23664 14962 23716 14968
rect 23676 14550 23704 14962
rect 23664 14544 23716 14550
rect 23664 14486 23716 14492
rect 23662 14240 23718 14249
rect 23662 14175 23718 14184
rect 23676 14074 23704 14175
rect 23664 14068 23716 14074
rect 23664 14010 23716 14016
rect 23662 13560 23718 13569
rect 23662 13495 23718 13504
rect 23572 12708 23624 12714
rect 23572 12650 23624 12656
rect 23676 12594 23704 13495
rect 23584 12566 23704 12594
rect 23388 12300 23440 12306
rect 23388 12242 23440 12248
rect 23584 12209 23612 12566
rect 23662 12472 23718 12481
rect 23662 12407 23718 12416
rect 23570 12200 23626 12209
rect 23570 12135 23626 12144
rect 23386 11928 23442 11937
rect 23386 11863 23442 11872
rect 23572 11892 23624 11898
rect 23400 11286 23428 11863
rect 23572 11834 23624 11840
rect 23388 11280 23440 11286
rect 23388 11222 23440 11228
rect 23480 11144 23532 11150
rect 23400 11092 23480 11098
rect 23400 11086 23532 11092
rect 23296 11076 23348 11082
rect 23296 11018 23348 11024
rect 23400 11070 23520 11086
rect 23296 10668 23348 10674
rect 23296 10610 23348 10616
rect 23204 10124 23256 10130
rect 23204 10066 23256 10072
rect 23202 9752 23258 9761
rect 23202 9687 23258 9696
rect 23216 6798 23244 9687
rect 23308 7954 23336 10610
rect 23400 10418 23428 11070
rect 23480 11008 23532 11014
rect 23478 10976 23480 10985
rect 23532 10976 23534 10985
rect 23478 10911 23534 10920
rect 23492 10606 23520 10911
rect 23584 10810 23612 11834
rect 23572 10804 23624 10810
rect 23572 10746 23624 10752
rect 23480 10600 23532 10606
rect 23480 10542 23532 10548
rect 23400 10390 23612 10418
rect 23584 10130 23612 10390
rect 23572 10124 23624 10130
rect 23572 10066 23624 10072
rect 23388 9988 23440 9994
rect 23388 9930 23440 9936
rect 23400 9602 23428 9930
rect 23400 9574 23520 9602
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 23296 7948 23348 7954
rect 23296 7890 23348 7896
rect 23296 7404 23348 7410
rect 23296 7346 23348 7352
rect 23204 6792 23256 6798
rect 23204 6734 23256 6740
rect 23202 5944 23258 5953
rect 23202 5879 23258 5888
rect 23112 4752 23164 4758
rect 23112 4694 23164 4700
rect 23124 4146 23152 4694
rect 23112 4140 23164 4146
rect 23112 4082 23164 4088
rect 23020 3732 23072 3738
rect 23020 3674 23072 3680
rect 22928 3664 22980 3670
rect 22848 3632 22928 3652
rect 22980 3632 22982 3641
rect 22848 3624 22926 3632
rect 22926 3567 22982 3576
rect 22928 3528 22980 3534
rect 22928 3470 22980 3476
rect 22940 3058 22968 3470
rect 23124 3097 23152 4082
rect 23110 3088 23166 3097
rect 22928 3052 22980 3058
rect 22928 2994 22980 3000
rect 23020 3052 23072 3058
rect 23110 3023 23166 3032
rect 23020 2994 23072 3000
rect 23032 2854 23060 2994
rect 23020 2848 23072 2854
rect 23020 2790 23072 2796
rect 22744 2644 22796 2650
rect 22744 2586 22796 2592
rect 23032 2446 23060 2790
rect 23020 2440 23072 2446
rect 23020 2382 23072 2388
rect 23020 2304 23072 2310
rect 23020 2246 23072 2252
rect 22742 1864 22798 1873
rect 22742 1799 22798 1808
rect 22756 610 22784 1799
rect 23032 1465 23060 2246
rect 23018 1456 23074 1465
rect 23018 1391 23074 1400
rect 22652 604 22704 610
rect 22652 546 22704 552
rect 22744 604 22796 610
rect 22744 546 22796 552
rect 22664 480 22692 546
rect 23216 480 23244 5879
rect 23308 4690 23336 7346
rect 23400 5710 23428 9454
rect 23492 7546 23520 9574
rect 23584 9518 23612 10066
rect 23572 9512 23624 9518
rect 23572 9454 23624 9460
rect 23584 9042 23612 9454
rect 23572 9036 23624 9042
rect 23572 8978 23624 8984
rect 23676 8634 23704 12407
rect 23664 8628 23716 8634
rect 23664 8570 23716 8576
rect 23662 8528 23718 8537
rect 23662 8463 23718 8472
rect 23572 8356 23624 8362
rect 23572 8298 23624 8304
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 23480 7200 23532 7206
rect 23478 7168 23480 7177
rect 23532 7168 23534 7177
rect 23478 7103 23534 7112
rect 23478 6216 23534 6225
rect 23478 6151 23480 6160
rect 23532 6151 23534 6160
rect 23480 6122 23532 6128
rect 23478 5808 23534 5817
rect 23584 5794 23612 8298
rect 23676 6254 23704 8463
rect 23768 8022 23796 16934
rect 23860 16590 23888 17734
rect 23952 17678 23980 17983
rect 24044 17921 24072 19858
rect 24136 18970 24164 20402
rect 24216 20256 24268 20262
rect 24216 20198 24268 20204
rect 24228 20058 24256 20198
rect 24216 20052 24268 20058
rect 24216 19994 24268 20000
rect 24320 19802 24348 20488
rect 24584 20470 24636 20476
rect 24596 19922 24624 20470
rect 24584 19916 24636 19922
rect 24584 19858 24636 19864
rect 24492 19848 24544 19854
rect 24228 19774 24348 19802
rect 24490 19816 24492 19825
rect 24544 19816 24546 19825
rect 24124 18964 24176 18970
rect 24124 18906 24176 18912
rect 24030 17912 24086 17921
rect 24030 17847 24086 17856
rect 24228 17864 24256 19774
rect 24490 19751 24546 19760
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24584 19440 24636 19446
rect 24582 19408 24584 19417
rect 24636 19408 24638 19417
rect 24582 19343 24638 19352
rect 24490 19000 24546 19009
rect 24490 18935 24492 18944
rect 24544 18935 24546 18944
rect 24492 18906 24544 18912
rect 24596 18748 24624 19343
rect 24688 19310 24716 21626
rect 24780 21162 24808 22471
rect 24872 22098 24900 22630
rect 24860 22092 24912 22098
rect 24860 22034 24912 22040
rect 24780 21146 24900 21162
rect 24780 21140 24912 21146
rect 24780 21134 24860 21140
rect 24964 21128 24992 22732
rect 25044 22714 25096 22720
rect 25044 21548 25096 21554
rect 25044 21490 25096 21496
rect 25056 21350 25084 21490
rect 25228 21480 25280 21486
rect 25228 21422 25280 21428
rect 25044 21344 25096 21350
rect 25042 21312 25044 21321
rect 25096 21312 25098 21321
rect 25042 21247 25098 21256
rect 24964 21100 25084 21128
rect 24860 21082 24912 21088
rect 24952 21004 25004 21010
rect 24952 20946 25004 20952
rect 24860 20936 24912 20942
rect 24860 20878 24912 20884
rect 24872 20534 24900 20878
rect 24964 20602 24992 20946
rect 24952 20596 25004 20602
rect 24952 20538 25004 20544
rect 24860 20528 24912 20534
rect 24860 20470 24912 20476
rect 24768 20460 24820 20466
rect 24768 20402 24820 20408
rect 24780 19854 24808 20402
rect 24952 20392 25004 20398
rect 24952 20334 25004 20340
rect 24860 19984 24912 19990
rect 24860 19926 24912 19932
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 24676 19304 24728 19310
rect 24676 19246 24728 19252
rect 24688 18902 24716 19246
rect 24780 19174 24808 19790
rect 24872 19310 24900 19926
rect 24860 19304 24912 19310
rect 24860 19246 24912 19252
rect 24768 19168 24820 19174
rect 24768 19110 24820 19116
rect 24858 19136 24914 19145
rect 24676 18896 24728 18902
rect 24676 18838 24728 18844
rect 24676 18760 24728 18766
rect 24596 18720 24676 18748
rect 24676 18702 24728 18708
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24688 18358 24716 18702
rect 24676 18352 24728 18358
rect 24676 18294 24728 18300
rect 24308 17876 24360 17882
rect 24228 17836 24308 17864
rect 24308 17818 24360 17824
rect 24032 17808 24084 17814
rect 24032 17750 24084 17756
rect 23940 17672 23992 17678
rect 23940 17614 23992 17620
rect 23848 16584 23900 16590
rect 23848 16526 23900 16532
rect 23952 16522 23980 17614
rect 24044 17270 24072 17750
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24216 17536 24268 17542
rect 24216 17478 24268 17484
rect 24032 17264 24084 17270
rect 24032 17206 24084 17212
rect 24228 17202 24256 17478
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24688 17338 24716 17682
rect 24780 17513 24808 19110
rect 24858 19071 24914 19080
rect 24766 17504 24822 17513
rect 24766 17439 24822 17448
rect 24676 17332 24728 17338
rect 24872 17320 24900 19071
rect 24964 18630 24992 20334
rect 25056 19922 25084 21100
rect 25136 21004 25188 21010
rect 25136 20946 25188 20952
rect 25044 19916 25096 19922
rect 25044 19858 25096 19864
rect 25056 19174 25084 19858
rect 25044 19168 25096 19174
rect 25044 19110 25096 19116
rect 25044 18828 25096 18834
rect 25044 18770 25096 18776
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 24952 18420 25004 18426
rect 24952 18362 25004 18368
rect 24676 17274 24728 17280
rect 24780 17292 24900 17320
rect 24780 17218 24808 17292
rect 24216 17196 24268 17202
rect 24216 17138 24268 17144
rect 24688 17190 24808 17218
rect 24858 17232 24914 17241
rect 24688 16998 24716 17190
rect 24858 17167 24914 17176
rect 24768 17128 24820 17134
rect 24768 17070 24820 17076
rect 24032 16992 24084 16998
rect 24032 16934 24084 16940
rect 24216 16992 24268 16998
rect 24216 16934 24268 16940
rect 24676 16992 24728 16998
rect 24676 16934 24728 16940
rect 23940 16516 23992 16522
rect 23940 16458 23992 16464
rect 23848 16448 23900 16454
rect 23848 16390 23900 16396
rect 23860 15910 23888 16390
rect 24044 16114 24072 16934
rect 24032 16108 24084 16114
rect 24032 16050 24084 16056
rect 23848 15904 23900 15910
rect 23848 15846 23900 15852
rect 23860 14278 23888 15846
rect 24030 15736 24086 15745
rect 24030 15671 24032 15680
rect 24084 15671 24086 15680
rect 24032 15642 24084 15648
rect 23940 15564 23992 15570
rect 23940 15506 23992 15512
rect 23952 14890 23980 15506
rect 24044 15162 24072 15642
rect 24032 15156 24084 15162
rect 24032 15098 24084 15104
rect 23940 14884 23992 14890
rect 23940 14826 23992 14832
rect 23952 14618 23980 14826
rect 24228 14618 24256 16934
rect 24676 16652 24728 16658
rect 24676 16594 24728 16600
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24688 16250 24716 16594
rect 24676 16244 24728 16250
rect 24676 16186 24728 16192
rect 24676 16108 24728 16114
rect 24676 16050 24728 16056
rect 24688 15638 24716 16050
rect 24676 15632 24728 15638
rect 24676 15574 24728 15580
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24306 15056 24362 15065
rect 24688 15026 24716 15574
rect 24780 15348 24808 17070
rect 24872 16794 24900 17167
rect 24964 17134 24992 18362
rect 25056 17882 25084 18770
rect 25044 17876 25096 17882
rect 25044 17818 25096 17824
rect 25044 17672 25096 17678
rect 25044 17614 25096 17620
rect 24952 17128 25004 17134
rect 24952 17070 25004 17076
rect 24860 16788 24912 16794
rect 24860 16730 24912 16736
rect 25056 16726 25084 17614
rect 25044 16720 25096 16726
rect 25044 16662 25096 16668
rect 25148 16658 25176 20946
rect 25240 20233 25268 21422
rect 25226 20224 25282 20233
rect 25226 20159 25282 20168
rect 25228 19712 25280 19718
rect 25228 19654 25280 19660
rect 25240 18630 25268 19654
rect 25228 18624 25280 18630
rect 25228 18566 25280 18572
rect 25228 18216 25280 18222
rect 25226 18184 25228 18193
rect 25280 18184 25282 18193
rect 25226 18119 25282 18128
rect 25228 18080 25280 18086
rect 25228 18022 25280 18028
rect 25240 17542 25268 18022
rect 25228 17536 25280 17542
rect 25228 17478 25280 17484
rect 25332 17270 25360 23174
rect 25410 22672 25466 22681
rect 25410 22607 25466 22616
rect 25424 22574 25452 22607
rect 25412 22568 25464 22574
rect 25412 22510 25464 22516
rect 25410 21856 25466 21865
rect 25410 21791 25466 21800
rect 25424 20602 25452 21791
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25516 19394 25544 25350
rect 25594 25327 25650 25336
rect 25608 24954 25636 25327
rect 25596 24948 25648 24954
rect 25596 24890 25648 24896
rect 25594 23624 25650 23633
rect 25594 23559 25650 23568
rect 25608 22778 25636 23559
rect 25686 23080 25742 23089
rect 25686 23015 25742 23024
rect 25596 22772 25648 22778
rect 25596 22714 25648 22720
rect 25700 21690 25728 23015
rect 25688 21684 25740 21690
rect 25688 21626 25740 21632
rect 25688 21344 25740 21350
rect 25594 21312 25650 21321
rect 25688 21286 25740 21292
rect 25594 21247 25650 21256
rect 25424 19366 25544 19394
rect 25424 17377 25452 19366
rect 25504 19304 25556 19310
rect 25504 19246 25556 19252
rect 25516 18290 25544 19246
rect 25608 19174 25636 21247
rect 25596 19168 25648 19174
rect 25596 19110 25648 19116
rect 25700 18986 25728 21286
rect 25608 18958 25728 18986
rect 25504 18284 25556 18290
rect 25504 18226 25556 18232
rect 25410 17368 25466 17377
rect 25410 17303 25466 17312
rect 25320 17264 25372 17270
rect 25320 17206 25372 17212
rect 25412 17196 25464 17202
rect 25412 17138 25464 17144
rect 25424 17105 25452 17138
rect 25410 17096 25466 17105
rect 25410 17031 25466 17040
rect 25318 16688 25374 16697
rect 25136 16652 25188 16658
rect 25318 16623 25374 16632
rect 25412 16652 25464 16658
rect 25136 16594 25188 16600
rect 25136 16516 25188 16522
rect 25136 16458 25188 16464
rect 24858 16144 24914 16153
rect 24858 16079 24914 16088
rect 24872 15473 24900 16079
rect 25044 15904 25096 15910
rect 25044 15846 25096 15852
rect 24858 15464 24914 15473
rect 24858 15399 24914 15408
rect 24780 15320 24900 15348
rect 24306 14991 24362 15000
rect 24676 15020 24728 15026
rect 24320 14822 24348 14991
rect 24676 14962 24728 14968
rect 24308 14816 24360 14822
rect 24308 14758 24360 14764
rect 24320 14618 24348 14758
rect 23940 14612 23992 14618
rect 23940 14554 23992 14560
rect 24032 14612 24084 14618
rect 24032 14554 24084 14560
rect 24216 14612 24268 14618
rect 24216 14554 24268 14560
rect 24308 14612 24360 14618
rect 24308 14554 24360 14560
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 23940 13728 23992 13734
rect 23940 13670 23992 13676
rect 23848 12708 23900 12714
rect 23848 12650 23900 12656
rect 23860 12442 23888 12650
rect 23848 12436 23900 12442
rect 23848 12378 23900 12384
rect 23848 12300 23900 12306
rect 23848 12242 23900 12248
rect 23756 8016 23808 8022
rect 23756 7958 23808 7964
rect 23860 7410 23888 12242
rect 23952 12186 23980 13670
rect 24044 13394 24072 14554
rect 24214 14512 24270 14521
rect 24214 14447 24216 14456
rect 24268 14447 24270 14456
rect 24216 14418 24268 14424
rect 24228 14074 24256 14418
rect 24688 14414 24716 14962
rect 24768 14476 24820 14482
rect 24768 14418 24820 14424
rect 24676 14408 24728 14414
rect 24676 14350 24728 14356
rect 24676 14272 24728 14278
rect 24676 14214 24728 14220
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24216 14068 24268 14074
rect 24216 14010 24268 14016
rect 24032 13388 24084 13394
rect 24032 13330 24084 13336
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24122 12472 24178 12481
rect 24688 12458 24716 14214
rect 24780 13326 24808 14418
rect 24768 13320 24820 13326
rect 24766 13288 24768 13297
rect 24820 13288 24822 13297
rect 24766 13223 24822 13232
rect 24766 13016 24822 13025
rect 24766 12951 24822 12960
rect 24780 12646 24808 12951
rect 24872 12889 24900 15320
rect 25056 14618 25084 15846
rect 25148 15706 25176 16458
rect 25228 16040 25280 16046
rect 25228 15982 25280 15988
rect 25136 15700 25188 15706
rect 25136 15642 25188 15648
rect 25240 15609 25268 15982
rect 25332 15706 25360 16623
rect 25412 16594 25464 16600
rect 25504 16652 25556 16658
rect 25504 16594 25556 16600
rect 25320 15700 25372 15706
rect 25320 15642 25372 15648
rect 25226 15600 25282 15609
rect 25136 15564 25188 15570
rect 25226 15535 25282 15544
rect 25320 15564 25372 15570
rect 25136 15506 25188 15512
rect 25320 15506 25372 15512
rect 25148 15162 25176 15506
rect 25136 15156 25188 15162
rect 25136 15098 25188 15104
rect 25044 14612 25096 14618
rect 25044 14554 25096 14560
rect 25044 14476 25096 14482
rect 25044 14418 25096 14424
rect 24858 12880 24914 12889
rect 24858 12815 24914 12824
rect 24768 12640 24820 12646
rect 24768 12582 24820 12588
rect 24688 12430 24808 12458
rect 24122 12407 24124 12416
rect 24176 12407 24178 12416
rect 24124 12378 24176 12384
rect 23952 12158 24072 12186
rect 23940 12096 23992 12102
rect 23940 12038 23992 12044
rect 23952 11121 23980 12038
rect 24044 11354 24072 12158
rect 24136 11762 24164 12378
rect 24676 12096 24728 12102
rect 24676 12038 24728 12044
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24688 11898 24716 12038
rect 24676 11892 24728 11898
rect 24676 11834 24728 11840
rect 24124 11756 24176 11762
rect 24124 11698 24176 11704
rect 24216 11620 24268 11626
rect 24216 11562 24268 11568
rect 24032 11348 24084 11354
rect 24032 11290 24084 11296
rect 23938 11112 23994 11121
rect 23938 11047 23994 11056
rect 24228 10810 24256 11562
rect 24676 11280 24728 11286
rect 24676 11222 24728 11228
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24688 10810 24716 11222
rect 24216 10804 24268 10810
rect 24216 10746 24268 10752
rect 24676 10804 24728 10810
rect 24676 10746 24728 10752
rect 23938 10704 23994 10713
rect 23938 10639 23994 10648
rect 23952 9518 23980 10639
rect 24674 10568 24730 10577
rect 24674 10503 24730 10512
rect 24032 10464 24084 10470
rect 24032 10406 24084 10412
rect 23940 9512 23992 9518
rect 23940 9454 23992 9460
rect 23952 9178 23980 9454
rect 23940 9172 23992 9178
rect 23940 9114 23992 9120
rect 24044 8090 24072 10406
rect 24214 10296 24270 10305
rect 24214 10231 24270 10240
rect 24228 10198 24256 10231
rect 24216 10192 24268 10198
rect 24122 10160 24178 10169
rect 24216 10134 24268 10140
rect 24122 10095 24178 10104
rect 24136 8430 24164 10095
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24214 9616 24270 9625
rect 24214 9551 24270 9560
rect 24228 8537 24256 9551
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24214 8528 24270 8537
rect 24214 8463 24270 8472
rect 24124 8424 24176 8430
rect 24124 8366 24176 8372
rect 24032 8084 24084 8090
rect 24032 8026 24084 8032
rect 24136 7886 24164 8366
rect 24688 8242 24716 10503
rect 24780 8362 24808 12430
rect 24952 12368 25004 12374
rect 24952 12310 25004 12316
rect 24964 11778 24992 12310
rect 24872 11750 24992 11778
rect 24872 11626 24900 11750
rect 24950 11656 25006 11665
rect 24860 11620 24912 11626
rect 24950 11591 25006 11600
rect 24860 11562 24912 11568
rect 24964 11354 24992 11591
rect 24952 11348 25004 11354
rect 24952 11290 25004 11296
rect 24860 10804 24912 10810
rect 24860 10746 24912 10752
rect 24872 10266 24900 10746
rect 24950 10296 25006 10305
rect 24860 10260 24912 10266
rect 24950 10231 25006 10240
rect 24860 10202 24912 10208
rect 24964 9722 24992 10231
rect 24952 9716 25004 9722
rect 24952 9658 25004 9664
rect 24952 9376 25004 9382
rect 24952 9318 25004 9324
rect 24964 9042 24992 9318
rect 24952 9036 25004 9042
rect 24952 8978 25004 8984
rect 24964 8634 24992 8978
rect 24952 8628 25004 8634
rect 24952 8570 25004 8576
rect 24768 8356 24820 8362
rect 24768 8298 24820 8304
rect 24688 8214 24808 8242
rect 24214 7984 24270 7993
rect 24780 7970 24808 8214
rect 24214 7919 24270 7928
rect 24676 7948 24728 7954
rect 24124 7880 24176 7886
rect 24030 7848 24086 7857
rect 24124 7822 24176 7828
rect 24030 7783 24086 7792
rect 23940 7744 23992 7750
rect 23940 7686 23992 7692
rect 23848 7404 23900 7410
rect 23848 7346 23900 7352
rect 23756 7336 23808 7342
rect 23756 7278 23808 7284
rect 23768 6322 23796 7278
rect 23860 7002 23888 7346
rect 23848 6996 23900 7002
rect 23848 6938 23900 6944
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 23664 6248 23716 6254
rect 23664 6190 23716 6196
rect 23676 5914 23704 6190
rect 23664 5908 23716 5914
rect 23664 5850 23716 5856
rect 23584 5766 23704 5794
rect 23478 5743 23534 5752
rect 23388 5704 23440 5710
rect 23388 5646 23440 5652
rect 23492 5370 23520 5743
rect 23572 5568 23624 5574
rect 23572 5510 23624 5516
rect 23480 5364 23532 5370
rect 23480 5306 23532 5312
rect 23296 4684 23348 4690
rect 23296 4626 23348 4632
rect 23584 4298 23612 5510
rect 23676 5302 23704 5766
rect 23664 5296 23716 5302
rect 23664 5238 23716 5244
rect 23664 5024 23716 5030
rect 23664 4966 23716 4972
rect 23676 4729 23704 4966
rect 23662 4720 23718 4729
rect 23662 4655 23718 4664
rect 23664 4480 23716 4486
rect 23662 4448 23664 4457
rect 23716 4448 23718 4457
rect 23662 4383 23718 4392
rect 23400 4270 23612 4298
rect 23400 2122 23428 4270
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 23492 3942 23520 4082
rect 23480 3936 23532 3942
rect 23480 3878 23532 3884
rect 23572 3936 23624 3942
rect 23572 3878 23624 3884
rect 23492 3058 23520 3878
rect 23480 3052 23532 3058
rect 23480 2994 23532 3000
rect 23584 2553 23612 3878
rect 23756 3392 23808 3398
rect 23952 3369 23980 7686
rect 24044 7290 24072 7783
rect 24228 7313 24256 7919
rect 24780 7942 24900 7970
rect 24676 7890 24728 7896
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24214 7304 24270 7313
rect 24044 7274 24164 7290
rect 24044 7268 24176 7274
rect 24044 7262 24124 7268
rect 24214 7239 24270 7248
rect 24124 7210 24176 7216
rect 24124 6860 24176 6866
rect 24124 6802 24176 6808
rect 24030 6760 24086 6769
rect 24030 6695 24032 6704
rect 24084 6695 24086 6704
rect 24032 6666 24084 6672
rect 24030 6080 24086 6089
rect 24030 6015 24086 6024
rect 24044 4010 24072 6015
rect 24136 5914 24164 6802
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24688 6458 24716 7890
rect 24768 7880 24820 7886
rect 24768 7822 24820 7828
rect 24780 7546 24808 7822
rect 24768 7540 24820 7546
rect 24768 7482 24820 7488
rect 24872 7426 24900 7942
rect 24780 7410 24900 7426
rect 24768 7404 24900 7410
rect 24820 7398 24900 7404
rect 24768 7346 24820 7352
rect 25056 7018 25084 14418
rect 25148 13938 25176 15098
rect 25228 14952 25280 14958
rect 25228 14894 25280 14900
rect 25240 14278 25268 14894
rect 25332 14550 25360 15506
rect 25320 14544 25372 14550
rect 25320 14486 25372 14492
rect 25228 14272 25280 14278
rect 25226 14240 25228 14249
rect 25280 14240 25282 14249
rect 25226 14175 25282 14184
rect 25226 13968 25282 13977
rect 25136 13932 25188 13938
rect 25226 13903 25282 13912
rect 25136 13874 25188 13880
rect 25240 13870 25268 13903
rect 25228 13864 25280 13870
rect 25228 13806 25280 13812
rect 25332 12986 25360 14486
rect 25320 12980 25372 12986
rect 25320 12922 25372 12928
rect 25228 12300 25280 12306
rect 25228 12242 25280 12248
rect 25134 11928 25190 11937
rect 25134 11863 25190 11872
rect 25148 11257 25176 11863
rect 25240 11830 25268 12242
rect 25228 11824 25280 11830
rect 25228 11766 25280 11772
rect 25240 11354 25268 11766
rect 25332 11354 25360 12922
rect 25424 12442 25452 16594
rect 25412 12436 25464 12442
rect 25412 12378 25464 12384
rect 25424 11694 25452 12378
rect 25412 11688 25464 11694
rect 25412 11630 25464 11636
rect 25410 11520 25466 11529
rect 25410 11455 25466 11464
rect 25228 11348 25280 11354
rect 25228 11290 25280 11296
rect 25320 11348 25372 11354
rect 25320 11290 25372 11296
rect 25134 11248 25190 11257
rect 25134 11183 25190 11192
rect 25318 11112 25374 11121
rect 25318 11047 25374 11056
rect 25134 10024 25190 10033
rect 25134 9959 25136 9968
rect 25188 9959 25190 9968
rect 25136 9930 25188 9936
rect 25148 9178 25176 9930
rect 25136 9172 25188 9178
rect 25188 9132 25268 9160
rect 25136 9114 25188 9120
rect 25136 8832 25188 8838
rect 25136 8774 25188 8780
rect 25148 8673 25176 8774
rect 25134 8664 25190 8673
rect 25134 8599 25190 8608
rect 25136 8424 25188 8430
rect 25136 8366 25188 8372
rect 25148 7177 25176 8366
rect 25240 8090 25268 9132
rect 25228 8084 25280 8090
rect 25228 8026 25280 8032
rect 25228 7200 25280 7206
rect 25134 7168 25190 7177
rect 25228 7142 25280 7148
rect 25134 7103 25190 7112
rect 24780 6990 25084 7018
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 24780 6338 24808 6990
rect 24952 6928 25004 6934
rect 24952 6870 25004 6876
rect 24860 6860 24912 6866
rect 24860 6802 24912 6808
rect 24872 6390 24900 6802
rect 24688 6310 24808 6338
rect 24860 6384 24912 6390
rect 24860 6326 24912 6332
rect 24688 5914 24716 6310
rect 24860 6248 24912 6254
rect 24860 6190 24912 6196
rect 24768 6180 24820 6186
rect 24768 6122 24820 6128
rect 24124 5908 24176 5914
rect 24124 5850 24176 5856
rect 24676 5908 24728 5914
rect 24676 5850 24728 5856
rect 24136 5574 24164 5850
rect 24214 5672 24270 5681
rect 24214 5607 24270 5616
rect 24124 5568 24176 5574
rect 24124 5510 24176 5516
rect 24122 5400 24178 5409
rect 24122 5335 24178 5344
rect 24136 4826 24164 5335
rect 24124 4820 24176 4826
rect 24124 4762 24176 4768
rect 24122 4312 24178 4321
rect 24122 4247 24178 4256
rect 24136 4078 24164 4247
rect 24124 4072 24176 4078
rect 24124 4014 24176 4020
rect 24032 4004 24084 4010
rect 24032 3946 24084 3952
rect 24136 3738 24164 4014
rect 24124 3732 24176 3738
rect 24124 3674 24176 3680
rect 24032 3392 24084 3398
rect 23756 3334 23808 3340
rect 23938 3360 23994 3369
rect 23768 2990 23796 3334
rect 24032 3334 24084 3340
rect 23938 3295 23994 3304
rect 23756 2984 23808 2990
rect 23756 2926 23808 2932
rect 23952 2922 23980 3295
rect 24044 3233 24072 3334
rect 24030 3224 24086 3233
rect 24030 3159 24086 3168
rect 24032 2984 24084 2990
rect 24032 2926 24084 2932
rect 23940 2916 23992 2922
rect 23940 2858 23992 2864
rect 23664 2848 23716 2854
rect 23662 2816 23664 2825
rect 23716 2816 23718 2825
rect 23662 2751 23718 2760
rect 23938 2680 23994 2689
rect 23938 2615 23940 2624
rect 23992 2615 23994 2624
rect 23940 2586 23992 2592
rect 23570 2544 23626 2553
rect 23480 2508 23532 2514
rect 23570 2479 23626 2488
rect 23480 2450 23532 2456
rect 23492 2310 23520 2450
rect 23664 2440 23716 2446
rect 23662 2408 23664 2417
rect 23716 2408 23718 2417
rect 23662 2343 23718 2352
rect 23480 2304 23532 2310
rect 23478 2272 23480 2281
rect 23532 2272 23534 2281
rect 23478 2207 23534 2216
rect 23400 2094 23520 2122
rect 23492 921 23520 2094
rect 24044 1193 24072 2926
rect 24228 1986 24256 5607
rect 24780 5545 24808 6122
rect 24766 5536 24822 5545
rect 24289 5468 24585 5488
rect 24766 5471 24822 5480
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24872 5386 24900 6190
rect 24688 5358 24900 5386
rect 24308 5296 24360 5302
rect 24308 5238 24360 5244
rect 24320 5001 24348 5238
rect 24492 5160 24544 5166
rect 24492 5102 24544 5108
rect 24306 4992 24362 5001
rect 24306 4927 24362 4936
rect 24504 4554 24532 5102
rect 24688 4826 24716 5358
rect 24676 4820 24728 4826
rect 24676 4762 24728 4768
rect 24492 4548 24544 4554
rect 24492 4490 24544 4496
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24688 4282 24716 4762
rect 24860 4480 24912 4486
rect 24780 4440 24860 4468
rect 24676 4276 24728 4282
rect 24676 4218 24728 4224
rect 24780 4010 24808 4440
rect 24860 4422 24912 4428
rect 24964 4298 24992 6870
rect 25136 6724 25188 6730
rect 25136 6666 25188 6672
rect 25044 5772 25096 5778
rect 25044 5714 25096 5720
rect 25056 5098 25084 5714
rect 25148 5710 25176 6666
rect 25136 5704 25188 5710
rect 25240 5681 25268 7142
rect 25136 5646 25188 5652
rect 25226 5672 25282 5681
rect 25044 5092 25096 5098
rect 25044 5034 25096 5040
rect 25148 4826 25176 5646
rect 25226 5607 25282 5616
rect 25228 5568 25280 5574
rect 25228 5510 25280 5516
rect 25240 5302 25268 5510
rect 25228 5296 25280 5302
rect 25228 5238 25280 5244
rect 25136 4820 25188 4826
rect 25136 4762 25188 4768
rect 25148 4622 25176 4762
rect 25136 4616 25188 4622
rect 25136 4558 25188 4564
rect 25042 4448 25098 4457
rect 25042 4383 25098 4392
rect 24872 4270 24992 4298
rect 24768 4004 24820 4010
rect 24768 3946 24820 3952
rect 24490 3768 24546 3777
rect 24490 3703 24546 3712
rect 24504 3670 24532 3703
rect 24492 3664 24544 3670
rect 24492 3606 24544 3612
rect 24768 3664 24820 3670
rect 24768 3606 24820 3612
rect 24676 3528 24728 3534
rect 24676 3470 24728 3476
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24688 3058 24716 3470
rect 24676 3052 24728 3058
rect 24676 2994 24728 3000
rect 24780 2650 24808 3606
rect 24768 2644 24820 2650
rect 24768 2586 24820 2592
rect 24676 2440 24728 2446
rect 24676 2382 24728 2388
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24228 1958 24348 1986
rect 24030 1184 24086 1193
rect 24030 1119 24086 1128
rect 23478 912 23534 921
rect 23478 847 23534 856
rect 23756 604 23808 610
rect 23756 546 23808 552
rect 23768 480 23796 546
rect 24320 480 24348 1958
rect 24688 1601 24716 2382
rect 24674 1592 24730 1601
rect 24674 1527 24730 1536
rect 24872 480 24900 4270
rect 25056 4214 25084 4383
rect 25148 4282 25176 4558
rect 25136 4276 25188 4282
rect 25136 4218 25188 4224
rect 25044 4208 25096 4214
rect 25044 4150 25096 4156
rect 25228 4072 25280 4078
rect 25228 4014 25280 4020
rect 24952 4004 25004 4010
rect 24952 3946 25004 3952
rect 24964 1329 24992 3946
rect 25042 3632 25098 3641
rect 25042 3567 25098 3576
rect 25056 3194 25084 3567
rect 25044 3188 25096 3194
rect 25044 3130 25096 3136
rect 25240 2961 25268 4014
rect 25332 2990 25360 11047
rect 25424 10674 25452 11455
rect 25412 10668 25464 10674
rect 25412 10610 25464 10616
rect 25412 6656 25464 6662
rect 25412 6598 25464 6604
rect 25424 6458 25452 6598
rect 25412 6452 25464 6458
rect 25412 6394 25464 6400
rect 25412 6112 25464 6118
rect 25412 6054 25464 6060
rect 25320 2984 25372 2990
rect 25226 2952 25282 2961
rect 25320 2926 25372 2932
rect 25226 2887 25282 2896
rect 24950 1320 25006 1329
rect 24950 1255 25006 1264
rect 25424 480 25452 6054
rect 25516 4758 25544 16594
rect 25608 14482 25636 18958
rect 25792 17490 25820 26143
rect 25884 25498 25912 27520
rect 25872 25492 25924 25498
rect 25872 25434 25924 25440
rect 25872 23724 25924 23730
rect 25872 23666 25924 23672
rect 25884 21729 25912 23666
rect 25962 22400 26018 22409
rect 25962 22335 26018 22344
rect 25870 21720 25926 21729
rect 25870 21655 25926 21664
rect 25870 21584 25926 21593
rect 25870 21519 25926 21528
rect 25700 17462 25820 17490
rect 25596 14476 25648 14482
rect 25596 14418 25648 14424
rect 25596 12096 25648 12102
rect 25596 12038 25648 12044
rect 25608 11014 25636 12038
rect 25596 11008 25648 11014
rect 25596 10950 25648 10956
rect 25608 10470 25636 10950
rect 25596 10464 25648 10470
rect 25596 10406 25648 10412
rect 25608 9926 25636 10406
rect 25596 9920 25648 9926
rect 25596 9862 25648 9868
rect 25608 9450 25636 9862
rect 25596 9444 25648 9450
rect 25596 9386 25648 9392
rect 25608 9178 25636 9386
rect 25596 9172 25648 9178
rect 25596 9114 25648 9120
rect 25596 8900 25648 8906
rect 25596 8842 25648 8848
rect 25608 6458 25636 8842
rect 25596 6452 25648 6458
rect 25596 6394 25648 6400
rect 25608 5914 25636 6394
rect 25700 6100 25728 17462
rect 25884 17354 25912 21519
rect 25792 17326 25912 17354
rect 25792 16658 25820 17326
rect 25872 17264 25924 17270
rect 25872 17206 25924 17212
rect 25780 16652 25832 16658
rect 25780 16594 25832 16600
rect 25778 16552 25834 16561
rect 25778 16487 25834 16496
rect 25792 10810 25820 16487
rect 25884 11762 25912 17206
rect 25976 13530 26004 22335
rect 26068 16250 26096 27639
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 26528 25702 26556 27520
rect 26516 25696 26568 25702
rect 26516 25638 26568 25644
rect 27080 25226 27108 27520
rect 27632 25673 27660 27520
rect 27618 25664 27674 25673
rect 27618 25599 27674 25608
rect 27068 25220 27120 25226
rect 27068 25162 27120 25168
rect 26148 23520 26200 23526
rect 26148 23462 26200 23468
rect 26056 16244 26108 16250
rect 26056 16186 26108 16192
rect 26056 14816 26108 14822
rect 26056 14758 26108 14764
rect 26068 14278 26096 14758
rect 26056 14272 26108 14278
rect 26056 14214 26108 14220
rect 26068 13734 26096 14214
rect 26056 13728 26108 13734
rect 26056 13670 26108 13676
rect 25964 13524 26016 13530
rect 25964 13466 26016 13472
rect 26068 13462 26096 13670
rect 26056 13456 26108 13462
rect 26056 13398 26108 13404
rect 26068 12986 26096 13398
rect 26056 12980 26108 12986
rect 26056 12922 26108 12928
rect 26068 12442 26096 12922
rect 26056 12436 26108 12442
rect 26056 12378 26108 12384
rect 25962 11792 26018 11801
rect 25872 11756 25924 11762
rect 25962 11727 26018 11736
rect 25872 11698 25924 11704
rect 25780 10804 25832 10810
rect 25780 10746 25832 10752
rect 25792 10606 25820 10746
rect 25780 10600 25832 10606
rect 25780 10542 25832 10548
rect 25872 8288 25924 8294
rect 25872 8230 25924 8236
rect 25700 6072 25820 6100
rect 25596 5908 25648 5914
rect 25648 5868 25728 5896
rect 25596 5850 25648 5856
rect 25700 5370 25728 5868
rect 25688 5364 25740 5370
rect 25688 5306 25740 5312
rect 25596 5296 25648 5302
rect 25596 5238 25648 5244
rect 25504 4752 25556 4758
rect 25504 4694 25556 4700
rect 25504 2916 25556 2922
rect 25504 2858 25556 2864
rect 25516 1057 25544 2858
rect 25608 2530 25636 5238
rect 25688 5024 25740 5030
rect 25688 4966 25740 4972
rect 25700 4185 25728 4966
rect 25686 4176 25742 4185
rect 25686 4111 25742 4120
rect 25792 3738 25820 6072
rect 25884 5302 25912 8230
rect 25976 6089 26004 11727
rect 26056 10192 26108 10198
rect 26056 10134 26108 10140
rect 25962 6080 26018 6089
rect 25962 6015 26018 6024
rect 25872 5296 25924 5302
rect 25872 5238 25924 5244
rect 26068 5166 26096 10134
rect 26160 9330 26188 23462
rect 26238 19816 26294 19825
rect 26238 19751 26294 19760
rect 26252 19310 26280 19751
rect 26240 19304 26292 19310
rect 26240 19246 26292 19252
rect 26422 19000 26478 19009
rect 26422 18935 26478 18944
rect 26240 18624 26292 18630
rect 26240 18566 26292 18572
rect 26252 17542 26280 18566
rect 26330 18320 26386 18329
rect 26330 18255 26332 18264
rect 26384 18255 26386 18264
rect 26332 18226 26384 18232
rect 26330 17640 26386 17649
rect 26330 17575 26386 17584
rect 26240 17536 26292 17542
rect 26240 17478 26292 17484
rect 26252 16810 26280 17478
rect 26344 17338 26372 17575
rect 26332 17332 26384 17338
rect 26332 17274 26384 17280
rect 26252 16782 26372 16810
rect 26240 16720 26292 16726
rect 26240 16662 26292 16668
rect 26252 16250 26280 16662
rect 26344 16590 26372 16782
rect 26332 16584 26384 16590
rect 26332 16526 26384 16532
rect 26240 16244 26292 16250
rect 26240 16186 26292 16192
rect 26332 16108 26384 16114
rect 26332 16050 26384 16056
rect 26240 11552 26292 11558
rect 26240 11494 26292 11500
rect 26252 9994 26280 11494
rect 26344 10849 26372 16050
rect 26436 11898 26464 18935
rect 26424 11892 26476 11898
rect 26424 11834 26476 11840
rect 26330 10840 26386 10849
rect 26330 10775 26386 10784
rect 26240 9988 26292 9994
rect 26240 9930 26292 9936
rect 26160 9302 26280 9330
rect 26148 9172 26200 9178
rect 26148 9114 26200 9120
rect 26160 8634 26188 9114
rect 26148 8628 26200 8634
rect 26148 8570 26200 8576
rect 26148 8084 26200 8090
rect 26148 8026 26200 8032
rect 26160 7546 26188 8026
rect 26252 7750 26280 9302
rect 26240 7744 26292 7750
rect 26240 7686 26292 7692
rect 26148 7540 26200 7546
rect 26148 7482 26200 7488
rect 26160 7002 26188 7482
rect 26608 7472 26660 7478
rect 26608 7414 26660 7420
rect 26148 6996 26200 7002
rect 26148 6938 26200 6944
rect 26160 5846 26188 6938
rect 26240 6384 26292 6390
rect 26240 6326 26292 6332
rect 26148 5840 26200 5846
rect 26148 5782 26200 5788
rect 26148 5364 26200 5370
rect 26148 5306 26200 5312
rect 26056 5160 26108 5166
rect 25962 5128 26018 5137
rect 25872 5092 25924 5098
rect 26056 5102 26108 5108
rect 25962 5063 26018 5072
rect 25872 5034 25924 5040
rect 25780 3732 25832 3738
rect 25780 3674 25832 3680
rect 25608 2502 25728 2530
rect 25596 2440 25648 2446
rect 25596 2382 25648 2388
rect 25608 2009 25636 2382
rect 25594 2000 25650 2009
rect 25594 1935 25650 1944
rect 25502 1048 25558 1057
rect 25502 983 25558 992
rect 25700 610 25728 2502
rect 25884 2009 25912 5034
rect 25870 2000 25926 2009
rect 25870 1935 25926 1944
rect 25688 604 25740 610
rect 25688 546 25740 552
rect 25976 480 26004 5063
rect 26160 3738 26188 5306
rect 26148 3732 26200 3738
rect 26148 3674 26200 3680
rect 21086 96 21142 105
rect 21086 31 21142 40
rect 21546 0 21602 480
rect 22098 0 22154 480
rect 22650 0 22706 480
rect 23202 0 23258 480
rect 23754 0 23810 480
rect 24306 0 24362 480
rect 24858 0 24914 480
rect 25410 0 25466 480
rect 25962 0 26018 480
rect 26252 377 26280 6326
rect 26332 5840 26384 5846
rect 26332 5782 26384 5788
rect 26344 4826 26372 5782
rect 26332 4820 26384 4826
rect 26332 4762 26384 4768
rect 26344 4706 26372 4762
rect 26344 4678 26464 4706
rect 26332 4072 26384 4078
rect 26330 4040 26332 4049
rect 26384 4040 26386 4049
rect 26330 3975 26386 3984
rect 26330 3496 26386 3505
rect 26330 3431 26386 3440
rect 26344 3194 26372 3431
rect 26332 3188 26384 3194
rect 26332 3130 26384 3136
rect 26436 2650 26464 4678
rect 26620 2689 26648 7414
rect 27160 5228 27212 5234
rect 27160 5170 27212 5176
rect 26606 2680 26662 2689
rect 26424 2644 26476 2650
rect 26606 2615 26662 2624
rect 26424 2586 26476 2592
rect 26514 1728 26570 1737
rect 26514 1663 26570 1672
rect 26528 480 26556 1663
rect 27172 1465 27200 5170
rect 27618 4176 27674 4185
rect 27618 4111 27674 4120
rect 26790 1456 26846 1465
rect 27158 1456 27214 1465
rect 26846 1414 27108 1442
rect 26790 1391 26846 1400
rect 27080 480 27108 1414
rect 27158 1391 27214 1400
rect 27632 480 27660 4111
rect 26238 368 26294 377
rect 26238 303 26294 312
rect 26514 0 26570 480
rect 27066 0 27122 480
rect 27618 0 27674 480
<< via2 >>
rect 3514 27648 3570 27704
rect 1674 27104 1730 27160
rect 1490 26560 1546 26616
rect 1582 25336 1638 25392
rect 1582 24792 1638 24848
rect 1398 24112 1454 24168
rect 846 23296 902 23352
rect 294 22208 350 22264
rect 1490 23024 1546 23080
rect 1674 23060 1676 23080
rect 1676 23060 1728 23080
rect 1728 23060 1730 23080
rect 1674 23024 1730 23060
rect 1582 22480 1638 22536
rect 2042 23160 2098 23216
rect 2134 22480 2190 22536
rect 2042 21548 2098 21584
rect 2042 21528 2044 21548
rect 2044 21528 2096 21548
rect 2096 21528 2098 21548
rect 1950 20712 2006 20768
rect 1858 20576 1914 20632
rect 1030 17176 1086 17232
rect 846 13096 902 13152
rect 938 11872 994 11928
rect 846 11192 902 11248
rect 2042 20476 2044 20496
rect 2044 20476 2096 20496
rect 2096 20476 2098 20496
rect 2042 20440 2098 20476
rect 2410 22380 2412 22400
rect 2412 22380 2464 22400
rect 2464 22380 2466 22400
rect 2410 22344 2466 22380
rect 2686 25880 2742 25936
rect 2686 22480 2742 22536
rect 2962 22208 3018 22264
rect 2686 22072 2742 22128
rect 2594 21800 2650 21856
rect 2686 21256 2742 21312
rect 2410 20204 2412 20224
rect 2412 20204 2464 20224
rect 2464 20204 2466 20224
rect 2410 20168 2466 20204
rect 2318 19760 2374 19816
rect 1398 16632 1454 16688
rect 1122 13640 1178 13696
rect 2778 19488 2834 19544
rect 2778 19352 2834 19408
rect 2042 18028 2044 18048
rect 2044 18028 2096 18048
rect 2096 18028 2098 18048
rect 2042 17992 2098 18028
rect 1766 16632 1822 16688
rect 2410 17876 2466 17912
rect 2410 17856 2412 17876
rect 2412 17856 2464 17876
rect 2464 17856 2466 17876
rect 3146 21664 3202 21720
rect 3054 20848 3110 20904
rect 3146 20324 3202 20360
rect 3146 20304 3148 20324
rect 3148 20304 3200 20324
rect 3200 20304 3202 20324
rect 2870 18264 2926 18320
rect 3054 18128 3110 18184
rect 2594 17992 2650 18048
rect 2502 17040 2558 17096
rect 1858 15852 1860 15872
rect 1860 15852 1912 15872
rect 1912 15852 1914 15872
rect 1858 15816 1914 15852
rect 1490 12416 1546 12472
rect 1214 3576 1270 3632
rect 202 1672 258 1728
rect 1306 3168 1362 3224
rect 1766 13132 1768 13152
rect 1768 13132 1820 13152
rect 1820 13132 1822 13152
rect 1766 13096 1822 13132
rect 2134 13796 2190 13832
rect 2134 13776 2136 13796
rect 2136 13776 2188 13796
rect 2188 13776 2190 13796
rect 1950 12416 2006 12472
rect 1766 8356 1822 8392
rect 1766 8336 1768 8356
rect 1768 8336 1820 8356
rect 1820 8336 1822 8356
rect 1674 4392 1730 4448
rect 2134 11056 2190 11112
rect 2962 16904 3018 16960
rect 2870 13796 2926 13832
rect 2870 13776 2872 13796
rect 2872 13776 2924 13796
rect 2924 13776 2926 13796
rect 2686 12960 2742 13016
rect 2778 12860 2780 12880
rect 2780 12860 2832 12880
rect 2832 12860 2834 12880
rect 4066 23568 4122 23624
rect 3790 20032 3846 20088
rect 3698 19216 3754 19272
rect 3790 19080 3846 19136
rect 3698 17720 3754 17776
rect 3238 15680 3294 15736
rect 3422 15308 3424 15328
rect 3424 15308 3476 15328
rect 3476 15308 3478 15328
rect 3422 15272 3478 15308
rect 3238 13912 3294 13968
rect 2778 12824 2834 12860
rect 2686 11620 2742 11656
rect 2686 11600 2688 11620
rect 2688 11600 2740 11620
rect 2740 11600 2742 11620
rect 2686 11464 2742 11520
rect 1858 3848 1914 3904
rect 1766 3712 1822 3768
rect 1674 3168 1730 3224
rect 1398 1944 1454 2000
rect 1674 2624 1730 2680
rect 1582 856 1638 912
rect 2410 9988 2466 10024
rect 2410 9968 2412 9988
rect 2412 9968 2464 9988
rect 2464 9968 2466 9988
rect 3514 13268 3516 13288
rect 3516 13268 3568 13288
rect 3568 13268 3570 13288
rect 2962 8356 3018 8392
rect 2962 8336 2964 8356
rect 2964 8336 3016 8356
rect 3016 8336 3018 8356
rect 2870 8064 2926 8120
rect 2318 2896 2374 2952
rect 2870 7792 2926 7848
rect 3514 13232 3570 13268
rect 3422 11736 3478 11792
rect 3238 11600 3294 11656
rect 3330 10512 3386 10568
rect 3146 7928 3202 7984
rect 3698 16088 3754 16144
rect 4250 20168 4306 20224
rect 3790 14864 3846 14920
rect 3974 15272 4030 15328
rect 4066 13368 4122 13424
rect 3882 13096 3938 13152
rect 3698 11736 3754 11792
rect 3606 11056 3662 11112
rect 3698 10240 3754 10296
rect 3698 8472 3754 8528
rect 4066 13096 4122 13152
rect 4342 19252 4344 19272
rect 4344 19252 4396 19272
rect 4396 19252 4398 19272
rect 4342 19216 4398 19252
rect 3974 11600 4030 11656
rect 3974 10376 4030 10432
rect 3974 9560 4030 9616
rect 4066 8472 4122 8528
rect 6090 26016 6146 26072
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 6458 23160 6514 23216
rect 6642 23160 6698 23216
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 4710 22480 4766 22536
rect 5262 22344 5318 22400
rect 4710 22072 4766 22128
rect 4894 21684 4950 21720
rect 4894 21664 4896 21684
rect 4896 21664 4948 21684
rect 4948 21664 4950 21684
rect 4894 21140 4950 21176
rect 4894 21120 4896 21140
rect 4896 21120 4948 21140
rect 4948 21120 4950 21140
rect 4618 16768 4674 16824
rect 4986 20576 5042 20632
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5538 21292 5540 21312
rect 5540 21292 5592 21312
rect 5592 21292 5594 21312
rect 5538 21256 5594 21292
rect 5262 19896 5318 19952
rect 5538 21004 5594 21040
rect 5538 20984 5540 21004
rect 5540 20984 5592 21004
rect 5592 20984 5594 21004
rect 6090 20984 6146 21040
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5538 19760 5594 19816
rect 5722 19760 5778 19816
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 4986 18672 5042 18728
rect 5538 18808 5594 18864
rect 8114 25880 8170 25936
rect 7930 25744 7986 25800
rect 7746 24656 7802 24712
rect 7194 23316 7250 23352
rect 7194 23296 7196 23316
rect 7196 23296 7248 23316
rect 7248 23296 7250 23316
rect 7378 22888 7434 22944
rect 7286 22616 7342 22672
rect 7102 22208 7158 22264
rect 6918 21120 6974 21176
rect 6826 20712 6882 20768
rect 7470 22344 7526 22400
rect 7194 20984 7250 21040
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5538 17856 5594 17912
rect 5630 17720 5686 17776
rect 5170 17312 5226 17368
rect 4986 17176 5042 17232
rect 4986 16496 5042 16552
rect 4066 7792 4122 7848
rect 4434 7792 4490 7848
rect 3974 7148 3976 7168
rect 3976 7148 4028 7168
rect 4028 7148 4030 7168
rect 3974 7112 4030 7148
rect 3882 6024 3938 6080
rect 3514 5480 3570 5536
rect 3422 3168 3478 3224
rect 2042 1536 2098 1592
rect 2870 2760 2926 2816
rect 2962 2388 2964 2408
rect 2964 2388 3016 2408
rect 3016 2388 3018 2408
rect 2962 2352 3018 2388
rect 3790 3440 3846 3496
rect 4066 3732 4122 3768
rect 4066 3712 4068 3732
rect 4068 3712 4120 3732
rect 4120 3712 4122 3732
rect 3974 3032 4030 3088
rect 3882 1400 3938 1456
rect 3514 856 3570 912
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5630 15816 5686 15872
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 6458 17448 6514 17504
rect 6274 16904 6330 16960
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5630 13912 5686 13968
rect 5170 12844 5226 12880
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5170 12824 5172 12844
rect 5172 12824 5224 12844
rect 5224 12824 5226 12844
rect 5078 8880 5134 8936
rect 4894 7828 4896 7848
rect 4896 7828 4948 7848
rect 4948 7828 4950 7848
rect 4894 7792 4950 7828
rect 5446 12416 5502 12472
rect 6090 12044 6092 12064
rect 6092 12044 6144 12064
rect 6144 12044 6146 12064
rect 6090 12008 6146 12044
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5538 11620 5594 11656
rect 5538 11600 5540 11620
rect 5540 11600 5592 11620
rect 5592 11600 5594 11620
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 6734 18944 6790 19000
rect 6642 17584 6698 17640
rect 7194 20204 7196 20224
rect 7196 20204 7248 20224
rect 7248 20204 7250 20224
rect 7194 20168 7250 20204
rect 7010 18808 7066 18864
rect 6642 16652 6698 16688
rect 6642 16632 6644 16652
rect 6644 16632 6696 16652
rect 6696 16632 6698 16652
rect 6642 15816 6698 15872
rect 6366 13504 6422 13560
rect 6366 13096 6422 13152
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5446 9560 5502 9616
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5998 8200 6054 8256
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5998 7520 6054 7576
rect 5630 6860 5686 6896
rect 5630 6840 5632 6860
rect 5632 6840 5684 6860
rect 5684 6840 5686 6860
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5262 4528 5318 4584
rect 5078 1944 5134 2000
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5538 3984 5594 4040
rect 6182 8200 6238 8256
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6642 14184 6698 14240
rect 7286 18944 7342 19000
rect 7194 16632 7250 16688
rect 7010 14592 7066 14648
rect 6734 12980 6790 13016
rect 6734 12960 6736 12980
rect 6736 12960 6788 12980
rect 6788 12960 6790 12980
rect 7194 12416 7250 12472
rect 6734 12280 6790 12336
rect 6550 9832 6606 9888
rect 6458 9424 6514 9480
rect 6642 7928 6698 7984
rect 6642 7656 6698 7712
rect 6366 6840 6422 6896
rect 6642 2916 6698 2952
rect 6642 2896 6644 2916
rect 6644 2896 6696 2916
rect 6696 2896 6698 2916
rect 6274 1128 6330 1184
rect 6826 11500 6828 11520
rect 6828 11500 6880 11520
rect 6880 11500 6882 11520
rect 6826 11464 6882 11500
rect 7654 22752 7710 22808
rect 7562 18672 7618 18728
rect 8666 24248 8722 24304
rect 7654 15544 7710 15600
rect 7654 15308 7656 15328
rect 7656 15308 7708 15328
rect 7708 15308 7710 15328
rect 7654 15272 7710 15308
rect 7378 11348 7434 11384
rect 7378 11328 7380 11348
rect 7380 11328 7432 11348
rect 7432 11328 7434 11348
rect 7378 10784 7434 10840
rect 7562 12144 7618 12200
rect 7654 10920 7710 10976
rect 7102 8336 7158 8392
rect 6918 7948 6974 7984
rect 6918 7928 6920 7948
rect 6920 7928 6972 7948
rect 6972 7928 6974 7948
rect 7010 7812 7066 7848
rect 7010 7792 7012 7812
rect 7012 7792 7064 7812
rect 7064 7792 7066 7812
rect 7010 7384 7066 7440
rect 6826 6568 6882 6624
rect 8666 23160 8722 23216
rect 8206 22380 8208 22400
rect 8208 22380 8260 22400
rect 8260 22380 8262 22400
rect 8206 22344 8262 22380
rect 8390 21936 8446 21992
rect 8114 20576 8170 20632
rect 7930 18128 7986 18184
rect 8482 21256 8538 21312
rect 8298 19760 8354 19816
rect 8114 18944 8170 19000
rect 8574 20032 8630 20088
rect 8482 18264 8538 18320
rect 8390 17740 8446 17776
rect 8390 17720 8392 17740
rect 8392 17720 8444 17740
rect 8444 17720 8446 17740
rect 8114 17040 8170 17096
rect 8482 16768 8538 16824
rect 8022 15952 8078 16008
rect 8390 15988 8392 16008
rect 8392 15988 8444 16008
rect 8444 15988 8446 16008
rect 8390 15952 8446 15988
rect 9034 24792 9090 24848
rect 8850 23432 8906 23488
rect 26054 27648 26110 27704
rect 9494 24928 9550 24984
rect 9218 22072 9274 22128
rect 8942 20324 8998 20360
rect 8942 20304 8944 20324
rect 8944 20304 8996 20324
rect 8996 20304 8998 20324
rect 9126 19660 9128 19680
rect 9128 19660 9180 19680
rect 9180 19660 9182 19680
rect 9126 19624 9182 19660
rect 9034 18536 9090 18592
rect 8850 17876 8906 17912
rect 8850 17856 8852 17876
rect 8852 17856 8904 17876
rect 8904 17856 8906 17876
rect 9034 17176 9090 17232
rect 8942 17040 8998 17096
rect 9034 15816 9090 15872
rect 8022 13776 8078 13832
rect 8850 14884 8906 14920
rect 8850 14864 8852 14884
rect 8852 14864 8904 14884
rect 8904 14864 8906 14884
rect 8942 14456 8998 14512
rect 8942 14220 8944 14240
rect 8944 14220 8996 14240
rect 8996 14220 8998 14240
rect 8942 14184 8998 14220
rect 8206 12960 8262 13016
rect 8022 12588 8024 12608
rect 8024 12588 8076 12608
rect 8076 12588 8078 12608
rect 8022 12552 8078 12588
rect 8114 12280 8170 12336
rect 7838 11056 7894 11112
rect 7654 10104 7710 10160
rect 7930 10532 7986 10568
rect 7930 10512 7932 10532
rect 7932 10512 7984 10532
rect 7984 10512 7986 10532
rect 7654 8744 7710 8800
rect 7930 8628 7986 8664
rect 7930 8608 7932 8628
rect 7932 8608 7984 8628
rect 7984 8608 7986 8628
rect 7286 7520 7342 7576
rect 6826 4664 6882 4720
rect 6826 2080 6882 2136
rect 6918 1264 6974 1320
rect 4250 312 4306 368
rect 7194 6160 7250 6216
rect 7654 8084 7710 8120
rect 7654 8064 7656 8084
rect 7656 8064 7708 8084
rect 7708 8064 7710 8084
rect 7562 6724 7618 6760
rect 7562 6704 7564 6724
rect 7564 6704 7616 6724
rect 7616 6704 7618 6724
rect 8390 12688 8446 12744
rect 8298 10804 8354 10840
rect 8298 10784 8300 10804
rect 8300 10784 8352 10804
rect 8352 10784 8354 10804
rect 8298 9016 8354 9072
rect 8482 11872 8538 11928
rect 8482 8336 8538 8392
rect 7746 6568 7802 6624
rect 7562 5788 7564 5808
rect 7564 5788 7616 5808
rect 7616 5788 7618 5808
rect 7562 5752 7618 5788
rect 7286 5344 7342 5400
rect 7286 3460 7342 3496
rect 7286 3440 7288 3460
rect 7288 3440 7340 3460
rect 7340 3440 7342 3460
rect 7194 3168 7250 3224
rect 7194 2760 7250 2816
rect 7102 312 7158 368
rect 7654 2760 7710 2816
rect 7746 2624 7802 2680
rect 8022 5888 8078 5944
rect 8022 5636 8078 5672
rect 8022 5616 8024 5636
rect 8024 5616 8076 5636
rect 8076 5616 8078 5636
rect 9034 13368 9090 13424
rect 8942 11192 8998 11248
rect 8482 6568 8538 6624
rect 7930 5480 7986 5536
rect 8666 4548 8722 4584
rect 8666 4528 8668 4548
rect 8668 4528 8720 4548
rect 8720 4528 8722 4548
rect 9494 21936 9550 21992
rect 9678 25064 9734 25120
rect 9310 20440 9366 20496
rect 9770 24792 9826 24848
rect 9678 20440 9734 20496
rect 9494 20304 9550 20360
rect 9586 20204 9588 20224
rect 9588 20204 9640 20224
rect 9640 20204 9642 20224
rect 9586 20168 9642 20204
rect 9494 19488 9550 19544
rect 9402 17584 9458 17640
rect 9310 16496 9366 16552
rect 9402 15700 9458 15736
rect 9402 15680 9404 15700
rect 9404 15680 9456 15700
rect 9456 15680 9458 15700
rect 9402 15136 9458 15192
rect 9586 18808 9642 18864
rect 10046 23568 10102 23624
rect 10874 26152 10930 26208
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10414 24132 10470 24168
rect 10414 24112 10416 24132
rect 10416 24112 10468 24132
rect 10468 24112 10470 24132
rect 10230 23704 10286 23760
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10690 21936 10746 21992
rect 9862 19080 9918 19136
rect 9862 18944 9918 19000
rect 9678 17756 9680 17776
rect 9680 17756 9732 17776
rect 9732 17756 9734 17776
rect 9678 17720 9734 17756
rect 9770 17584 9826 17640
rect 9678 16088 9734 16144
rect 9770 14456 9826 14512
rect 9770 13640 9826 13696
rect 9402 12960 9458 13016
rect 9310 12280 9366 12336
rect 9494 11056 9550 11112
rect 9678 11600 9734 11656
rect 9678 9696 9734 9752
rect 9310 8744 9366 8800
rect 9218 8064 9274 8120
rect 9218 7792 9274 7848
rect 8022 2932 8024 2952
rect 8024 2932 8076 2952
rect 8076 2932 8078 2952
rect 8022 2896 8078 2932
rect 8850 2760 8906 2816
rect 8758 2488 8814 2544
rect 7562 176 7618 232
rect 9218 3168 9274 3224
rect 9126 992 9182 1048
rect 8482 40 8538 96
rect 9586 8608 9642 8664
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10598 20848 10654 20904
rect 10782 20440 10838 20496
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10230 19252 10232 19272
rect 10232 19252 10284 19272
rect 10284 19252 10286 19272
rect 10230 19216 10286 19252
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10322 18400 10378 18456
rect 11794 26288 11850 26344
rect 11518 25608 11574 25664
rect 11426 24656 11482 24712
rect 11242 22344 11298 22400
rect 10966 19760 11022 19816
rect 11058 19624 11114 19680
rect 10966 18944 11022 19000
rect 11334 20032 11390 20088
rect 11334 19896 11390 19952
rect 11242 19236 11298 19272
rect 11242 19216 11244 19236
rect 11244 19216 11296 19236
rect 11296 19216 11298 19236
rect 11242 19080 11298 19136
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 9954 15272 10010 15328
rect 9862 12552 9918 12608
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10506 16244 10562 16280
rect 10506 16224 10508 16244
rect 10508 16224 10560 16244
rect 10560 16224 10562 16244
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10966 18672 11022 18728
rect 11058 17992 11114 18048
rect 11058 17856 11114 17912
rect 10966 15952 11022 16008
rect 10874 15852 10876 15872
rect 10876 15852 10928 15872
rect 10928 15852 10930 15872
rect 10874 15816 10930 15852
rect 10414 15000 10470 15056
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10138 13640 10194 13696
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 9770 8356 9826 8392
rect 9770 8336 9772 8356
rect 9772 8336 9824 8356
rect 9824 8336 9826 8356
rect 9678 7792 9734 7848
rect 9862 7792 9918 7848
rect 9862 7112 9918 7168
rect 10874 15272 10930 15328
rect 11242 16496 11298 16552
rect 11610 22888 11666 22944
rect 11518 22480 11574 22536
rect 11518 20712 11574 20768
rect 11518 19896 11574 19952
rect 11886 22072 11942 22128
rect 11702 20440 11758 20496
rect 11610 19760 11666 19816
rect 11886 20168 11942 20224
rect 11886 19760 11942 19816
rect 12346 23468 12348 23488
rect 12348 23468 12400 23488
rect 12400 23468 12402 23488
rect 12346 23432 12402 23468
rect 12346 22480 12402 22536
rect 12346 20576 12402 20632
rect 12530 22480 12586 22536
rect 12898 24928 12954 24984
rect 12898 24384 12954 24440
rect 12990 23432 13046 23488
rect 12254 20032 12310 20088
rect 12438 20304 12494 20360
rect 11794 19216 11850 19272
rect 11978 19116 11980 19136
rect 11980 19116 12032 19136
rect 12032 19116 12034 19136
rect 11978 19080 12034 19116
rect 11426 15952 11482 16008
rect 11426 15680 11482 15736
rect 11334 15272 11390 15328
rect 11058 14320 11114 14376
rect 10966 14048 11022 14104
rect 10874 13640 10930 13696
rect 10782 13524 10838 13560
rect 10782 13504 10784 13524
rect 10784 13504 10836 13524
rect 10836 13504 10838 13524
rect 10874 12960 10930 13016
rect 10782 12824 10838 12880
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10414 12280 10470 12336
rect 10690 12280 10746 12336
rect 10230 12008 10286 12064
rect 10138 11736 10194 11792
rect 11242 14456 11298 14512
rect 11242 13912 11298 13968
rect 11426 13776 11482 13832
rect 11794 18672 11850 18728
rect 11702 17856 11758 17912
rect 11702 17448 11758 17504
rect 11610 15156 11666 15192
rect 11610 15136 11612 15156
rect 11612 15136 11664 15156
rect 11664 15136 11666 15156
rect 11150 12552 11206 12608
rect 10414 12008 10470 12064
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10598 10668 10654 10704
rect 10598 10648 10600 10668
rect 10600 10648 10652 10668
rect 10652 10648 10654 10668
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10046 7656 10102 7712
rect 10782 9152 10838 9208
rect 11334 11872 11390 11928
rect 11242 11600 11298 11656
rect 10966 9696 11022 9752
rect 11610 13368 11666 13424
rect 11518 12144 11574 12200
rect 11334 10412 11336 10432
rect 11336 10412 11388 10432
rect 11388 10412 11390 10432
rect 11334 10376 11390 10412
rect 11242 9832 11298 9888
rect 11242 9560 11298 9616
rect 11058 9288 11114 9344
rect 10782 7656 10838 7712
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10138 6740 10140 6760
rect 10140 6740 10192 6760
rect 10192 6740 10194 6760
rect 10138 6704 10194 6740
rect 9586 4120 9642 4176
rect 10046 5888 10102 5944
rect 9954 5072 10010 5128
rect 10046 3884 10048 3904
rect 10048 3884 10100 3904
rect 10100 3884 10102 3904
rect 10046 3848 10102 3884
rect 9862 3712 9918 3768
rect 9954 2760 10010 2816
rect 9862 2624 9918 2680
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10690 5616 10746 5672
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 11150 8608 11206 8664
rect 11334 9016 11390 9072
rect 11058 7520 11114 7576
rect 11058 7420 11060 7440
rect 11060 7420 11112 7440
rect 11112 7420 11114 7440
rect 11058 7384 11114 7420
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 11886 15816 11942 15872
rect 12162 18808 12218 18864
rect 12162 18536 12218 18592
rect 12162 17856 12218 17912
rect 12346 18264 12402 18320
rect 12806 20712 12862 20768
rect 12806 20052 12862 20088
rect 12806 20032 12808 20052
rect 12808 20032 12860 20052
rect 12860 20032 12862 20052
rect 12622 19760 12678 19816
rect 12622 19352 12678 19408
rect 12806 19488 12862 19544
rect 12530 18708 12532 18728
rect 12532 18708 12584 18728
rect 12584 18708 12586 18728
rect 12530 18672 12586 18708
rect 12714 19080 12770 19136
rect 12990 18944 13046 19000
rect 12162 14864 12218 14920
rect 11886 12688 11942 12744
rect 11702 11872 11758 11928
rect 11794 11736 11850 11792
rect 11978 11600 12034 11656
rect 11702 10140 11704 10160
rect 11704 10140 11756 10160
rect 11756 10140 11758 10160
rect 11702 10104 11758 10140
rect 11610 9832 11666 9888
rect 11518 6452 11574 6488
rect 11518 6432 11520 6452
rect 11520 6432 11572 6452
rect 11572 6432 11574 6452
rect 11242 5480 11298 5536
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10598 2216 10654 2272
rect 11334 4120 11390 4176
rect 11886 9696 11942 9752
rect 12070 11092 12072 11112
rect 12072 11092 12124 11112
rect 12124 11092 12126 11112
rect 12070 11056 12126 11092
rect 12714 18536 12770 18592
rect 12622 17584 12678 17640
rect 12346 13776 12402 13832
rect 12530 16224 12586 16280
rect 13542 25064 13598 25120
rect 13542 23704 13598 23760
rect 13450 23160 13506 23216
rect 13450 22072 13506 22128
rect 13174 19216 13230 19272
rect 12806 15680 12862 15736
rect 12714 15544 12770 15600
rect 11978 8744 12034 8800
rect 11702 7792 11758 7848
rect 11702 5480 11758 5536
rect 11518 3712 11574 3768
rect 11518 3068 11520 3088
rect 11520 3068 11572 3088
rect 11572 3068 11574 3088
rect 11518 3032 11574 3068
rect 11518 1672 11574 1728
rect 11610 1400 11666 1456
rect 11794 4800 11850 4856
rect 11794 4256 11850 4312
rect 11794 2624 11850 2680
rect 12990 15544 13046 15600
rect 12806 13252 12862 13288
rect 12806 13232 12808 13252
rect 12808 13232 12860 13252
rect 12860 13232 12862 13252
rect 12346 11212 12402 11248
rect 12346 11192 12348 11212
rect 12348 11192 12400 11212
rect 12400 11192 12402 11212
rect 12346 11076 12402 11112
rect 12346 11056 12348 11076
rect 12348 11056 12400 11076
rect 12400 11056 12402 11076
rect 12438 9716 12494 9752
rect 12438 9696 12440 9716
rect 12440 9696 12492 9716
rect 12492 9696 12494 9716
rect 12438 9016 12494 9072
rect 12070 6024 12126 6080
rect 11978 4936 12034 4992
rect 12806 10920 12862 10976
rect 12622 7692 12624 7712
rect 12624 7692 12676 7712
rect 12676 7692 12678 7712
rect 12622 7656 12678 7692
rect 13266 16768 13322 16824
rect 13450 18808 13506 18864
rect 13450 14900 13452 14920
rect 13452 14900 13504 14920
rect 13504 14900 13506 14920
rect 13450 14864 13506 14900
rect 13450 14592 13506 14648
rect 13450 13948 13452 13968
rect 13452 13948 13504 13968
rect 13504 13948 13506 13968
rect 13450 13912 13506 13948
rect 13450 13404 13452 13424
rect 13452 13404 13504 13424
rect 13504 13404 13506 13424
rect 13450 13368 13506 13404
rect 13174 9152 13230 9208
rect 12622 5344 12678 5400
rect 12622 5072 12678 5128
rect 12254 4256 12310 4312
rect 12070 1944 12126 2000
rect 11886 1672 11942 1728
rect 12438 3984 12494 4040
rect 12438 3304 12494 3360
rect 12990 6024 13046 6080
rect 12898 5752 12954 5808
rect 12806 5616 12862 5672
rect 12990 5208 13046 5264
rect 13174 5772 13230 5808
rect 13174 5752 13176 5772
rect 13176 5752 13228 5772
rect 13228 5752 13230 5772
rect 12990 4664 13046 4720
rect 14462 25880 14518 25936
rect 14278 24928 14334 24984
rect 13818 22616 13874 22672
rect 13726 18536 13782 18592
rect 13726 17856 13782 17912
rect 14186 22752 14242 22808
rect 14094 21120 14150 21176
rect 14462 24520 14518 24576
rect 14186 20596 14242 20632
rect 14186 20576 14188 20596
rect 14188 20576 14240 20596
rect 14240 20576 14242 20596
rect 13634 17176 13690 17232
rect 13634 16224 13690 16280
rect 13634 15408 13690 15464
rect 13634 13776 13690 13832
rect 14186 18264 14242 18320
rect 14094 17448 14150 17504
rect 13910 16632 13966 16688
rect 13818 13504 13874 13560
rect 13910 13388 13966 13424
rect 13910 13368 13912 13388
rect 13912 13368 13964 13388
rect 13964 13368 13966 13388
rect 13726 13096 13782 13152
rect 13634 12280 13690 12336
rect 14186 17176 14242 17232
rect 14094 13404 14096 13424
rect 14096 13404 14148 13424
rect 14148 13404 14150 13424
rect 14094 13368 14150 13404
rect 13818 11600 13874 11656
rect 13542 10512 13598 10568
rect 13358 4936 13414 4992
rect 13358 4120 13414 4176
rect 12990 2216 13046 2272
rect 13634 6976 13690 7032
rect 13726 5480 13782 5536
rect 13542 4800 13598 4856
rect 13634 4548 13690 4584
rect 13634 4528 13636 4548
rect 13636 4528 13688 4548
rect 13688 4528 13690 4548
rect 13542 3984 13598 4040
rect 13542 3440 13598 3496
rect 14370 18944 14426 19000
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14922 24792 14978 24848
rect 15106 24556 15108 24576
rect 15108 24556 15160 24576
rect 15160 24556 15162 24576
rect 15106 24520 15162 24556
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14830 23296 14886 23352
rect 15290 23160 15346 23216
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14646 19932 14648 19952
rect 14648 19932 14700 19952
rect 14700 19932 14702 19952
rect 14646 19896 14702 19932
rect 14462 17076 14464 17096
rect 14464 17076 14516 17096
rect 14516 17076 14518 17096
rect 14462 17040 14518 17076
rect 14278 16904 14334 16960
rect 14370 16788 14426 16824
rect 14370 16768 14372 16788
rect 14372 16768 14424 16788
rect 14424 16768 14426 16788
rect 14370 16088 14426 16144
rect 15106 22208 15162 22264
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 15106 20440 15162 20496
rect 14830 20304 14886 20360
rect 14830 19896 14886 19952
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 15934 26016 15990 26072
rect 15934 24928 15990 24984
rect 15566 24404 15622 24440
rect 15566 24384 15568 24404
rect 15568 24384 15620 24404
rect 15620 24384 15622 24404
rect 15474 23860 15530 23896
rect 15474 23840 15476 23860
rect 15476 23840 15528 23860
rect 15528 23840 15530 23860
rect 15474 23568 15530 23624
rect 15658 23432 15714 23488
rect 15658 22888 15714 22944
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 15106 17876 15162 17912
rect 15106 17856 15108 17876
rect 15108 17856 15160 17876
rect 15160 17856 15162 17876
rect 14830 17584 14886 17640
rect 14646 17076 14648 17096
rect 14648 17076 14700 17096
rect 14700 17076 14702 17096
rect 14646 17040 14702 17076
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14738 16904 14794 16960
rect 15198 16652 15254 16688
rect 15198 16632 15200 16652
rect 15200 16632 15252 16652
rect 15252 16632 15254 16652
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14738 16224 14794 16280
rect 14462 13912 14518 13968
rect 14462 13812 14464 13832
rect 14464 13812 14516 13832
rect 14516 13812 14518 13832
rect 14462 13776 14518 13812
rect 14646 15136 14702 15192
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 15106 15000 15162 15056
rect 14830 14728 14886 14784
rect 14738 14184 14794 14240
rect 14646 13932 14702 13968
rect 14646 13912 14648 13932
rect 14648 13912 14700 13932
rect 14700 13912 14702 13932
rect 14646 12960 14702 13016
rect 14370 12416 14426 12472
rect 14462 12008 14518 12064
rect 14646 11872 14702 11928
rect 14370 9832 14426 9888
rect 14186 8608 14242 8664
rect 14370 8508 14372 8528
rect 14372 8508 14424 8528
rect 14424 8508 14426 8528
rect 14370 8472 14426 8508
rect 14278 8064 14334 8120
rect 14646 10784 14702 10840
rect 15106 14456 15162 14512
rect 15290 14340 15346 14376
rect 15290 14320 15292 14340
rect 15292 14320 15344 14340
rect 15344 14320 15346 14340
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 15290 13912 15346 13968
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14922 12416 14978 12472
rect 15566 20576 15622 20632
rect 15382 12552 15438 12608
rect 15382 12280 15438 12336
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14830 10684 14832 10704
rect 14832 10684 14884 10704
rect 14884 10684 14886 10704
rect 14830 10648 14886 10684
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 15106 9560 15162 9616
rect 14646 9460 14648 9480
rect 14648 9460 14700 9480
rect 14700 9460 14702 9480
rect 14646 9424 14702 9460
rect 14830 9424 14886 9480
rect 15014 9152 15070 9208
rect 14830 8880 14886 8936
rect 14646 8608 14702 8664
rect 14370 6976 14426 7032
rect 14094 4564 14096 4584
rect 14096 4564 14148 4584
rect 14148 4564 14150 4584
rect 14094 4528 14150 4564
rect 14370 2760 14426 2816
rect 14002 2488 14058 2544
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 15106 8472 15162 8528
rect 15106 7792 15162 7848
rect 15290 7812 15346 7848
rect 15290 7792 15292 7812
rect 15292 7792 15344 7812
rect 15344 7792 15346 7812
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14646 6568 14702 6624
rect 15290 6840 15346 6896
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 15290 5752 15346 5808
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14646 4800 14702 4856
rect 14554 3712 14610 3768
rect 15014 4936 15070 4992
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14922 2896 14978 2952
rect 15658 15680 15714 15736
rect 15658 14612 15714 14648
rect 15658 14592 15660 14612
rect 15660 14592 15712 14612
rect 15712 14592 15714 14612
rect 16118 26016 16174 26072
rect 17038 25472 17094 25528
rect 16026 24792 16082 24848
rect 15934 23704 15990 23760
rect 15934 23604 15936 23624
rect 15936 23604 15988 23624
rect 15988 23604 15990 23624
rect 15934 23568 15990 23604
rect 15934 23060 15936 23080
rect 15936 23060 15988 23080
rect 15988 23060 15990 23080
rect 15934 23024 15990 23060
rect 15842 22380 15844 22400
rect 15844 22380 15896 22400
rect 15896 22380 15898 22400
rect 15842 22344 15898 22380
rect 16302 23704 16358 23760
rect 16026 21936 16082 21992
rect 15842 20576 15898 20632
rect 15842 17584 15898 17640
rect 15934 16224 15990 16280
rect 15934 15852 15936 15872
rect 15936 15852 15988 15872
rect 15988 15852 15990 15872
rect 15934 15816 15990 15852
rect 15658 12688 15714 12744
rect 16026 13232 16082 13288
rect 15934 12280 15990 12336
rect 15750 11872 15806 11928
rect 15658 11464 15714 11520
rect 15566 10240 15622 10296
rect 15750 11056 15806 11112
rect 15658 9968 15714 10024
rect 15842 10412 15844 10432
rect 15844 10412 15896 10432
rect 15896 10412 15898 10432
rect 15842 10376 15898 10412
rect 15750 8916 15752 8936
rect 15752 8916 15804 8936
rect 15804 8916 15806 8936
rect 15750 8880 15806 8916
rect 15474 7248 15530 7304
rect 15658 7248 15714 7304
rect 15658 6296 15714 6352
rect 15566 6160 15622 6216
rect 14554 2524 14556 2544
rect 14556 2524 14608 2544
rect 14608 2524 14610 2544
rect 14554 2488 14610 2524
rect 14462 2388 14464 2408
rect 14464 2388 14516 2408
rect 14516 2388 14518 2408
rect 14462 2352 14518 2388
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 15290 1944 15346 2000
rect 15658 4820 15714 4856
rect 15658 4800 15660 4820
rect 15660 4800 15712 4820
rect 15712 4800 15714 4820
rect 16026 9968 16082 10024
rect 16026 9016 16082 9072
rect 15934 7928 15990 7984
rect 16026 7540 16082 7576
rect 16026 7520 16028 7540
rect 16028 7520 16080 7540
rect 16080 7520 16082 7540
rect 16026 7248 16082 7304
rect 15934 6060 15936 6080
rect 15936 6060 15988 6080
rect 15988 6060 15990 6080
rect 15934 6024 15990 6060
rect 17038 24792 17094 24848
rect 16854 24520 16910 24576
rect 17130 23976 17186 24032
rect 16394 22480 16450 22536
rect 16302 21800 16358 21856
rect 16302 21664 16358 21720
rect 16578 21392 16634 21448
rect 16854 23160 16910 23216
rect 16394 21256 16450 21312
rect 16394 20712 16450 20768
rect 16302 19216 16358 19272
rect 16670 19352 16726 19408
rect 16302 18128 16358 18184
rect 16486 18808 16542 18864
rect 16578 18128 16634 18184
rect 16394 16632 16450 16688
rect 16210 15564 16266 15600
rect 16210 15544 16212 15564
rect 16212 15544 16264 15564
rect 16264 15544 16266 15564
rect 16394 14864 16450 14920
rect 16394 14456 16450 14512
rect 16394 12144 16450 12200
rect 16394 10240 16450 10296
rect 17866 26288 17922 26344
rect 18050 24928 18106 24984
rect 17130 22380 17132 22400
rect 17132 22380 17184 22400
rect 17184 22380 17186 22400
rect 17130 22344 17186 22380
rect 17130 21564 17132 21584
rect 17132 21564 17184 21584
rect 17184 21564 17186 21584
rect 17130 21528 17186 21564
rect 17038 20440 17094 20496
rect 16946 17176 17002 17232
rect 16762 16224 16818 16280
rect 16762 15020 16818 15056
rect 16762 15000 16764 15020
rect 16764 15000 16816 15020
rect 16816 15000 16818 15020
rect 16762 14728 16818 14784
rect 16670 13504 16726 13560
rect 17130 15680 17186 15736
rect 16762 12280 16818 12336
rect 16210 7520 16266 7576
rect 17130 13796 17186 13832
rect 17130 13776 17132 13796
rect 17132 13776 17184 13796
rect 17184 13776 17186 13796
rect 17038 13368 17094 13424
rect 17682 24248 17738 24304
rect 17314 21528 17370 21584
rect 17222 13232 17278 13288
rect 17038 12416 17094 12472
rect 17130 11872 17186 11928
rect 16394 8780 16396 8800
rect 16396 8780 16448 8800
rect 16448 8780 16450 8800
rect 16394 8744 16450 8780
rect 16302 6704 16358 6760
rect 16394 3440 16450 3496
rect 17314 12436 17370 12472
rect 17314 12416 17316 12436
rect 17316 12416 17368 12436
rect 17368 12416 17370 12436
rect 18050 24248 18106 24304
rect 17682 19116 17684 19136
rect 17684 19116 17736 19136
rect 17736 19116 17738 19136
rect 17682 19080 17738 19116
rect 17682 17720 17738 17776
rect 17590 17176 17646 17232
rect 17590 13368 17646 13424
rect 17866 20576 17922 20632
rect 17866 20476 17868 20496
rect 17868 20476 17920 20496
rect 17920 20476 17922 20496
rect 17866 20440 17922 20476
rect 17866 19760 17922 19816
rect 18142 23024 18198 23080
rect 19062 24384 19118 24440
rect 18418 23316 18474 23352
rect 18418 23296 18420 23316
rect 18420 23296 18472 23316
rect 18472 23296 18474 23316
rect 18234 22480 18290 22536
rect 18142 22072 18198 22128
rect 18142 21256 18198 21312
rect 18050 21120 18106 21176
rect 18234 20984 18290 21040
rect 18142 20168 18198 20224
rect 18234 19660 18236 19680
rect 18236 19660 18288 19680
rect 18288 19660 18290 19680
rect 18234 19624 18290 19660
rect 17866 18128 17922 18184
rect 18050 17448 18106 17504
rect 18050 17176 18106 17232
rect 18142 16632 18198 16688
rect 17958 16360 18014 16416
rect 18050 15272 18106 15328
rect 18050 14592 18106 14648
rect 17958 13504 18014 13560
rect 17958 12824 18014 12880
rect 17406 11736 17462 11792
rect 17314 11500 17316 11520
rect 17316 11500 17368 11520
rect 17368 11500 17370 11520
rect 17314 11464 17370 11500
rect 17130 7964 17132 7984
rect 17132 7964 17184 7984
rect 17184 7964 17186 7984
rect 17130 7928 17186 7964
rect 16762 7268 16818 7304
rect 16762 7248 16764 7268
rect 16764 7248 16816 7268
rect 16816 7248 16818 7268
rect 16854 6976 16910 7032
rect 17498 10104 17554 10160
rect 17498 9172 17554 9208
rect 17498 9152 17500 9172
rect 17500 9152 17552 9172
rect 17552 9152 17554 9172
rect 17406 8608 17462 8664
rect 17406 7792 17462 7848
rect 17038 6704 17094 6760
rect 17222 6704 17278 6760
rect 17406 6604 17408 6624
rect 17408 6604 17460 6624
rect 17460 6604 17462 6624
rect 17406 6568 17462 6604
rect 17038 5208 17094 5264
rect 16670 3304 16726 3360
rect 17406 4664 17462 4720
rect 17314 4120 17370 4176
rect 17682 11192 17738 11248
rect 17682 10920 17738 10976
rect 17774 10648 17830 10704
rect 17958 12416 18014 12472
rect 18234 15136 18290 15192
rect 18234 13912 18290 13968
rect 18050 10920 18106 10976
rect 18050 10784 18106 10840
rect 18142 10648 18198 10704
rect 17958 9832 18014 9888
rect 18418 22344 18474 22400
rect 18602 23432 18658 23488
rect 18510 21392 18566 21448
rect 18418 20984 18474 21040
rect 18418 20712 18474 20768
rect 18694 19760 18750 19816
rect 18602 18536 18658 18592
rect 18510 18264 18566 18320
rect 18510 17176 18566 17232
rect 18694 18264 18750 18320
rect 18694 17584 18750 17640
rect 18510 16904 18566 16960
rect 18418 15988 18420 16008
rect 18420 15988 18472 16008
rect 18472 15988 18474 16008
rect 18418 15952 18474 15988
rect 18602 16768 18658 16824
rect 18510 13232 18566 13288
rect 17866 9016 17922 9072
rect 17866 7112 17922 7168
rect 17774 4684 17830 4720
rect 17774 4664 17776 4684
rect 17776 4664 17828 4684
rect 17828 4664 17830 4684
rect 18050 4528 18106 4584
rect 17406 3984 17462 4040
rect 16854 3476 16856 3496
rect 16856 3476 16908 3496
rect 16908 3476 16910 3496
rect 16854 3440 16910 3476
rect 17038 3440 17094 3496
rect 16578 2760 16634 2816
rect 16118 856 16174 912
rect 17590 3984 17646 4040
rect 17774 3576 17830 3632
rect 17406 2896 17462 2952
rect 17498 2796 17500 2816
rect 17500 2796 17552 2816
rect 17552 2796 17554 2816
rect 17498 2760 17554 2796
rect 18142 4120 18198 4176
rect 18510 9832 18566 9888
rect 18326 9716 18382 9752
rect 18326 9696 18328 9716
rect 18328 9696 18380 9716
rect 18380 9696 18382 9716
rect 18418 9288 18474 9344
rect 18326 6160 18382 6216
rect 18234 3712 18290 3768
rect 18326 3304 18382 3360
rect 17590 1808 17646 1864
rect 9310 40 9366 96
rect 18326 2508 18382 2544
rect 18326 2488 18328 2508
rect 18328 2488 18380 2508
rect 18380 2488 18382 2508
rect 19062 22752 19118 22808
rect 18878 20440 18934 20496
rect 19062 21800 19118 21856
rect 18970 18400 19026 18456
rect 19062 18028 19064 18048
rect 19064 18028 19116 18048
rect 19116 18028 19118 18048
rect 19062 17992 19118 18028
rect 18878 16668 18880 16688
rect 18880 16668 18932 16688
rect 18932 16668 18934 16688
rect 18878 16632 18934 16668
rect 18878 12844 18934 12880
rect 18878 12824 18880 12844
rect 18880 12824 18932 12844
rect 18932 12824 18934 12844
rect 19430 22380 19432 22400
rect 19432 22380 19484 22400
rect 19484 22380 19486 22400
rect 19430 22344 19486 22380
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19614 23160 19670 23216
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19338 21528 19394 21584
rect 19522 21392 19578 21448
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19706 21004 19762 21040
rect 19706 20984 19708 21004
rect 19708 20984 19760 21004
rect 19760 20984 19762 21004
rect 19890 20868 19946 20904
rect 19890 20848 19892 20868
rect 19892 20848 19944 20868
rect 19944 20848 19946 20868
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19614 19896 19670 19952
rect 19522 19352 19578 19408
rect 19430 18828 19486 18864
rect 19430 18808 19432 18828
rect 19432 18808 19484 18828
rect 19484 18808 19486 18828
rect 19706 19216 19762 19272
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19430 17856 19486 17912
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 20350 25200 20406 25256
rect 20074 24112 20130 24168
rect 20626 24656 20682 24712
rect 21086 24248 21142 24304
rect 20074 21684 20130 21720
rect 20074 21664 20076 21684
rect 20076 21664 20128 21684
rect 20128 21664 20130 21684
rect 20074 20304 20130 20360
rect 20074 17756 20076 17776
rect 20076 17756 20128 17776
rect 20128 17756 20130 17776
rect 20074 17720 20130 17756
rect 19154 15408 19210 15464
rect 18694 3576 18750 3632
rect 18694 3440 18750 3496
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19430 16088 19486 16144
rect 19338 14356 19340 14376
rect 19340 14356 19392 14376
rect 19392 14356 19394 14376
rect 19338 14320 19394 14356
rect 19338 13504 19394 13560
rect 19614 16088 19670 16144
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 20074 15544 20130 15600
rect 21086 22208 21142 22264
rect 20442 19896 20498 19952
rect 20534 19760 20590 19816
rect 20442 18808 20498 18864
rect 20350 17740 20406 17776
rect 20350 17720 20352 17740
rect 20352 17720 20404 17740
rect 20404 17720 20406 17740
rect 20258 15952 20314 16008
rect 20074 14884 20130 14920
rect 20074 14864 20076 14884
rect 20076 14864 20128 14884
rect 20128 14864 20130 14884
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19982 14456 20038 14512
rect 19706 14068 19762 14104
rect 19706 14048 19708 14068
rect 19708 14048 19760 14068
rect 19760 14048 19762 14068
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 20994 20712 21050 20768
rect 20718 20460 20774 20496
rect 20718 20440 20720 20460
rect 20720 20440 20772 20460
rect 20772 20440 20774 20460
rect 20718 20168 20774 20224
rect 20810 19896 20866 19952
rect 21178 19624 21234 19680
rect 20902 19352 20958 19408
rect 20534 16632 20590 16688
rect 20718 18672 20774 18728
rect 20718 18148 20774 18184
rect 20718 18128 20720 18148
rect 20720 18128 20772 18148
rect 20772 18128 20774 18148
rect 20718 17992 20774 18048
rect 20626 15680 20682 15736
rect 20626 15564 20682 15600
rect 20626 15544 20628 15564
rect 20628 15544 20680 15564
rect 20680 15544 20682 15564
rect 20626 14456 20682 14512
rect 20258 12980 20314 13016
rect 20258 12960 20260 12980
rect 20260 12960 20312 12980
rect 20312 12960 20314 12980
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19154 10260 19210 10296
rect 19154 10240 19156 10260
rect 19156 10240 19208 10260
rect 19208 10240 19210 10260
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19522 10124 19578 10160
rect 19522 10104 19524 10124
rect 19524 10104 19576 10124
rect 19576 10104 19578 10124
rect 19338 9560 19394 9616
rect 19890 9460 19892 9480
rect 19892 9460 19944 9480
rect 19944 9460 19946 9480
rect 19890 9424 19946 9460
rect 19430 9324 19432 9344
rect 19432 9324 19484 9344
rect 19484 9324 19486 9344
rect 19430 9288 19486 9324
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19430 9016 19486 9072
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19430 6876 19432 6896
rect 19432 6876 19484 6896
rect 19484 6876 19486 6896
rect 19430 6840 19486 6876
rect 19522 6740 19524 6760
rect 19524 6740 19576 6760
rect 19576 6740 19578 6760
rect 19522 6704 19578 6740
rect 19154 6452 19210 6488
rect 19154 6432 19156 6452
rect 19156 6432 19208 6452
rect 19208 6432 19210 6452
rect 18970 5616 19026 5672
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19982 4528 20038 4584
rect 19430 3848 19486 3904
rect 19338 3712 19394 3768
rect 18786 3304 18842 3360
rect 18694 3168 18750 3224
rect 18510 1944 18566 2000
rect 18326 1672 18382 1728
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19614 3068 19616 3088
rect 19616 3068 19668 3088
rect 19668 3068 19670 3088
rect 19614 3032 19670 3068
rect 20626 14048 20682 14104
rect 20626 13912 20682 13968
rect 20718 13812 20720 13832
rect 20720 13812 20772 13832
rect 20772 13812 20774 13832
rect 20718 13776 20774 13812
rect 20994 15952 21050 16008
rect 20994 15408 21050 15464
rect 20994 15136 21050 15192
rect 20994 14592 21050 14648
rect 20994 12708 21050 12744
rect 20994 12688 20996 12708
rect 20996 12688 21048 12708
rect 21048 12688 21050 12708
rect 20810 12144 20866 12200
rect 20718 11192 20774 11248
rect 20902 11464 20958 11520
rect 20902 10920 20958 10976
rect 20350 8064 20406 8120
rect 20350 7520 20406 7576
rect 20534 9172 20590 9208
rect 20534 9152 20536 9172
rect 20536 9152 20588 9172
rect 20588 9152 20590 9172
rect 21178 17992 21234 18048
rect 21178 15036 21180 15056
rect 21180 15036 21232 15056
rect 21232 15036 21234 15056
rect 21178 15000 21234 15036
rect 21178 13232 21234 13288
rect 21086 12164 21142 12200
rect 21086 12144 21088 12164
rect 21088 12144 21140 12164
rect 21140 12144 21142 12164
rect 21086 11600 21142 11656
rect 20534 8608 20590 8664
rect 20810 7928 20866 7984
rect 20810 7792 20866 7848
rect 20442 5888 20498 5944
rect 20350 5208 20406 5264
rect 20074 2796 20076 2816
rect 20076 2796 20128 2816
rect 20128 2796 20130 2816
rect 20074 2760 20130 2796
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20810 6296 20866 6352
rect 21822 23432 21878 23488
rect 21362 18708 21364 18728
rect 21364 18708 21416 18728
rect 21416 18708 21418 18728
rect 21362 18672 21418 18708
rect 21362 18264 21418 18320
rect 21362 11600 21418 11656
rect 21362 11192 21418 11248
rect 22190 23840 22246 23896
rect 21822 22616 21878 22672
rect 21638 21392 21694 21448
rect 21638 20576 21694 20632
rect 21546 17584 21602 17640
rect 21638 15680 21694 15736
rect 21546 15272 21602 15328
rect 21546 14220 21548 14240
rect 21548 14220 21600 14240
rect 21600 14220 21602 14240
rect 21546 14184 21602 14220
rect 21638 14048 21694 14104
rect 21546 12008 21602 12064
rect 21362 6568 21418 6624
rect 21822 21936 21878 21992
rect 22098 21428 22100 21448
rect 22100 21428 22152 21448
rect 22152 21428 22154 21448
rect 22098 21392 22154 21428
rect 21914 18944 21970 19000
rect 22650 25064 22706 25120
rect 22374 22072 22430 22128
rect 22282 21972 22284 21992
rect 22284 21972 22336 21992
rect 22336 21972 22338 21992
rect 22282 21936 22338 21972
rect 22282 21392 22338 21448
rect 22282 20748 22284 20768
rect 22284 20748 22336 20768
rect 22336 20748 22338 20768
rect 22282 20712 22338 20748
rect 21914 18264 21970 18320
rect 21914 18128 21970 18184
rect 21822 17992 21878 18048
rect 21822 17856 21878 17912
rect 22006 17720 22062 17776
rect 22374 18536 22430 18592
rect 22374 17448 22430 17504
rect 21822 12824 21878 12880
rect 22006 12280 22062 12336
rect 22006 10920 22062 10976
rect 21730 8336 21786 8392
rect 21178 5616 21234 5672
rect 20442 3984 20498 4040
rect 19982 1808 20038 1864
rect 20166 1672 20222 1728
rect 17590 312 17646 368
rect 21454 5208 21510 5264
rect 20902 3984 20958 4040
rect 21178 4392 21234 4448
rect 20994 3440 21050 3496
rect 19430 176 19486 232
rect 21270 3440 21326 3496
rect 22282 12280 22338 12336
rect 22282 9696 22338 9752
rect 22190 8780 22192 8800
rect 22192 8780 22244 8800
rect 22244 8780 22246 8800
rect 22190 8744 22246 8780
rect 22190 8628 22246 8664
rect 22190 8608 22192 8628
rect 22192 8608 22244 8628
rect 22244 8608 22246 8628
rect 22006 7520 22062 7576
rect 21914 6432 21970 6488
rect 22466 15136 22522 15192
rect 23386 27104 23442 27160
rect 23202 26560 23258 26616
rect 22742 21392 22798 21448
rect 23018 22208 23074 22264
rect 23018 21936 23074 21992
rect 22742 16904 22798 16960
rect 22742 15000 22798 15056
rect 22650 12960 22706 13016
rect 22650 12824 22706 12880
rect 22926 18536 22982 18592
rect 22926 16360 22982 16416
rect 22926 16224 22982 16280
rect 23570 25880 23626 25936
rect 23110 21528 23166 21584
rect 23110 20032 23166 20088
rect 23386 23568 23442 23624
rect 23478 22208 23534 22264
rect 23478 20984 23534 21040
rect 23386 20304 23442 20360
rect 23202 19080 23258 19136
rect 23294 18536 23350 18592
rect 23478 19624 23534 19680
rect 23294 18264 23350 18320
rect 23202 17584 23258 17640
rect 23110 17196 23166 17232
rect 23110 17176 23112 17196
rect 23112 17176 23164 17196
rect 23164 17176 23166 17196
rect 23110 16904 23166 16960
rect 23110 14048 23166 14104
rect 23294 17176 23350 17232
rect 23386 16788 23442 16824
rect 23386 16768 23388 16788
rect 23388 16768 23440 16788
rect 23440 16768 23442 16788
rect 23386 16360 23442 16416
rect 23846 24112 23902 24168
rect 24674 25880 24730 25936
rect 24122 24792 24178 24848
rect 24122 24012 24124 24032
rect 24124 24012 24176 24032
rect 24176 24012 24178 24032
rect 24122 23976 24178 24012
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24858 24556 24860 24576
rect 24860 24556 24912 24576
rect 24912 24556 24914 24576
rect 24858 24520 24914 24556
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24306 23568 24362 23624
rect 24122 23432 24178 23488
rect 23846 22480 23902 22536
rect 23754 18420 23810 18456
rect 23754 18400 23756 18420
rect 23756 18400 23808 18420
rect 23808 18400 23810 18420
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24398 22344 24454 22400
rect 24122 22108 24124 22128
rect 24124 22108 24176 22128
rect 24176 22108 24178 22128
rect 24122 22072 24178 22108
rect 24398 22072 24454 22128
rect 25778 26152 25834 26208
rect 25410 25336 25466 25392
rect 25410 24792 25466 24848
rect 25318 24656 25374 24712
rect 25226 24112 25282 24168
rect 25042 23024 25098 23080
rect 24766 22480 24822 22536
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 23938 21392 23994 21448
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 23938 17992 23994 18048
rect 23754 17332 23810 17368
rect 23754 17312 23756 17332
rect 23756 17312 23808 17332
rect 23808 17312 23810 17332
rect 23662 16632 23718 16688
rect 23570 16496 23626 16552
rect 23478 14864 23534 14920
rect 23202 13504 23258 13560
rect 22926 12824 22982 12880
rect 23202 13096 23258 13152
rect 22834 12688 22890 12744
rect 22742 10684 22744 10704
rect 22744 10684 22796 10704
rect 22796 10684 22798 10704
rect 22742 10648 22798 10684
rect 22742 10260 22798 10296
rect 22742 10240 22744 10260
rect 22744 10240 22796 10260
rect 22796 10240 22798 10260
rect 22834 9152 22890 9208
rect 23018 11600 23074 11656
rect 23018 10004 23020 10024
rect 23020 10004 23072 10024
rect 23072 10004 23074 10024
rect 23018 9968 23074 10004
rect 22834 8064 22890 8120
rect 22466 6840 22522 6896
rect 22098 4120 22154 4176
rect 21546 3032 21602 3088
rect 21638 2644 21694 2680
rect 21638 2624 21640 2644
rect 21640 2624 21692 2644
rect 21692 2624 21694 2644
rect 21730 2388 21732 2408
rect 21732 2388 21784 2408
rect 21784 2388 21786 2408
rect 21730 2352 21786 2388
rect 23202 11636 23204 11656
rect 23204 11636 23256 11656
rect 23256 11636 23258 11656
rect 23202 11600 23258 11636
rect 23662 14184 23718 14240
rect 23662 13504 23718 13560
rect 23662 12416 23718 12472
rect 23570 12144 23626 12200
rect 23386 11872 23442 11928
rect 23202 9696 23258 9752
rect 23478 10956 23480 10976
rect 23480 10956 23532 10976
rect 23532 10956 23534 10976
rect 23478 10920 23534 10956
rect 23202 5888 23258 5944
rect 22926 3612 22928 3632
rect 22928 3612 22980 3632
rect 22980 3612 22982 3632
rect 22926 3576 22982 3612
rect 23110 3032 23166 3088
rect 22742 1808 22798 1864
rect 23018 1400 23074 1456
rect 23662 8472 23718 8528
rect 23478 7148 23480 7168
rect 23480 7148 23532 7168
rect 23532 7148 23534 7168
rect 23478 7112 23534 7148
rect 23478 6180 23534 6216
rect 23478 6160 23480 6180
rect 23480 6160 23532 6180
rect 23532 6160 23534 6180
rect 23478 5752 23534 5808
rect 24490 19796 24492 19816
rect 24492 19796 24544 19816
rect 24544 19796 24546 19816
rect 24030 17856 24086 17912
rect 24490 19760 24546 19796
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24582 19388 24584 19408
rect 24584 19388 24636 19408
rect 24636 19388 24638 19408
rect 24582 19352 24638 19388
rect 24490 18964 24546 19000
rect 24490 18944 24492 18964
rect 24492 18944 24544 18964
rect 24544 18944 24546 18964
rect 25042 21292 25044 21312
rect 25044 21292 25096 21312
rect 25096 21292 25098 21312
rect 25042 21256 25098 21292
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24858 19080 24914 19136
rect 24766 17448 24822 17504
rect 24858 17176 24914 17232
rect 24030 15700 24086 15736
rect 24030 15680 24032 15700
rect 24032 15680 24084 15700
rect 24084 15680 24086 15700
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24306 15000 24362 15056
rect 25226 20168 25282 20224
rect 25226 18164 25228 18184
rect 25228 18164 25280 18184
rect 25280 18164 25282 18184
rect 25226 18128 25282 18164
rect 25410 22616 25466 22672
rect 25410 21800 25466 21856
rect 25594 25336 25650 25392
rect 25594 23568 25650 23624
rect 25686 23024 25742 23080
rect 25594 21256 25650 21312
rect 25410 17312 25466 17368
rect 25410 17040 25466 17096
rect 25318 16632 25374 16688
rect 24858 16088 24914 16144
rect 24858 15408 24914 15464
rect 24214 14476 24270 14512
rect 24214 14456 24216 14476
rect 24216 14456 24268 14476
rect 24268 14456 24270 14476
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24122 12436 24178 12472
rect 24122 12416 24124 12436
rect 24124 12416 24176 12436
rect 24176 12416 24178 12436
rect 24766 13268 24768 13288
rect 24768 13268 24820 13288
rect 24820 13268 24822 13288
rect 24766 13232 24822 13268
rect 24766 12960 24822 13016
rect 25226 15544 25282 15600
rect 24858 12824 24914 12880
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 23938 11056 23994 11112
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 23938 10648 23994 10704
rect 24674 10512 24730 10568
rect 24214 10240 24270 10296
rect 24122 10104 24178 10160
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24214 9560 24270 9616
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24214 8472 24270 8528
rect 24950 11600 25006 11656
rect 24950 10240 25006 10296
rect 24214 7928 24270 7984
rect 24030 7792 24086 7848
rect 23662 4664 23718 4720
rect 23662 4428 23664 4448
rect 23664 4428 23716 4448
rect 23716 4428 23718 4448
rect 23662 4392 23718 4428
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24214 7248 24270 7304
rect 24030 6724 24086 6760
rect 24030 6704 24032 6724
rect 24032 6704 24084 6724
rect 24084 6704 24086 6724
rect 24030 6024 24086 6080
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 25226 14220 25228 14240
rect 25228 14220 25280 14240
rect 25280 14220 25282 14240
rect 25226 14184 25282 14220
rect 25226 13912 25282 13968
rect 25134 11872 25190 11928
rect 25410 11464 25466 11520
rect 25134 11192 25190 11248
rect 25318 11056 25374 11112
rect 25134 9988 25190 10024
rect 25134 9968 25136 9988
rect 25136 9968 25188 9988
rect 25188 9968 25190 9988
rect 25134 8608 25190 8664
rect 25134 7112 25190 7168
rect 24214 5616 24270 5672
rect 24122 5344 24178 5400
rect 24122 4256 24178 4312
rect 23938 3304 23994 3360
rect 24030 3168 24086 3224
rect 23662 2796 23664 2816
rect 23664 2796 23716 2816
rect 23716 2796 23718 2816
rect 23662 2760 23718 2796
rect 23938 2644 23994 2680
rect 23938 2624 23940 2644
rect 23940 2624 23992 2644
rect 23992 2624 23994 2644
rect 23570 2488 23626 2544
rect 23662 2388 23664 2408
rect 23664 2388 23716 2408
rect 23716 2388 23718 2408
rect 23662 2352 23718 2388
rect 23478 2252 23480 2272
rect 23480 2252 23532 2272
rect 23532 2252 23534 2272
rect 23478 2216 23534 2252
rect 24766 5480 24822 5536
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24306 4936 24362 4992
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 25226 5616 25282 5672
rect 25042 4392 25098 4448
rect 24490 3712 24546 3768
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 24030 1128 24086 1184
rect 23478 856 23534 912
rect 24674 1536 24730 1592
rect 25042 3576 25098 3632
rect 25226 2896 25282 2952
rect 24950 1264 25006 1320
rect 25962 22344 26018 22400
rect 25870 21664 25926 21720
rect 25870 21528 25926 21584
rect 25778 16496 25834 16552
rect 27618 25608 27674 25664
rect 25962 11736 26018 11792
rect 25686 4120 25742 4176
rect 25962 6024 26018 6080
rect 26238 19760 26294 19816
rect 26422 18944 26478 19000
rect 26330 18284 26386 18320
rect 26330 18264 26332 18284
rect 26332 18264 26384 18284
rect 26384 18264 26386 18284
rect 26330 17584 26386 17640
rect 26330 10784 26386 10840
rect 25962 5072 26018 5128
rect 25594 1944 25650 2000
rect 25502 992 25558 1048
rect 25870 1944 25926 2000
rect 21086 40 21142 96
rect 26330 4020 26332 4040
rect 26332 4020 26384 4040
rect 26384 4020 26386 4040
rect 26330 3984 26386 4020
rect 26330 3440 26386 3496
rect 26606 2624 26662 2680
rect 26514 1672 26570 1728
rect 27618 4120 27674 4176
rect 26790 1400 26846 1456
rect 27158 1400 27214 1456
rect 26238 312 26294 368
<< metal3 >>
rect 0 27706 480 27736
rect 3509 27706 3575 27709
rect 0 27704 3575 27706
rect 0 27648 3514 27704
rect 3570 27648 3575 27704
rect 0 27646 3575 27648
rect 0 27616 480 27646
rect 3509 27643 3575 27646
rect 26049 27706 26115 27709
rect 27520 27706 28000 27736
rect 26049 27704 28000 27706
rect 26049 27648 26054 27704
rect 26110 27648 28000 27704
rect 26049 27646 28000 27648
rect 26049 27643 26115 27646
rect 27520 27616 28000 27646
rect 0 27162 480 27192
rect 1669 27162 1735 27165
rect 0 27160 1735 27162
rect 0 27104 1674 27160
rect 1730 27104 1735 27160
rect 0 27102 1735 27104
rect 0 27072 480 27102
rect 1669 27099 1735 27102
rect 23381 27162 23447 27165
rect 27520 27162 28000 27192
rect 23381 27160 28000 27162
rect 23381 27104 23386 27160
rect 23442 27104 28000 27160
rect 23381 27102 28000 27104
rect 23381 27099 23447 27102
rect 27520 27072 28000 27102
rect 0 26618 480 26648
rect 1485 26618 1551 26621
rect 0 26616 1551 26618
rect 0 26560 1490 26616
rect 1546 26560 1551 26616
rect 0 26558 1551 26560
rect 0 26528 480 26558
rect 1485 26555 1551 26558
rect 23197 26618 23263 26621
rect 27520 26618 28000 26648
rect 23197 26616 28000 26618
rect 23197 26560 23202 26616
rect 23258 26560 28000 26616
rect 23197 26558 28000 26560
rect 23197 26555 23263 26558
rect 27520 26528 28000 26558
rect 11789 26346 11855 26349
rect 17861 26346 17927 26349
rect 11789 26344 17927 26346
rect 11789 26288 11794 26344
rect 11850 26288 17866 26344
rect 17922 26288 17927 26344
rect 11789 26286 17927 26288
rect 11789 26283 11855 26286
rect 17861 26283 17927 26286
rect 10869 26210 10935 26213
rect 25773 26210 25839 26213
rect 10869 26208 25839 26210
rect 10869 26152 10874 26208
rect 10930 26152 25778 26208
rect 25834 26152 25839 26208
rect 10869 26150 25839 26152
rect 10869 26147 10935 26150
rect 25773 26147 25839 26150
rect 6085 26074 6151 26077
rect 15929 26074 15995 26077
rect 6085 26072 15995 26074
rect 6085 26016 6090 26072
rect 6146 26016 15934 26072
rect 15990 26016 15995 26072
rect 6085 26014 15995 26016
rect 6085 26011 6151 26014
rect 15929 26011 15995 26014
rect 16113 26074 16179 26077
rect 20110 26074 20116 26076
rect 16113 26072 20116 26074
rect 16113 26016 16118 26072
rect 16174 26016 20116 26072
rect 16113 26014 20116 26016
rect 16113 26011 16179 26014
rect 20110 26012 20116 26014
rect 20180 26012 20186 26076
rect 0 25938 480 25968
rect 2681 25938 2747 25941
rect 0 25936 2747 25938
rect 0 25880 2686 25936
rect 2742 25880 2747 25936
rect 0 25878 2747 25880
rect 0 25848 480 25878
rect 2681 25875 2747 25878
rect 8109 25938 8175 25941
rect 14457 25938 14523 25941
rect 8109 25936 14523 25938
rect 8109 25880 8114 25936
rect 8170 25880 14462 25936
rect 14518 25880 14523 25936
rect 8109 25878 14523 25880
rect 8109 25875 8175 25878
rect 14457 25875 14523 25878
rect 14590 25876 14596 25940
rect 14660 25938 14666 25940
rect 23565 25938 23631 25941
rect 14660 25936 23631 25938
rect 14660 25880 23570 25936
rect 23626 25880 23631 25936
rect 14660 25878 23631 25880
rect 14660 25876 14666 25878
rect 23565 25875 23631 25878
rect 24669 25938 24735 25941
rect 27520 25938 28000 25968
rect 24669 25936 28000 25938
rect 24669 25880 24674 25936
rect 24730 25880 28000 25936
rect 24669 25878 28000 25880
rect 24669 25875 24735 25878
rect 27520 25848 28000 25878
rect 7925 25802 7991 25805
rect 7925 25800 24962 25802
rect 7925 25744 7930 25800
rect 7986 25744 24962 25800
rect 7925 25742 24962 25744
rect 7925 25739 7991 25742
rect 11513 25666 11579 25669
rect 24902 25666 24962 25742
rect 27613 25666 27679 25669
rect 11513 25664 17234 25666
rect 11513 25608 11518 25664
rect 11574 25608 17234 25664
rect 11513 25606 17234 25608
rect 24902 25664 27679 25666
rect 24902 25608 27618 25664
rect 27674 25608 27679 25664
rect 24902 25606 27679 25608
rect 11513 25603 11579 25606
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 14038 25468 14044 25532
rect 14108 25530 14114 25532
rect 17033 25530 17099 25533
rect 14108 25528 17099 25530
rect 14108 25472 17038 25528
rect 17094 25472 17099 25528
rect 14108 25470 17099 25472
rect 14108 25468 14114 25470
rect 17033 25467 17099 25470
rect 0 25394 480 25424
rect 1577 25394 1643 25397
rect 0 25392 1643 25394
rect 0 25336 1582 25392
rect 1638 25336 1643 25392
rect 0 25334 1643 25336
rect 17174 25394 17234 25606
rect 27613 25603 27679 25606
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 25405 25394 25471 25397
rect 17174 25392 25471 25394
rect 17174 25336 25410 25392
rect 25466 25336 25471 25392
rect 17174 25334 25471 25336
rect 0 25304 480 25334
rect 1577 25331 1643 25334
rect 25405 25331 25471 25334
rect 25589 25394 25655 25397
rect 27520 25394 28000 25424
rect 25589 25392 28000 25394
rect 25589 25336 25594 25392
rect 25650 25336 28000 25392
rect 25589 25334 28000 25336
rect 25589 25331 25655 25334
rect 27520 25304 28000 25334
rect 11278 25196 11284 25260
rect 11348 25258 11354 25260
rect 20345 25258 20411 25261
rect 11348 25256 20411 25258
rect 11348 25200 20350 25256
rect 20406 25200 20411 25256
rect 11348 25198 20411 25200
rect 11348 25196 11354 25198
rect 20345 25195 20411 25198
rect 9673 25122 9739 25125
rect 13537 25122 13603 25125
rect 22645 25122 22711 25125
rect 9673 25120 13603 25122
rect 9673 25064 9678 25120
rect 9734 25064 13542 25120
rect 13598 25064 13603 25120
rect 9673 25062 13603 25064
rect 9673 25059 9739 25062
rect 13537 25059 13603 25062
rect 15334 25120 22711 25122
rect 15334 25064 22650 25120
rect 22706 25064 22711 25120
rect 15334 25062 22711 25064
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 9489 24986 9555 24989
rect 12893 24986 12959 24989
rect 9489 24984 12959 24986
rect 9489 24928 9494 24984
rect 9550 24928 12898 24984
rect 12954 24928 12959 24984
rect 9489 24926 12959 24928
rect 9489 24923 9555 24926
rect 12893 24923 12959 24926
rect 13670 24924 13676 24988
rect 13740 24986 13746 24988
rect 14273 24986 14339 24989
rect 13740 24984 14339 24986
rect 13740 24928 14278 24984
rect 14334 24928 14339 24984
rect 13740 24926 14339 24928
rect 13740 24924 13746 24926
rect 14273 24923 14339 24926
rect 0 24850 480 24880
rect 1577 24850 1643 24853
rect 0 24848 1643 24850
rect 0 24792 1582 24848
rect 1638 24792 1643 24848
rect 0 24790 1643 24792
rect 0 24760 480 24790
rect 1577 24787 1643 24790
rect 9029 24850 9095 24853
rect 9765 24850 9831 24853
rect 9029 24848 9831 24850
rect 9029 24792 9034 24848
rect 9090 24792 9770 24848
rect 9826 24792 9831 24848
rect 9029 24790 9831 24792
rect 9029 24787 9095 24790
rect 9765 24787 9831 24790
rect 14917 24850 14983 24853
rect 15334 24850 15394 25062
rect 22645 25059 22711 25062
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 15929 24986 15995 24989
rect 18045 24986 18111 24989
rect 15929 24984 18111 24986
rect 15929 24928 15934 24984
rect 15990 24928 18050 24984
rect 18106 24928 18111 24984
rect 15929 24926 18111 24928
rect 15929 24923 15995 24926
rect 18045 24923 18111 24926
rect 14917 24848 15394 24850
rect 14917 24792 14922 24848
rect 14978 24792 15394 24848
rect 14917 24790 15394 24792
rect 14917 24787 14983 24790
rect 15510 24788 15516 24852
rect 15580 24850 15586 24852
rect 16021 24850 16087 24853
rect 15580 24848 16087 24850
rect 15580 24792 16026 24848
rect 16082 24792 16087 24848
rect 15580 24790 16087 24792
rect 15580 24788 15586 24790
rect 16021 24787 16087 24790
rect 17033 24850 17099 24853
rect 17033 24848 23490 24850
rect 17033 24792 17038 24848
rect 17094 24792 23490 24848
rect 17033 24790 23490 24792
rect 17033 24787 17099 24790
rect 7741 24714 7807 24717
rect 11421 24714 11487 24717
rect 20621 24714 20687 24717
rect 7741 24712 11346 24714
rect 7741 24656 7746 24712
rect 7802 24656 11346 24712
rect 7741 24654 11346 24656
rect 7741 24651 7807 24654
rect 11286 24578 11346 24654
rect 11421 24712 20687 24714
rect 11421 24656 11426 24712
rect 11482 24656 20626 24712
rect 20682 24656 20687 24712
rect 11421 24654 20687 24656
rect 23430 24714 23490 24790
rect 23606 24788 23612 24852
rect 23676 24850 23682 24852
rect 24117 24850 24183 24853
rect 23676 24848 24183 24850
rect 23676 24792 24122 24848
rect 24178 24792 24183 24848
rect 23676 24790 24183 24792
rect 23676 24788 23682 24790
rect 24117 24787 24183 24790
rect 25405 24850 25471 24853
rect 27520 24850 28000 24880
rect 25405 24848 28000 24850
rect 25405 24792 25410 24848
rect 25466 24792 28000 24848
rect 25405 24790 28000 24792
rect 25405 24787 25471 24790
rect 27520 24760 28000 24790
rect 25313 24714 25379 24717
rect 23430 24712 25379 24714
rect 23430 24656 25318 24712
rect 25374 24656 25379 24712
rect 23430 24654 25379 24656
rect 11421 24651 11487 24654
rect 20621 24651 20687 24654
rect 25313 24651 25379 24654
rect 14457 24578 14523 24581
rect 11286 24576 14523 24578
rect 11286 24520 14462 24576
rect 14518 24520 14523 24576
rect 11286 24518 14523 24520
rect 14457 24515 14523 24518
rect 15101 24578 15167 24581
rect 16849 24578 16915 24581
rect 15101 24576 16915 24578
rect 15101 24520 15106 24576
rect 15162 24520 16854 24576
rect 16910 24520 16915 24576
rect 15101 24518 16915 24520
rect 15101 24515 15167 24518
rect 16849 24515 16915 24518
rect 20662 24516 20668 24580
rect 20732 24578 20738 24580
rect 24853 24578 24919 24581
rect 20732 24576 24919 24578
rect 20732 24520 24858 24576
rect 24914 24520 24919 24576
rect 20732 24518 24919 24520
rect 20732 24516 20738 24518
rect 24853 24515 24919 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 12893 24442 12959 24445
rect 13486 24442 13492 24444
rect 12893 24440 13492 24442
rect 12893 24384 12898 24440
rect 12954 24384 13492 24440
rect 12893 24382 13492 24384
rect 12893 24379 12959 24382
rect 13486 24380 13492 24382
rect 13556 24442 13562 24444
rect 15561 24442 15627 24445
rect 13556 24440 15627 24442
rect 13556 24384 15566 24440
rect 15622 24384 15627 24440
rect 13556 24382 15627 24384
rect 13556 24380 13562 24382
rect 15561 24379 15627 24382
rect 15694 24380 15700 24444
rect 15764 24442 15770 24444
rect 19057 24442 19123 24445
rect 15764 24440 19123 24442
rect 15764 24384 19062 24440
rect 19118 24384 19123 24440
rect 15764 24382 19123 24384
rect 15764 24380 15770 24382
rect 19057 24379 19123 24382
rect 8661 24306 8727 24309
rect 17677 24306 17743 24309
rect 8661 24304 17743 24306
rect 8661 24248 8666 24304
rect 8722 24248 17682 24304
rect 17738 24248 17743 24304
rect 8661 24246 17743 24248
rect 8661 24243 8727 24246
rect 17677 24243 17743 24246
rect 18045 24306 18111 24309
rect 21081 24306 21147 24309
rect 18045 24304 21147 24306
rect 18045 24248 18050 24304
rect 18106 24248 21086 24304
rect 21142 24248 21147 24304
rect 18045 24246 21147 24248
rect 18045 24243 18111 24246
rect 21081 24243 21147 24246
rect 0 24170 480 24200
rect 1393 24170 1459 24173
rect 0 24168 1459 24170
rect 0 24112 1398 24168
rect 1454 24112 1459 24168
rect 0 24110 1459 24112
rect 0 24080 480 24110
rect 1393 24107 1459 24110
rect 10409 24170 10475 24173
rect 20069 24170 20135 24173
rect 10409 24168 20135 24170
rect 10409 24112 10414 24168
rect 10470 24112 20074 24168
rect 20130 24112 20135 24168
rect 10409 24110 20135 24112
rect 10409 24107 10475 24110
rect 20069 24107 20135 24110
rect 23841 24170 23907 24173
rect 23974 24170 23980 24172
rect 23841 24168 23980 24170
rect 23841 24112 23846 24168
rect 23902 24112 23980 24168
rect 23841 24110 23980 24112
rect 23841 24107 23907 24110
rect 23974 24108 23980 24110
rect 24044 24108 24050 24172
rect 25221 24170 25287 24173
rect 27520 24170 28000 24200
rect 25221 24168 28000 24170
rect 25221 24112 25226 24168
rect 25282 24112 28000 24168
rect 25221 24110 28000 24112
rect 25221 24107 25287 24110
rect 27520 24080 28000 24110
rect 17125 24034 17191 24037
rect 24117 24034 24183 24037
rect 17125 24032 24183 24034
rect 17125 23976 17130 24032
rect 17186 23976 24122 24032
rect 24178 23976 24183 24032
rect 17125 23974 24183 23976
rect 17125 23971 17191 23974
rect 24117 23971 24183 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 15469 23898 15535 23901
rect 22185 23898 22251 23901
rect 15469 23896 22251 23898
rect 15469 23840 15474 23896
rect 15530 23840 22190 23896
rect 22246 23840 22251 23896
rect 15469 23838 22251 23840
rect 15469 23835 15535 23838
rect 22185 23835 22251 23838
rect 10225 23762 10291 23765
rect 9860 23760 10291 23762
rect 9860 23704 10230 23760
rect 10286 23704 10291 23760
rect 9860 23702 10291 23704
rect 0 23626 480 23656
rect 4061 23626 4127 23629
rect 0 23624 4127 23626
rect 0 23568 4066 23624
rect 4122 23568 4127 23624
rect 0 23566 4127 23568
rect 0 23536 480 23566
rect 4061 23563 4127 23566
rect 8845 23490 8911 23493
rect 9860 23490 9920 23702
rect 10225 23699 10291 23702
rect 13537 23762 13603 23765
rect 15929 23764 15995 23765
rect 15326 23762 15332 23764
rect 13537 23760 15332 23762
rect 13537 23704 13542 23760
rect 13598 23704 15332 23760
rect 13537 23702 15332 23704
rect 13537 23699 13603 23702
rect 15326 23700 15332 23702
rect 15396 23700 15402 23764
rect 15878 23762 15884 23764
rect 15838 23702 15884 23762
rect 15948 23760 15995 23764
rect 15990 23704 15995 23760
rect 15878 23700 15884 23702
rect 15948 23700 15995 23704
rect 15929 23699 15995 23700
rect 16297 23762 16363 23765
rect 21398 23762 21404 23764
rect 16297 23760 21404 23762
rect 16297 23704 16302 23760
rect 16358 23704 21404 23760
rect 16297 23702 21404 23704
rect 16297 23699 16363 23702
rect 21398 23700 21404 23702
rect 21468 23700 21474 23764
rect 10041 23626 10107 23629
rect 15469 23626 15535 23629
rect 10041 23624 15535 23626
rect 10041 23568 10046 23624
rect 10102 23568 15474 23624
rect 15530 23568 15535 23624
rect 10041 23566 15535 23568
rect 10041 23563 10107 23566
rect 15469 23563 15535 23566
rect 15929 23626 15995 23629
rect 19006 23626 19012 23628
rect 15929 23624 19012 23626
rect 15929 23568 15934 23624
rect 15990 23568 19012 23624
rect 15929 23566 19012 23568
rect 15929 23563 15995 23566
rect 19006 23564 19012 23566
rect 19076 23564 19082 23628
rect 23054 23564 23060 23628
rect 23124 23626 23130 23628
rect 23381 23626 23447 23629
rect 23124 23624 23447 23626
rect 23124 23568 23386 23624
rect 23442 23568 23447 23624
rect 23124 23566 23447 23568
rect 23124 23564 23130 23566
rect 23381 23563 23447 23566
rect 24301 23626 24367 23629
rect 25262 23626 25268 23628
rect 24301 23624 25268 23626
rect 24301 23568 24306 23624
rect 24362 23568 25268 23624
rect 24301 23566 25268 23568
rect 24301 23563 24367 23566
rect 25262 23564 25268 23566
rect 25332 23564 25338 23628
rect 25589 23626 25655 23629
rect 27520 23626 28000 23656
rect 25589 23624 28000 23626
rect 25589 23568 25594 23624
rect 25650 23568 28000 23624
rect 25589 23566 28000 23568
rect 25589 23563 25655 23566
rect 27520 23536 28000 23566
rect 12341 23492 12407 23493
rect 12341 23490 12388 23492
rect 8845 23488 9920 23490
rect 8845 23432 8850 23488
rect 8906 23432 9920 23488
rect 8845 23430 9920 23432
rect 12296 23488 12388 23490
rect 12296 23432 12346 23488
rect 12296 23430 12388 23432
rect 8845 23427 8911 23430
rect 12341 23428 12388 23430
rect 12452 23428 12458 23492
rect 12985 23490 13051 23493
rect 14774 23490 14780 23492
rect 12985 23488 14780 23490
rect 12985 23432 12990 23488
rect 13046 23432 14780 23488
rect 12985 23430 14780 23432
rect 12341 23427 12407 23428
rect 12985 23427 13051 23430
rect 14774 23428 14780 23430
rect 14844 23428 14850 23492
rect 15653 23490 15719 23493
rect 18597 23490 18663 23493
rect 15653 23488 18663 23490
rect 15653 23432 15658 23488
rect 15714 23432 18602 23488
rect 18658 23432 18663 23488
rect 15653 23430 18663 23432
rect 15653 23427 15719 23430
rect 18597 23427 18663 23430
rect 21817 23490 21883 23493
rect 24117 23490 24183 23493
rect 21817 23488 24183 23490
rect 21817 23432 21822 23488
rect 21878 23432 24122 23488
rect 24178 23432 24183 23488
rect 21817 23430 24183 23432
rect 21817 23427 21883 23430
rect 24117 23427 24183 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 841 23354 907 23357
rect 7189 23354 7255 23357
rect 841 23352 7255 23354
rect 841 23296 846 23352
rect 902 23296 7194 23352
rect 7250 23296 7255 23352
rect 841 23294 7255 23296
rect 841 23291 907 23294
rect 7189 23291 7255 23294
rect 14825 23354 14891 23357
rect 18413 23354 18479 23357
rect 14825 23352 18479 23354
rect 14825 23296 14830 23352
rect 14886 23296 18418 23352
rect 18474 23296 18479 23352
rect 14825 23294 18479 23296
rect 14825 23291 14891 23294
rect 18413 23291 18479 23294
rect 2037 23218 2103 23221
rect 6453 23218 6519 23221
rect 2037 23216 6519 23218
rect 2037 23160 2042 23216
rect 2098 23160 6458 23216
rect 6514 23160 6519 23216
rect 2037 23158 6519 23160
rect 2037 23155 2103 23158
rect 6453 23155 6519 23158
rect 6637 23218 6703 23221
rect 8661 23218 8727 23221
rect 6637 23216 8727 23218
rect 6637 23160 6642 23216
rect 6698 23160 8666 23216
rect 8722 23160 8727 23216
rect 6637 23158 8727 23160
rect 6637 23155 6703 23158
rect 8661 23155 8727 23158
rect 13445 23218 13511 23221
rect 15285 23218 15351 23221
rect 13445 23216 15351 23218
rect 13445 23160 13450 23216
rect 13506 23160 15290 23216
rect 15346 23160 15351 23216
rect 13445 23158 15351 23160
rect 13445 23155 13511 23158
rect 15285 23155 15351 23158
rect 16849 23218 16915 23221
rect 19609 23218 19675 23221
rect 16849 23216 19675 23218
rect 16849 23160 16854 23216
rect 16910 23160 19614 23216
rect 19670 23160 19675 23216
rect 16849 23158 19675 23160
rect 16849 23155 16915 23158
rect 19609 23155 19675 23158
rect 0 23082 480 23112
rect 1485 23082 1551 23085
rect 0 23080 1551 23082
rect 0 23024 1490 23080
rect 1546 23024 1551 23080
rect 0 23022 1551 23024
rect 0 22992 480 23022
rect 1485 23019 1551 23022
rect 1669 23082 1735 23085
rect 10910 23082 10916 23084
rect 1669 23080 10916 23082
rect 1669 23024 1674 23080
rect 1730 23024 10916 23080
rect 1669 23022 10916 23024
rect 1669 23019 1735 23022
rect 10910 23020 10916 23022
rect 10980 23020 10986 23084
rect 15929 23082 15995 23085
rect 18137 23082 18203 23085
rect 25037 23082 25103 23085
rect 15929 23080 18203 23082
rect 15929 23024 15934 23080
rect 15990 23024 18142 23080
rect 18198 23024 18203 23080
rect 15929 23022 18203 23024
rect 15929 23019 15995 23022
rect 18137 23019 18203 23022
rect 23982 23080 25103 23082
rect 23982 23024 25042 23080
rect 25098 23024 25103 23080
rect 23982 23022 25103 23024
rect 7373 22946 7439 22949
rect 11605 22946 11671 22949
rect 7373 22944 11671 22946
rect 7373 22888 7378 22944
rect 7434 22888 11610 22944
rect 11666 22888 11671 22944
rect 7373 22886 11671 22888
rect 7373 22883 7439 22886
rect 11605 22883 11671 22886
rect 15653 22946 15719 22949
rect 23982 22946 24042 23022
rect 25037 23019 25103 23022
rect 25681 23082 25747 23085
rect 27520 23082 28000 23112
rect 25681 23080 28000 23082
rect 25681 23024 25686 23080
rect 25742 23024 28000 23080
rect 25681 23022 28000 23024
rect 25681 23019 25747 23022
rect 27520 22992 28000 23022
rect 15653 22944 24042 22946
rect 15653 22888 15658 22944
rect 15714 22888 24042 22944
rect 15653 22886 24042 22888
rect 15653 22883 15719 22886
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 7649 22810 7715 22813
rect 14181 22810 14247 22813
rect 7649 22808 14247 22810
rect 7649 22752 7654 22808
rect 7710 22752 14186 22808
rect 14242 22752 14247 22808
rect 7649 22750 14247 22752
rect 7649 22747 7715 22750
rect 14181 22747 14247 22750
rect 19057 22810 19123 22813
rect 19057 22808 24042 22810
rect 19057 22752 19062 22808
rect 19118 22752 24042 22808
rect 19057 22750 24042 22752
rect 19057 22747 19123 22750
rect 7281 22674 7347 22677
rect 7281 22672 11898 22674
rect 7281 22616 7286 22672
rect 7342 22616 11898 22672
rect 7281 22614 11898 22616
rect 7281 22611 7347 22614
rect 0 22538 480 22568
rect 1577 22538 1643 22541
rect 0 22536 1643 22538
rect 0 22480 1582 22536
rect 1638 22480 1643 22536
rect 0 22478 1643 22480
rect 0 22448 480 22478
rect 1577 22475 1643 22478
rect 2129 22538 2195 22541
rect 2681 22538 2747 22541
rect 2129 22536 2747 22538
rect 2129 22480 2134 22536
rect 2190 22480 2686 22536
rect 2742 22480 2747 22536
rect 2129 22478 2747 22480
rect 2129 22475 2195 22478
rect 2681 22475 2747 22478
rect 4705 22538 4771 22541
rect 11513 22538 11579 22541
rect 4705 22536 11579 22538
rect 4705 22480 4710 22536
rect 4766 22480 11518 22536
rect 11574 22480 11579 22536
rect 4705 22478 11579 22480
rect 11838 22538 11898 22614
rect 12014 22612 12020 22676
rect 12084 22674 12090 22676
rect 13813 22674 13879 22677
rect 21817 22674 21883 22677
rect 12084 22614 13186 22674
rect 12084 22612 12090 22614
rect 12341 22538 12407 22541
rect 11838 22536 12407 22538
rect 11838 22480 12346 22536
rect 12402 22480 12407 22536
rect 11838 22478 12407 22480
rect 4705 22475 4771 22478
rect 11513 22475 11579 22478
rect 12341 22475 12407 22478
rect 12525 22538 12591 22541
rect 12750 22538 12756 22540
rect 12525 22536 12756 22538
rect 12525 22480 12530 22536
rect 12586 22480 12756 22536
rect 12525 22478 12756 22480
rect 12525 22475 12591 22478
rect 12750 22476 12756 22478
rect 12820 22476 12826 22540
rect 13126 22538 13186 22614
rect 13813 22672 21883 22674
rect 13813 22616 13818 22672
rect 13874 22616 21822 22672
rect 21878 22616 21883 22672
rect 13813 22614 21883 22616
rect 23982 22674 24042 22750
rect 25405 22674 25471 22677
rect 23982 22672 25471 22674
rect 23982 22616 25410 22672
rect 25466 22616 25471 22672
rect 23982 22614 25471 22616
rect 13813 22611 13879 22614
rect 21817 22611 21883 22614
rect 25405 22611 25471 22614
rect 16389 22538 16455 22541
rect 18229 22538 18295 22541
rect 23841 22538 23907 22541
rect 13126 22536 18154 22538
rect 13126 22480 16394 22536
rect 16450 22480 18154 22536
rect 13126 22478 18154 22480
rect 16389 22475 16455 22478
rect 2405 22402 2471 22405
rect 3918 22402 3924 22404
rect 2405 22400 3924 22402
rect 2405 22344 2410 22400
rect 2466 22344 3924 22400
rect 2405 22342 3924 22344
rect 2405 22339 2471 22342
rect 3918 22340 3924 22342
rect 3988 22340 3994 22404
rect 5257 22402 5323 22405
rect 7465 22402 7531 22405
rect 8201 22402 8267 22405
rect 5257 22400 8267 22402
rect 5257 22344 5262 22400
rect 5318 22344 7470 22400
rect 7526 22344 8206 22400
rect 8262 22344 8267 22400
rect 5257 22342 8267 22344
rect 5257 22339 5323 22342
rect 7465 22339 7531 22342
rect 8201 22339 8267 22342
rect 11237 22402 11303 22405
rect 15837 22402 15903 22405
rect 11237 22400 15903 22402
rect 11237 22344 11242 22400
rect 11298 22344 15842 22400
rect 15898 22344 15903 22400
rect 11237 22342 15903 22344
rect 11237 22339 11303 22342
rect 15837 22339 15903 22342
rect 17125 22402 17191 22405
rect 17534 22402 17540 22404
rect 17125 22400 17540 22402
rect 17125 22344 17130 22400
rect 17186 22344 17540 22400
rect 17125 22342 17540 22344
rect 17125 22339 17191 22342
rect 17534 22340 17540 22342
rect 17604 22340 17610 22404
rect 18094 22402 18154 22478
rect 18229 22536 23907 22538
rect 18229 22480 18234 22536
rect 18290 22480 23846 22536
rect 23902 22480 23907 22536
rect 18229 22478 23907 22480
rect 18229 22475 18295 22478
rect 23841 22475 23907 22478
rect 24761 22538 24827 22541
rect 27520 22538 28000 22568
rect 24761 22536 28000 22538
rect 24761 22480 24766 22536
rect 24822 22480 28000 22536
rect 24761 22478 28000 22480
rect 24761 22475 24827 22478
rect 27520 22448 28000 22478
rect 18413 22402 18479 22405
rect 19425 22404 19491 22405
rect 18094 22400 18479 22402
rect 18094 22344 18418 22400
rect 18474 22344 18479 22400
rect 18094 22342 18479 22344
rect 18413 22339 18479 22342
rect 19374 22340 19380 22404
rect 19444 22402 19491 22404
rect 24393 22402 24459 22405
rect 25957 22402 26023 22405
rect 19444 22400 19536 22402
rect 19486 22344 19536 22400
rect 19444 22342 19536 22344
rect 24393 22400 26023 22402
rect 24393 22344 24398 22400
rect 24454 22344 25962 22400
rect 26018 22344 26023 22400
rect 24393 22342 26023 22344
rect 19444 22340 19491 22342
rect 19425 22339 19491 22340
rect 24393 22339 24459 22342
rect 25957 22339 26023 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 289 22266 355 22269
rect 2957 22266 3023 22269
rect 7097 22266 7163 22269
rect 289 22264 7163 22266
rect 289 22208 294 22264
rect 350 22208 2962 22264
rect 3018 22208 7102 22264
rect 7158 22208 7163 22264
rect 289 22206 7163 22208
rect 289 22203 355 22206
rect 2957 22203 3023 22206
rect 7097 22203 7163 22206
rect 15101 22266 15167 22269
rect 21081 22266 21147 22269
rect 23013 22266 23079 22269
rect 23473 22266 23539 22269
rect 15101 22264 18706 22266
rect 15101 22208 15106 22264
rect 15162 22208 18706 22264
rect 15101 22206 18706 22208
rect 15101 22203 15167 22206
rect 2681 22130 2747 22133
rect 4705 22130 4771 22133
rect 2681 22128 4771 22130
rect 2681 22072 2686 22128
rect 2742 22072 4710 22128
rect 4766 22072 4771 22128
rect 2681 22070 4771 22072
rect 2681 22067 2747 22070
rect 4705 22067 4771 22070
rect 9213 22130 9279 22133
rect 11881 22130 11947 22133
rect 13445 22132 13511 22133
rect 13445 22130 13492 22132
rect 9213 22128 11947 22130
rect 9213 22072 9218 22128
rect 9274 22072 11886 22128
rect 11942 22072 11947 22128
rect 9213 22070 11947 22072
rect 13400 22128 13492 22130
rect 13400 22072 13450 22128
rect 13400 22070 13492 22072
rect 9213 22067 9279 22070
rect 11881 22067 11947 22070
rect 13445 22068 13492 22070
rect 13556 22068 13562 22132
rect 18137 22130 18203 22133
rect 15104 22128 18203 22130
rect 15104 22072 18142 22128
rect 18198 22072 18203 22128
rect 15104 22070 18203 22072
rect 18646 22130 18706 22206
rect 21081 22264 23539 22266
rect 21081 22208 21086 22264
rect 21142 22208 23018 22264
rect 23074 22208 23478 22264
rect 23534 22208 23539 22264
rect 21081 22206 23539 22208
rect 21081 22203 21147 22206
rect 23013 22203 23079 22206
rect 23473 22203 23539 22206
rect 22369 22130 22435 22133
rect 18646 22128 22435 22130
rect 18646 22072 22374 22128
rect 22430 22072 22435 22128
rect 18646 22070 22435 22072
rect 13445 22067 13511 22068
rect 8385 21994 8451 21997
rect 9070 21994 9076 21996
rect 8385 21992 9076 21994
rect 8385 21936 8390 21992
rect 8446 21936 9076 21992
rect 8385 21934 9076 21936
rect 8385 21931 8451 21934
rect 9070 21932 9076 21934
rect 9140 21932 9146 21996
rect 9489 21994 9555 21997
rect 10685 21994 10751 21997
rect 9489 21992 10751 21994
rect 9489 21936 9494 21992
rect 9550 21936 10690 21992
rect 10746 21936 10751 21992
rect 9489 21934 10751 21936
rect 9489 21931 9555 21934
rect 10685 21931 10751 21934
rect 11094 21932 11100 21996
rect 11164 21994 11170 21996
rect 15104 21994 15164 22070
rect 18137 22067 18203 22070
rect 22369 22067 22435 22070
rect 24117 22130 24183 22133
rect 24393 22130 24459 22133
rect 24117 22128 24459 22130
rect 24117 22072 24122 22128
rect 24178 22072 24398 22128
rect 24454 22072 24459 22128
rect 24117 22070 24459 22072
rect 24117 22067 24183 22070
rect 24393 22067 24459 22070
rect 11164 21934 15164 21994
rect 11164 21932 11170 21934
rect 15878 21932 15884 21996
rect 15948 21994 15954 21996
rect 16021 21994 16087 21997
rect 15948 21992 16087 21994
rect 15948 21936 16026 21992
rect 16082 21936 16087 21992
rect 15948 21934 16087 21936
rect 15948 21932 15954 21934
rect 16021 21931 16087 21934
rect 19006 21932 19012 21996
rect 19076 21994 19082 21996
rect 21817 21994 21883 21997
rect 22277 21996 22343 21997
rect 23013 21996 23079 21997
rect 22277 21994 22324 21996
rect 19076 21992 21883 21994
rect 19076 21936 21822 21992
rect 21878 21936 21883 21992
rect 19076 21934 21883 21936
rect 22232 21992 22324 21994
rect 22232 21936 22282 21992
rect 22232 21934 22324 21936
rect 19076 21932 19082 21934
rect 21817 21931 21883 21934
rect 22277 21932 22324 21934
rect 22388 21932 22394 21996
rect 23013 21994 23060 21996
rect 22968 21992 23060 21994
rect 22968 21936 23018 21992
rect 22968 21934 23060 21936
rect 23013 21932 23060 21934
rect 23124 21932 23130 21996
rect 22277 21931 22343 21932
rect 23013 21931 23079 21932
rect 0 21858 480 21888
rect 2589 21858 2655 21861
rect 0 21856 2655 21858
rect 0 21800 2594 21856
rect 2650 21800 2655 21856
rect 0 21798 2655 21800
rect 0 21768 480 21798
rect 2589 21795 2655 21798
rect 16297 21858 16363 21861
rect 16430 21858 16436 21860
rect 16297 21856 16436 21858
rect 16297 21800 16302 21856
rect 16358 21800 16436 21856
rect 16297 21798 16436 21800
rect 16297 21795 16363 21798
rect 16430 21796 16436 21798
rect 16500 21796 16506 21860
rect 19057 21858 19123 21861
rect 20294 21858 20300 21860
rect 19057 21856 20300 21858
rect 19057 21800 19062 21856
rect 19118 21800 20300 21856
rect 19057 21798 20300 21800
rect 19057 21795 19123 21798
rect 20294 21796 20300 21798
rect 20364 21796 20370 21860
rect 25405 21858 25471 21861
rect 27520 21858 28000 21888
rect 25405 21856 28000 21858
rect 25405 21800 25410 21856
rect 25466 21800 28000 21856
rect 25405 21798 28000 21800
rect 25405 21795 25471 21798
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 27520 21768 28000 21798
rect 24277 21727 24597 21728
rect 3141 21722 3207 21725
rect 4889 21722 4955 21725
rect 3141 21720 4955 21722
rect 3141 21664 3146 21720
rect 3202 21664 4894 21720
rect 4950 21664 4955 21720
rect 3141 21662 4955 21664
rect 3141 21659 3207 21662
rect 4889 21659 4955 21662
rect 16297 21722 16363 21725
rect 20069 21722 20135 21725
rect 25865 21724 25931 21725
rect 25814 21722 25820 21724
rect 16297 21720 20135 21722
rect 16297 21664 16302 21720
rect 16358 21664 20074 21720
rect 20130 21664 20135 21720
rect 16297 21662 20135 21664
rect 25774 21662 25820 21722
rect 25884 21720 25931 21724
rect 25926 21664 25931 21720
rect 16297 21659 16363 21662
rect 20069 21659 20135 21662
rect 25814 21660 25820 21662
rect 25884 21660 25931 21664
rect 25865 21659 25931 21660
rect 2037 21586 2103 21589
rect 13302 21586 13308 21588
rect 2037 21584 13308 21586
rect 2037 21528 2042 21584
rect 2098 21528 13308 21584
rect 2037 21526 13308 21528
rect 2037 21523 2103 21526
rect 13302 21524 13308 21526
rect 13372 21524 13378 21588
rect 17125 21586 17191 21589
rect 15196 21584 17191 21586
rect 15196 21528 17130 21584
rect 17186 21528 17191 21584
rect 15196 21526 17191 21528
rect 10910 21388 10916 21452
rect 10980 21450 10986 21452
rect 15196 21450 15256 21526
rect 17125 21523 17191 21526
rect 17309 21586 17375 21589
rect 19333 21586 19399 21589
rect 17309 21584 19399 21586
rect 17309 21528 17314 21584
rect 17370 21528 19338 21584
rect 19394 21528 19399 21584
rect 17309 21526 19399 21528
rect 17309 21523 17375 21526
rect 19333 21523 19399 21526
rect 23105 21586 23171 21589
rect 25865 21586 25931 21589
rect 23105 21584 25931 21586
rect 23105 21528 23110 21584
rect 23166 21528 25870 21584
rect 25926 21528 25931 21584
rect 23105 21526 25931 21528
rect 23105 21523 23171 21526
rect 25865 21523 25931 21526
rect 10980 21390 15256 21450
rect 16573 21450 16639 21453
rect 18505 21450 18571 21453
rect 19517 21450 19583 21453
rect 16573 21448 19583 21450
rect 16573 21392 16578 21448
rect 16634 21392 18510 21448
rect 18566 21392 19522 21448
rect 19578 21392 19583 21448
rect 16573 21390 19583 21392
rect 10980 21388 10986 21390
rect 16573 21387 16639 21390
rect 18505 21387 18571 21390
rect 19517 21387 19583 21390
rect 21030 21388 21036 21452
rect 21100 21450 21106 21452
rect 21633 21450 21699 21453
rect 22093 21450 22159 21453
rect 21100 21448 22159 21450
rect 21100 21392 21638 21448
rect 21694 21392 22098 21448
rect 22154 21392 22159 21448
rect 21100 21390 22159 21392
rect 21100 21388 21106 21390
rect 21633 21387 21699 21390
rect 22093 21387 22159 21390
rect 22277 21450 22343 21453
rect 22737 21450 22803 21453
rect 23933 21450 23999 21453
rect 24710 21450 24716 21452
rect 22277 21448 22938 21450
rect 22277 21392 22282 21448
rect 22338 21392 22742 21448
rect 22798 21392 22938 21448
rect 22277 21390 22938 21392
rect 22277 21387 22343 21390
rect 22737 21387 22803 21390
rect 0 21314 480 21344
rect 2681 21314 2747 21317
rect 0 21312 2747 21314
rect 0 21256 2686 21312
rect 2742 21256 2747 21312
rect 0 21254 2747 21256
rect 0 21224 480 21254
rect 2681 21251 2747 21254
rect 5533 21314 5599 21317
rect 8477 21314 8543 21317
rect 5533 21312 8543 21314
rect 5533 21256 5538 21312
rect 5594 21256 8482 21312
rect 8538 21256 8543 21312
rect 5533 21254 8543 21256
rect 5533 21251 5599 21254
rect 8477 21251 8543 21254
rect 16389 21314 16455 21317
rect 18137 21314 18203 21317
rect 16389 21312 18203 21314
rect 16389 21256 16394 21312
rect 16450 21256 18142 21312
rect 18198 21256 18203 21312
rect 16389 21254 18203 21256
rect 22878 21314 22938 21390
rect 23933 21448 24716 21450
rect 23933 21392 23938 21448
rect 23994 21392 24716 21448
rect 23933 21390 24716 21392
rect 23933 21387 23999 21390
rect 24710 21388 24716 21390
rect 24780 21388 24786 21452
rect 25037 21316 25103 21317
rect 24710 21314 24716 21316
rect 22878 21254 24716 21314
rect 16389 21251 16455 21254
rect 18137 21251 18203 21254
rect 24710 21252 24716 21254
rect 24780 21252 24786 21316
rect 25037 21314 25084 21316
rect 24992 21312 25084 21314
rect 24992 21256 25042 21312
rect 24992 21254 25084 21256
rect 25037 21252 25084 21254
rect 25148 21252 25154 21316
rect 25589 21314 25655 21317
rect 27520 21314 28000 21344
rect 25589 21312 28000 21314
rect 25589 21256 25594 21312
rect 25650 21256 28000 21312
rect 25589 21254 28000 21256
rect 25037 21251 25103 21252
rect 25589 21251 25655 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 27520 21224 28000 21254
rect 19610 21183 19930 21184
rect 4889 21178 4955 21181
rect 6913 21178 6979 21181
rect 4889 21176 6979 21178
rect 4889 21120 4894 21176
rect 4950 21120 6918 21176
rect 6974 21120 6979 21176
rect 4889 21118 6979 21120
rect 4889 21115 4955 21118
rect 6913 21115 6979 21118
rect 14089 21178 14155 21181
rect 18045 21178 18111 21181
rect 14089 21176 18111 21178
rect 14089 21120 14094 21176
rect 14150 21120 18050 21176
rect 18106 21120 18111 21176
rect 14089 21118 18111 21120
rect 14089 21115 14155 21118
rect 18045 21115 18111 21118
rect 5533 21042 5599 21045
rect 6085 21042 6151 21045
rect 7189 21042 7255 21045
rect 5533 21040 7255 21042
rect 5533 20984 5538 21040
rect 5594 20984 6090 21040
rect 6146 20984 7194 21040
rect 7250 20984 7255 21040
rect 5533 20982 7255 20984
rect 5533 20979 5599 20982
rect 6085 20979 6151 20982
rect 7189 20979 7255 20982
rect 15326 20980 15332 21044
rect 15396 21042 15402 21044
rect 18229 21042 18295 21045
rect 18413 21044 18479 21045
rect 18413 21042 18460 21044
rect 15396 21040 18295 21042
rect 15396 20984 18234 21040
rect 18290 20984 18295 21040
rect 15396 20982 18295 20984
rect 18368 21040 18460 21042
rect 18368 20984 18418 21040
rect 18368 20982 18460 20984
rect 15396 20980 15402 20982
rect 18229 20979 18295 20982
rect 18413 20980 18460 20982
rect 18524 20980 18530 21044
rect 19701 21042 19767 21045
rect 23473 21042 23539 21045
rect 19701 21040 23539 21042
rect 19701 20984 19706 21040
rect 19762 20984 23478 21040
rect 23534 20984 23539 21040
rect 19701 20982 23539 20984
rect 18413 20979 18479 20980
rect 19701 20979 19767 20982
rect 23473 20979 23539 20982
rect 3049 20906 3115 20909
rect 10593 20906 10659 20909
rect 19885 20906 19951 20909
rect 3049 20904 6148 20906
rect 3049 20848 3054 20904
rect 3110 20848 6148 20904
rect 3049 20846 6148 20848
rect 3049 20843 3115 20846
rect 0 20770 480 20800
rect 1945 20770 2011 20773
rect 0 20768 2011 20770
rect 0 20712 1950 20768
rect 2006 20712 2011 20768
rect 0 20710 2011 20712
rect 0 20680 480 20710
rect 1945 20707 2011 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 1853 20634 1919 20637
rect 4981 20634 5047 20637
rect 1853 20632 5047 20634
rect 1853 20576 1858 20632
rect 1914 20576 4986 20632
rect 5042 20576 5047 20632
rect 1853 20574 5047 20576
rect 6088 20634 6148 20846
rect 10593 20904 19810 20906
rect 10593 20848 10598 20904
rect 10654 20848 19810 20904
rect 10593 20846 19810 20848
rect 10593 20843 10659 20846
rect 6821 20770 6887 20773
rect 11513 20770 11579 20773
rect 6821 20768 11579 20770
rect 6821 20712 6826 20768
rect 6882 20712 11518 20768
rect 11574 20712 11579 20768
rect 6821 20710 11579 20712
rect 6821 20707 6887 20710
rect 11513 20707 11579 20710
rect 12801 20770 12867 20773
rect 14406 20770 14412 20772
rect 12801 20768 14412 20770
rect 12801 20712 12806 20768
rect 12862 20712 14412 20768
rect 12801 20710 14412 20712
rect 12801 20707 12867 20710
rect 14406 20708 14412 20710
rect 14476 20708 14482 20772
rect 16389 20770 16455 20773
rect 18413 20770 18479 20773
rect 16389 20768 18479 20770
rect 16389 20712 16394 20768
rect 16450 20712 18418 20768
rect 18474 20712 18479 20768
rect 16389 20710 18479 20712
rect 19750 20770 19810 20846
rect 19885 20904 24962 20906
rect 19885 20848 19890 20904
rect 19946 20848 24962 20904
rect 19885 20846 24962 20848
rect 19885 20843 19951 20846
rect 20989 20770 21055 20773
rect 22277 20772 22343 20773
rect 22277 20770 22324 20772
rect 19750 20768 21055 20770
rect 19750 20712 20994 20768
rect 21050 20712 21055 20768
rect 19750 20710 21055 20712
rect 22232 20768 22324 20770
rect 22232 20712 22282 20768
rect 22232 20710 22324 20712
rect 16389 20707 16455 20710
rect 18413 20707 18479 20710
rect 20989 20707 21055 20710
rect 22277 20708 22324 20710
rect 22388 20708 22394 20772
rect 24902 20770 24962 20846
rect 27520 20770 28000 20800
rect 24902 20710 28000 20770
rect 22277 20707 22343 20708
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 27520 20680 28000 20710
rect 24277 20639 24597 20640
rect 8109 20634 8175 20637
rect 6088 20632 8175 20634
rect 6088 20576 8114 20632
rect 8170 20576 8175 20632
rect 6088 20574 8175 20576
rect 1853 20571 1919 20574
rect 4981 20571 5047 20574
rect 8109 20571 8175 20574
rect 12341 20634 12407 20637
rect 14181 20634 14247 20637
rect 12341 20632 14247 20634
rect 12341 20576 12346 20632
rect 12402 20576 14186 20632
rect 14242 20576 14247 20632
rect 12341 20574 14247 20576
rect 12341 20571 12407 20574
rect 14181 20571 14247 20574
rect 15561 20634 15627 20637
rect 15837 20634 15903 20637
rect 15561 20632 15903 20634
rect 15561 20576 15566 20632
rect 15622 20576 15842 20632
rect 15898 20576 15903 20632
rect 15561 20574 15903 20576
rect 15561 20571 15627 20574
rect 15837 20571 15903 20574
rect 17861 20634 17927 20637
rect 21633 20634 21699 20637
rect 17861 20632 21699 20634
rect 17861 20576 17866 20632
rect 17922 20576 21638 20632
rect 21694 20576 21699 20632
rect 17861 20574 21699 20576
rect 17861 20571 17927 20574
rect 21633 20571 21699 20574
rect 2037 20498 2103 20501
rect 9305 20498 9371 20501
rect 2037 20496 9371 20498
rect 2037 20440 2042 20496
rect 2098 20440 9310 20496
rect 9366 20440 9371 20496
rect 2037 20438 9371 20440
rect 2037 20435 2103 20438
rect 9305 20435 9371 20438
rect 9673 20498 9739 20501
rect 10777 20498 10843 20501
rect 9673 20496 10843 20498
rect 9673 20440 9678 20496
rect 9734 20440 10782 20496
rect 10838 20440 10843 20496
rect 9673 20438 10843 20440
rect 9673 20435 9739 20438
rect 10777 20435 10843 20438
rect 11697 20498 11763 20501
rect 11830 20498 11836 20500
rect 11697 20496 11836 20498
rect 11697 20440 11702 20496
rect 11758 20440 11836 20496
rect 11697 20438 11836 20440
rect 11697 20435 11763 20438
rect 11830 20436 11836 20438
rect 11900 20498 11906 20500
rect 15101 20498 15167 20501
rect 17033 20498 17099 20501
rect 17861 20498 17927 20501
rect 11900 20438 15026 20498
rect 11900 20436 11906 20438
rect 3141 20362 3207 20365
rect 8937 20362 9003 20365
rect 9489 20362 9555 20365
rect 12433 20362 12499 20365
rect 3141 20360 8770 20362
rect 3141 20304 3146 20360
rect 3202 20304 8770 20360
rect 3141 20302 8770 20304
rect 3141 20299 3207 20302
rect 2405 20226 2471 20229
rect 4245 20226 4311 20229
rect 7189 20226 7255 20229
rect 2405 20224 4170 20226
rect 2405 20168 2410 20224
rect 2466 20168 4170 20224
rect 2405 20166 4170 20168
rect 2405 20163 2471 20166
rect 0 20090 480 20120
rect 3785 20090 3851 20093
rect 0 20088 3851 20090
rect 0 20032 3790 20088
rect 3846 20032 3851 20088
rect 0 20030 3851 20032
rect 4110 20090 4170 20166
rect 4245 20224 7255 20226
rect 4245 20168 4250 20224
rect 4306 20168 7194 20224
rect 7250 20168 7255 20224
rect 4245 20166 7255 20168
rect 4245 20163 4311 20166
rect 7189 20163 7255 20166
rect 8569 20090 8635 20093
rect 4110 20088 8635 20090
rect 4110 20032 8574 20088
rect 8630 20032 8635 20088
rect 4110 20030 8635 20032
rect 8710 20090 8770 20302
rect 8937 20360 12499 20362
rect 8937 20304 8942 20360
rect 8998 20304 9494 20360
rect 9550 20304 12438 20360
rect 12494 20304 12499 20360
rect 8937 20302 12499 20304
rect 8937 20299 9003 20302
rect 9489 20299 9555 20302
rect 12433 20299 12499 20302
rect 13302 20300 13308 20364
rect 13372 20362 13378 20364
rect 14825 20362 14891 20365
rect 13372 20360 14891 20362
rect 13372 20304 14830 20360
rect 14886 20304 14891 20360
rect 13372 20302 14891 20304
rect 14966 20362 15026 20438
rect 15101 20496 17927 20498
rect 15101 20440 15106 20496
rect 15162 20440 17038 20496
rect 17094 20440 17866 20496
rect 17922 20440 17927 20496
rect 15101 20438 17927 20440
rect 15101 20435 15167 20438
rect 17033 20435 17099 20438
rect 17861 20435 17927 20438
rect 18873 20498 18939 20501
rect 20713 20498 20779 20501
rect 18873 20496 20779 20498
rect 18873 20440 18878 20496
rect 18934 20440 20718 20496
rect 20774 20440 20779 20496
rect 18873 20438 20779 20440
rect 18873 20435 18939 20438
rect 20713 20435 20779 20438
rect 20069 20362 20135 20365
rect 14966 20360 20135 20362
rect 14966 20304 20074 20360
rect 20130 20304 20135 20360
rect 14966 20302 20135 20304
rect 13372 20300 13378 20302
rect 14825 20299 14891 20302
rect 20069 20299 20135 20302
rect 23381 20362 23447 20365
rect 23790 20362 23796 20364
rect 23381 20360 23796 20362
rect 23381 20304 23386 20360
rect 23442 20304 23796 20360
rect 23381 20302 23796 20304
rect 23381 20299 23447 20302
rect 23790 20300 23796 20302
rect 23860 20300 23866 20364
rect 9581 20228 9647 20229
rect 9581 20226 9628 20228
rect 9536 20224 9628 20226
rect 9536 20168 9586 20224
rect 9536 20166 9628 20168
rect 9581 20164 9628 20166
rect 9692 20164 9698 20228
rect 11881 20226 11947 20229
rect 18137 20226 18203 20229
rect 11881 20224 18203 20226
rect 11881 20168 11886 20224
rect 11942 20168 18142 20224
rect 18198 20168 18203 20224
rect 11881 20166 18203 20168
rect 9581 20163 9647 20164
rect 11881 20163 11947 20166
rect 18137 20163 18203 20166
rect 20713 20226 20779 20229
rect 25221 20226 25287 20229
rect 20713 20224 25287 20226
rect 20713 20168 20718 20224
rect 20774 20168 25226 20224
rect 25282 20168 25287 20224
rect 20713 20166 25287 20168
rect 20713 20163 20779 20166
rect 25221 20163 25287 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 9990 20090 9996 20092
rect 8710 20030 9996 20090
rect 0 20000 480 20030
rect 3785 20027 3851 20030
rect 8569 20027 8635 20030
rect 9990 20028 9996 20030
rect 10060 20028 10066 20092
rect 11329 20090 11395 20093
rect 11462 20090 11468 20092
rect 11329 20088 11468 20090
rect 11329 20032 11334 20088
rect 11390 20032 11468 20088
rect 11329 20030 11468 20032
rect 11329 20027 11395 20030
rect 11462 20028 11468 20030
rect 11532 20028 11538 20092
rect 12249 20090 12315 20093
rect 12801 20090 12867 20093
rect 12249 20088 12867 20090
rect 12249 20032 12254 20088
rect 12310 20032 12806 20088
rect 12862 20032 12867 20088
rect 12249 20030 12867 20032
rect 12249 20027 12315 20030
rect 12801 20027 12867 20030
rect 14406 20028 14412 20092
rect 14476 20090 14482 20092
rect 14476 20030 19442 20090
rect 14476 20028 14482 20030
rect 5257 19954 5323 19957
rect 11329 19954 11395 19957
rect 5257 19952 11395 19954
rect 5257 19896 5262 19952
rect 5318 19896 11334 19952
rect 11390 19896 11395 19952
rect 5257 19894 11395 19896
rect 5257 19891 5323 19894
rect 11329 19891 11395 19894
rect 11513 19954 11579 19957
rect 14641 19954 14707 19957
rect 11513 19952 14707 19954
rect 11513 19896 11518 19952
rect 11574 19896 14646 19952
rect 14702 19896 14707 19952
rect 11513 19894 14707 19896
rect 11513 19891 11579 19894
rect 14641 19891 14707 19894
rect 14825 19954 14891 19957
rect 17534 19954 17540 19956
rect 14825 19952 17540 19954
rect 14825 19896 14830 19952
rect 14886 19896 17540 19952
rect 14825 19894 17540 19896
rect 14825 19891 14891 19894
rect 17534 19892 17540 19894
rect 17604 19892 17610 19956
rect 19382 19954 19442 20030
rect 20662 20028 20668 20092
rect 20732 20090 20738 20092
rect 21766 20090 21772 20092
rect 20732 20030 21772 20090
rect 20732 20028 20738 20030
rect 21766 20028 21772 20030
rect 21836 20028 21842 20092
rect 23105 20090 23171 20093
rect 23422 20090 23428 20092
rect 23105 20088 23428 20090
rect 23105 20032 23110 20088
rect 23166 20032 23428 20088
rect 23105 20030 23428 20032
rect 23105 20027 23171 20030
rect 23422 20028 23428 20030
rect 23492 20028 23498 20092
rect 27520 20090 28000 20120
rect 23568 20030 28000 20090
rect 19609 19954 19675 19957
rect 20437 19956 20503 19957
rect 20805 19956 20871 19957
rect 20437 19954 20484 19956
rect 19382 19952 19675 19954
rect 19382 19896 19614 19952
rect 19670 19896 19675 19952
rect 19382 19894 19675 19896
rect 20392 19952 20484 19954
rect 20392 19896 20442 19952
rect 20392 19894 20484 19896
rect 19609 19891 19675 19894
rect 20437 19892 20484 19894
rect 20548 19892 20554 19956
rect 20805 19954 20852 19956
rect 20760 19952 20852 19954
rect 20760 19896 20810 19952
rect 20760 19894 20852 19896
rect 20805 19892 20852 19894
rect 20916 19892 20922 19956
rect 23054 19892 23060 19956
rect 23124 19954 23130 19956
rect 23568 19954 23628 20030
rect 27520 20000 28000 20030
rect 23124 19894 23628 19954
rect 23798 19894 26434 19954
rect 23124 19892 23130 19894
rect 20437 19891 20503 19892
rect 20805 19891 20871 19892
rect 2313 19818 2379 19821
rect 5533 19818 5599 19821
rect 2313 19816 5599 19818
rect 2313 19760 2318 19816
rect 2374 19760 5538 19816
rect 5594 19760 5599 19816
rect 2313 19758 5599 19760
rect 2313 19755 2379 19758
rect 5533 19755 5599 19758
rect 5717 19818 5783 19821
rect 8293 19818 8359 19821
rect 10961 19820 11027 19821
rect 5717 19816 8359 19818
rect 5717 19760 5722 19816
rect 5778 19760 8298 19816
rect 8354 19760 8359 19816
rect 5717 19758 8359 19760
rect 5717 19755 5783 19758
rect 8293 19755 8359 19758
rect 10910 19756 10916 19820
rect 10980 19818 11027 19820
rect 11605 19818 11671 19821
rect 11881 19818 11947 19821
rect 10980 19816 11072 19818
rect 11022 19760 11072 19816
rect 10980 19758 11072 19760
rect 11605 19816 11947 19818
rect 11605 19760 11610 19816
rect 11666 19760 11886 19816
rect 11942 19760 11947 19816
rect 11605 19758 11947 19760
rect 10980 19756 11027 19758
rect 10961 19755 11027 19756
rect 11605 19755 11671 19758
rect 11881 19755 11947 19758
rect 12617 19818 12683 19821
rect 16062 19818 16068 19820
rect 12617 19816 16068 19818
rect 12617 19760 12622 19816
rect 12678 19760 16068 19816
rect 12617 19758 16068 19760
rect 12617 19755 12683 19758
rect 16062 19756 16068 19758
rect 16132 19756 16138 19820
rect 17861 19818 17927 19821
rect 18689 19818 18755 19821
rect 20529 19818 20595 19821
rect 23798 19818 23858 19894
rect 17861 19816 20595 19818
rect 17861 19760 17866 19816
rect 17922 19760 18694 19816
rect 18750 19760 20534 19816
rect 20590 19760 20595 19816
rect 17861 19758 20595 19760
rect 17861 19755 17927 19758
rect 18689 19755 18755 19758
rect 20529 19755 20595 19758
rect 21038 19758 23858 19818
rect 24485 19818 24551 19821
rect 26233 19818 26299 19821
rect 24485 19816 26299 19818
rect 24485 19760 24490 19816
rect 24546 19760 26238 19816
rect 26294 19760 26299 19816
rect 24485 19758 26299 19760
rect 9121 19682 9187 19685
rect 11053 19682 11119 19685
rect 9121 19680 11119 19682
rect 9121 19624 9126 19680
rect 9182 19624 11058 19680
rect 11114 19624 11119 19680
rect 9121 19622 11119 19624
rect 9121 19619 9187 19622
rect 11053 19619 11119 19622
rect 17902 19620 17908 19684
rect 17972 19682 17978 19684
rect 18229 19682 18295 19685
rect 20662 19682 20668 19684
rect 17972 19680 20668 19682
rect 17972 19624 18234 19680
rect 18290 19624 20668 19680
rect 17972 19622 20668 19624
rect 17972 19620 17978 19622
rect 18229 19619 18295 19622
rect 20662 19620 20668 19622
rect 20732 19620 20738 19684
rect 5610 19616 5930 19617
rect 0 19546 480 19576
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 2773 19546 2839 19549
rect 0 19544 2839 19546
rect 0 19488 2778 19544
rect 2834 19488 2839 19544
rect 0 19486 2839 19488
rect 0 19456 480 19486
rect 2773 19483 2839 19486
rect 9489 19546 9555 19549
rect 12801 19546 12867 19549
rect 21038 19546 21098 19758
rect 24485 19755 24551 19758
rect 26233 19755 26299 19758
rect 21173 19682 21239 19685
rect 23473 19682 23539 19685
rect 21173 19680 23539 19682
rect 21173 19624 21178 19680
rect 21234 19624 23478 19680
rect 23534 19624 23539 19680
rect 21173 19622 23539 19624
rect 21173 19619 21239 19622
rect 23473 19619 23539 19622
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 9489 19544 12867 19546
rect 9489 19488 9494 19544
rect 9550 19488 12806 19544
rect 12862 19488 12867 19544
rect 9489 19486 12867 19488
rect 9489 19483 9555 19486
rect 12801 19483 12867 19486
rect 16806 19486 21098 19546
rect 26374 19546 26434 19894
rect 27520 19546 28000 19576
rect 26374 19486 28000 19546
rect 2773 19410 2839 19413
rect 12617 19410 12683 19413
rect 16665 19412 16731 19413
rect 16614 19410 16620 19412
rect 2773 19408 12683 19410
rect 2773 19352 2778 19408
rect 2834 19352 12622 19408
rect 12678 19352 12683 19408
rect 2773 19350 12683 19352
rect 2773 19347 2839 19350
rect 12617 19347 12683 19350
rect 16070 19350 16620 19410
rect 16684 19408 16731 19412
rect 16726 19352 16731 19408
rect 3693 19274 3759 19277
rect 4337 19274 4403 19277
rect 10225 19274 10291 19277
rect 3693 19272 10291 19274
rect 3693 19216 3698 19272
rect 3754 19216 4342 19272
rect 4398 19216 10230 19272
rect 10286 19216 10291 19272
rect 3693 19214 10291 19216
rect 3693 19211 3759 19214
rect 4337 19211 4403 19214
rect 10225 19211 10291 19214
rect 10910 19212 10916 19276
rect 10980 19274 10986 19276
rect 11237 19274 11303 19277
rect 10980 19272 11303 19274
rect 10980 19216 11242 19272
rect 11298 19216 11303 19272
rect 10980 19214 11303 19216
rect 10980 19212 10986 19214
rect 11237 19211 11303 19214
rect 11646 19212 11652 19276
rect 11716 19274 11722 19276
rect 11789 19274 11855 19277
rect 11716 19272 11855 19274
rect 11716 19216 11794 19272
rect 11850 19216 11855 19272
rect 11716 19214 11855 19216
rect 11716 19212 11722 19214
rect 11789 19211 11855 19214
rect 13169 19274 13235 19277
rect 16070 19274 16130 19350
rect 16614 19348 16620 19350
rect 16684 19348 16731 19352
rect 16665 19347 16731 19348
rect 13169 19272 16130 19274
rect 13169 19216 13174 19272
rect 13230 19216 16130 19272
rect 13169 19214 16130 19216
rect 16297 19274 16363 19277
rect 16806 19274 16866 19486
rect 27520 19456 28000 19486
rect 19517 19410 19583 19413
rect 20662 19410 20668 19412
rect 19517 19408 20668 19410
rect 19517 19352 19522 19408
rect 19578 19352 20668 19408
rect 19517 19350 20668 19352
rect 19517 19347 19583 19350
rect 20662 19348 20668 19350
rect 20732 19348 20738 19412
rect 20897 19410 20963 19413
rect 21030 19410 21036 19412
rect 20897 19408 21036 19410
rect 20897 19352 20902 19408
rect 20958 19352 21036 19408
rect 20897 19350 21036 19352
rect 20897 19347 20963 19350
rect 21030 19348 21036 19350
rect 21100 19348 21106 19412
rect 24577 19410 24643 19413
rect 25078 19410 25084 19412
rect 24577 19408 25084 19410
rect 24577 19352 24582 19408
rect 24638 19352 25084 19408
rect 24577 19350 25084 19352
rect 24577 19347 24643 19350
rect 25078 19348 25084 19350
rect 25148 19348 25154 19412
rect 19701 19274 19767 19277
rect 21950 19274 21956 19276
rect 16297 19272 16866 19274
rect 16297 19216 16302 19272
rect 16358 19216 16866 19272
rect 16297 19214 16866 19216
rect 17864 19272 21956 19274
rect 17864 19216 19706 19272
rect 19762 19216 21956 19272
rect 17864 19214 21956 19216
rect 13169 19211 13235 19214
rect 16297 19211 16363 19214
rect 3785 19138 3851 19141
rect 9857 19138 9923 19141
rect 3785 19136 9923 19138
rect 3785 19080 3790 19136
rect 3846 19080 9862 19136
rect 9918 19080 9923 19136
rect 3785 19078 9923 19080
rect 3785 19075 3851 19078
rect 9857 19075 9923 19078
rect 11237 19138 11303 19141
rect 11973 19138 12039 19141
rect 11237 19136 12039 19138
rect 11237 19080 11242 19136
rect 11298 19080 11978 19136
rect 12034 19080 12039 19136
rect 11237 19078 12039 19080
rect 11237 19075 11303 19078
rect 11973 19075 12039 19078
rect 12709 19138 12775 19141
rect 17677 19138 17743 19141
rect 12709 19136 17743 19138
rect 12709 19080 12714 19136
rect 12770 19080 17682 19136
rect 17738 19080 17743 19136
rect 12709 19078 17743 19080
rect 12709 19075 12775 19078
rect 17677 19075 17743 19078
rect 10277 19072 10597 19073
rect 0 19002 480 19032
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 6729 19002 6795 19005
rect 0 19000 6795 19002
rect 0 18944 6734 19000
rect 6790 18944 6795 19000
rect 0 18942 6795 18944
rect 0 18912 480 18942
rect 6729 18939 6795 18942
rect 7281 19002 7347 19005
rect 8109 19002 8175 19005
rect 9857 19002 9923 19005
rect 7281 19000 9923 19002
rect 7281 18944 7286 19000
rect 7342 18944 8114 19000
rect 8170 18944 9862 19000
rect 9918 18944 9923 19000
rect 7281 18942 9923 18944
rect 7281 18939 7347 18942
rect 8109 18939 8175 18942
rect 9857 18939 9923 18942
rect 10961 19002 11027 19005
rect 12985 19002 13051 19005
rect 10961 19000 13051 19002
rect 10961 18944 10966 19000
rect 11022 18944 12990 19000
rect 13046 18944 13051 19000
rect 10961 18942 13051 18944
rect 10961 18939 11027 18942
rect 12985 18939 13051 18942
rect 14365 19002 14431 19005
rect 17864 19002 17924 19214
rect 19701 19211 19767 19214
rect 21950 19212 21956 19214
rect 22020 19212 22026 19276
rect 22870 19076 22876 19140
rect 22940 19138 22946 19140
rect 23197 19138 23263 19141
rect 22940 19136 23263 19138
rect 22940 19080 23202 19136
rect 23258 19080 23263 19136
rect 22940 19078 23263 19080
rect 22940 19076 22946 19078
rect 23197 19075 23263 19078
rect 24853 19138 24919 19141
rect 25262 19138 25268 19140
rect 24853 19136 25268 19138
rect 24853 19080 24858 19136
rect 24914 19080 25268 19136
rect 24853 19078 25268 19080
rect 24853 19075 24919 19078
rect 25262 19076 25268 19078
rect 25332 19076 25338 19140
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 14365 19000 17924 19002
rect 14365 18944 14370 19000
rect 14426 18944 17924 19000
rect 14365 18942 17924 18944
rect 21909 19002 21975 19005
rect 24485 19002 24551 19005
rect 21909 19000 24551 19002
rect 21909 18944 21914 19000
rect 21970 18944 24490 19000
rect 24546 18944 24551 19000
rect 21909 18942 24551 18944
rect 14365 18939 14431 18942
rect 21909 18939 21975 18942
rect 24485 18939 24551 18942
rect 26417 19002 26483 19005
rect 27520 19002 28000 19032
rect 26417 19000 28000 19002
rect 26417 18944 26422 19000
rect 26478 18944 28000 19000
rect 26417 18942 28000 18944
rect 26417 18939 26483 18942
rect 27520 18912 28000 18942
rect 5533 18866 5599 18869
rect 6310 18866 6316 18868
rect 5533 18864 6316 18866
rect 5533 18808 5538 18864
rect 5594 18808 6316 18864
rect 5533 18806 6316 18808
rect 5533 18803 5599 18806
rect 6310 18804 6316 18806
rect 6380 18804 6386 18868
rect 7005 18866 7071 18869
rect 9581 18866 9647 18869
rect 7005 18864 9647 18866
rect 7005 18808 7010 18864
rect 7066 18808 9586 18864
rect 9642 18808 9647 18864
rect 7005 18806 9647 18808
rect 7005 18803 7071 18806
rect 9581 18803 9647 18806
rect 12157 18866 12223 18869
rect 13445 18866 13511 18869
rect 15694 18866 15700 18868
rect 12157 18864 13511 18866
rect 12157 18808 12162 18864
rect 12218 18808 13450 18864
rect 13506 18808 13511 18864
rect 12157 18806 13511 18808
rect 12157 18803 12223 18806
rect 13445 18803 13511 18806
rect 14644 18806 15700 18866
rect 4981 18730 5047 18733
rect 7557 18730 7623 18733
rect 10961 18732 11027 18733
rect 9806 18730 9812 18732
rect 4981 18728 6148 18730
rect 4981 18672 4986 18728
rect 5042 18672 6148 18728
rect 4981 18670 6148 18672
rect 4981 18667 5047 18670
rect 6088 18594 6148 18670
rect 7557 18728 9812 18730
rect 7557 18672 7562 18728
rect 7618 18672 9812 18728
rect 7557 18670 9812 18672
rect 7557 18667 7623 18670
rect 9806 18668 9812 18670
rect 9876 18668 9882 18732
rect 10910 18730 10916 18732
rect 10870 18670 10916 18730
rect 10980 18728 11027 18732
rect 11022 18672 11027 18728
rect 10910 18668 10916 18670
rect 10980 18668 11027 18672
rect 11646 18668 11652 18732
rect 11716 18730 11722 18732
rect 11789 18730 11855 18733
rect 11716 18728 11855 18730
rect 11716 18672 11794 18728
rect 11850 18672 11855 18728
rect 11716 18670 11855 18672
rect 11716 18668 11722 18670
rect 10961 18667 11027 18668
rect 11789 18667 11855 18670
rect 12525 18730 12591 18733
rect 14644 18730 14704 18806
rect 15694 18804 15700 18806
rect 15764 18804 15770 18868
rect 16481 18866 16547 18869
rect 19425 18866 19491 18869
rect 16481 18864 19491 18866
rect 16481 18808 16486 18864
rect 16542 18808 19430 18864
rect 19486 18808 19491 18864
rect 16481 18806 19491 18808
rect 16481 18803 16547 18806
rect 19425 18803 19491 18806
rect 20437 18866 20503 18869
rect 20437 18864 24962 18866
rect 20437 18808 20442 18864
rect 20498 18808 24962 18864
rect 20437 18806 24962 18808
rect 20437 18803 20503 18806
rect 12525 18728 14704 18730
rect 12525 18672 12530 18728
rect 12586 18672 14704 18728
rect 12525 18670 14704 18672
rect 12525 18667 12591 18670
rect 17166 18668 17172 18732
rect 17236 18730 17242 18732
rect 20713 18730 20779 18733
rect 17236 18728 20779 18730
rect 17236 18672 20718 18728
rect 20774 18672 20779 18728
rect 17236 18670 20779 18672
rect 17236 18668 17242 18670
rect 20713 18667 20779 18670
rect 21357 18730 21423 18733
rect 21357 18728 24042 18730
rect 21357 18672 21362 18728
rect 21418 18672 24042 18728
rect 21357 18670 24042 18672
rect 21357 18667 21423 18670
rect 9029 18594 9095 18597
rect 12157 18594 12223 18597
rect 6088 18592 12223 18594
rect 6088 18536 9034 18592
rect 9090 18536 12162 18592
rect 12218 18536 12223 18592
rect 6088 18534 12223 18536
rect 9029 18531 9095 18534
rect 12157 18531 12223 18534
rect 12709 18594 12775 18597
rect 13721 18594 13787 18597
rect 12709 18592 13787 18594
rect 12709 18536 12714 18592
rect 12770 18536 13726 18592
rect 13782 18536 13787 18592
rect 12709 18534 13787 18536
rect 12709 18531 12775 18534
rect 13721 18531 13787 18534
rect 18597 18594 18663 18597
rect 22369 18594 22435 18597
rect 22921 18594 22987 18597
rect 23289 18596 23355 18597
rect 18597 18592 22987 18594
rect 18597 18536 18602 18592
rect 18658 18536 22374 18592
rect 22430 18536 22926 18592
rect 22982 18536 22987 18592
rect 18597 18534 22987 18536
rect 18597 18531 18663 18534
rect 22369 18531 22435 18534
rect 22921 18531 22987 18534
rect 23238 18532 23244 18596
rect 23308 18594 23355 18596
rect 23308 18592 23400 18594
rect 23350 18536 23400 18592
rect 23308 18534 23400 18536
rect 23308 18532 23355 18534
rect 23289 18531 23355 18532
rect 5610 18528 5930 18529
rect 0 18458 480 18488
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 10317 18458 10383 18461
rect 10910 18458 10916 18460
rect 0 18398 4722 18458
rect 0 18368 480 18398
rect 2865 18322 2931 18325
rect 2998 18322 3004 18324
rect 2865 18320 3004 18322
rect 2865 18264 2870 18320
rect 2926 18264 3004 18320
rect 2865 18262 3004 18264
rect 2865 18259 2931 18262
rect 2998 18260 3004 18262
rect 3068 18260 3074 18324
rect 4662 18322 4722 18398
rect 10317 18456 10916 18458
rect 10317 18400 10322 18456
rect 10378 18400 10916 18456
rect 10317 18398 10916 18400
rect 10317 18395 10383 18398
rect 10910 18396 10916 18398
rect 10980 18396 10986 18460
rect 12382 18458 12388 18460
rect 11056 18398 12388 18458
rect 8477 18322 8543 18325
rect 4662 18320 8543 18322
rect 4662 18264 8482 18320
rect 8538 18264 8543 18320
rect 4662 18262 8543 18264
rect 8477 18259 8543 18262
rect 10726 18260 10732 18324
rect 10796 18288 10802 18324
rect 11056 18288 11116 18398
rect 12382 18396 12388 18398
rect 12452 18458 12458 18460
rect 18965 18458 19031 18461
rect 23749 18458 23815 18461
rect 12452 18398 14106 18458
rect 12452 18396 12458 18398
rect 10796 18260 11116 18288
rect 10734 18228 11116 18260
rect 12341 18320 12407 18325
rect 12341 18264 12346 18320
rect 12402 18264 12407 18320
rect 12341 18259 12407 18264
rect 3049 18186 3115 18189
rect 7925 18186 7991 18189
rect 3049 18184 7991 18186
rect 3049 18128 3054 18184
rect 3110 18128 7930 18184
rect 7986 18128 7991 18184
rect 3049 18126 7991 18128
rect 3049 18123 3115 18126
rect 7925 18123 7991 18126
rect 2037 18052 2103 18053
rect 2037 18048 2084 18052
rect 2148 18050 2154 18052
rect 2589 18050 2655 18053
rect 3550 18050 3556 18052
rect 2037 17992 2042 18048
rect 2037 17988 2084 17992
rect 2148 17990 2194 18050
rect 2589 18048 3556 18050
rect 2589 17992 2594 18048
rect 2650 17992 3556 18048
rect 2589 17990 3556 17992
rect 2148 17988 2154 17990
rect 2037 17987 2103 17988
rect 2589 17987 2655 17990
rect 3550 17988 3556 17990
rect 3620 17988 3626 18052
rect 11053 18050 11119 18053
rect 12344 18050 12404 18259
rect 14046 18186 14106 18398
rect 18965 18456 23815 18458
rect 18965 18400 18970 18456
rect 19026 18400 23754 18456
rect 23810 18400 23815 18456
rect 18965 18398 23815 18400
rect 18965 18395 19031 18398
rect 23749 18395 23815 18398
rect 14181 18322 14247 18325
rect 18505 18322 18571 18325
rect 14181 18320 18571 18322
rect 14181 18264 14186 18320
rect 14242 18264 18510 18320
rect 18566 18264 18571 18320
rect 14181 18262 18571 18264
rect 14181 18259 14247 18262
rect 18505 18259 18571 18262
rect 18689 18322 18755 18325
rect 21357 18322 21423 18325
rect 18689 18320 21423 18322
rect 18689 18264 18694 18320
rect 18750 18264 21362 18320
rect 21418 18264 21423 18320
rect 18689 18262 21423 18264
rect 18689 18259 18755 18262
rect 21357 18259 21423 18262
rect 21909 18322 21975 18325
rect 23289 18322 23355 18325
rect 21909 18320 23355 18322
rect 21909 18264 21914 18320
rect 21970 18264 23294 18320
rect 23350 18264 23355 18320
rect 21909 18262 23355 18264
rect 23982 18322 24042 18670
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 24902 18458 24962 18806
rect 27520 18458 28000 18488
rect 24902 18398 28000 18458
rect 27520 18368 28000 18398
rect 26325 18322 26391 18325
rect 23982 18320 26391 18322
rect 23982 18264 26330 18320
rect 26386 18264 26391 18320
rect 23982 18262 26391 18264
rect 21909 18259 21975 18262
rect 23289 18259 23355 18262
rect 26325 18259 26391 18262
rect 16297 18186 16363 18189
rect 16573 18186 16639 18189
rect 14046 18184 16639 18186
rect 14046 18128 16302 18184
rect 16358 18128 16578 18184
rect 16634 18128 16639 18184
rect 14046 18126 16639 18128
rect 16297 18123 16363 18126
rect 16573 18123 16639 18126
rect 17861 18186 17927 18189
rect 20713 18186 20779 18189
rect 17861 18184 20779 18186
rect 17861 18128 17866 18184
rect 17922 18128 20718 18184
rect 20774 18128 20779 18184
rect 17861 18126 20779 18128
rect 17861 18123 17927 18126
rect 20713 18123 20779 18126
rect 21909 18186 21975 18189
rect 25221 18186 25287 18189
rect 21909 18184 25287 18186
rect 21909 18128 21914 18184
rect 21970 18128 25226 18184
rect 25282 18128 25287 18184
rect 21909 18126 25287 18128
rect 21909 18123 21975 18126
rect 25221 18123 25287 18126
rect 19057 18050 19123 18053
rect 11053 18048 11162 18050
rect 11053 17992 11058 18048
rect 11114 17992 11162 18048
rect 11053 17987 11162 17992
rect 12344 18048 19123 18050
rect 12344 17992 19062 18048
rect 19118 17992 19123 18048
rect 12344 17990 19123 17992
rect 19057 17987 19123 17990
rect 20713 18050 20779 18053
rect 21173 18052 21239 18053
rect 20846 18050 20852 18052
rect 20713 18048 20852 18050
rect 20713 17992 20718 18048
rect 20774 17992 20852 18048
rect 20713 17990 20852 17992
rect 20713 17987 20779 17990
rect 20846 17988 20852 17990
rect 20916 17988 20922 18052
rect 21173 18048 21220 18052
rect 21284 18050 21290 18052
rect 21817 18050 21883 18053
rect 23933 18050 23999 18053
rect 21173 17992 21178 18048
rect 21173 17988 21220 17992
rect 21284 17990 21330 18050
rect 21817 18048 23999 18050
rect 21817 17992 21822 18048
rect 21878 17992 23938 18048
rect 23994 17992 23999 18048
rect 21817 17990 23999 17992
rect 21284 17988 21290 17990
rect 21173 17987 21239 17988
rect 21817 17987 21883 17990
rect 23933 17987 23999 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 11102 17917 11162 17987
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 2405 17914 2471 17917
rect 5533 17914 5599 17917
rect 8845 17914 8911 17917
rect 2405 17912 5458 17914
rect 2405 17856 2410 17912
rect 2466 17856 5458 17912
rect 2405 17854 5458 17856
rect 2405 17851 2471 17854
rect 0 17778 480 17808
rect 3693 17778 3759 17781
rect 0 17776 3759 17778
rect 0 17720 3698 17776
rect 3754 17720 3759 17776
rect 0 17718 3759 17720
rect 5398 17778 5458 17854
rect 5533 17912 8911 17914
rect 5533 17856 5538 17912
rect 5594 17856 8850 17912
rect 8906 17856 8911 17912
rect 5533 17854 8911 17856
rect 5533 17851 5599 17854
rect 8845 17851 8911 17854
rect 11053 17912 11162 17917
rect 11053 17856 11058 17912
rect 11114 17856 11162 17912
rect 11053 17854 11162 17856
rect 11697 17914 11763 17917
rect 12157 17914 12223 17917
rect 11697 17912 12223 17914
rect 11697 17856 11702 17912
rect 11758 17856 12162 17912
rect 12218 17856 12223 17912
rect 11697 17854 12223 17856
rect 11053 17851 11119 17854
rect 11697 17851 11763 17854
rect 12157 17851 12223 17854
rect 12750 17852 12756 17916
rect 12820 17914 12826 17916
rect 13721 17914 13787 17917
rect 12820 17912 13787 17914
rect 12820 17856 13726 17912
rect 13782 17856 13787 17912
rect 12820 17854 13787 17856
rect 12820 17852 12826 17854
rect 13721 17851 13787 17854
rect 15101 17914 15167 17917
rect 19425 17914 19491 17917
rect 15101 17912 19491 17914
rect 15101 17856 15106 17912
rect 15162 17856 19430 17912
rect 19486 17856 19491 17912
rect 15101 17854 19491 17856
rect 15101 17851 15167 17854
rect 19425 17851 19491 17854
rect 20110 17852 20116 17916
rect 20180 17914 20186 17916
rect 21817 17914 21883 17917
rect 20180 17912 21883 17914
rect 20180 17856 21822 17912
rect 21878 17856 21883 17912
rect 20180 17854 21883 17856
rect 20180 17852 20186 17854
rect 21817 17851 21883 17854
rect 24025 17914 24091 17917
rect 25630 17914 25636 17916
rect 24025 17912 25636 17914
rect 24025 17856 24030 17912
rect 24086 17856 25636 17912
rect 24025 17854 25636 17856
rect 24025 17851 24091 17854
rect 25630 17852 25636 17854
rect 25700 17852 25706 17916
rect 5625 17778 5691 17781
rect 8385 17778 8451 17781
rect 5398 17776 8451 17778
rect 5398 17720 5630 17776
rect 5686 17720 8390 17776
rect 8446 17720 8451 17776
rect 5398 17718 8451 17720
rect 0 17688 480 17718
rect 3693 17715 3759 17718
rect 5625 17715 5691 17718
rect 8385 17715 8451 17718
rect 9673 17778 9739 17781
rect 17677 17778 17743 17781
rect 20069 17778 20135 17781
rect 9673 17776 17234 17778
rect 9673 17720 9678 17776
rect 9734 17720 17234 17776
rect 9673 17718 17234 17720
rect 9673 17715 9739 17718
rect 6637 17642 6703 17645
rect 9397 17642 9463 17645
rect 6637 17640 9463 17642
rect 6637 17584 6642 17640
rect 6698 17584 9402 17640
rect 9458 17584 9463 17640
rect 6637 17582 9463 17584
rect 6637 17579 6703 17582
rect 9397 17579 9463 17582
rect 9765 17642 9831 17645
rect 12617 17642 12683 17645
rect 9765 17640 12683 17642
rect 9765 17584 9770 17640
rect 9826 17584 12622 17640
rect 12678 17584 12683 17640
rect 9765 17582 12683 17584
rect 9765 17579 9831 17582
rect 12617 17579 12683 17582
rect 14590 17580 14596 17644
rect 14660 17642 14666 17644
rect 14825 17642 14891 17645
rect 14660 17640 14891 17642
rect 14660 17584 14830 17640
rect 14886 17584 14891 17640
rect 14660 17582 14891 17584
rect 14660 17580 14666 17582
rect 14825 17579 14891 17582
rect 15694 17580 15700 17644
rect 15764 17642 15770 17644
rect 15837 17642 15903 17645
rect 15764 17640 15903 17642
rect 15764 17584 15842 17640
rect 15898 17584 15903 17640
rect 15764 17582 15903 17584
rect 15764 17580 15770 17582
rect 15837 17579 15903 17582
rect 6453 17506 6519 17509
rect 11697 17506 11763 17509
rect 6453 17504 11763 17506
rect 6453 17448 6458 17504
rect 6514 17448 11702 17504
rect 11758 17448 11763 17504
rect 6453 17446 11763 17448
rect 6453 17443 6519 17446
rect 11697 17443 11763 17446
rect 13670 17444 13676 17508
rect 13740 17506 13746 17508
rect 14089 17506 14155 17509
rect 13740 17504 14155 17506
rect 13740 17448 14094 17504
rect 14150 17448 14155 17504
rect 13740 17446 14155 17448
rect 13740 17444 13746 17446
rect 14089 17443 14155 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 5165 17372 5231 17373
rect 5165 17370 5212 17372
rect 5120 17368 5212 17370
rect 5120 17312 5170 17368
rect 5120 17310 5212 17312
rect 5165 17308 5212 17310
rect 5276 17308 5282 17372
rect 17174 17370 17234 17718
rect 17677 17776 20135 17778
rect 17677 17720 17682 17776
rect 17738 17720 20074 17776
rect 20130 17720 20135 17776
rect 17677 17718 20135 17720
rect 17677 17715 17743 17718
rect 20069 17715 20135 17718
rect 20345 17778 20411 17781
rect 22001 17778 22067 17781
rect 20345 17776 22067 17778
rect 20345 17720 20350 17776
rect 20406 17720 22006 17776
rect 22062 17720 22067 17776
rect 20345 17718 22067 17720
rect 20345 17715 20411 17718
rect 22001 17715 22067 17718
rect 25078 17716 25084 17780
rect 25148 17778 25154 17780
rect 27520 17778 28000 17808
rect 25148 17718 28000 17778
rect 25148 17716 25154 17718
rect 27520 17688 28000 17718
rect 18689 17642 18755 17645
rect 21541 17642 21607 17645
rect 18689 17640 21607 17642
rect 18689 17584 18694 17640
rect 18750 17584 21546 17640
rect 21602 17584 21607 17640
rect 18689 17582 21607 17584
rect 18689 17579 18755 17582
rect 21541 17579 21607 17582
rect 23197 17642 23263 17645
rect 26325 17642 26391 17645
rect 23197 17640 26391 17642
rect 23197 17584 23202 17640
rect 23258 17584 26330 17640
rect 26386 17584 26391 17640
rect 23197 17582 26391 17584
rect 23197 17579 23263 17582
rect 26325 17579 26391 17582
rect 18045 17506 18111 17509
rect 22369 17506 22435 17509
rect 18045 17504 22435 17506
rect 18045 17448 18050 17504
rect 18106 17448 22374 17504
rect 22430 17448 22435 17504
rect 18045 17446 22435 17448
rect 18045 17443 18111 17446
rect 22369 17443 22435 17446
rect 24761 17506 24827 17509
rect 25262 17506 25268 17508
rect 24761 17504 25268 17506
rect 24761 17448 24766 17504
rect 24822 17448 25268 17504
rect 24761 17446 25268 17448
rect 24761 17443 24827 17446
rect 25262 17444 25268 17446
rect 25332 17444 25338 17508
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 23749 17370 23815 17373
rect 17174 17368 23815 17370
rect 17174 17312 23754 17368
rect 23810 17312 23815 17368
rect 17174 17310 23815 17312
rect 5165 17307 5231 17308
rect 23749 17307 23815 17310
rect 25405 17372 25471 17373
rect 25405 17368 25452 17372
rect 25516 17370 25522 17372
rect 25405 17312 25410 17368
rect 25405 17308 25452 17312
rect 25516 17310 25562 17370
rect 25516 17308 25522 17310
rect 25405 17307 25471 17308
rect 0 17234 480 17264
rect 1025 17234 1091 17237
rect 0 17232 1091 17234
rect 0 17176 1030 17232
rect 1086 17176 1091 17232
rect 0 17174 1091 17176
rect 0 17144 480 17174
rect 1025 17171 1091 17174
rect 4981 17234 5047 17237
rect 9029 17234 9095 17237
rect 4981 17232 9095 17234
rect 4981 17176 4986 17232
rect 5042 17176 9034 17232
rect 9090 17176 9095 17232
rect 4981 17174 9095 17176
rect 4981 17171 5047 17174
rect 9029 17171 9095 17174
rect 13629 17234 13695 17237
rect 14181 17234 14247 17237
rect 13629 17232 14247 17234
rect 13629 17176 13634 17232
rect 13690 17176 14186 17232
rect 14242 17176 14247 17232
rect 13629 17174 14247 17176
rect 13629 17171 13695 17174
rect 14181 17171 14247 17174
rect 15878 17172 15884 17236
rect 15948 17234 15954 17236
rect 16941 17234 17007 17237
rect 17585 17236 17651 17237
rect 17534 17234 17540 17236
rect 15948 17232 17007 17234
rect 15948 17176 16946 17232
rect 17002 17176 17007 17232
rect 15948 17174 17007 17176
rect 17494 17174 17540 17234
rect 17604 17232 17651 17236
rect 17646 17176 17651 17232
rect 15948 17172 15954 17174
rect 16941 17171 17007 17174
rect 17534 17172 17540 17174
rect 17604 17172 17651 17176
rect 17585 17171 17651 17172
rect 18045 17234 18111 17237
rect 18505 17234 18571 17237
rect 23105 17234 23171 17237
rect 18045 17232 23171 17234
rect 18045 17176 18050 17232
rect 18106 17176 18510 17232
rect 18566 17176 23110 17232
rect 23166 17176 23171 17232
rect 18045 17174 23171 17176
rect 18045 17171 18111 17174
rect 18505 17171 18571 17174
rect 23105 17171 23171 17174
rect 23289 17234 23355 17237
rect 24853 17234 24919 17237
rect 27520 17234 28000 17264
rect 23289 17232 24919 17234
rect 23289 17176 23294 17232
rect 23350 17176 24858 17232
rect 24914 17176 24919 17232
rect 23289 17174 24919 17176
rect 23289 17171 23355 17174
rect 24853 17171 24919 17174
rect 25638 17174 28000 17234
rect 2497 17098 2563 17101
rect 8109 17098 8175 17101
rect 2497 17096 8175 17098
rect 2497 17040 2502 17096
rect 2558 17040 8114 17096
rect 8170 17040 8175 17096
rect 2497 17038 8175 17040
rect 2497 17035 2563 17038
rect 8109 17035 8175 17038
rect 8937 17098 9003 17101
rect 11462 17098 11468 17100
rect 8937 17096 11468 17098
rect 8937 17040 8942 17096
rect 8998 17040 11468 17096
rect 8937 17038 11468 17040
rect 8937 17035 9003 17038
rect 11462 17036 11468 17038
rect 11532 17098 11538 17100
rect 14457 17098 14523 17101
rect 11532 17096 14523 17098
rect 11532 17040 14462 17096
rect 14518 17040 14523 17096
rect 11532 17038 14523 17040
rect 11532 17036 11538 17038
rect 14457 17035 14523 17038
rect 14641 17098 14707 17101
rect 25405 17098 25471 17101
rect 14641 17096 25471 17098
rect 14641 17040 14646 17096
rect 14702 17040 25410 17096
rect 25466 17040 25471 17096
rect 14641 17038 25471 17040
rect 14641 17035 14707 17038
rect 25405 17035 25471 17038
rect 2957 16962 3023 16965
rect 6269 16962 6335 16965
rect 2957 16960 6335 16962
rect 2957 16904 2962 16960
rect 3018 16904 6274 16960
rect 6330 16904 6335 16960
rect 2957 16902 6335 16904
rect 2957 16899 3023 16902
rect 6269 16899 6335 16902
rect 14273 16962 14339 16965
rect 14590 16962 14596 16964
rect 14273 16960 14596 16962
rect 14273 16904 14278 16960
rect 14334 16904 14596 16960
rect 14273 16902 14596 16904
rect 14273 16899 14339 16902
rect 14590 16900 14596 16902
rect 14660 16900 14666 16964
rect 14733 16962 14799 16965
rect 18505 16962 18571 16965
rect 22737 16964 22803 16965
rect 22686 16962 22692 16964
rect 14733 16960 18571 16962
rect 14733 16904 14738 16960
rect 14794 16904 18510 16960
rect 18566 16904 18571 16960
rect 14733 16902 18571 16904
rect 22646 16902 22692 16962
rect 22756 16960 22803 16964
rect 22798 16904 22803 16960
rect 14733 16899 14799 16902
rect 18505 16899 18571 16902
rect 22686 16900 22692 16902
rect 22756 16900 22803 16904
rect 22737 16899 22803 16900
rect 23105 16962 23171 16965
rect 25638 16962 25698 17174
rect 27520 17144 28000 17174
rect 23105 16960 25698 16962
rect 23105 16904 23110 16960
rect 23166 16904 25698 16960
rect 23105 16902 25698 16904
rect 23105 16899 23171 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 4613 16826 4679 16829
rect 8477 16826 8543 16829
rect 13261 16826 13327 16829
rect 14365 16826 14431 16829
rect 18597 16826 18663 16829
rect 23381 16826 23447 16829
rect 4613 16824 8586 16826
rect 4613 16768 4618 16824
rect 4674 16768 8482 16824
rect 8538 16768 8586 16824
rect 4613 16766 8586 16768
rect 4613 16763 4679 16766
rect 8477 16763 8586 16766
rect 13261 16824 14106 16826
rect 13261 16768 13266 16824
rect 13322 16768 14106 16824
rect 13261 16766 14106 16768
rect 13261 16763 13327 16766
rect 0 16690 480 16720
rect 1393 16690 1459 16693
rect 0 16688 1459 16690
rect 0 16632 1398 16688
rect 1454 16632 1459 16688
rect 0 16630 1459 16632
rect 0 16600 480 16630
rect 1393 16627 1459 16630
rect 1761 16690 1827 16693
rect 6637 16690 6703 16693
rect 1761 16688 6703 16690
rect 1761 16632 1766 16688
rect 1822 16632 6642 16688
rect 6698 16632 6703 16688
rect 1761 16630 6703 16632
rect 1761 16627 1827 16630
rect 6637 16627 6703 16630
rect 7189 16690 7255 16693
rect 8150 16690 8156 16692
rect 7189 16688 8156 16690
rect 7189 16632 7194 16688
rect 7250 16632 8156 16688
rect 7189 16630 8156 16632
rect 7189 16627 7255 16630
rect 8150 16628 8156 16630
rect 8220 16628 8226 16692
rect 8526 16690 8586 16763
rect 13905 16690 13971 16693
rect 8526 16688 13971 16690
rect 8526 16632 13910 16688
rect 13966 16632 13971 16688
rect 8526 16630 13971 16632
rect 13905 16627 13971 16630
rect 4981 16554 5047 16557
rect 9305 16554 9371 16557
rect 11237 16554 11303 16557
rect 4981 16552 6148 16554
rect 4981 16496 4986 16552
rect 5042 16496 6148 16552
rect 4981 16494 6148 16496
rect 4981 16491 5047 16494
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 6088 16282 6148 16494
rect 9305 16552 11303 16554
rect 9305 16496 9310 16552
rect 9366 16496 11242 16552
rect 11298 16496 11303 16552
rect 9305 16494 11303 16496
rect 9305 16491 9371 16494
rect 11237 16491 11303 16494
rect 14046 16554 14106 16766
rect 14365 16824 18663 16826
rect 14365 16768 14370 16824
rect 14426 16768 18602 16824
rect 18658 16768 18663 16824
rect 14365 16766 18663 16768
rect 14365 16763 14431 16766
rect 18597 16763 18663 16766
rect 20072 16824 23447 16826
rect 20072 16768 23386 16824
rect 23442 16768 23447 16824
rect 20072 16766 23447 16768
rect 15193 16690 15259 16693
rect 15326 16690 15332 16692
rect 15193 16688 15332 16690
rect 15193 16632 15198 16688
rect 15254 16632 15332 16688
rect 15193 16630 15332 16632
rect 15193 16627 15259 16630
rect 15326 16628 15332 16630
rect 15396 16628 15402 16692
rect 16389 16690 16455 16693
rect 18137 16690 18203 16693
rect 16389 16688 18203 16690
rect 16389 16632 16394 16688
rect 16450 16632 18142 16688
rect 18198 16632 18203 16688
rect 16389 16630 18203 16632
rect 16389 16627 16455 16630
rect 18137 16627 18203 16630
rect 18873 16690 18939 16693
rect 20072 16690 20132 16766
rect 23381 16763 23447 16766
rect 23606 16764 23612 16828
rect 23676 16764 23682 16828
rect 23790 16764 23796 16828
rect 23860 16764 23866 16828
rect 23614 16693 23674 16764
rect 18873 16688 20132 16690
rect 18873 16632 18878 16688
rect 18934 16632 20132 16688
rect 18873 16630 20132 16632
rect 20529 16690 20595 16693
rect 22686 16690 22692 16692
rect 20529 16688 22692 16690
rect 20529 16632 20534 16688
rect 20590 16632 22692 16688
rect 20529 16630 22692 16632
rect 18873 16627 18939 16630
rect 20529 16627 20595 16630
rect 22686 16628 22692 16630
rect 22756 16628 22762 16692
rect 23614 16688 23723 16693
rect 23614 16632 23662 16688
rect 23718 16632 23723 16688
rect 23614 16630 23723 16632
rect 23657 16627 23723 16630
rect 22502 16554 22508 16556
rect 14046 16494 22508 16554
rect 14046 16418 14106 16494
rect 22502 16492 22508 16494
rect 22572 16492 22578 16556
rect 23422 16492 23428 16556
rect 23492 16554 23498 16556
rect 23565 16554 23631 16557
rect 23492 16552 23631 16554
rect 23492 16496 23570 16552
rect 23626 16496 23631 16552
rect 23492 16494 23631 16496
rect 23798 16554 23858 16764
rect 25313 16690 25379 16693
rect 27520 16690 28000 16720
rect 25313 16688 28000 16690
rect 25313 16632 25318 16688
rect 25374 16632 28000 16688
rect 25313 16630 28000 16632
rect 25313 16627 25379 16630
rect 27520 16600 28000 16630
rect 25773 16554 25839 16557
rect 23798 16552 25839 16554
rect 23798 16496 25778 16552
rect 25834 16496 25839 16552
rect 23798 16494 25839 16496
rect 23492 16492 23498 16494
rect 23565 16491 23631 16494
rect 25773 16491 25839 16494
rect 10366 16358 14106 16418
rect 10366 16282 10426 16358
rect 16430 16356 16436 16420
rect 16500 16418 16506 16420
rect 17953 16418 18019 16421
rect 21582 16418 21588 16420
rect 16500 16416 21588 16418
rect 16500 16360 17958 16416
rect 18014 16360 21588 16416
rect 16500 16358 21588 16360
rect 16500 16356 16506 16358
rect 17953 16355 18019 16358
rect 21582 16356 21588 16358
rect 21652 16356 21658 16420
rect 22921 16418 22987 16421
rect 23381 16418 23447 16421
rect 22921 16416 23447 16418
rect 22921 16360 22926 16416
rect 22982 16360 23386 16416
rect 23442 16360 23447 16416
rect 22921 16358 23447 16360
rect 22921 16355 22987 16358
rect 23381 16355 23447 16358
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 6088 16222 10426 16282
rect 10501 16282 10567 16285
rect 12525 16282 12591 16285
rect 10501 16280 12591 16282
rect 10501 16224 10506 16280
rect 10562 16224 12530 16280
rect 12586 16224 12591 16280
rect 10501 16222 12591 16224
rect 10501 16219 10567 16222
rect 12525 16219 12591 16222
rect 12750 16220 12756 16284
rect 12820 16282 12826 16284
rect 13629 16282 13695 16285
rect 12820 16280 13695 16282
rect 12820 16224 13634 16280
rect 13690 16224 13695 16280
rect 12820 16222 13695 16224
rect 12820 16220 12826 16222
rect 13629 16219 13695 16222
rect 14038 16220 14044 16284
rect 14108 16282 14114 16284
rect 14733 16282 14799 16285
rect 14108 16280 14799 16282
rect 14108 16224 14738 16280
rect 14794 16224 14799 16280
rect 14108 16222 14799 16224
rect 14108 16220 14114 16222
rect 14733 16219 14799 16222
rect 15929 16282 15995 16285
rect 16246 16282 16252 16284
rect 15929 16280 16252 16282
rect 15929 16224 15934 16280
rect 15990 16224 16252 16280
rect 15929 16222 16252 16224
rect 15929 16219 15995 16222
rect 16246 16220 16252 16222
rect 16316 16220 16322 16284
rect 16757 16282 16823 16285
rect 22921 16282 22987 16285
rect 16757 16280 22987 16282
rect 16757 16224 16762 16280
rect 16818 16224 22926 16280
rect 22982 16224 22987 16280
rect 16757 16222 22987 16224
rect 16757 16219 16823 16222
rect 22921 16219 22987 16222
rect 3693 16146 3759 16149
rect 9673 16146 9739 16149
rect 3693 16144 9739 16146
rect 3693 16088 3698 16144
rect 3754 16088 9678 16144
rect 9734 16088 9739 16144
rect 3693 16086 9739 16088
rect 3693 16083 3759 16086
rect 9673 16083 9739 16086
rect 9806 16084 9812 16148
rect 9876 16146 9882 16148
rect 12382 16146 12388 16148
rect 9876 16086 12388 16146
rect 9876 16084 9882 16086
rect 12382 16084 12388 16086
rect 12452 16084 12458 16148
rect 14365 16146 14431 16149
rect 19425 16146 19491 16149
rect 14365 16144 19491 16146
rect 14365 16088 14370 16144
rect 14426 16088 19430 16144
rect 19486 16088 19491 16144
rect 14365 16086 19491 16088
rect 14365 16083 14431 16086
rect 19425 16083 19491 16086
rect 19609 16146 19675 16149
rect 24853 16146 24919 16149
rect 19609 16144 24919 16146
rect 19609 16088 19614 16144
rect 19670 16088 24858 16144
rect 24914 16088 24919 16144
rect 19609 16086 24919 16088
rect 19609 16083 19675 16086
rect 24853 16083 24919 16086
rect 0 16010 480 16040
rect 8017 16010 8083 16013
rect 0 16008 8083 16010
rect 0 15952 8022 16008
rect 8078 15952 8083 16008
rect 0 15950 8083 15952
rect 0 15920 480 15950
rect 8017 15947 8083 15950
rect 8385 16010 8451 16013
rect 10961 16010 11027 16013
rect 11421 16010 11487 16013
rect 18413 16010 18479 16013
rect 20253 16010 20319 16013
rect 8385 16008 10794 16010
rect 8385 15952 8390 16008
rect 8446 15952 10794 16008
rect 8385 15950 10794 15952
rect 8385 15947 8451 15950
rect 1853 15874 1919 15877
rect 5625 15874 5691 15877
rect 1853 15872 5691 15874
rect 1853 15816 1858 15872
rect 1914 15816 5630 15872
rect 5686 15816 5691 15872
rect 1853 15814 5691 15816
rect 1853 15811 1919 15814
rect 5625 15811 5691 15814
rect 6637 15874 6703 15877
rect 9029 15874 9095 15877
rect 6637 15872 9095 15874
rect 6637 15816 6642 15872
rect 6698 15816 9034 15872
rect 9090 15816 9095 15872
rect 6637 15814 9095 15816
rect 6637 15811 6703 15814
rect 9029 15811 9095 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 3233 15738 3299 15741
rect 9397 15738 9463 15741
rect 3233 15736 9463 15738
rect 3233 15680 3238 15736
rect 3294 15680 9402 15736
rect 9458 15680 9463 15736
rect 3233 15678 9463 15680
rect 10734 15738 10794 15950
rect 10961 16008 18479 16010
rect 10961 15952 10966 16008
rect 11022 15952 11426 16008
rect 11482 15952 18418 16008
rect 18474 15952 18479 16008
rect 10961 15950 18479 15952
rect 10961 15947 11027 15950
rect 11421 15947 11487 15950
rect 18413 15947 18479 15950
rect 18600 16008 20776 16010
rect 18600 15952 20258 16008
rect 20314 15952 20776 16008
rect 18600 15950 20776 15952
rect 10869 15874 10935 15877
rect 11881 15874 11947 15877
rect 15929 15874 15995 15877
rect 10869 15872 15995 15874
rect 10869 15816 10874 15872
rect 10930 15816 11886 15872
rect 11942 15816 15934 15872
rect 15990 15816 15995 15872
rect 10869 15814 15995 15816
rect 10869 15811 10935 15814
rect 11881 15811 11947 15814
rect 15929 15811 15995 15814
rect 11421 15738 11487 15741
rect 10734 15736 11487 15738
rect 10734 15680 11426 15736
rect 11482 15680 11487 15736
rect 10734 15678 11487 15680
rect 3233 15675 3299 15678
rect 9397 15675 9463 15678
rect 11421 15675 11487 15678
rect 11830 15676 11836 15740
rect 11900 15738 11906 15740
rect 12198 15738 12204 15740
rect 11900 15678 12204 15738
rect 11900 15676 11906 15678
rect 12198 15676 12204 15678
rect 12268 15676 12274 15740
rect 12801 15738 12867 15741
rect 15653 15738 15719 15741
rect 17125 15738 17191 15741
rect 18600 15738 18660 15950
rect 20253 15947 20319 15950
rect 20716 15874 20776 15950
rect 20846 15948 20852 16012
rect 20916 16010 20922 16012
rect 20989 16010 21055 16013
rect 20916 16008 21055 16010
rect 20916 15952 20994 16008
rect 21050 15952 21055 16008
rect 20916 15950 21055 15952
rect 20916 15948 20922 15950
rect 20989 15947 21055 15950
rect 21950 15948 21956 16012
rect 22020 16010 22026 16012
rect 22134 16010 22140 16012
rect 22020 15950 22140 16010
rect 22020 15948 22026 15950
rect 22134 15948 22140 15950
rect 22204 15948 22210 16012
rect 27520 16010 28000 16040
rect 22280 15950 28000 16010
rect 22280 15874 22340 15950
rect 27520 15920 28000 15950
rect 20716 15814 22340 15874
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 12801 15736 15719 15738
rect 12801 15680 12806 15736
rect 12862 15680 15658 15736
rect 15714 15680 15719 15736
rect 12801 15678 15719 15680
rect 12801 15675 12867 15678
rect 15653 15675 15719 15678
rect 16070 15736 17191 15738
rect 16070 15680 17130 15736
rect 17186 15680 17191 15736
rect 16070 15678 17191 15680
rect 7649 15602 7715 15605
rect 12709 15602 12775 15605
rect 12985 15602 13051 15605
rect 16070 15602 16130 15678
rect 17125 15675 17191 15678
rect 18094 15678 18660 15738
rect 20621 15738 20687 15741
rect 21633 15738 21699 15741
rect 24025 15738 24091 15741
rect 20621 15736 21282 15738
rect 20621 15680 20626 15736
rect 20682 15680 21282 15736
rect 20621 15678 21282 15680
rect 7649 15600 13051 15602
rect 7649 15544 7654 15600
rect 7710 15544 12714 15600
rect 12770 15544 12990 15600
rect 13046 15544 13051 15600
rect 7649 15542 13051 15544
rect 7649 15539 7715 15542
rect 12709 15539 12775 15542
rect 12985 15539 13051 15542
rect 14598 15542 16130 15602
rect 16205 15602 16271 15605
rect 18094 15602 18154 15678
rect 20621 15675 20687 15678
rect 20069 15602 20135 15605
rect 20621 15602 20687 15605
rect 16205 15600 18154 15602
rect 16205 15544 16210 15600
rect 16266 15544 18154 15600
rect 16205 15542 18154 15544
rect 18232 15600 20687 15602
rect 18232 15544 20074 15600
rect 20130 15544 20626 15600
rect 20682 15544 20687 15600
rect 18232 15542 20687 15544
rect 0 15466 480 15496
rect 13629 15466 13695 15469
rect 0 15464 13695 15466
rect 0 15408 13634 15464
rect 13690 15408 13695 15464
rect 0 15406 13695 15408
rect 0 15376 480 15406
rect 13629 15403 13695 15406
rect 3417 15330 3483 15333
rect 3969 15330 4035 15333
rect 7649 15330 7715 15333
rect 9949 15330 10015 15333
rect 3417 15328 5458 15330
rect 3417 15272 3422 15328
rect 3478 15272 3974 15328
rect 4030 15272 5458 15328
rect 3417 15270 5458 15272
rect 3417 15267 3483 15270
rect 3969 15267 4035 15270
rect 5398 15058 5458 15270
rect 7649 15328 10015 15330
rect 7649 15272 7654 15328
rect 7710 15272 9954 15328
rect 10010 15272 10015 15328
rect 7649 15270 10015 15272
rect 7649 15267 7715 15270
rect 9949 15267 10015 15270
rect 10869 15330 10935 15333
rect 11329 15330 11395 15333
rect 14598 15330 14658 15542
rect 16205 15539 16271 15542
rect 18232 15466 18292 15542
rect 20069 15539 20135 15542
rect 20621 15539 20687 15542
rect 10869 15328 14658 15330
rect 10869 15272 10874 15328
rect 10930 15272 11334 15328
rect 11390 15272 14658 15328
rect 10869 15270 14658 15272
rect 14782 15406 18292 15466
rect 19149 15466 19215 15469
rect 20989 15466 21055 15469
rect 19149 15464 21055 15466
rect 19149 15408 19154 15464
rect 19210 15408 20994 15464
rect 21050 15408 21055 15464
rect 19149 15406 21055 15408
rect 21222 15466 21282 15678
rect 21633 15736 24091 15738
rect 21633 15680 21638 15736
rect 21694 15680 24030 15736
rect 24086 15680 24091 15736
rect 21633 15678 24091 15680
rect 21633 15675 21699 15678
rect 24025 15675 24091 15678
rect 21582 15540 21588 15604
rect 21652 15602 21658 15604
rect 25221 15602 25287 15605
rect 21652 15600 25287 15602
rect 21652 15544 25226 15600
rect 25282 15544 25287 15600
rect 21652 15542 25287 15544
rect 21652 15540 21658 15542
rect 25221 15539 25287 15542
rect 21582 15466 21588 15468
rect 21222 15406 21588 15466
rect 10869 15267 10935 15270
rect 11329 15267 11395 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 9397 15194 9463 15197
rect 11605 15196 11671 15197
rect 9990 15194 9996 15196
rect 9397 15192 9996 15194
rect 9397 15136 9402 15192
rect 9458 15136 9996 15192
rect 9397 15134 9996 15136
rect 9397 15131 9463 15134
rect 9990 15132 9996 15134
rect 10060 15132 10066 15196
rect 11605 15194 11652 15196
rect 11560 15192 11652 15194
rect 11560 15136 11610 15192
rect 11560 15134 11652 15136
rect 11605 15132 11652 15134
rect 11716 15132 11722 15196
rect 14641 15194 14707 15197
rect 14782 15194 14842 15406
rect 19149 15403 19215 15406
rect 20989 15403 21055 15406
rect 21582 15404 21588 15406
rect 21652 15404 21658 15468
rect 24853 15466 24919 15469
rect 27520 15466 28000 15496
rect 24853 15464 28000 15466
rect 24853 15408 24858 15464
rect 24914 15408 28000 15464
rect 24853 15406 28000 15408
rect 24853 15403 24919 15406
rect 27520 15376 28000 15406
rect 18045 15330 18111 15333
rect 21541 15330 21607 15333
rect 18045 15328 21607 15330
rect 18045 15272 18050 15328
rect 18106 15272 21546 15328
rect 21602 15272 21607 15328
rect 18045 15270 21607 15272
rect 18045 15267 18111 15270
rect 21541 15267 21607 15270
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 14641 15192 14842 15194
rect 14641 15136 14646 15192
rect 14702 15136 14842 15192
rect 14641 15134 14842 15136
rect 18229 15194 18295 15197
rect 18454 15194 18460 15196
rect 18229 15192 18460 15194
rect 18229 15136 18234 15192
rect 18290 15136 18460 15192
rect 18229 15134 18460 15136
rect 11605 15131 11671 15132
rect 14641 15131 14707 15134
rect 18229 15131 18295 15134
rect 18454 15132 18460 15134
rect 18524 15132 18530 15196
rect 20989 15194 21055 15197
rect 22461 15194 22527 15197
rect 20989 15192 22527 15194
rect 20989 15136 20994 15192
rect 21050 15136 22466 15192
rect 22522 15136 22527 15192
rect 20989 15134 22527 15136
rect 20989 15131 21055 15134
rect 22461 15131 22527 15134
rect 9806 15058 9812 15060
rect 5398 14998 9812 15058
rect 9806 14996 9812 14998
rect 9876 14996 9882 15060
rect 9990 14996 9996 15060
rect 10060 15058 10066 15060
rect 10409 15058 10475 15061
rect 13486 15058 13492 15060
rect 10060 15056 10475 15058
rect 10060 15000 10414 15056
rect 10470 15000 10475 15056
rect 10060 14998 10475 15000
rect 10060 14996 10066 14998
rect 10409 14995 10475 14998
rect 11792 14998 13492 15058
rect 0 14922 480 14952
rect 3785 14922 3851 14925
rect 0 14920 3851 14922
rect 0 14864 3790 14920
rect 3846 14864 3851 14920
rect 0 14862 3851 14864
rect 0 14832 480 14862
rect 3785 14859 3851 14862
rect 8845 14922 8911 14925
rect 11792 14922 11852 14998
rect 13486 14996 13492 14998
rect 13556 14996 13562 15060
rect 15101 15058 15167 15061
rect 16757 15058 16823 15061
rect 21173 15058 21239 15061
rect 15101 15056 21239 15058
rect 15101 15000 15106 15056
rect 15162 15000 16762 15056
rect 16818 15000 21178 15056
rect 21234 15000 21239 15056
rect 15101 14998 21239 15000
rect 15101 14995 15167 14998
rect 16757 14995 16823 14998
rect 21173 14995 21239 14998
rect 22737 15058 22803 15061
rect 23054 15058 23060 15060
rect 22737 15056 23060 15058
rect 22737 15000 22742 15056
rect 22798 15000 23060 15056
rect 22737 14998 23060 15000
rect 22737 14995 22803 14998
rect 23054 14996 23060 14998
rect 23124 14996 23130 15060
rect 24301 15058 24367 15061
rect 24710 15058 24716 15060
rect 24301 15056 24716 15058
rect 24301 15000 24306 15056
rect 24362 15000 24716 15056
rect 24301 14998 24716 15000
rect 24301 14995 24367 14998
rect 24710 14996 24716 14998
rect 24780 14996 24786 15060
rect 12157 14922 12223 14925
rect 8845 14920 12223 14922
rect 8845 14864 8850 14920
rect 8906 14864 12162 14920
rect 12218 14864 12223 14920
rect 8845 14862 12223 14864
rect 8845 14859 8911 14862
rect 12157 14859 12223 14862
rect 12382 14860 12388 14924
rect 12452 14922 12458 14924
rect 13445 14922 13511 14925
rect 12452 14920 13511 14922
rect 12452 14864 13450 14920
rect 13506 14864 13511 14920
rect 12452 14862 13511 14864
rect 12452 14860 12458 14862
rect 13445 14859 13511 14862
rect 16389 14922 16455 14925
rect 20069 14922 20135 14925
rect 16389 14920 20135 14922
rect 16389 14864 16394 14920
rect 16450 14864 20074 14920
rect 20130 14864 20135 14920
rect 16389 14862 20135 14864
rect 16389 14859 16455 14862
rect 20069 14859 20135 14862
rect 20294 14860 20300 14924
rect 20364 14922 20370 14924
rect 23473 14922 23539 14925
rect 27520 14922 28000 14952
rect 20364 14920 28000 14922
rect 20364 14864 23478 14920
rect 23534 14864 28000 14920
rect 20364 14862 28000 14864
rect 20364 14860 20370 14862
rect 23473 14859 23539 14862
rect 27520 14832 28000 14862
rect 14825 14786 14891 14789
rect 16757 14786 16823 14789
rect 14825 14784 16823 14786
rect 14825 14728 14830 14784
rect 14886 14728 16762 14784
rect 16818 14728 16823 14784
rect 14825 14726 16823 14728
rect 14825 14723 14891 14726
rect 16757 14723 16823 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 7005 14652 7071 14653
rect 7005 14648 7052 14652
rect 7116 14650 7122 14652
rect 13445 14650 13511 14653
rect 15653 14650 15719 14653
rect 18045 14650 18111 14653
rect 19006 14650 19012 14652
rect 7005 14592 7010 14648
rect 7005 14588 7052 14592
rect 7116 14590 7162 14650
rect 13445 14648 15719 14650
rect 13445 14592 13450 14648
rect 13506 14592 15658 14648
rect 15714 14592 15719 14648
rect 13445 14590 15719 14592
rect 7116 14588 7122 14590
rect 7005 14587 7071 14588
rect 13445 14587 13511 14590
rect 15653 14587 15719 14590
rect 16254 14648 19012 14650
rect 16254 14592 18050 14648
rect 18106 14592 19012 14648
rect 16254 14590 19012 14592
rect 8937 14514 9003 14517
rect 9765 14514 9831 14517
rect 11237 14514 11303 14517
rect 8937 14512 11303 14514
rect 8937 14456 8942 14512
rect 8998 14456 9770 14512
rect 9826 14456 11242 14512
rect 11298 14456 11303 14512
rect 8937 14454 11303 14456
rect 8937 14451 9003 14454
rect 9765 14451 9831 14454
rect 11237 14451 11303 14454
rect 15101 14514 15167 14517
rect 16254 14514 16314 14590
rect 18045 14587 18111 14590
rect 19006 14588 19012 14590
rect 19076 14588 19082 14652
rect 20989 14650 21055 14653
rect 25814 14650 25820 14652
rect 20989 14648 25820 14650
rect 20989 14592 20994 14648
rect 21050 14592 25820 14648
rect 20989 14590 25820 14592
rect 20989 14587 21055 14590
rect 25814 14588 25820 14590
rect 25884 14588 25890 14652
rect 15101 14512 16314 14514
rect 15101 14456 15106 14512
rect 15162 14456 16314 14512
rect 15101 14454 16314 14456
rect 16389 14514 16455 14517
rect 19977 14514 20043 14517
rect 16389 14512 20043 14514
rect 16389 14456 16394 14512
rect 16450 14456 19982 14512
rect 20038 14456 20043 14512
rect 16389 14454 20043 14456
rect 15101 14451 15167 14454
rect 16389 14451 16455 14454
rect 19977 14451 20043 14454
rect 20621 14514 20687 14517
rect 24209 14514 24275 14517
rect 20621 14512 24275 14514
rect 20621 14456 20626 14512
rect 20682 14456 24214 14512
rect 24270 14456 24275 14512
rect 20621 14454 24275 14456
rect 20621 14451 20687 14454
rect 24209 14451 24275 14454
rect 0 14378 480 14408
rect 11053 14378 11119 14381
rect 0 14376 11119 14378
rect 0 14320 11058 14376
rect 11114 14320 11119 14376
rect 0 14318 11119 14320
rect 0 14288 480 14318
rect 11053 14315 11119 14318
rect 15285 14378 15351 14381
rect 19333 14378 19399 14381
rect 27520 14378 28000 14408
rect 15285 14376 19399 14378
rect 15285 14320 15290 14376
rect 15346 14320 19338 14376
rect 19394 14320 19399 14376
rect 15285 14318 19399 14320
rect 15285 14315 15351 14318
rect 19333 14315 19399 14318
rect 19566 14318 28000 14378
rect 6637 14242 6703 14245
rect 8937 14242 9003 14245
rect 6637 14240 9003 14242
rect 6637 14184 6642 14240
rect 6698 14184 8942 14240
rect 8998 14184 9003 14240
rect 6637 14182 9003 14184
rect 6637 14179 6703 14182
rect 8937 14179 9003 14182
rect 9806 14180 9812 14244
rect 9876 14242 9882 14244
rect 14733 14242 14799 14245
rect 9876 14240 14799 14242
rect 9876 14184 14738 14240
rect 14794 14184 14799 14240
rect 9876 14182 14799 14184
rect 9876 14180 9882 14182
rect 14733 14179 14799 14182
rect 16246 14180 16252 14244
rect 16316 14242 16322 14244
rect 19566 14242 19626 14318
rect 27520 14288 28000 14318
rect 16316 14182 19626 14242
rect 21541 14242 21607 14245
rect 23657 14242 23723 14245
rect 21541 14240 23723 14242
rect 21541 14184 21546 14240
rect 21602 14184 23662 14240
rect 23718 14184 23723 14240
rect 21541 14182 23723 14184
rect 16316 14180 16322 14182
rect 21541 14179 21607 14182
rect 23657 14179 23723 14182
rect 24710 14180 24716 14244
rect 24780 14242 24786 14244
rect 25221 14242 25287 14245
rect 24780 14240 25287 14242
rect 24780 14184 25226 14240
rect 25282 14184 25287 14240
rect 24780 14182 25287 14184
rect 24780 14180 24786 14182
rect 25221 14179 25287 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 10961 14106 11027 14109
rect 10961 14104 14842 14106
rect 10961 14048 10966 14104
rect 11022 14048 14842 14104
rect 10961 14046 14842 14048
rect 10961 14043 11027 14046
rect 3233 13970 3299 13973
rect 5625 13970 5691 13973
rect 3233 13968 5691 13970
rect 3233 13912 3238 13968
rect 3294 13912 5630 13968
rect 5686 13912 5691 13968
rect 3233 13910 5691 13912
rect 3233 13907 3299 13910
rect 5625 13907 5691 13910
rect 6862 13908 6868 13972
rect 6932 13970 6938 13972
rect 11237 13970 11303 13973
rect 6932 13968 11303 13970
rect 6932 13912 11242 13968
rect 11298 13912 11303 13968
rect 6932 13910 11303 13912
rect 6932 13908 6938 13910
rect 11237 13907 11303 13910
rect 11646 13908 11652 13972
rect 11716 13970 11722 13972
rect 13445 13970 13511 13973
rect 11716 13968 13511 13970
rect 11716 13912 13450 13968
rect 13506 13912 13511 13968
rect 11716 13910 13511 13912
rect 11716 13908 11722 13910
rect 13445 13907 13511 13910
rect 14457 13970 14523 13973
rect 14641 13970 14707 13973
rect 14457 13968 14707 13970
rect 14457 13912 14462 13968
rect 14518 13912 14646 13968
rect 14702 13912 14707 13968
rect 14457 13910 14707 13912
rect 14457 13907 14523 13910
rect 14641 13907 14707 13910
rect 2129 13834 2195 13837
rect 2865 13834 2931 13837
rect 2129 13832 2931 13834
rect 2129 13776 2134 13832
rect 2190 13776 2870 13832
rect 2926 13776 2931 13832
rect 2129 13774 2931 13776
rect 2129 13771 2195 13774
rect 2865 13771 2931 13774
rect 8017 13834 8083 13837
rect 11421 13834 11487 13837
rect 8017 13832 11487 13834
rect 8017 13776 8022 13832
rect 8078 13776 11426 13832
rect 11482 13776 11487 13832
rect 8017 13774 11487 13776
rect 8017 13771 8083 13774
rect 11421 13771 11487 13774
rect 12341 13836 12407 13837
rect 12341 13832 12388 13836
rect 12452 13834 12458 13836
rect 12341 13776 12346 13832
rect 12341 13772 12388 13776
rect 12452 13774 12498 13834
rect 12452 13772 12458 13774
rect 13302 13772 13308 13836
rect 13372 13834 13378 13836
rect 13629 13834 13695 13837
rect 14457 13836 14523 13837
rect 13372 13832 13695 13834
rect 13372 13776 13634 13832
rect 13690 13776 13695 13832
rect 13372 13774 13695 13776
rect 13372 13772 13378 13774
rect 12341 13771 12407 13772
rect 13629 13771 13695 13774
rect 14406 13772 14412 13836
rect 14476 13834 14523 13836
rect 14782 13834 14842 14046
rect 16798 14044 16804 14108
rect 16868 14106 16874 14108
rect 19701 14106 19767 14109
rect 20621 14106 20687 14109
rect 16868 14104 19767 14106
rect 16868 14048 19706 14104
rect 19762 14048 19767 14104
rect 16868 14046 19767 14048
rect 16868 14044 16874 14046
rect 19701 14043 19767 14046
rect 20486 14104 20687 14106
rect 20486 14048 20626 14104
rect 20682 14048 20687 14104
rect 20486 14046 20687 14048
rect 15285 13972 15351 13973
rect 15285 13970 15332 13972
rect 15240 13968 15332 13970
rect 15240 13912 15290 13968
rect 15240 13910 15332 13912
rect 15285 13908 15332 13910
rect 15396 13908 15402 13972
rect 18229 13970 18295 13973
rect 20486 13970 20546 14046
rect 20621 14043 20687 14046
rect 21633 14106 21699 14109
rect 23105 14106 23171 14109
rect 21633 14104 23171 14106
rect 21633 14048 21638 14104
rect 21694 14048 23110 14104
rect 23166 14048 23171 14104
rect 21633 14046 23171 14048
rect 21633 14043 21699 14046
rect 23105 14043 23171 14046
rect 18229 13968 20546 13970
rect 18229 13912 18234 13968
rect 18290 13912 20546 13968
rect 18229 13910 20546 13912
rect 20621 13970 20687 13973
rect 25221 13970 25287 13973
rect 20621 13968 25287 13970
rect 20621 13912 20626 13968
rect 20682 13912 25226 13968
rect 25282 13912 25287 13968
rect 20621 13910 25287 13912
rect 15285 13907 15351 13908
rect 18229 13907 18295 13910
rect 20621 13907 20687 13910
rect 25221 13907 25287 13910
rect 17125 13834 17191 13837
rect 20713 13834 20779 13837
rect 14476 13832 14568 13834
rect 14518 13776 14568 13832
rect 14476 13774 14568 13776
rect 14782 13832 17191 13834
rect 14782 13776 17130 13832
rect 17186 13776 17191 13832
rect 14782 13774 17191 13776
rect 14476 13772 14523 13774
rect 14457 13771 14523 13772
rect 17125 13771 17191 13774
rect 18094 13832 20779 13834
rect 18094 13776 20718 13832
rect 20774 13776 20779 13832
rect 18094 13774 20779 13776
rect 0 13698 480 13728
rect 1117 13698 1183 13701
rect 0 13696 1183 13698
rect 0 13640 1122 13696
rect 1178 13640 1183 13696
rect 0 13638 1183 13640
rect 0 13608 480 13638
rect 1117 13635 1183 13638
rect 9765 13698 9831 13701
rect 10133 13698 10199 13701
rect 9765 13696 10199 13698
rect 9765 13640 9770 13696
rect 9826 13640 10138 13696
rect 10194 13640 10199 13696
rect 9765 13638 10199 13640
rect 9765 13635 9831 13638
rect 10133 13635 10199 13638
rect 10869 13698 10935 13701
rect 18094 13698 18154 13774
rect 20713 13771 20779 13774
rect 10869 13696 18154 13698
rect 10869 13640 10874 13696
rect 10930 13640 18154 13696
rect 10869 13638 18154 13640
rect 10869 13635 10935 13638
rect 22686 13636 22692 13700
rect 22756 13698 22762 13700
rect 27520 13698 28000 13728
rect 22756 13638 28000 13698
rect 22756 13636 22762 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 27520 13608 28000 13638
rect 19610 13567 19930 13568
rect 6361 13562 6427 13565
rect 6318 13560 6427 13562
rect 6318 13504 6366 13560
rect 6422 13504 6427 13560
rect 6318 13499 6427 13504
rect 10777 13562 10843 13565
rect 13670 13562 13676 13564
rect 10777 13560 13676 13562
rect 10777 13504 10782 13560
rect 10838 13504 13676 13560
rect 10777 13502 13676 13504
rect 10777 13499 10843 13502
rect 13670 13500 13676 13502
rect 13740 13500 13746 13564
rect 13813 13562 13879 13565
rect 16665 13562 16731 13565
rect 13813 13560 16731 13562
rect 13813 13504 13818 13560
rect 13874 13504 16670 13560
rect 16726 13504 16731 13560
rect 13813 13502 16731 13504
rect 4061 13426 4127 13429
rect 6318 13426 6378 13499
rect 4061 13424 6378 13426
rect 4061 13368 4066 13424
rect 4122 13368 6378 13424
rect 4061 13366 6378 13368
rect 9029 13426 9095 13429
rect 11605 13426 11671 13429
rect 13445 13426 13511 13429
rect 9029 13424 13511 13426
rect 9029 13368 9034 13424
rect 9090 13368 11610 13424
rect 11666 13368 13450 13424
rect 13506 13368 13511 13424
rect 9029 13366 13511 13368
rect 13678 13426 13738 13500
rect 13813 13499 13879 13502
rect 16665 13499 16731 13502
rect 17953 13562 18019 13565
rect 19333 13562 19399 13565
rect 23197 13562 23263 13565
rect 17953 13560 19399 13562
rect 17953 13504 17958 13560
rect 18014 13504 19338 13560
rect 19394 13504 19399 13560
rect 17953 13502 19399 13504
rect 17953 13499 18019 13502
rect 19333 13499 19399 13502
rect 20072 13560 23263 13562
rect 20072 13504 23202 13560
rect 23258 13504 23263 13560
rect 20072 13502 23263 13504
rect 13905 13426 13971 13429
rect 13678 13424 13971 13426
rect 13678 13368 13910 13424
rect 13966 13368 13971 13424
rect 13678 13366 13971 13368
rect 4061 13363 4127 13366
rect 9029 13363 9095 13366
rect 11605 13363 11671 13366
rect 13445 13363 13511 13366
rect 13905 13363 13971 13366
rect 14089 13426 14155 13429
rect 17033 13426 17099 13429
rect 14089 13424 17099 13426
rect 14089 13368 14094 13424
rect 14150 13368 17038 13424
rect 17094 13368 17099 13424
rect 14089 13366 17099 13368
rect 14089 13363 14155 13366
rect 17033 13363 17099 13366
rect 17585 13426 17651 13429
rect 20072 13426 20132 13502
rect 23197 13499 23263 13502
rect 23657 13562 23723 13565
rect 25078 13562 25084 13564
rect 23657 13560 25084 13562
rect 23657 13504 23662 13560
rect 23718 13504 25084 13560
rect 23657 13502 25084 13504
rect 23657 13499 23723 13502
rect 25078 13500 25084 13502
rect 25148 13500 25154 13564
rect 17585 13424 20132 13426
rect 17585 13368 17590 13424
rect 17646 13368 20132 13424
rect 17585 13366 20132 13368
rect 20302 13366 24962 13426
rect 17585 13363 17651 13366
rect 3509 13290 3575 13293
rect 12801 13290 12867 13293
rect 16021 13290 16087 13293
rect 16246 13290 16252 13292
rect 3509 13288 12220 13290
rect 3509 13232 3514 13288
rect 3570 13232 12220 13288
rect 3509 13230 12220 13232
rect 3509 13227 3575 13230
rect 0 13154 480 13184
rect 841 13154 907 13157
rect 0 13152 907 13154
rect 0 13096 846 13152
rect 902 13096 907 13152
rect 0 13094 907 13096
rect 0 13064 480 13094
rect 841 13091 907 13094
rect 1761 13154 1827 13157
rect 2446 13154 2452 13156
rect 1761 13152 2452 13154
rect 1761 13096 1766 13152
rect 1822 13096 2452 13152
rect 1761 13094 2452 13096
rect 1761 13091 1827 13094
rect 2446 13092 2452 13094
rect 2516 13092 2522 13156
rect 3877 13154 3943 13157
rect 4061 13154 4127 13157
rect 6361 13156 6427 13157
rect 3877 13152 4127 13154
rect 3877 13096 3882 13152
rect 3938 13096 4066 13152
rect 4122 13096 4127 13152
rect 3877 13094 4127 13096
rect 3877 13091 3943 13094
rect 4061 13091 4127 13094
rect 6310 13092 6316 13156
rect 6380 13154 6427 13156
rect 12160 13154 12220 13230
rect 12801 13288 15394 13290
rect 12801 13232 12806 13288
rect 12862 13232 15394 13288
rect 12801 13230 15394 13232
rect 12801 13227 12867 13230
rect 13721 13154 13787 13157
rect 6380 13152 6472 13154
rect 6422 13096 6472 13152
rect 6380 13094 6472 13096
rect 12160 13152 13787 13154
rect 12160 13096 13726 13152
rect 13782 13096 13787 13152
rect 12160 13094 13787 13096
rect 15334 13154 15394 13230
rect 16021 13288 16252 13290
rect 16021 13232 16026 13288
rect 16082 13232 16252 13288
rect 16021 13230 16252 13232
rect 16021 13227 16087 13230
rect 16246 13228 16252 13230
rect 16316 13228 16322 13292
rect 17217 13290 17283 13293
rect 17718 13290 17724 13292
rect 17217 13288 17724 13290
rect 17217 13232 17222 13288
rect 17278 13232 17724 13288
rect 17217 13230 17724 13232
rect 17217 13227 17283 13230
rect 17718 13228 17724 13230
rect 17788 13228 17794 13292
rect 18505 13290 18571 13293
rect 20302 13290 20362 13366
rect 18505 13288 20362 13290
rect 18505 13232 18510 13288
rect 18566 13232 20362 13288
rect 18505 13230 20362 13232
rect 21173 13290 21239 13293
rect 24761 13290 24827 13293
rect 21173 13288 24827 13290
rect 21173 13232 21178 13288
rect 21234 13232 24766 13288
rect 24822 13232 24827 13288
rect 21173 13230 24827 13232
rect 18505 13227 18571 13230
rect 21173 13227 21239 13230
rect 24761 13227 24827 13230
rect 23197 13154 23263 13157
rect 15334 13152 23263 13154
rect 15334 13096 23202 13152
rect 23258 13096 23263 13152
rect 15334 13094 23263 13096
rect 24902 13154 24962 13366
rect 27520 13154 28000 13184
rect 24902 13094 28000 13154
rect 6380 13092 6427 13094
rect 6361 13091 6427 13092
rect 13721 13091 13787 13094
rect 23197 13091 23263 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 27520 13064 28000 13094
rect 24277 13023 24597 13024
rect 2681 13018 2747 13021
rect 3366 13018 3372 13020
rect 2681 13016 3372 13018
rect 2681 12960 2686 13016
rect 2742 12960 3372 13016
rect 2681 12958 3372 12960
rect 2681 12955 2747 12958
rect 3366 12956 3372 12958
rect 3436 12956 3442 13020
rect 6729 13018 6795 13021
rect 8201 13018 8267 13021
rect 6729 13016 8267 13018
rect 6729 12960 6734 13016
rect 6790 12960 8206 13016
rect 8262 12960 8267 13016
rect 6729 12958 8267 12960
rect 6729 12955 6795 12958
rect 8201 12955 8267 12958
rect 9397 13018 9463 13021
rect 10869 13018 10935 13021
rect 14641 13020 14707 13021
rect 9397 13016 10935 13018
rect 9397 12960 9402 13016
rect 9458 12960 10874 13016
rect 10930 12960 10935 13016
rect 9397 12958 10935 12960
rect 9397 12955 9463 12958
rect 10869 12955 10935 12958
rect 14590 12956 14596 13020
rect 14660 13018 14707 13020
rect 20253 13018 20319 13021
rect 22645 13018 22711 13021
rect 14660 13016 14752 13018
rect 14702 12960 14752 13016
rect 14660 12958 14752 12960
rect 20253 13016 22711 13018
rect 20253 12960 20258 13016
rect 20314 12960 22650 13016
rect 22706 12960 22711 13016
rect 20253 12958 22711 12960
rect 14660 12956 14707 12958
rect 14641 12955 14707 12956
rect 20253 12955 20319 12958
rect 22645 12955 22711 12958
rect 24761 13018 24827 13021
rect 24894 13018 24900 13020
rect 24761 13016 24900 13018
rect 24761 12960 24766 13016
rect 24822 12960 24900 13016
rect 24761 12958 24900 12960
rect 24761 12955 24827 12958
rect 24894 12956 24900 12958
rect 24964 12956 24970 13020
rect 2773 12882 2839 12885
rect 5165 12882 5231 12885
rect 10777 12882 10843 12885
rect 17953 12882 18019 12885
rect 2773 12880 3250 12882
rect 2773 12824 2778 12880
rect 2834 12824 3250 12880
rect 2773 12822 3250 12824
rect 2773 12819 2839 12822
rect 3190 12746 3250 12822
rect 5165 12880 10843 12882
rect 5165 12824 5170 12880
rect 5226 12824 10782 12880
rect 10838 12824 10843 12880
rect 5165 12822 10843 12824
rect 5165 12819 5231 12822
rect 10777 12819 10843 12822
rect 12022 12880 18019 12882
rect 12022 12824 17958 12880
rect 18014 12824 18019 12880
rect 12022 12822 18019 12824
rect 8385 12746 8451 12749
rect 11881 12746 11947 12749
rect 3190 12744 8451 12746
rect 3190 12688 8390 12744
rect 8446 12688 8451 12744
rect 3190 12686 8451 12688
rect 8385 12683 8451 12686
rect 8526 12744 11947 12746
rect 8526 12688 11886 12744
rect 11942 12688 11947 12744
rect 8526 12686 11947 12688
rect 0 12610 480 12640
rect 4838 12610 4844 12612
rect 0 12550 4844 12610
rect 0 12520 480 12550
rect 4838 12548 4844 12550
rect 4908 12548 4914 12612
rect 8017 12610 8083 12613
rect 8526 12610 8586 12686
rect 11881 12683 11947 12686
rect 8017 12608 8586 12610
rect 8017 12552 8022 12608
rect 8078 12552 8586 12608
rect 8017 12550 8586 12552
rect 9857 12610 9923 12613
rect 9990 12610 9996 12612
rect 9857 12608 9996 12610
rect 9857 12552 9862 12608
rect 9918 12552 9996 12608
rect 9857 12550 9996 12552
rect 8017 12547 8083 12550
rect 9857 12547 9923 12550
rect 9990 12548 9996 12550
rect 10060 12548 10066 12612
rect 11145 12610 11211 12613
rect 12022 12610 12082 12822
rect 17953 12819 18019 12822
rect 18873 12882 18939 12885
rect 21817 12882 21883 12885
rect 18873 12880 21883 12882
rect 18873 12824 18878 12880
rect 18934 12824 21822 12880
rect 21878 12824 21883 12880
rect 18873 12822 21883 12824
rect 18873 12819 18939 12822
rect 21817 12819 21883 12822
rect 22318 12820 22324 12884
rect 22388 12882 22394 12884
rect 22645 12882 22711 12885
rect 22388 12880 22711 12882
rect 22388 12824 22650 12880
rect 22706 12824 22711 12880
rect 22388 12822 22711 12824
rect 22388 12820 22394 12822
rect 22645 12819 22711 12822
rect 22921 12882 22987 12885
rect 24853 12884 24919 12885
rect 23238 12882 23244 12884
rect 22921 12880 23244 12882
rect 22921 12824 22926 12880
rect 22982 12824 23244 12880
rect 22921 12822 23244 12824
rect 22921 12819 22987 12822
rect 23238 12820 23244 12822
rect 23308 12820 23314 12884
rect 24853 12882 24900 12884
rect 24808 12880 24900 12882
rect 24808 12824 24858 12880
rect 24808 12822 24900 12824
rect 24853 12820 24900 12822
rect 24964 12820 24970 12884
rect 24853 12819 24919 12820
rect 15653 12746 15719 12749
rect 20989 12746 21055 12749
rect 22829 12748 22895 12749
rect 22829 12746 22876 12748
rect 15653 12744 21055 12746
rect 15653 12688 15658 12744
rect 15714 12688 20994 12744
rect 21050 12688 21055 12744
rect 15653 12686 21055 12688
rect 22784 12744 22876 12746
rect 22784 12688 22834 12744
rect 22784 12686 22876 12688
rect 15653 12683 15719 12686
rect 20989 12683 21055 12686
rect 22829 12684 22876 12686
rect 22940 12684 22946 12748
rect 22829 12683 22895 12684
rect 15377 12610 15443 12613
rect 11145 12608 12082 12610
rect 11145 12552 11150 12608
rect 11206 12552 12082 12608
rect 11145 12550 12082 12552
rect 14230 12608 15443 12610
rect 14230 12552 15382 12608
rect 15438 12552 15443 12608
rect 14230 12550 15443 12552
rect 11145 12547 11211 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 1485 12474 1551 12477
rect 1945 12474 2011 12477
rect 1485 12472 2011 12474
rect 1485 12416 1490 12472
rect 1546 12416 1950 12472
rect 2006 12416 2011 12472
rect 1485 12414 2011 12416
rect 1485 12411 1551 12414
rect 1945 12411 2011 12414
rect 5441 12474 5507 12477
rect 6862 12474 6868 12476
rect 5441 12472 6868 12474
rect 5441 12416 5446 12472
rect 5502 12416 6868 12472
rect 5441 12414 6868 12416
rect 5441 12411 5507 12414
rect 6862 12412 6868 12414
rect 6932 12412 6938 12476
rect 7189 12474 7255 12477
rect 9990 12474 9996 12476
rect 7008 12472 9996 12474
rect 7008 12416 7194 12472
rect 7250 12416 9996 12472
rect 7008 12414 9996 12416
rect 6729 12338 6795 12341
rect 7008 12338 7068 12414
rect 7189 12411 7255 12414
rect 9990 12412 9996 12414
rect 10060 12412 10066 12476
rect 13302 12412 13308 12476
rect 13372 12474 13378 12476
rect 14230 12474 14290 12550
rect 15377 12547 15443 12550
rect 15518 12550 19488 12610
rect 13372 12414 14290 12474
rect 14365 12474 14431 12477
rect 14590 12474 14596 12476
rect 14365 12472 14596 12474
rect 14365 12416 14370 12472
rect 14426 12416 14596 12472
rect 14365 12414 14596 12416
rect 13372 12412 13378 12414
rect 14365 12411 14431 12414
rect 14590 12412 14596 12414
rect 14660 12412 14666 12476
rect 14917 12474 14983 12477
rect 15518 12474 15578 12550
rect 14917 12472 15578 12474
rect 14917 12416 14922 12472
rect 14978 12416 15578 12472
rect 14917 12414 15578 12416
rect 17033 12474 17099 12477
rect 17309 12474 17375 12477
rect 17033 12472 17375 12474
rect 17033 12416 17038 12472
rect 17094 12416 17314 12472
rect 17370 12416 17375 12472
rect 17033 12414 17375 12416
rect 14917 12411 14983 12414
rect 17033 12411 17099 12414
rect 17309 12411 17375 12414
rect 17953 12474 18019 12477
rect 17953 12472 19258 12474
rect 17953 12416 17958 12472
rect 18014 12416 19258 12472
rect 17953 12414 19258 12416
rect 17953 12411 18019 12414
rect 6729 12336 7068 12338
rect 6729 12280 6734 12336
rect 6790 12280 7068 12336
rect 6729 12278 7068 12280
rect 8109 12338 8175 12341
rect 9305 12338 9371 12341
rect 10409 12338 10475 12341
rect 8109 12336 10475 12338
rect 8109 12280 8114 12336
rect 8170 12280 9310 12336
rect 9366 12280 10414 12336
rect 10470 12280 10475 12336
rect 8109 12278 10475 12280
rect 6729 12275 6795 12278
rect 8109 12275 8175 12278
rect 9305 12275 9371 12278
rect 10409 12275 10475 12278
rect 10685 12338 10751 12341
rect 13629 12338 13695 12341
rect 10685 12336 13695 12338
rect 10685 12280 10690 12336
rect 10746 12280 13634 12336
rect 13690 12280 13695 12336
rect 10685 12278 13695 12280
rect 10685 12275 10751 12278
rect 13629 12275 13695 12278
rect 13854 12276 13860 12340
rect 13924 12338 13930 12340
rect 15377 12338 15443 12341
rect 13924 12336 15443 12338
rect 13924 12280 15382 12336
rect 15438 12280 15443 12336
rect 13924 12278 15443 12280
rect 13924 12276 13930 12278
rect 15377 12275 15443 12278
rect 15929 12338 15995 12341
rect 16757 12340 16823 12341
rect 16246 12338 16252 12340
rect 15929 12336 16252 12338
rect 15929 12280 15934 12336
rect 15990 12280 16252 12336
rect 15929 12278 16252 12280
rect 15929 12275 15995 12278
rect 16246 12276 16252 12278
rect 16316 12276 16322 12340
rect 16757 12338 16804 12340
rect 16712 12336 16804 12338
rect 16712 12280 16762 12336
rect 16712 12278 16804 12280
rect 16757 12276 16804 12278
rect 16868 12276 16874 12340
rect 16757 12275 16823 12276
rect 7557 12202 7623 12205
rect 11513 12202 11579 12205
rect 7557 12200 11579 12202
rect 7557 12144 7562 12200
rect 7618 12144 11518 12200
rect 11574 12144 11579 12200
rect 7557 12142 11579 12144
rect 7557 12139 7623 12142
rect 11513 12139 11579 12142
rect 11830 12140 11836 12204
rect 11900 12202 11906 12204
rect 16389 12202 16455 12205
rect 11900 12200 16455 12202
rect 11900 12144 16394 12200
rect 16450 12144 16455 12200
rect 11900 12142 16455 12144
rect 19198 12202 19258 12414
rect 19428 12338 19488 12550
rect 22502 12548 22508 12612
rect 22572 12610 22578 12612
rect 27520 12610 28000 12640
rect 22572 12550 28000 12610
rect 22572 12548 22578 12550
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 27520 12520 28000 12550
rect 19610 12479 19930 12480
rect 23657 12476 23723 12477
rect 23606 12474 23612 12476
rect 23566 12414 23612 12474
rect 23676 12472 23723 12476
rect 23718 12416 23723 12472
rect 23606 12412 23612 12414
rect 23676 12412 23723 12416
rect 23657 12411 23723 12412
rect 24117 12474 24183 12477
rect 25446 12474 25452 12476
rect 24117 12472 25452 12474
rect 24117 12416 24122 12472
rect 24178 12416 25452 12472
rect 24117 12414 25452 12416
rect 24117 12411 24183 12414
rect 25446 12412 25452 12414
rect 25516 12412 25522 12476
rect 22001 12338 22067 12341
rect 19428 12336 22067 12338
rect 19428 12280 22006 12336
rect 22062 12280 22067 12336
rect 19428 12278 22067 12280
rect 22001 12275 22067 12278
rect 22277 12338 22343 12341
rect 22870 12338 22876 12340
rect 22277 12336 22876 12338
rect 22277 12280 22282 12336
rect 22338 12280 22876 12336
rect 22277 12278 22876 12280
rect 22277 12275 22343 12278
rect 22870 12276 22876 12278
rect 22940 12276 22946 12340
rect 20805 12202 20871 12205
rect 19198 12200 20871 12202
rect 19198 12144 20810 12200
rect 20866 12144 20871 12200
rect 19198 12142 20871 12144
rect 11900 12140 11906 12142
rect 16389 12139 16455 12142
rect 20805 12139 20871 12142
rect 21081 12202 21147 12205
rect 23565 12202 23631 12205
rect 21081 12200 23631 12202
rect 21081 12144 21086 12200
rect 21142 12144 23570 12200
rect 23626 12144 23631 12200
rect 21081 12142 23631 12144
rect 21081 12139 21147 12142
rect 23565 12139 23631 12142
rect 6085 12066 6151 12069
rect 10225 12066 10291 12069
rect 6085 12064 10291 12066
rect 6085 12008 6090 12064
rect 6146 12008 10230 12064
rect 10286 12008 10291 12064
rect 6085 12006 10291 12008
rect 6085 12003 6151 12006
rect 10225 12003 10291 12006
rect 10409 12066 10475 12069
rect 14457 12066 14523 12069
rect 21541 12066 21607 12069
rect 10409 12064 14842 12066
rect 10409 12008 10414 12064
rect 10470 12008 14462 12064
rect 14518 12008 14842 12064
rect 10409 12006 14842 12008
rect 10409 12003 10475 12006
rect 14457 12003 14523 12006
rect 5610 12000 5930 12001
rect 0 11930 480 11960
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 933 11930 999 11933
rect 0 11928 999 11930
rect 0 11872 938 11928
rect 994 11872 999 11928
rect 0 11870 999 11872
rect 0 11840 480 11870
rect 933 11867 999 11870
rect 8477 11930 8543 11933
rect 11329 11930 11395 11933
rect 8477 11928 11395 11930
rect 8477 11872 8482 11928
rect 8538 11872 11334 11928
rect 11390 11872 11395 11928
rect 8477 11870 11395 11872
rect 8477 11867 8543 11870
rect 11329 11867 11395 11870
rect 11697 11930 11763 11933
rect 12566 11930 12572 11932
rect 11697 11928 12572 11930
rect 11697 11872 11702 11928
rect 11758 11872 12572 11928
rect 11697 11870 12572 11872
rect 11697 11867 11763 11870
rect 12566 11868 12572 11870
rect 12636 11868 12642 11932
rect 13670 11868 13676 11932
rect 13740 11930 13746 11932
rect 14641 11930 14707 11933
rect 13740 11928 14707 11930
rect 13740 11872 14646 11928
rect 14702 11872 14707 11928
rect 13740 11870 14707 11872
rect 13740 11868 13746 11870
rect 14641 11867 14707 11870
rect 3417 11794 3483 11797
rect 3693 11794 3759 11797
rect 10133 11794 10199 11797
rect 11789 11796 11855 11797
rect 11789 11794 11836 11796
rect 3417 11792 10199 11794
rect 3417 11736 3422 11792
rect 3478 11736 3698 11792
rect 3754 11736 10138 11792
rect 10194 11736 10199 11792
rect 3417 11734 10199 11736
rect 3417 11731 3483 11734
rect 3693 11731 3759 11734
rect 10133 11731 10199 11734
rect 11102 11792 11836 11794
rect 11102 11736 11794 11792
rect 11102 11734 11836 11736
rect 2681 11658 2747 11661
rect 3233 11658 3299 11661
rect 3969 11658 4035 11661
rect 2681 11656 4035 11658
rect 2681 11600 2686 11656
rect 2742 11600 3238 11656
rect 3294 11600 3974 11656
rect 4030 11600 4035 11656
rect 2681 11598 4035 11600
rect 2681 11595 2747 11598
rect 3233 11595 3299 11598
rect 3969 11595 4035 11598
rect 5533 11658 5599 11661
rect 9673 11658 9739 11661
rect 11102 11658 11162 11734
rect 11789 11732 11836 11734
rect 11900 11732 11906 11796
rect 14782 11794 14842 12006
rect 16990 12064 21607 12066
rect 16990 12008 21546 12064
rect 21602 12008 21607 12064
rect 16990 12006 21607 12008
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 15745 11930 15811 11933
rect 16990 11930 17050 12006
rect 21541 12003 21607 12006
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 15745 11928 17050 11930
rect 15745 11872 15750 11928
rect 15806 11872 17050 11928
rect 15745 11870 17050 11872
rect 17125 11930 17191 11933
rect 21030 11930 21036 11932
rect 17125 11928 21036 11930
rect 17125 11872 17130 11928
rect 17186 11872 21036 11928
rect 17125 11870 21036 11872
rect 15745 11867 15811 11870
rect 17125 11867 17191 11870
rect 21030 11868 21036 11870
rect 21100 11868 21106 11932
rect 23054 11868 23060 11932
rect 23124 11930 23130 11932
rect 23381 11930 23447 11933
rect 23124 11928 23447 11930
rect 23124 11872 23386 11928
rect 23442 11872 23447 11928
rect 23124 11870 23447 11872
rect 23124 11868 23130 11870
rect 23381 11867 23447 11870
rect 25129 11930 25195 11933
rect 27520 11930 28000 11960
rect 25129 11928 28000 11930
rect 25129 11872 25134 11928
rect 25190 11872 28000 11928
rect 25129 11870 28000 11872
rect 25129 11867 25195 11870
rect 27520 11840 28000 11870
rect 17401 11794 17467 11797
rect 14782 11792 17467 11794
rect 14782 11736 17406 11792
rect 17462 11736 17467 11792
rect 14782 11734 17467 11736
rect 11789 11731 11855 11732
rect 17401 11731 17467 11734
rect 20478 11732 20484 11796
rect 20548 11794 20554 11796
rect 25957 11794 26023 11797
rect 20548 11792 26023 11794
rect 20548 11736 25962 11792
rect 26018 11736 26023 11792
rect 20548 11734 26023 11736
rect 20548 11732 20554 11734
rect 25957 11731 26023 11734
rect 5533 11656 9739 11658
rect 5533 11600 5538 11656
rect 5594 11600 9678 11656
rect 9734 11600 9739 11656
rect 5533 11598 9739 11600
rect 5533 11595 5599 11598
rect 9673 11595 9739 11598
rect 9998 11598 11162 11658
rect 11237 11660 11303 11661
rect 11237 11656 11284 11660
rect 11348 11658 11354 11660
rect 11973 11658 12039 11661
rect 13813 11658 13879 11661
rect 21081 11658 21147 11661
rect 11237 11600 11242 11656
rect 2681 11522 2747 11525
rect 6821 11522 6887 11525
rect 9998 11522 10058 11598
rect 11237 11596 11284 11600
rect 11348 11598 11394 11658
rect 11973 11656 21147 11658
rect 11973 11600 11978 11656
rect 12034 11600 13818 11656
rect 13874 11600 21086 11656
rect 21142 11600 21147 11656
rect 11973 11598 21147 11600
rect 11348 11596 11354 11598
rect 11237 11595 11303 11596
rect 11973 11595 12039 11598
rect 13813 11595 13879 11598
rect 21081 11595 21147 11598
rect 21357 11658 21423 11661
rect 23013 11658 23079 11661
rect 21357 11656 23079 11658
rect 21357 11600 21362 11656
rect 21418 11600 23018 11656
rect 23074 11600 23079 11656
rect 21357 11598 23079 11600
rect 21357 11595 21423 11598
rect 23013 11595 23079 11598
rect 23197 11658 23263 11661
rect 24945 11658 25011 11661
rect 23197 11656 25011 11658
rect 23197 11600 23202 11656
rect 23258 11600 24950 11656
rect 25006 11600 25011 11656
rect 23197 11598 25011 11600
rect 23197 11595 23263 11598
rect 24945 11595 25011 11598
rect 15653 11522 15719 11525
rect 2681 11520 6887 11522
rect 2681 11464 2686 11520
rect 2742 11464 6826 11520
rect 6882 11464 6887 11520
rect 2681 11462 6887 11464
rect 2681 11459 2747 11462
rect 6821 11459 6887 11462
rect 7054 11462 10058 11522
rect 10688 11520 15719 11522
rect 10688 11464 15658 11520
rect 15714 11464 15719 11520
rect 10688 11462 15719 11464
rect 0 11386 480 11416
rect 7054 11386 7114 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 7373 11388 7439 11389
rect 7373 11386 7420 11388
rect 0 11326 7114 11386
rect 7328 11384 7420 11386
rect 7328 11328 7378 11384
rect 7328 11326 7420 11328
rect 0 11296 480 11326
rect 7373 11324 7420 11326
rect 7484 11324 7490 11388
rect 7373 11323 7439 11324
rect 841 11250 907 11253
rect 8937 11250 9003 11253
rect 841 11248 9003 11250
rect 841 11192 846 11248
rect 902 11192 8942 11248
rect 8998 11192 9003 11248
rect 841 11190 9003 11192
rect 841 11187 907 11190
rect 8937 11187 9003 11190
rect 9990 11188 9996 11252
rect 10060 11250 10066 11252
rect 10688 11250 10748 11462
rect 15653 11459 15719 11462
rect 17309 11522 17375 11525
rect 17718 11522 17724 11524
rect 17309 11520 17724 11522
rect 17309 11464 17314 11520
rect 17370 11464 17724 11520
rect 17309 11462 17724 11464
rect 17309 11459 17375 11462
rect 17718 11460 17724 11462
rect 17788 11460 17794 11524
rect 20897 11522 20963 11525
rect 25405 11522 25471 11525
rect 20897 11520 25471 11522
rect 20897 11464 20902 11520
rect 20958 11464 25410 11520
rect 25466 11464 25471 11520
rect 20897 11462 25471 11464
rect 20897 11459 20963 11462
rect 25405 11459 25471 11462
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 10910 11324 10916 11388
rect 10980 11386 10986 11388
rect 10980 11326 19488 11386
rect 10980 11324 10986 11326
rect 10060 11190 10748 11250
rect 12341 11250 12407 11253
rect 17677 11250 17743 11253
rect 12341 11248 17743 11250
rect 12341 11192 12346 11248
rect 12402 11192 17682 11248
rect 17738 11192 17743 11248
rect 12341 11190 17743 11192
rect 19428 11250 19488 11326
rect 21950 11324 21956 11388
rect 22020 11386 22026 11388
rect 27520 11386 28000 11416
rect 22020 11326 28000 11386
rect 22020 11324 22026 11326
rect 27520 11296 28000 11326
rect 20713 11250 20779 11253
rect 21357 11250 21423 11253
rect 25129 11250 25195 11253
rect 19428 11248 21423 11250
rect 19428 11192 20718 11248
rect 20774 11192 21362 11248
rect 21418 11192 21423 11248
rect 19428 11190 21423 11192
rect 10060 11188 10066 11190
rect 12341 11187 12407 11190
rect 17677 11187 17743 11190
rect 20713 11187 20779 11190
rect 21357 11187 21423 11190
rect 21590 11248 25195 11250
rect 21590 11192 25134 11248
rect 25190 11192 25195 11248
rect 21590 11190 25195 11192
rect 2129 11114 2195 11117
rect 3366 11114 3372 11116
rect 2129 11112 3372 11114
rect 2129 11056 2134 11112
rect 2190 11056 3372 11112
rect 2129 11054 3372 11056
rect 2129 11051 2195 11054
rect 3366 11052 3372 11054
rect 3436 11052 3442 11116
rect 3601 11114 3667 11117
rect 7833 11114 7899 11117
rect 3601 11112 7899 11114
rect 3601 11056 3606 11112
rect 3662 11056 7838 11112
rect 7894 11056 7899 11112
rect 3601 11054 7899 11056
rect 3601 11051 3667 11054
rect 7833 11051 7899 11054
rect 9489 11114 9555 11117
rect 12065 11114 12131 11117
rect 12341 11114 12407 11117
rect 15745 11116 15811 11117
rect 15694 11114 15700 11116
rect 9489 11112 12407 11114
rect 9489 11056 9494 11112
rect 9550 11056 12070 11112
rect 12126 11056 12346 11112
rect 12402 11056 12407 11112
rect 9489 11054 12407 11056
rect 9489 11051 9555 11054
rect 12065 11051 12131 11054
rect 12341 11051 12407 11054
rect 14782 11054 15394 11114
rect 15654 11054 15700 11114
rect 15764 11112 15811 11116
rect 15806 11056 15811 11112
rect 7649 10978 7715 10981
rect 12801 10978 12867 10981
rect 7649 10976 12867 10978
rect 7649 10920 7654 10976
rect 7710 10920 12806 10976
rect 12862 10920 12867 10976
rect 7649 10918 12867 10920
rect 7649 10915 7715 10918
rect 12801 10915 12867 10918
rect 5610 10912 5930 10913
rect 0 10842 480 10872
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 4838 10842 4844 10844
rect 0 10782 4844 10842
rect 0 10752 480 10782
rect 4838 10780 4844 10782
rect 4908 10780 4914 10844
rect 7373 10842 7439 10845
rect 8293 10842 8359 10845
rect 14641 10842 14707 10845
rect 14782 10842 14842 11054
rect 15334 10978 15394 11054
rect 15694 11052 15700 11054
rect 15764 11052 15811 11056
rect 19374 11052 19380 11116
rect 19444 11114 19450 11116
rect 21590 11114 21650 11190
rect 25129 11187 25195 11190
rect 19444 11054 21650 11114
rect 23933 11114 23999 11117
rect 25313 11114 25379 11117
rect 23933 11112 25379 11114
rect 23933 11056 23938 11112
rect 23994 11056 25318 11112
rect 25374 11056 25379 11112
rect 23933 11054 25379 11056
rect 19444 11052 19450 11054
rect 15745 11051 15811 11052
rect 23933 11051 23999 11054
rect 25313 11051 25379 11054
rect 17166 10978 17172 10980
rect 15334 10918 17172 10978
rect 17166 10916 17172 10918
rect 17236 10978 17242 10980
rect 17677 10978 17743 10981
rect 17236 10976 17743 10978
rect 17236 10920 17682 10976
rect 17738 10920 17743 10976
rect 17236 10918 17743 10920
rect 17236 10916 17242 10918
rect 17677 10915 17743 10918
rect 18045 10978 18111 10981
rect 20897 10978 20963 10981
rect 18045 10976 20963 10978
rect 18045 10920 18050 10976
rect 18106 10920 20902 10976
rect 20958 10920 20963 10976
rect 18045 10918 20963 10920
rect 18045 10915 18111 10918
rect 20897 10915 20963 10918
rect 22001 10978 22067 10981
rect 23473 10978 23539 10981
rect 22001 10976 23539 10978
rect 22001 10920 22006 10976
rect 22062 10920 23478 10976
rect 23534 10920 23539 10976
rect 22001 10918 23539 10920
rect 22001 10915 22067 10918
rect 23473 10915 23539 10918
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 7373 10840 14842 10842
rect 7373 10784 7378 10840
rect 7434 10784 8298 10840
rect 8354 10784 14646 10840
rect 14702 10784 14842 10840
rect 7373 10782 14842 10784
rect 7373 10779 7439 10782
rect 8293 10779 8359 10782
rect 14641 10779 14707 10782
rect 15510 10780 15516 10844
rect 15580 10842 15586 10844
rect 18045 10842 18111 10845
rect 15580 10840 18111 10842
rect 15580 10784 18050 10840
rect 18106 10784 18111 10840
rect 15580 10782 18111 10784
rect 15580 10780 15586 10782
rect 18045 10779 18111 10782
rect 26325 10842 26391 10845
rect 27520 10842 28000 10872
rect 26325 10840 28000 10842
rect 26325 10784 26330 10840
rect 26386 10784 28000 10840
rect 26325 10782 28000 10784
rect 26325 10779 26391 10782
rect 27520 10752 28000 10782
rect 10593 10706 10659 10709
rect 6870 10704 10659 10706
rect 6870 10648 10598 10704
rect 10654 10648 10659 10704
rect 6870 10646 10659 10648
rect 3325 10570 3391 10573
rect 6870 10570 6930 10646
rect 10593 10643 10659 10646
rect 14825 10706 14891 10709
rect 17769 10706 17835 10709
rect 14825 10704 17835 10706
rect 14825 10648 14830 10704
rect 14886 10648 17774 10704
rect 17830 10648 17835 10704
rect 14825 10646 17835 10648
rect 14825 10643 14891 10646
rect 17769 10643 17835 10646
rect 18137 10706 18203 10709
rect 22737 10706 22803 10709
rect 18137 10704 22803 10706
rect 18137 10648 18142 10704
rect 18198 10648 22742 10704
rect 22798 10648 22803 10704
rect 18137 10646 22803 10648
rect 18137 10643 18203 10646
rect 22737 10643 22803 10646
rect 23933 10706 23999 10709
rect 25262 10706 25268 10708
rect 23933 10704 25268 10706
rect 23933 10648 23938 10704
rect 23994 10648 25268 10704
rect 23933 10646 25268 10648
rect 23933 10643 23999 10646
rect 25262 10644 25268 10646
rect 25332 10644 25338 10708
rect 7925 10572 7991 10573
rect 7925 10570 7972 10572
rect 3325 10568 6930 10570
rect 3325 10512 3330 10568
rect 3386 10512 6930 10568
rect 3325 10510 6930 10512
rect 7880 10568 7972 10570
rect 7880 10512 7930 10568
rect 7880 10510 7972 10512
rect 3325 10507 3391 10510
rect 7925 10508 7972 10510
rect 8036 10508 8042 10572
rect 10726 10570 10732 10572
rect 8158 10510 10732 10570
rect 7925 10507 7991 10508
rect 3969 10434 4035 10437
rect 8158 10434 8218 10510
rect 10726 10508 10732 10510
rect 10796 10508 10802 10572
rect 10910 10508 10916 10572
rect 10980 10570 10986 10572
rect 13302 10570 13308 10572
rect 10980 10510 13308 10570
rect 10980 10508 10986 10510
rect 13302 10508 13308 10510
rect 13372 10508 13378 10572
rect 13537 10570 13603 10573
rect 24669 10570 24735 10573
rect 24894 10570 24900 10572
rect 13537 10568 24900 10570
rect 13537 10512 13542 10568
rect 13598 10512 24674 10568
rect 24730 10512 24900 10568
rect 13537 10510 24900 10512
rect 13537 10507 13603 10510
rect 24669 10507 24735 10510
rect 24894 10508 24900 10510
rect 24964 10508 24970 10572
rect 3969 10432 8218 10434
rect 3969 10376 3974 10432
rect 4030 10376 8218 10432
rect 3969 10374 8218 10376
rect 11329 10434 11395 10437
rect 15837 10434 15903 10437
rect 11329 10432 15903 10434
rect 11329 10376 11334 10432
rect 11390 10376 15842 10432
rect 15898 10376 15903 10432
rect 11329 10374 15903 10376
rect 3969 10371 4035 10374
rect 11329 10371 11395 10374
rect 15837 10371 15903 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 3693 10298 3759 10301
rect 3693 10296 9874 10298
rect 3693 10240 3698 10296
rect 3754 10240 9874 10296
rect 3693 10238 9874 10240
rect 3693 10235 3759 10238
rect 0 10162 480 10192
rect 7649 10162 7715 10165
rect 0 10160 7715 10162
rect 0 10104 7654 10160
rect 7710 10104 7715 10160
rect 0 10102 7715 10104
rect 9814 10162 9874 10238
rect 12566 10236 12572 10300
rect 12636 10298 12642 10300
rect 15561 10298 15627 10301
rect 12636 10296 15627 10298
rect 12636 10240 15566 10296
rect 15622 10240 15627 10296
rect 12636 10238 15627 10240
rect 12636 10236 12642 10238
rect 15561 10235 15627 10238
rect 16389 10298 16455 10301
rect 19149 10298 19215 10301
rect 16389 10296 19215 10298
rect 16389 10240 16394 10296
rect 16450 10240 19154 10296
rect 19210 10240 19215 10296
rect 16389 10238 19215 10240
rect 16389 10235 16455 10238
rect 19149 10235 19215 10238
rect 22737 10298 22803 10301
rect 23422 10298 23428 10300
rect 22737 10296 23428 10298
rect 22737 10240 22742 10296
rect 22798 10240 23428 10296
rect 22737 10238 23428 10240
rect 22737 10235 22803 10238
rect 23422 10236 23428 10238
rect 23492 10236 23498 10300
rect 24209 10298 24275 10301
rect 24945 10298 25011 10301
rect 25630 10298 25636 10300
rect 24209 10296 25636 10298
rect 24209 10240 24214 10296
rect 24270 10240 24950 10296
rect 25006 10240 25636 10296
rect 24209 10238 25636 10240
rect 24209 10235 24275 10238
rect 24945 10235 25011 10238
rect 25630 10236 25636 10238
rect 25700 10236 25706 10300
rect 11697 10162 11763 10165
rect 9814 10160 11763 10162
rect 9814 10104 11702 10160
rect 11758 10104 11763 10160
rect 9814 10102 11763 10104
rect 0 10072 480 10102
rect 7649 10099 7715 10102
rect 11697 10099 11763 10102
rect 17493 10162 17559 10165
rect 19517 10162 19583 10165
rect 24117 10162 24183 10165
rect 27520 10162 28000 10192
rect 17493 10160 19583 10162
rect 17493 10104 17498 10160
rect 17554 10104 19522 10160
rect 19578 10104 19583 10160
rect 17493 10102 19583 10104
rect 17493 10099 17559 10102
rect 19517 10099 19583 10102
rect 22372 10160 28000 10162
rect 22372 10104 24122 10160
rect 24178 10104 28000 10160
rect 22372 10102 28000 10104
rect 2405 10026 2471 10029
rect 15653 10026 15719 10029
rect 2405 10024 15719 10026
rect 2405 9968 2410 10024
rect 2466 9968 15658 10024
rect 15714 9968 15719 10024
rect 2405 9966 15719 9968
rect 2405 9963 2471 9966
rect 15653 9963 15719 9966
rect 16021 10026 16087 10029
rect 22372 10026 22432 10102
rect 24117 10099 24183 10102
rect 27520 10072 28000 10102
rect 23013 10026 23079 10029
rect 25129 10026 25195 10029
rect 16021 10024 22432 10026
rect 16021 9968 16026 10024
rect 16082 9968 22432 10024
rect 16021 9966 22432 9968
rect 22510 10024 25195 10026
rect 22510 9968 23018 10024
rect 23074 9968 25134 10024
rect 25190 9968 25195 10024
rect 22510 9966 25195 9968
rect 16021 9963 16087 9966
rect 6545 9890 6611 9893
rect 11237 9890 11303 9893
rect 6545 9888 11303 9890
rect 6545 9832 6550 9888
rect 6606 9832 11242 9888
rect 11298 9832 11303 9888
rect 6545 9830 11303 9832
rect 6545 9827 6611 9830
rect 11237 9827 11303 9830
rect 11605 9890 11671 9893
rect 14365 9890 14431 9893
rect 11605 9888 14431 9890
rect 11605 9832 11610 9888
rect 11666 9832 14370 9888
rect 14426 9832 14431 9888
rect 11605 9830 14431 9832
rect 11605 9827 11671 9830
rect 14365 9827 14431 9830
rect 17953 9890 18019 9893
rect 18505 9890 18571 9893
rect 22510 9890 22570 9966
rect 23013 9963 23079 9966
rect 25129 9963 25195 9966
rect 17953 9888 22570 9890
rect 17953 9832 17958 9888
rect 18014 9832 18510 9888
rect 18566 9832 22570 9888
rect 17953 9830 22570 9832
rect 17953 9827 18019 9830
rect 18505 9827 18571 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 9673 9754 9739 9757
rect 6088 9752 9739 9754
rect 6088 9696 9678 9752
rect 9734 9696 9739 9752
rect 6088 9694 9739 9696
rect 0 9618 480 9648
rect 3969 9618 4035 9621
rect 0 9616 4035 9618
rect 0 9560 3974 9616
rect 4030 9560 4035 9616
rect 0 9558 4035 9560
rect 0 9528 480 9558
rect 3969 9555 4035 9558
rect 5441 9618 5507 9621
rect 6088 9618 6148 9694
rect 9673 9691 9739 9694
rect 10961 9754 11027 9757
rect 11881 9754 11947 9757
rect 12433 9754 12499 9757
rect 10961 9752 12499 9754
rect 10961 9696 10966 9752
rect 11022 9696 11886 9752
rect 11942 9696 12438 9752
rect 12494 9696 12499 9752
rect 10961 9694 12499 9696
rect 10961 9691 11027 9694
rect 11881 9691 11947 9694
rect 12433 9691 12499 9694
rect 18321 9754 18387 9757
rect 22277 9754 22343 9757
rect 23197 9754 23263 9757
rect 18321 9752 23263 9754
rect 18321 9696 18326 9752
rect 18382 9696 22282 9752
rect 22338 9696 23202 9752
rect 23258 9696 23263 9752
rect 18321 9694 23263 9696
rect 18321 9691 18387 9694
rect 22277 9691 22343 9694
rect 23197 9691 23263 9694
rect 5441 9616 6148 9618
rect 5441 9560 5446 9616
rect 5502 9560 6148 9616
rect 5441 9558 6148 9560
rect 11237 9618 11303 9621
rect 12750 9618 12756 9620
rect 11237 9616 12756 9618
rect 11237 9560 11242 9616
rect 11298 9560 12756 9616
rect 11237 9558 12756 9560
rect 5441 9555 5507 9558
rect 11237 9555 11303 9558
rect 12750 9556 12756 9558
rect 12820 9556 12826 9620
rect 14222 9556 14228 9620
rect 14292 9618 14298 9620
rect 15101 9618 15167 9621
rect 19333 9618 19399 9621
rect 20846 9618 20852 9620
rect 14292 9616 15167 9618
rect 14292 9560 15106 9616
rect 15162 9560 15167 9616
rect 14292 9558 15167 9560
rect 14292 9556 14298 9558
rect 15101 9555 15167 9558
rect 16070 9616 20852 9618
rect 16070 9560 19338 9616
rect 19394 9560 20852 9616
rect 16070 9558 20852 9560
rect 6453 9482 6519 9485
rect 14641 9482 14707 9485
rect 6453 9480 14707 9482
rect 6453 9424 6458 9480
rect 6514 9424 14646 9480
rect 14702 9424 14707 9480
rect 6453 9422 14707 9424
rect 6453 9419 6519 9422
rect 14641 9419 14707 9422
rect 14825 9482 14891 9485
rect 16070 9482 16130 9558
rect 19333 9555 19399 9558
rect 20846 9556 20852 9558
rect 20916 9556 20922 9620
rect 21766 9556 21772 9620
rect 21836 9618 21842 9620
rect 24209 9618 24275 9621
rect 27520 9618 28000 9648
rect 21836 9616 28000 9618
rect 21836 9560 24214 9616
rect 24270 9560 28000 9616
rect 21836 9558 28000 9560
rect 21836 9556 21842 9558
rect 24209 9555 24275 9558
rect 27520 9528 28000 9558
rect 19885 9482 19951 9485
rect 14825 9480 16130 9482
rect 14825 9424 14830 9480
rect 14886 9424 16130 9480
rect 14825 9422 16130 9424
rect 16254 9480 19951 9482
rect 16254 9424 19890 9480
rect 19946 9424 19951 9480
rect 16254 9422 19951 9424
rect 14825 9419 14891 9422
rect 11053 9346 11119 9349
rect 12382 9346 12388 9348
rect 11053 9344 12388 9346
rect 11053 9288 11058 9344
rect 11114 9288 12388 9344
rect 11053 9286 12388 9288
rect 11053 9283 11119 9286
rect 12382 9284 12388 9286
rect 12452 9346 12458 9348
rect 16254 9346 16314 9422
rect 19885 9419 19951 9422
rect 12452 9286 16314 9346
rect 18413 9346 18479 9349
rect 19425 9346 19491 9349
rect 18413 9344 19491 9346
rect 18413 9288 18418 9344
rect 18474 9288 19430 9344
rect 19486 9288 19491 9344
rect 18413 9286 19491 9288
rect 12452 9284 12458 9286
rect 18413 9283 18479 9286
rect 19425 9283 19491 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 10777 9210 10843 9213
rect 13169 9210 13235 9213
rect 10777 9208 13235 9210
rect 10777 9152 10782 9208
rect 10838 9152 13174 9208
rect 13230 9152 13235 9208
rect 10777 9150 13235 9152
rect 10777 9147 10843 9150
rect 13169 9147 13235 9150
rect 15009 9210 15075 9213
rect 17493 9210 17559 9213
rect 15009 9208 17559 9210
rect 15009 9152 15014 9208
rect 15070 9152 17498 9208
rect 17554 9152 17559 9208
rect 15009 9150 17559 9152
rect 15009 9147 15075 9150
rect 17493 9147 17559 9150
rect 20529 9210 20595 9213
rect 22829 9210 22895 9213
rect 23054 9210 23060 9212
rect 20529 9208 23060 9210
rect 20529 9152 20534 9208
rect 20590 9152 22834 9208
rect 22890 9152 23060 9208
rect 20529 9150 23060 9152
rect 20529 9147 20595 9150
rect 22829 9147 22895 9150
rect 23054 9148 23060 9150
rect 23124 9148 23130 9212
rect 0 9074 480 9104
rect 8293 9074 8359 9077
rect 0 9072 8359 9074
rect 0 9016 8298 9072
rect 8354 9016 8359 9072
rect 0 9014 8359 9016
rect 0 8984 480 9014
rect 8293 9011 8359 9014
rect 11329 9074 11395 9077
rect 12433 9074 12499 9077
rect 15878 9074 15884 9076
rect 11329 9072 15884 9074
rect 11329 9016 11334 9072
rect 11390 9016 12438 9072
rect 12494 9016 15884 9072
rect 11329 9014 15884 9016
rect 11329 9011 11395 9014
rect 12433 9011 12499 9014
rect 15878 9012 15884 9014
rect 15948 9012 15954 9076
rect 16021 9074 16087 9077
rect 17861 9074 17927 9077
rect 19425 9074 19491 9077
rect 16021 9072 19491 9074
rect 16021 9016 16026 9072
rect 16082 9016 17866 9072
rect 17922 9016 19430 9072
rect 19486 9016 19491 9072
rect 16021 9014 19491 9016
rect 16021 9011 16087 9014
rect 17861 9011 17927 9014
rect 19425 9011 19491 9014
rect 23606 9012 23612 9076
rect 23676 9074 23682 9076
rect 27520 9074 28000 9104
rect 23676 9014 28000 9074
rect 23676 9012 23682 9014
rect 27520 8984 28000 9014
rect 5073 8938 5139 8941
rect 14825 8938 14891 8941
rect 15745 8938 15811 8941
rect 5073 8936 15811 8938
rect 5073 8880 5078 8936
rect 5134 8880 14830 8936
rect 14886 8880 15750 8936
rect 15806 8880 15811 8936
rect 5073 8878 15811 8880
rect 5073 8875 5139 8878
rect 14825 8875 14891 8878
rect 15745 8875 15811 8878
rect 15886 8878 24962 8938
rect 7649 8802 7715 8805
rect 9305 8802 9371 8805
rect 11973 8802 12039 8805
rect 7649 8800 9371 8802
rect 7649 8744 7654 8800
rect 7710 8744 9310 8800
rect 9366 8744 9371 8800
rect 7649 8742 9371 8744
rect 7649 8739 7715 8742
rect 9305 8739 9371 8742
rect 9446 8800 12039 8802
rect 9446 8744 11978 8800
rect 12034 8744 12039 8800
rect 9446 8742 12039 8744
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 7925 8666 7991 8669
rect 9446 8666 9506 8742
rect 11973 8739 12039 8742
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 7925 8664 9506 8666
rect 7925 8608 7930 8664
rect 7986 8608 9506 8664
rect 7925 8606 9506 8608
rect 9581 8666 9647 8669
rect 11145 8668 11211 8669
rect 10910 8666 10916 8668
rect 9581 8664 10916 8666
rect 9581 8608 9586 8664
rect 9642 8608 10916 8664
rect 9581 8606 10916 8608
rect 7925 8603 7991 8606
rect 9581 8603 9647 8606
rect 10910 8604 10916 8606
rect 10980 8604 10986 8668
rect 11094 8604 11100 8668
rect 11164 8666 11211 8668
rect 11164 8664 11256 8666
rect 11206 8608 11256 8664
rect 11164 8606 11256 8608
rect 11164 8604 11211 8606
rect 13854 8604 13860 8668
rect 13924 8666 13930 8668
rect 14181 8666 14247 8669
rect 14641 8666 14707 8669
rect 13924 8664 14707 8666
rect 13924 8608 14186 8664
rect 14242 8608 14646 8664
rect 14702 8608 14707 8664
rect 13924 8606 14707 8608
rect 13924 8604 13930 8606
rect 11145 8603 11211 8604
rect 14181 8603 14247 8606
rect 14641 8603 14707 8606
rect 0 8530 480 8560
rect 3693 8530 3759 8533
rect 0 8528 3759 8530
rect 0 8472 3698 8528
rect 3754 8472 3759 8528
rect 0 8470 3759 8472
rect 0 8440 480 8470
rect 3693 8467 3759 8470
rect 4061 8530 4127 8533
rect 14365 8530 14431 8533
rect 4061 8528 14431 8530
rect 4061 8472 4066 8528
rect 4122 8472 14370 8528
rect 14426 8472 14431 8528
rect 4061 8470 14431 8472
rect 4061 8467 4127 8470
rect 14365 8467 14431 8470
rect 14590 8468 14596 8532
rect 14660 8530 14666 8532
rect 15101 8530 15167 8533
rect 15886 8530 15946 8878
rect 16389 8802 16455 8805
rect 22185 8802 22251 8805
rect 16389 8800 22251 8802
rect 16389 8744 16394 8800
rect 16450 8744 22190 8800
rect 22246 8744 22251 8800
rect 16389 8742 22251 8744
rect 16389 8739 16455 8742
rect 22185 8739 22251 8742
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 17401 8666 17467 8669
rect 20529 8666 20595 8669
rect 22185 8666 22251 8669
rect 17401 8664 22251 8666
rect 17401 8608 17406 8664
rect 17462 8608 20534 8664
rect 20590 8608 22190 8664
rect 22246 8608 22251 8664
rect 17401 8606 22251 8608
rect 17401 8603 17467 8606
rect 20529 8603 20595 8606
rect 22185 8603 22251 8606
rect 14660 8528 15946 8530
rect 14660 8472 15106 8528
rect 15162 8472 15946 8528
rect 14660 8470 15946 8472
rect 23657 8530 23723 8533
rect 24209 8530 24275 8533
rect 23657 8528 24275 8530
rect 23657 8472 23662 8528
rect 23718 8472 24214 8528
rect 24270 8472 24275 8528
rect 23657 8470 24275 8472
rect 24902 8530 24962 8878
rect 25129 8668 25195 8669
rect 25078 8666 25084 8668
rect 25038 8606 25084 8666
rect 25148 8664 25195 8668
rect 25190 8608 25195 8664
rect 25078 8604 25084 8606
rect 25148 8604 25195 8608
rect 25129 8603 25195 8604
rect 27520 8530 28000 8560
rect 24902 8470 28000 8530
rect 14660 8468 14666 8470
rect 15101 8467 15167 8470
rect 23657 8467 23723 8470
rect 24209 8467 24275 8470
rect 27520 8440 28000 8470
rect 1761 8394 1827 8397
rect 2957 8394 3023 8397
rect 1761 8392 3023 8394
rect 1761 8336 1766 8392
rect 1822 8336 2962 8392
rect 3018 8336 3023 8392
rect 1761 8334 3023 8336
rect 1761 8331 1827 8334
rect 2957 8331 3023 8334
rect 7097 8394 7163 8397
rect 8477 8394 8543 8397
rect 9765 8394 9831 8397
rect 7097 8392 9831 8394
rect 7097 8336 7102 8392
rect 7158 8336 8482 8392
rect 8538 8336 9770 8392
rect 9826 8336 9831 8392
rect 7097 8334 9831 8336
rect 7097 8331 7163 8334
rect 8477 8331 8543 8334
rect 9765 8331 9831 8334
rect 9998 8334 10794 8394
rect 5993 8258 6059 8261
rect 6177 8258 6243 8261
rect 9998 8258 10058 8334
rect 5993 8256 10058 8258
rect 5993 8200 5998 8256
rect 6054 8200 6182 8256
rect 6238 8200 10058 8256
rect 5993 8198 10058 8200
rect 10734 8258 10794 8334
rect 19428 8334 20132 8394
rect 10734 8198 14474 8258
rect 5993 8195 6059 8198
rect 6177 8195 6243 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 2865 8122 2931 8125
rect 7649 8122 7715 8125
rect 9213 8124 9279 8125
rect 9213 8122 9260 8124
rect 2865 8120 7715 8122
rect 2865 8064 2870 8120
rect 2926 8064 7654 8120
rect 7710 8064 7715 8120
rect 2865 8062 7715 8064
rect 9168 8120 9260 8122
rect 9168 8064 9218 8120
rect 9168 8062 9260 8064
rect 2865 8059 2931 8062
rect 7649 8059 7715 8062
rect 9213 8060 9260 8062
rect 9324 8060 9330 8124
rect 14273 8122 14339 8125
rect 10734 8120 14339 8122
rect 10734 8064 14278 8120
rect 14334 8064 14339 8120
rect 10734 8062 14339 8064
rect 14414 8122 14474 8198
rect 19428 8122 19488 8334
rect 20072 8258 20132 8334
rect 21725 8392 21791 8397
rect 21725 8336 21730 8392
rect 21786 8336 21791 8392
rect 21725 8331 21791 8336
rect 21728 8258 21788 8331
rect 20072 8198 21788 8258
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 14414 8062 19488 8122
rect 20345 8122 20411 8125
rect 20345 8120 21052 8122
rect 20345 8064 20350 8120
rect 20406 8064 21052 8120
rect 20345 8062 21052 8064
rect 9213 8059 9279 8060
rect 3141 7986 3207 7989
rect 6637 7986 6703 7989
rect 3141 7984 6703 7986
rect 3141 7928 3146 7984
rect 3202 7928 6642 7984
rect 6698 7928 6703 7984
rect 3141 7926 6703 7928
rect 3141 7923 3207 7926
rect 6637 7923 6703 7926
rect 6913 7986 6979 7989
rect 10734 7986 10794 8062
rect 14273 8059 14339 8062
rect 20345 8059 20411 8062
rect 15929 7986 15995 7989
rect 6913 7984 10794 7986
rect 6913 7928 6918 7984
rect 6974 7928 10794 7984
rect 6913 7926 10794 7928
rect 10918 7984 15995 7986
rect 10918 7928 15934 7984
rect 15990 7928 15995 7984
rect 10918 7926 15995 7928
rect 6913 7923 6979 7926
rect 0 7850 480 7880
rect 2865 7850 2931 7853
rect 0 7848 2931 7850
rect 0 7792 2870 7848
rect 2926 7792 2931 7848
rect 0 7790 2931 7792
rect 0 7760 480 7790
rect 2865 7787 2931 7790
rect 4061 7850 4127 7853
rect 4286 7850 4292 7852
rect 4061 7848 4292 7850
rect 4061 7792 4066 7848
rect 4122 7792 4292 7848
rect 4061 7790 4292 7792
rect 4061 7787 4127 7790
rect 4286 7788 4292 7790
rect 4356 7850 4362 7852
rect 4429 7850 4495 7853
rect 4356 7848 4495 7850
rect 4356 7792 4434 7848
rect 4490 7792 4495 7848
rect 4356 7790 4495 7792
rect 4356 7788 4362 7790
rect 4429 7787 4495 7790
rect 4889 7850 4955 7853
rect 7005 7850 7071 7853
rect 4889 7848 7071 7850
rect 4889 7792 4894 7848
rect 4950 7792 7010 7848
rect 7066 7792 7071 7848
rect 4889 7790 7071 7792
rect 4889 7787 4955 7790
rect 7005 7787 7071 7790
rect 9213 7850 9279 7853
rect 9673 7850 9739 7853
rect 9213 7848 9739 7850
rect 9213 7792 9218 7848
rect 9274 7792 9678 7848
rect 9734 7792 9739 7848
rect 9213 7790 9739 7792
rect 9213 7787 9279 7790
rect 9673 7787 9739 7790
rect 9857 7850 9923 7853
rect 10918 7850 10978 7926
rect 15929 7923 15995 7926
rect 17125 7986 17191 7989
rect 20805 7986 20871 7989
rect 17125 7984 20871 7986
rect 17125 7928 17130 7984
rect 17186 7928 20810 7984
rect 20866 7928 20871 7984
rect 17125 7926 20871 7928
rect 20992 7986 21052 8062
rect 21398 8060 21404 8124
rect 21468 8122 21474 8124
rect 22829 8122 22895 8125
rect 21468 8120 22895 8122
rect 21468 8064 22834 8120
rect 22890 8064 22895 8120
rect 21468 8062 22895 8064
rect 21468 8060 21474 8062
rect 22829 8059 22895 8062
rect 24209 7986 24275 7989
rect 20992 7984 24275 7986
rect 20992 7928 24214 7984
rect 24270 7928 24275 7984
rect 20992 7926 24275 7928
rect 17125 7923 17191 7926
rect 20805 7923 20871 7926
rect 24209 7923 24275 7926
rect 9857 7848 10978 7850
rect 9857 7792 9862 7848
rect 9918 7792 10978 7848
rect 9857 7790 10978 7792
rect 11697 7850 11763 7853
rect 15101 7850 15167 7853
rect 11697 7848 15167 7850
rect 11697 7792 11702 7848
rect 11758 7792 15106 7848
rect 15162 7792 15167 7848
rect 11697 7790 15167 7792
rect 9857 7787 9923 7790
rect 11697 7787 11763 7790
rect 15101 7787 15167 7790
rect 15285 7850 15351 7853
rect 17401 7850 17467 7853
rect 20805 7850 20871 7853
rect 24025 7850 24091 7853
rect 27520 7850 28000 7880
rect 15285 7848 15394 7850
rect 15285 7792 15290 7848
rect 15346 7792 15394 7848
rect 15285 7787 15394 7792
rect 17401 7848 20871 7850
rect 17401 7792 17406 7848
rect 17462 7792 20810 7848
rect 20866 7792 20871 7848
rect 17401 7790 20871 7792
rect 17401 7787 17467 7790
rect 20805 7787 20871 7790
rect 21912 7848 24091 7850
rect 21912 7792 24030 7848
rect 24086 7792 24091 7848
rect 21912 7790 24091 7792
rect 6637 7714 6703 7717
rect 10041 7714 10107 7717
rect 6637 7712 10107 7714
rect 6637 7656 6642 7712
rect 6698 7656 10046 7712
rect 10102 7656 10107 7712
rect 6637 7654 10107 7656
rect 6637 7651 6703 7654
rect 10041 7651 10107 7654
rect 10777 7714 10843 7717
rect 12617 7714 12683 7717
rect 10777 7712 12683 7714
rect 10777 7656 10782 7712
rect 10838 7656 12622 7712
rect 12678 7656 12683 7712
rect 10777 7654 12683 7656
rect 15334 7714 15394 7787
rect 17718 7714 17724 7716
rect 15334 7654 17724 7714
rect 10777 7651 10843 7654
rect 12617 7651 12683 7654
rect 17718 7652 17724 7654
rect 17788 7714 17794 7716
rect 21912 7714 21972 7790
rect 24025 7787 24091 7790
rect 24902 7790 28000 7850
rect 17788 7654 21972 7714
rect 17788 7652 17794 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 5993 7578 6059 7581
rect 7281 7578 7347 7581
rect 11053 7578 11119 7581
rect 16021 7580 16087 7581
rect 16021 7578 16068 7580
rect 5993 7576 11119 7578
rect 5993 7520 5998 7576
rect 6054 7520 7286 7576
rect 7342 7520 11058 7576
rect 11114 7520 11119 7576
rect 5993 7518 11119 7520
rect 15976 7576 16068 7578
rect 15976 7520 16026 7576
rect 15976 7518 16068 7520
rect 5993 7515 6059 7518
rect 7281 7515 7347 7518
rect 11053 7515 11119 7518
rect 16021 7516 16068 7518
rect 16132 7516 16138 7580
rect 16205 7578 16271 7581
rect 20345 7578 20411 7581
rect 16205 7576 20411 7578
rect 16205 7520 16210 7576
rect 16266 7520 20350 7576
rect 20406 7520 20411 7576
rect 16205 7518 20411 7520
rect 16021 7515 16087 7516
rect 16205 7515 16271 7518
rect 20345 7515 20411 7518
rect 21582 7516 21588 7580
rect 21652 7578 21658 7580
rect 22001 7578 22067 7581
rect 21652 7576 22067 7578
rect 21652 7520 22006 7576
rect 22062 7520 22067 7576
rect 21652 7518 22067 7520
rect 21652 7516 21658 7518
rect 22001 7515 22067 7518
rect 7005 7442 7071 7445
rect 11053 7442 11119 7445
rect 24902 7442 24962 7790
rect 27520 7760 28000 7790
rect 7005 7440 10978 7442
rect 7005 7384 7010 7440
rect 7066 7384 10978 7440
rect 7005 7382 10978 7384
rect 7005 7379 7071 7382
rect 0 7306 480 7336
rect 10918 7306 10978 7382
rect 11053 7440 24962 7442
rect 11053 7384 11058 7440
rect 11114 7384 24962 7440
rect 11053 7382 24962 7384
rect 11053 7379 11119 7382
rect 15469 7306 15535 7309
rect 0 7246 10794 7306
rect 10918 7304 15535 7306
rect 10918 7248 15474 7304
rect 15530 7248 15535 7304
rect 10918 7246 15535 7248
rect 0 7216 480 7246
rect 3969 7170 4035 7173
rect 9857 7170 9923 7173
rect 3969 7168 9923 7170
rect 3969 7112 3974 7168
rect 4030 7112 9862 7168
rect 9918 7112 9923 7168
rect 3969 7110 9923 7112
rect 3969 7107 4035 7110
rect 9857 7107 9923 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 10734 7034 10794 7246
rect 15469 7243 15535 7246
rect 15653 7306 15719 7309
rect 16021 7306 16087 7309
rect 15653 7304 16087 7306
rect 15653 7248 15658 7304
rect 15714 7248 16026 7304
rect 16082 7248 16087 7304
rect 15653 7246 16087 7248
rect 15653 7243 15719 7246
rect 16021 7243 16087 7246
rect 16757 7306 16823 7309
rect 24209 7306 24275 7309
rect 27520 7306 28000 7336
rect 16757 7304 24042 7306
rect 16757 7248 16762 7304
rect 16818 7248 24042 7304
rect 16757 7246 24042 7248
rect 16757 7243 16823 7246
rect 11094 7108 11100 7172
rect 11164 7170 11170 7172
rect 17861 7170 17927 7173
rect 23473 7172 23539 7173
rect 11164 7168 17927 7170
rect 11164 7112 17866 7168
rect 17922 7112 17927 7168
rect 11164 7110 17927 7112
rect 11164 7108 11170 7110
rect 17861 7107 17927 7110
rect 23422 7108 23428 7172
rect 23492 7170 23539 7172
rect 23982 7170 24042 7246
rect 24209 7304 28000 7306
rect 24209 7248 24214 7304
rect 24270 7248 28000 7304
rect 24209 7246 28000 7248
rect 24209 7243 24275 7246
rect 27520 7216 28000 7246
rect 25129 7170 25195 7173
rect 23492 7168 23584 7170
rect 23534 7112 23584 7168
rect 23492 7110 23584 7112
rect 23982 7168 25195 7170
rect 23982 7112 25134 7168
rect 25190 7112 25195 7168
rect 23982 7110 25195 7112
rect 23492 7108 23539 7110
rect 23473 7107 23539 7108
rect 25129 7107 25195 7110
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 13629 7034 13695 7037
rect 10734 7032 13695 7034
rect 10734 6976 13634 7032
rect 13690 6976 13695 7032
rect 10734 6974 13695 6976
rect 13629 6971 13695 6974
rect 14365 7034 14431 7037
rect 16849 7034 16915 7037
rect 17534 7034 17540 7036
rect 14365 7032 15532 7034
rect 14365 6976 14370 7032
rect 14426 6976 15532 7032
rect 14365 6974 15532 6976
rect 14365 6971 14431 6974
rect 5625 6898 5691 6901
rect 6361 6898 6427 6901
rect 15285 6898 15351 6901
rect 5625 6896 15351 6898
rect 5625 6840 5630 6896
rect 5686 6840 6366 6896
rect 6422 6840 15290 6896
rect 15346 6840 15351 6896
rect 5625 6838 15351 6840
rect 15472 6898 15532 6974
rect 16849 7032 17540 7034
rect 16849 6976 16854 7032
rect 16910 6976 17540 7032
rect 16849 6974 17540 6976
rect 16849 6971 16915 6974
rect 17534 6972 17540 6974
rect 17604 6972 17610 7036
rect 17902 6898 17908 6900
rect 15472 6838 17908 6898
rect 5625 6835 5691 6838
rect 6361 6835 6427 6838
rect 15285 6835 15351 6838
rect 17902 6836 17908 6838
rect 17972 6836 17978 6900
rect 19425 6898 19491 6901
rect 22461 6898 22527 6901
rect 19425 6896 22527 6898
rect 19425 6840 19430 6896
rect 19486 6840 22466 6896
rect 22522 6840 22527 6896
rect 19425 6838 22527 6840
rect 19425 6835 19491 6838
rect 22461 6835 22527 6838
rect 23790 6836 23796 6900
rect 23860 6898 23866 6900
rect 23860 6838 24410 6898
rect 23860 6836 23866 6838
rect 0 6762 480 6792
rect 3550 6762 3556 6764
rect 0 6702 3556 6762
rect 0 6672 480 6702
rect 3550 6700 3556 6702
rect 3620 6700 3626 6764
rect 7557 6762 7623 6765
rect 10133 6762 10199 6765
rect 10726 6762 10732 6764
rect 7557 6760 8770 6762
rect 7557 6704 7562 6760
rect 7618 6704 8770 6760
rect 7557 6702 8770 6704
rect 7557 6699 7623 6702
rect 6821 6626 6887 6629
rect 7741 6626 7807 6629
rect 8477 6626 8543 6629
rect 6821 6624 8543 6626
rect 6821 6568 6826 6624
rect 6882 6568 7746 6624
rect 7802 6568 8482 6624
rect 8538 6568 8543 6624
rect 6821 6566 8543 6568
rect 8710 6626 8770 6702
rect 10133 6760 10732 6762
rect 10133 6704 10138 6760
rect 10194 6704 10732 6760
rect 10133 6702 10732 6704
rect 10133 6699 10199 6702
rect 10726 6700 10732 6702
rect 10796 6700 10802 6764
rect 15326 6762 15332 6764
rect 14782 6702 15332 6762
rect 14641 6626 14707 6629
rect 8710 6624 14707 6626
rect 8710 6568 14646 6624
rect 14702 6568 14707 6624
rect 8710 6566 14707 6568
rect 6821 6563 6887 6566
rect 7741 6563 7807 6566
rect 8477 6563 8543 6566
rect 14641 6563 14707 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 11513 6490 11579 6493
rect 12382 6490 12388 6492
rect 11513 6488 12388 6490
rect 11513 6432 11518 6488
rect 11574 6432 12388 6488
rect 11513 6430 12388 6432
rect 11513 6427 11579 6430
rect 12382 6428 12388 6430
rect 12452 6428 12458 6492
rect 14406 6490 14412 6492
rect 12528 6430 14412 6490
rect 11646 6292 11652 6356
rect 11716 6354 11722 6356
rect 12528 6354 12588 6430
rect 14406 6428 14412 6430
rect 14476 6490 14482 6492
rect 14782 6490 14842 6702
rect 15326 6700 15332 6702
rect 15396 6700 15402 6764
rect 16297 6762 16363 6765
rect 17033 6762 17099 6765
rect 16297 6760 17099 6762
rect 16297 6704 16302 6760
rect 16358 6704 17038 6760
rect 17094 6704 17099 6760
rect 16297 6702 17099 6704
rect 16297 6699 16363 6702
rect 17033 6699 17099 6702
rect 17217 6762 17283 6765
rect 19517 6762 19583 6765
rect 24025 6764 24091 6765
rect 17217 6760 19583 6762
rect 17217 6704 17222 6760
rect 17278 6704 19522 6760
rect 19578 6704 19583 6760
rect 17217 6702 19583 6704
rect 17217 6699 17283 6702
rect 19517 6699 19583 6702
rect 23974 6700 23980 6764
rect 24044 6762 24091 6764
rect 24350 6762 24410 6838
rect 27520 6762 28000 6792
rect 24044 6760 24136 6762
rect 24086 6704 24136 6760
rect 24044 6702 24136 6704
rect 24350 6702 28000 6762
rect 24044 6700 24091 6702
rect 24025 6699 24091 6700
rect 27520 6672 28000 6702
rect 17401 6626 17467 6629
rect 21357 6626 21423 6629
rect 17401 6624 21423 6626
rect 17401 6568 17406 6624
rect 17462 6568 21362 6624
rect 21418 6568 21423 6624
rect 17401 6566 21423 6568
rect 17401 6563 17467 6566
rect 21357 6563 21423 6566
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 14476 6430 14842 6490
rect 19149 6490 19215 6493
rect 21909 6490 21975 6493
rect 19149 6488 21975 6490
rect 19149 6432 19154 6488
rect 19210 6432 21914 6488
rect 21970 6432 21975 6488
rect 19149 6430 21975 6432
rect 14476 6428 14482 6430
rect 19149 6427 19215 6430
rect 21909 6427 21975 6430
rect 11716 6294 12588 6354
rect 15653 6354 15719 6357
rect 20805 6354 20871 6357
rect 15653 6352 20871 6354
rect 15653 6296 15658 6352
rect 15714 6296 20810 6352
rect 20866 6296 20871 6352
rect 15653 6294 20871 6296
rect 11716 6292 11722 6294
rect 15653 6291 15719 6294
rect 20805 6291 20871 6294
rect 7189 6218 7255 6221
rect 15561 6218 15627 6221
rect 7189 6216 15627 6218
rect 7189 6160 7194 6216
rect 7250 6160 15566 6216
rect 15622 6160 15627 6216
rect 7189 6158 15627 6160
rect 7189 6155 7255 6158
rect 15561 6155 15627 6158
rect 18321 6218 18387 6221
rect 23473 6218 23539 6221
rect 18321 6216 23539 6218
rect 18321 6160 18326 6216
rect 18382 6160 23478 6216
rect 23534 6160 23539 6216
rect 18321 6158 23539 6160
rect 18321 6155 18387 6158
rect 23473 6155 23539 6158
rect 0 6082 480 6112
rect 3877 6082 3943 6085
rect 12065 6084 12131 6085
rect 0 6080 3943 6082
rect 0 6024 3882 6080
rect 3938 6024 3943 6080
rect 0 6022 3943 6024
rect 0 5992 480 6022
rect 3877 6019 3943 6022
rect 12014 6020 12020 6084
rect 12084 6082 12131 6084
rect 12985 6082 13051 6085
rect 15929 6082 15995 6085
rect 12084 6080 12176 6082
rect 12126 6024 12176 6080
rect 12084 6022 12176 6024
rect 12985 6080 15995 6082
rect 12985 6024 12990 6080
rect 13046 6024 15934 6080
rect 15990 6024 15995 6080
rect 12985 6022 15995 6024
rect 12084 6020 12131 6022
rect 12065 6019 12131 6020
rect 12985 6019 13051 6022
rect 15929 6019 15995 6022
rect 20662 6020 20668 6084
rect 20732 6082 20738 6084
rect 24025 6082 24091 6085
rect 20732 6080 24091 6082
rect 20732 6024 24030 6080
rect 24086 6024 24091 6080
rect 20732 6022 24091 6024
rect 20732 6020 20738 6022
rect 24025 6019 24091 6022
rect 25957 6082 26023 6085
rect 27520 6082 28000 6112
rect 25957 6080 28000 6082
rect 25957 6024 25962 6080
rect 26018 6024 28000 6080
rect 25957 6022 28000 6024
rect 25957 6019 26023 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 27520 5992 28000 6022
rect 19610 5951 19930 5952
rect 8017 5946 8083 5949
rect 10041 5946 10107 5949
rect 8017 5944 10107 5946
rect 8017 5888 8022 5944
rect 8078 5888 10046 5944
rect 10102 5888 10107 5944
rect 8017 5886 10107 5888
rect 8017 5883 8083 5886
rect 10041 5883 10107 5886
rect 11094 5884 11100 5948
rect 11164 5946 11170 5948
rect 14590 5946 14596 5948
rect 11164 5886 14596 5946
rect 11164 5884 11170 5886
rect 14590 5884 14596 5886
rect 14660 5884 14666 5948
rect 20437 5946 20503 5949
rect 23197 5946 23263 5949
rect 20437 5944 23263 5946
rect 20437 5888 20442 5944
rect 20498 5888 23202 5944
rect 23258 5888 23263 5944
rect 20437 5886 23263 5888
rect 20437 5883 20503 5886
rect 23197 5883 23263 5886
rect 7557 5810 7623 5813
rect 12893 5810 12959 5813
rect 7557 5808 12959 5810
rect 7557 5752 7562 5808
rect 7618 5752 12898 5808
rect 12954 5752 12959 5808
rect 7557 5750 12959 5752
rect 7557 5747 7623 5750
rect 12893 5747 12959 5750
rect 13169 5810 13235 5813
rect 15285 5810 15351 5813
rect 23473 5810 23539 5813
rect 13169 5808 23539 5810
rect 13169 5752 13174 5808
rect 13230 5752 15290 5808
rect 15346 5752 23478 5808
rect 23534 5752 23539 5808
rect 13169 5750 23539 5752
rect 13169 5747 13235 5750
rect 15285 5747 15351 5750
rect 23473 5747 23539 5750
rect 8017 5674 8083 5677
rect 10685 5674 10751 5677
rect 8017 5672 10751 5674
rect 8017 5616 8022 5672
rect 8078 5616 10690 5672
rect 10746 5616 10751 5672
rect 8017 5614 10751 5616
rect 8017 5611 8083 5614
rect 10685 5611 10751 5614
rect 12801 5674 12867 5677
rect 18965 5674 19031 5677
rect 21173 5674 21239 5677
rect 12801 5672 15394 5674
rect 12801 5616 12806 5672
rect 12862 5616 15394 5672
rect 12801 5614 15394 5616
rect 12801 5611 12867 5614
rect 0 5538 480 5568
rect 3509 5538 3575 5541
rect 0 5536 3575 5538
rect 0 5480 3514 5536
rect 3570 5480 3575 5536
rect 0 5478 3575 5480
rect 0 5448 480 5478
rect 3509 5475 3575 5478
rect 7925 5538 7991 5541
rect 11237 5538 11303 5541
rect 7925 5536 11303 5538
rect 7925 5480 7930 5536
rect 7986 5480 11242 5536
rect 11298 5480 11303 5536
rect 7925 5478 11303 5480
rect 7925 5475 7991 5478
rect 11237 5475 11303 5478
rect 11697 5538 11763 5541
rect 13721 5538 13787 5541
rect 11697 5536 13787 5538
rect 11697 5480 11702 5536
rect 11758 5480 13726 5536
rect 13782 5480 13787 5536
rect 11697 5478 13787 5480
rect 11697 5475 11763 5478
rect 13721 5475 13787 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 7281 5402 7347 5405
rect 12617 5402 12683 5405
rect 7281 5400 12683 5402
rect 7281 5344 7286 5400
rect 7342 5344 12622 5400
rect 12678 5344 12683 5400
rect 7281 5342 12683 5344
rect 15334 5402 15394 5614
rect 18965 5672 21239 5674
rect 18965 5616 18970 5672
rect 19026 5616 21178 5672
rect 21234 5616 21239 5672
rect 18965 5614 21239 5616
rect 18965 5611 19031 5614
rect 21173 5611 21239 5614
rect 24209 5674 24275 5677
rect 25221 5674 25287 5677
rect 24209 5672 25287 5674
rect 24209 5616 24214 5672
rect 24270 5616 25226 5672
rect 25282 5616 25287 5672
rect 24209 5614 25287 5616
rect 24209 5611 24275 5614
rect 25221 5611 25287 5614
rect 24761 5538 24827 5541
rect 27520 5538 28000 5568
rect 24761 5536 28000 5538
rect 24761 5480 24766 5536
rect 24822 5480 28000 5536
rect 24761 5478 28000 5480
rect 24761 5475 24827 5478
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 27520 5448 28000 5478
rect 24277 5407 24597 5408
rect 24117 5402 24183 5405
rect 15334 5400 24183 5402
rect 15334 5344 24122 5400
rect 24178 5344 24183 5400
rect 15334 5342 24183 5344
rect 7281 5339 7347 5342
rect 12617 5339 12683 5342
rect 24117 5339 24183 5342
rect 12985 5266 13051 5269
rect 4892 5264 13051 5266
rect 4892 5208 12990 5264
rect 13046 5208 13051 5264
rect 4892 5206 13051 5208
rect 0 4994 480 5024
rect 4892 4994 4952 5206
rect 12985 5203 13051 5206
rect 17033 5266 17099 5269
rect 20345 5266 20411 5269
rect 21449 5266 21515 5269
rect 17033 5264 21515 5266
rect 17033 5208 17038 5264
rect 17094 5208 20350 5264
rect 20406 5208 21454 5264
rect 21510 5208 21515 5264
rect 17033 5206 21515 5208
rect 17033 5203 17099 5206
rect 20345 5203 20411 5206
rect 21449 5203 21515 5206
rect 23422 5204 23428 5268
rect 23492 5266 23498 5268
rect 24710 5266 24716 5268
rect 23492 5206 24716 5266
rect 23492 5204 23498 5206
rect 24710 5204 24716 5206
rect 24780 5204 24786 5268
rect 9949 5130 10015 5133
rect 12617 5130 12683 5133
rect 25957 5130 26023 5133
rect 9949 5128 11898 5130
rect 9949 5072 9954 5128
rect 10010 5072 11898 5128
rect 9949 5070 11898 5072
rect 9949 5067 10015 5070
rect 0 4934 4952 4994
rect 0 4904 480 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 11838 4861 11898 5070
rect 12617 5128 26023 5130
rect 12617 5072 12622 5128
rect 12678 5072 25962 5128
rect 26018 5072 26023 5128
rect 12617 5070 26023 5072
rect 12617 5067 12683 5070
rect 25957 5067 26023 5070
rect 11973 4994 12039 4997
rect 13353 4994 13419 4997
rect 11973 4992 13419 4994
rect 11973 4936 11978 4992
rect 12034 4936 13358 4992
rect 13414 4936 13419 4992
rect 11973 4934 13419 4936
rect 11973 4931 12039 4934
rect 13353 4931 13419 4934
rect 14774 4932 14780 4996
rect 14844 4994 14850 4996
rect 15009 4994 15075 4997
rect 14844 4992 15075 4994
rect 14844 4936 15014 4992
rect 15070 4936 15075 4992
rect 14844 4934 15075 4936
rect 14844 4932 14850 4934
rect 15009 4931 15075 4934
rect 24301 4994 24367 4997
rect 27520 4994 28000 5024
rect 24301 4992 28000 4994
rect 24301 4936 24306 4992
rect 24362 4936 28000 4992
rect 24301 4934 28000 4936
rect 24301 4931 24367 4934
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 27520 4904 28000 4934
rect 19610 4863 19930 4864
rect 11789 4858 11898 4861
rect 13537 4858 13603 4861
rect 14641 4858 14707 4861
rect 15653 4858 15719 4861
rect 11708 4856 13370 4858
rect 11708 4800 11794 4856
rect 11850 4800 13370 4856
rect 11708 4798 13370 4800
rect 11789 4795 11855 4798
rect 6821 4722 6887 4725
rect 12985 4722 13051 4725
rect 6821 4720 13051 4722
rect 6821 4664 6826 4720
rect 6882 4664 12990 4720
rect 13046 4664 13051 4720
rect 6821 4662 13051 4664
rect 13310 4722 13370 4798
rect 13537 4856 15719 4858
rect 13537 4800 13542 4856
rect 13598 4800 14646 4856
rect 14702 4800 15658 4856
rect 15714 4800 15719 4856
rect 13537 4798 15719 4800
rect 13537 4795 13603 4798
rect 14641 4795 14707 4798
rect 15653 4795 15719 4798
rect 17401 4722 17467 4725
rect 13310 4720 17467 4722
rect 13310 4664 17406 4720
rect 17462 4664 17467 4720
rect 13310 4662 17467 4664
rect 6821 4659 6887 4662
rect 12985 4659 13051 4662
rect 17401 4659 17467 4662
rect 17769 4722 17835 4725
rect 23657 4722 23723 4725
rect 17769 4720 23723 4722
rect 17769 4664 17774 4720
rect 17830 4664 23662 4720
rect 23718 4664 23723 4720
rect 17769 4662 23723 4664
rect 17769 4659 17835 4662
rect 23657 4659 23723 4662
rect 5257 4586 5323 4589
rect 8661 4588 8727 4589
rect 8661 4586 8708 4588
rect 5257 4584 6148 4586
rect 5257 4528 5262 4584
rect 5318 4528 6148 4584
rect 5257 4526 6148 4528
rect 8616 4584 8708 4586
rect 8616 4528 8666 4584
rect 8616 4526 8708 4528
rect 5257 4523 5323 4526
rect 0 4450 480 4480
rect 1669 4450 1735 4453
rect 0 4448 1735 4450
rect 0 4392 1674 4448
rect 1730 4392 1735 4448
rect 0 4390 1735 4392
rect 6088 4450 6148 4526
rect 8661 4524 8708 4526
rect 8772 4524 8778 4588
rect 13629 4586 13695 4589
rect 8894 4584 13695 4586
rect 8894 4528 13634 4584
rect 13690 4528 13695 4584
rect 8894 4526 13695 4528
rect 8661 4523 8727 4524
rect 8894 4450 8954 4526
rect 13629 4523 13695 4526
rect 14089 4586 14155 4589
rect 18045 4586 18111 4589
rect 14089 4584 18111 4586
rect 14089 4528 14094 4584
rect 14150 4528 18050 4584
rect 18106 4528 18111 4584
rect 14089 4526 18111 4528
rect 14089 4523 14155 4526
rect 18045 4523 18111 4526
rect 19977 4586 20043 4589
rect 23422 4586 23428 4588
rect 19977 4584 23428 4586
rect 19977 4528 19982 4584
rect 20038 4528 23428 4584
rect 19977 4526 23428 4528
rect 19977 4523 20043 4526
rect 23422 4524 23428 4526
rect 23492 4524 23498 4588
rect 6088 4390 8954 4450
rect 21173 4450 21239 4453
rect 23657 4450 23723 4453
rect 21173 4448 23723 4450
rect 21173 4392 21178 4448
rect 21234 4392 23662 4448
rect 23718 4392 23723 4448
rect 21173 4390 23723 4392
rect 0 4360 480 4390
rect 1669 4387 1735 4390
rect 21173 4387 21239 4390
rect 23657 4387 23723 4390
rect 25037 4450 25103 4453
rect 27520 4450 28000 4480
rect 25037 4448 28000 4450
rect 25037 4392 25042 4448
rect 25098 4392 28000 4448
rect 25037 4390 28000 4392
rect 25037 4387 25103 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 27520 4360 28000 4390
rect 24277 4319 24597 4320
rect 11789 4314 11855 4317
rect 12249 4314 12315 4317
rect 11789 4312 12315 4314
rect 11789 4256 11794 4312
rect 11850 4256 12254 4312
rect 12310 4256 12315 4312
rect 11789 4254 12315 4256
rect 11789 4251 11855 4254
rect 12249 4251 12315 4254
rect 21214 4252 21220 4316
rect 21284 4314 21290 4316
rect 24117 4314 24183 4317
rect 21284 4312 24183 4314
rect 21284 4256 24122 4312
rect 24178 4256 24183 4312
rect 21284 4254 24183 4256
rect 21284 4252 21290 4254
rect 24117 4251 24183 4254
rect 9581 4178 9647 4181
rect 11329 4178 11395 4181
rect 9581 4176 11395 4178
rect 9581 4120 9586 4176
rect 9642 4120 11334 4176
rect 11390 4120 11395 4176
rect 9581 4118 11395 4120
rect 9581 4115 9647 4118
rect 11329 4115 11395 4118
rect 13353 4178 13419 4181
rect 17309 4178 17375 4181
rect 13353 4176 17375 4178
rect 13353 4120 13358 4176
rect 13414 4120 17314 4176
rect 17370 4120 17375 4176
rect 13353 4118 17375 4120
rect 13353 4115 13419 4118
rect 17309 4115 17375 4118
rect 18137 4178 18203 4181
rect 22093 4178 22159 4181
rect 18137 4176 22159 4178
rect 18137 4120 18142 4176
rect 18198 4120 22098 4176
rect 22154 4120 22159 4176
rect 18137 4118 22159 4120
rect 18137 4115 18203 4118
rect 22093 4115 22159 4118
rect 25681 4178 25747 4181
rect 27613 4178 27679 4181
rect 25681 4176 27679 4178
rect 25681 4120 25686 4176
rect 25742 4120 27618 4176
rect 27674 4120 27679 4176
rect 25681 4118 27679 4120
rect 25681 4115 25747 4118
rect 27613 4115 27679 4118
rect 5533 4042 5599 4045
rect 12433 4042 12499 4045
rect 5533 4040 12499 4042
rect 5533 3984 5538 4040
rect 5594 3984 12438 4040
rect 12494 3984 12499 4040
rect 5533 3982 12499 3984
rect 5533 3979 5599 3982
rect 12433 3979 12499 3982
rect 13537 4042 13603 4045
rect 17401 4042 17467 4045
rect 13537 4040 17467 4042
rect 13537 3984 13542 4040
rect 13598 3984 17406 4040
rect 17462 3984 17467 4040
rect 13537 3982 17467 3984
rect 13537 3979 13603 3982
rect 17401 3979 17467 3982
rect 17585 4042 17651 4045
rect 20437 4042 20503 4045
rect 17585 4040 20503 4042
rect 17585 3984 17590 4040
rect 17646 3984 20442 4040
rect 20498 3984 20503 4040
rect 17585 3982 20503 3984
rect 17585 3979 17651 3982
rect 20437 3979 20503 3982
rect 20897 4042 20963 4045
rect 26325 4042 26391 4045
rect 20897 4040 26391 4042
rect 20897 3984 20902 4040
rect 20958 3984 26330 4040
rect 26386 3984 26391 4040
rect 20897 3982 26391 3984
rect 20897 3979 20963 3982
rect 26325 3979 26391 3982
rect 1853 3906 1919 3909
rect 10041 3906 10107 3909
rect 19425 3906 19491 3909
rect 1853 3904 10107 3906
rect 1853 3848 1858 3904
rect 1914 3848 10046 3904
rect 10102 3848 10107 3904
rect 1853 3846 10107 3848
rect 1853 3843 1919 3846
rect 10041 3843 10107 3846
rect 18094 3904 19491 3906
rect 18094 3848 19430 3904
rect 19486 3848 19491 3904
rect 18094 3846 19491 3848
rect 10277 3840 10597 3841
rect 0 3770 480 3800
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 1761 3770 1827 3773
rect 0 3768 1827 3770
rect 0 3712 1766 3768
rect 1822 3712 1827 3768
rect 0 3710 1827 3712
rect 0 3680 480 3710
rect 1761 3707 1827 3710
rect 3918 3708 3924 3772
rect 3988 3770 3994 3772
rect 4061 3770 4127 3773
rect 9857 3770 9923 3773
rect 3988 3768 4127 3770
rect 3988 3712 4066 3768
rect 4122 3712 4127 3768
rect 3988 3710 4127 3712
rect 3988 3708 3994 3710
rect 4061 3707 4127 3710
rect 4248 3768 9923 3770
rect 4248 3712 9862 3768
rect 9918 3712 9923 3768
rect 4248 3710 9923 3712
rect 1209 3634 1275 3637
rect 4248 3634 4308 3710
rect 9857 3707 9923 3710
rect 11513 3770 11579 3773
rect 11830 3770 11836 3772
rect 11513 3768 11836 3770
rect 11513 3712 11518 3768
rect 11574 3712 11836 3768
rect 11513 3710 11836 3712
rect 11513 3707 11579 3710
rect 11830 3708 11836 3710
rect 11900 3708 11906 3772
rect 14549 3770 14615 3773
rect 18094 3770 18154 3846
rect 19425 3843 19491 3846
rect 23054 3844 23060 3908
rect 23124 3906 23130 3908
rect 23124 3846 24732 3906
rect 23124 3844 23130 3846
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 14549 3768 18154 3770
rect 14549 3712 14554 3768
rect 14610 3712 18154 3768
rect 14549 3710 18154 3712
rect 18229 3770 18295 3773
rect 19333 3770 19399 3773
rect 18229 3768 19399 3770
rect 18229 3712 18234 3768
rect 18290 3712 19338 3768
rect 19394 3712 19399 3768
rect 18229 3710 19399 3712
rect 14549 3707 14615 3710
rect 18229 3707 18295 3710
rect 19333 3707 19399 3710
rect 23974 3708 23980 3772
rect 24044 3770 24050 3772
rect 24485 3770 24551 3773
rect 24044 3768 24551 3770
rect 24044 3712 24490 3768
rect 24546 3712 24551 3768
rect 24044 3710 24551 3712
rect 24672 3770 24732 3846
rect 27520 3770 28000 3800
rect 24672 3710 28000 3770
rect 24044 3708 24050 3710
rect 24485 3707 24551 3710
rect 27520 3680 28000 3710
rect 1209 3632 4308 3634
rect 1209 3576 1214 3632
rect 1270 3576 4308 3632
rect 1209 3574 4308 3576
rect 1209 3571 1275 3574
rect 9622 3572 9628 3636
rect 9692 3634 9698 3636
rect 17769 3634 17835 3637
rect 9692 3632 17835 3634
rect 9692 3576 17774 3632
rect 17830 3576 17835 3632
rect 9692 3574 17835 3576
rect 9692 3572 9698 3574
rect 17769 3571 17835 3574
rect 18689 3634 18755 3637
rect 22921 3634 22987 3637
rect 25037 3634 25103 3637
rect 18689 3632 21052 3634
rect 18689 3576 18694 3632
rect 18750 3576 21052 3632
rect 18689 3574 21052 3576
rect 18689 3571 18755 3574
rect 20992 3501 21052 3574
rect 22921 3632 25103 3634
rect 22921 3576 22926 3632
rect 22982 3576 25042 3632
rect 25098 3576 25103 3632
rect 22921 3574 25103 3576
rect 22921 3571 22987 3574
rect 25037 3571 25103 3574
rect 3785 3498 3851 3501
rect 7281 3498 7347 3501
rect 13537 3498 13603 3501
rect 16389 3498 16455 3501
rect 16849 3498 16915 3501
rect 3785 3496 16915 3498
rect 3785 3440 3790 3496
rect 3846 3440 7286 3496
rect 7342 3440 13542 3496
rect 13598 3440 16394 3496
rect 16450 3440 16854 3496
rect 16910 3440 16915 3496
rect 3785 3438 16915 3440
rect 3785 3435 3851 3438
rect 7281 3435 7347 3438
rect 13537 3435 13603 3438
rect 16389 3435 16455 3438
rect 16849 3435 16915 3438
rect 17033 3498 17099 3501
rect 18689 3498 18755 3501
rect 17033 3496 18755 3498
rect 17033 3440 17038 3496
rect 17094 3440 18694 3496
rect 18750 3440 18755 3496
rect 17033 3438 18755 3440
rect 17033 3435 17099 3438
rect 18689 3435 18755 3438
rect 20989 3496 21055 3501
rect 20989 3440 20994 3496
rect 21050 3440 21055 3496
rect 20989 3435 21055 3440
rect 21265 3498 21331 3501
rect 26325 3498 26391 3501
rect 21265 3496 26391 3498
rect 21265 3440 21270 3496
rect 21326 3440 26330 3496
rect 26386 3440 26391 3496
rect 21265 3438 26391 3440
rect 21265 3435 21331 3438
rect 26325 3435 26391 3438
rect 10726 3300 10732 3364
rect 10796 3362 10802 3364
rect 12433 3362 12499 3365
rect 10796 3360 12499 3362
rect 10796 3304 12438 3360
rect 12494 3304 12499 3360
rect 10796 3302 12499 3304
rect 10796 3300 10802 3302
rect 12433 3299 12499 3302
rect 16665 3362 16731 3365
rect 18321 3362 18387 3365
rect 16665 3360 18387 3362
rect 16665 3304 16670 3360
rect 16726 3304 18326 3360
rect 18382 3304 18387 3360
rect 16665 3302 18387 3304
rect 16665 3299 16731 3302
rect 18321 3299 18387 3302
rect 18781 3362 18847 3365
rect 23933 3362 23999 3365
rect 18781 3360 23999 3362
rect 18781 3304 18786 3360
rect 18842 3304 23938 3360
rect 23994 3304 23999 3360
rect 18781 3302 23999 3304
rect 18781 3299 18847 3302
rect 23933 3299 23999 3302
rect 5610 3296 5930 3297
rect 0 3226 480 3256
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 1301 3226 1367 3229
rect 1669 3226 1735 3229
rect 0 3224 1735 3226
rect 0 3168 1306 3224
rect 1362 3168 1674 3224
rect 1730 3168 1735 3224
rect 0 3166 1735 3168
rect 0 3136 480 3166
rect 1301 3163 1367 3166
rect 1669 3163 1735 3166
rect 3417 3226 3483 3229
rect 7189 3226 7255 3229
rect 9213 3226 9279 3229
rect 3417 3224 4354 3226
rect 3417 3168 3422 3224
rect 3478 3168 4354 3224
rect 3417 3166 4354 3168
rect 3417 3163 3483 3166
rect 3969 3092 4035 3093
rect 3918 3028 3924 3092
rect 3988 3090 4035 3092
rect 4294 3090 4354 3166
rect 7189 3224 9279 3226
rect 7189 3168 7194 3224
rect 7250 3168 9218 3224
rect 9274 3168 9279 3224
rect 7189 3166 9279 3168
rect 7189 3163 7255 3166
rect 9213 3163 9279 3166
rect 18689 3226 18755 3229
rect 24025 3226 24091 3229
rect 27520 3226 28000 3256
rect 18689 3224 24091 3226
rect 18689 3168 18694 3224
rect 18750 3168 24030 3224
rect 24086 3168 24091 3224
rect 18689 3166 24091 3168
rect 18689 3163 18755 3166
rect 24025 3163 24091 3166
rect 24672 3166 28000 3226
rect 11513 3090 11579 3093
rect 3988 3088 4080 3090
rect 4030 3032 4080 3088
rect 3988 3030 4080 3032
rect 4294 3088 11579 3090
rect 4294 3032 11518 3088
rect 11574 3032 11579 3088
rect 4294 3030 11579 3032
rect 3988 3028 4035 3030
rect 3969 3027 4035 3028
rect 11513 3027 11579 3030
rect 19374 3028 19380 3092
rect 19444 3090 19450 3092
rect 19609 3090 19675 3093
rect 19444 3088 19675 3090
rect 19444 3032 19614 3088
rect 19670 3032 19675 3088
rect 19444 3030 19675 3032
rect 19444 3028 19450 3030
rect 19609 3027 19675 3030
rect 20662 3028 20668 3092
rect 20732 3090 20738 3092
rect 21541 3090 21607 3093
rect 20732 3088 21607 3090
rect 20732 3032 21546 3088
rect 21602 3032 21607 3088
rect 20732 3030 21607 3032
rect 20732 3028 20738 3030
rect 21541 3027 21607 3030
rect 23105 3090 23171 3093
rect 24672 3090 24732 3166
rect 27520 3136 28000 3166
rect 23105 3088 24732 3090
rect 23105 3032 23110 3088
rect 23166 3032 24732 3088
rect 23105 3030 24732 3032
rect 23105 3027 23171 3030
rect 2313 2954 2379 2957
rect 6637 2954 6703 2957
rect 2313 2952 6703 2954
rect 2313 2896 2318 2952
rect 2374 2896 6642 2952
rect 6698 2896 6703 2952
rect 2313 2894 6703 2896
rect 2313 2891 2379 2894
rect 6637 2891 6703 2894
rect 8017 2954 8083 2957
rect 14917 2954 14983 2957
rect 8017 2952 14983 2954
rect 8017 2896 8022 2952
rect 8078 2896 14922 2952
rect 14978 2896 14983 2952
rect 8017 2894 14983 2896
rect 8017 2891 8083 2894
rect 14917 2891 14983 2894
rect 17401 2954 17467 2957
rect 25221 2954 25287 2957
rect 17401 2952 25287 2954
rect 17401 2896 17406 2952
rect 17462 2896 25226 2952
rect 25282 2896 25287 2952
rect 17401 2894 25287 2896
rect 17401 2891 17467 2894
rect 25221 2891 25287 2894
rect 2865 2818 2931 2821
rect 7189 2818 7255 2821
rect 2865 2816 7255 2818
rect 2865 2760 2870 2816
rect 2926 2760 7194 2816
rect 7250 2760 7255 2816
rect 2865 2758 7255 2760
rect 2865 2755 2931 2758
rect 7189 2755 7255 2758
rect 7649 2818 7715 2821
rect 8845 2818 8911 2821
rect 9949 2818 10015 2821
rect 7649 2816 10015 2818
rect 7649 2760 7654 2816
rect 7710 2760 8850 2816
rect 8906 2760 9954 2816
rect 10010 2760 10015 2816
rect 7649 2758 10015 2760
rect 7649 2755 7715 2758
rect 8845 2755 8911 2758
rect 9949 2755 10015 2758
rect 14365 2818 14431 2821
rect 16573 2818 16639 2821
rect 17493 2818 17559 2821
rect 14365 2816 17559 2818
rect 14365 2760 14370 2816
rect 14426 2760 16578 2816
rect 16634 2760 17498 2816
rect 17554 2760 17559 2816
rect 14365 2758 17559 2760
rect 14365 2755 14431 2758
rect 16573 2755 16639 2758
rect 17493 2755 17559 2758
rect 20069 2818 20135 2821
rect 23657 2818 23723 2821
rect 20069 2816 23723 2818
rect 20069 2760 20074 2816
rect 20130 2760 23662 2816
rect 23718 2760 23723 2816
rect 20069 2758 23723 2760
rect 20069 2755 20135 2758
rect 23657 2755 23723 2758
rect 10277 2752 10597 2753
rect 0 2682 480 2712
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 1669 2682 1735 2685
rect 0 2680 1735 2682
rect 0 2624 1674 2680
rect 1730 2624 1735 2680
rect 0 2622 1735 2624
rect 0 2592 480 2622
rect 1669 2619 1735 2622
rect 7741 2682 7807 2685
rect 9857 2682 9923 2685
rect 7741 2680 9923 2682
rect 7741 2624 7746 2680
rect 7802 2624 9862 2680
rect 9918 2624 9923 2680
rect 7741 2622 9923 2624
rect 7741 2619 7807 2622
rect 9857 2619 9923 2622
rect 11789 2682 11855 2685
rect 12382 2682 12388 2684
rect 11789 2680 12388 2682
rect 11789 2624 11794 2680
rect 11850 2624 12388 2680
rect 11789 2622 12388 2624
rect 11789 2619 11855 2622
rect 12382 2620 12388 2622
rect 12452 2620 12458 2684
rect 21633 2682 21699 2685
rect 23933 2682 23999 2685
rect 21633 2680 23999 2682
rect 21633 2624 21638 2680
rect 21694 2624 23938 2680
rect 23994 2624 23999 2680
rect 21633 2622 23999 2624
rect 21633 2619 21699 2622
rect 23933 2619 23999 2622
rect 26601 2682 26667 2685
rect 27520 2682 28000 2712
rect 26601 2680 28000 2682
rect 26601 2624 26606 2680
rect 26662 2624 28000 2680
rect 26601 2622 28000 2624
rect 26601 2619 26667 2622
rect 27520 2592 28000 2622
rect 8753 2546 8819 2549
rect 13997 2546 14063 2549
rect 8753 2544 14063 2546
rect 8753 2488 8758 2544
rect 8814 2488 14002 2544
rect 14058 2488 14063 2544
rect 8753 2486 14063 2488
rect 8753 2483 8819 2486
rect 13997 2483 14063 2486
rect 14549 2546 14615 2549
rect 18321 2546 18387 2549
rect 23565 2546 23631 2549
rect 14549 2544 23631 2546
rect 14549 2488 14554 2544
rect 14610 2488 18326 2544
rect 18382 2488 23570 2544
rect 23626 2488 23631 2544
rect 14549 2486 23631 2488
rect 14549 2483 14615 2486
rect 18321 2483 18387 2486
rect 23565 2483 23631 2486
rect 2957 2410 3023 2413
rect 14457 2410 14523 2413
rect 21725 2410 21791 2413
rect 23657 2412 23723 2413
rect 2957 2408 14523 2410
rect 2957 2352 2962 2408
rect 3018 2352 14462 2408
rect 14518 2352 14523 2408
rect 2957 2350 14523 2352
rect 2957 2347 3023 2350
rect 14457 2347 14523 2350
rect 14782 2408 21791 2410
rect 14782 2352 21730 2408
rect 21786 2352 21791 2408
rect 14782 2350 21791 2352
rect 10593 2274 10659 2277
rect 12985 2274 13051 2277
rect 14782 2274 14842 2350
rect 21725 2347 21791 2350
rect 23606 2348 23612 2412
rect 23676 2410 23723 2412
rect 23676 2408 23768 2410
rect 23718 2352 23768 2408
rect 23676 2350 23768 2352
rect 23676 2348 23723 2350
rect 23657 2347 23723 2348
rect 10593 2272 14842 2274
rect 10593 2216 10598 2272
rect 10654 2216 12990 2272
rect 13046 2216 14842 2272
rect 10593 2214 14842 2216
rect 10593 2211 10659 2214
rect 12985 2211 13051 2214
rect 15326 2212 15332 2276
rect 15396 2274 15402 2276
rect 23473 2274 23539 2277
rect 15396 2272 23539 2274
rect 15396 2216 23478 2272
rect 23534 2216 23539 2272
rect 15396 2214 23539 2216
rect 15396 2212 15402 2214
rect 23473 2211 23539 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 6821 2138 6887 2141
rect 6821 2136 12266 2138
rect 6821 2080 6826 2136
rect 6882 2080 12266 2136
rect 6821 2078 12266 2080
rect 6821 2075 6887 2078
rect 0 2002 480 2032
rect 1393 2002 1459 2005
rect 5073 2002 5139 2005
rect 12065 2002 12131 2005
rect 0 2000 1778 2002
rect 0 1944 1398 2000
rect 1454 1944 1778 2000
rect 0 1942 1778 1944
rect 0 1912 480 1942
rect 1393 1939 1459 1942
rect 1718 1866 1778 1942
rect 5073 2000 12131 2002
rect 5073 1944 5078 2000
rect 5134 1944 12070 2000
rect 12126 1944 12131 2000
rect 5073 1942 12131 1944
rect 12206 2002 12266 2078
rect 15285 2002 15351 2005
rect 12206 2000 15351 2002
rect 12206 1944 15290 2000
rect 15346 1944 15351 2000
rect 12206 1942 15351 1944
rect 5073 1939 5139 1942
rect 12065 1939 12131 1942
rect 15285 1939 15351 1942
rect 18505 2002 18571 2005
rect 25589 2002 25655 2005
rect 18505 2000 25655 2002
rect 18505 1944 18510 2000
rect 18566 1944 25594 2000
rect 25650 1944 25655 2000
rect 18505 1942 25655 1944
rect 18505 1939 18571 1942
rect 25589 1939 25655 1942
rect 25865 2002 25931 2005
rect 27520 2002 28000 2032
rect 25865 2000 28000 2002
rect 25865 1944 25870 2000
rect 25926 1944 28000 2000
rect 25865 1942 28000 1944
rect 25865 1939 25931 1942
rect 27520 1912 28000 1942
rect 17585 1866 17651 1869
rect 19977 1866 20043 1869
rect 1718 1864 17651 1866
rect 1718 1808 17590 1864
rect 17646 1808 17651 1864
rect 1718 1806 17651 1808
rect 17585 1803 17651 1806
rect 17726 1864 20043 1866
rect 17726 1808 19982 1864
rect 20038 1808 20043 1864
rect 17726 1806 20043 1808
rect 197 1730 263 1733
rect 11513 1730 11579 1733
rect 197 1728 11579 1730
rect 197 1672 202 1728
rect 258 1672 11518 1728
rect 11574 1672 11579 1728
rect 197 1670 11579 1672
rect 197 1667 263 1670
rect 11513 1667 11579 1670
rect 11881 1730 11947 1733
rect 17726 1730 17786 1806
rect 19977 1803 20043 1806
rect 22737 1866 22803 1869
rect 25078 1866 25084 1868
rect 22737 1864 25084 1866
rect 22737 1808 22742 1864
rect 22798 1808 25084 1864
rect 22737 1806 25084 1808
rect 22737 1803 22803 1806
rect 25078 1804 25084 1806
rect 25148 1804 25154 1868
rect 11881 1728 17786 1730
rect 11881 1672 11886 1728
rect 11942 1672 17786 1728
rect 11881 1670 17786 1672
rect 11881 1667 11947 1670
rect 17902 1668 17908 1732
rect 17972 1730 17978 1732
rect 18321 1730 18387 1733
rect 17972 1728 18387 1730
rect 17972 1672 18326 1728
rect 18382 1672 18387 1728
rect 17972 1670 18387 1672
rect 17972 1668 17978 1670
rect 18321 1667 18387 1670
rect 20161 1730 20227 1733
rect 26509 1730 26575 1733
rect 20161 1728 26575 1730
rect 20161 1672 20166 1728
rect 20222 1672 26514 1728
rect 26570 1672 26575 1728
rect 20161 1670 26575 1672
rect 20161 1667 20227 1670
rect 26509 1667 26575 1670
rect 2037 1594 2103 1597
rect 11646 1594 11652 1596
rect 2037 1592 11652 1594
rect 2037 1536 2042 1592
rect 2098 1536 11652 1592
rect 2037 1534 11652 1536
rect 2037 1531 2103 1534
rect 11646 1532 11652 1534
rect 11716 1532 11722 1596
rect 24669 1594 24735 1597
rect 22878 1592 24735 1594
rect 22878 1536 24674 1592
rect 24730 1536 24735 1592
rect 22878 1534 24735 1536
rect 0 1458 480 1488
rect 3877 1458 3943 1461
rect 0 1456 3943 1458
rect 0 1400 3882 1456
rect 3938 1400 3943 1456
rect 0 1398 3943 1400
rect 0 1368 480 1398
rect 3877 1395 3943 1398
rect 11605 1458 11671 1461
rect 22878 1458 22938 1534
rect 24669 1531 24735 1534
rect 11605 1456 22938 1458
rect 11605 1400 11610 1456
rect 11666 1400 22938 1456
rect 11605 1398 22938 1400
rect 23013 1458 23079 1461
rect 26785 1458 26851 1461
rect 23013 1456 26851 1458
rect 23013 1400 23018 1456
rect 23074 1400 26790 1456
rect 26846 1400 26851 1456
rect 23013 1398 26851 1400
rect 11605 1395 11671 1398
rect 23013 1395 23079 1398
rect 26785 1395 26851 1398
rect 27153 1458 27219 1461
rect 27520 1458 28000 1488
rect 27153 1456 28000 1458
rect 27153 1400 27158 1456
rect 27214 1400 28000 1456
rect 27153 1398 28000 1400
rect 27153 1395 27219 1398
rect 27520 1368 28000 1398
rect 6913 1322 6979 1325
rect 24945 1322 25011 1325
rect 6913 1320 25011 1322
rect 6913 1264 6918 1320
rect 6974 1264 24950 1320
rect 25006 1264 25011 1320
rect 6913 1262 25011 1264
rect 6913 1259 6979 1262
rect 24945 1259 25011 1262
rect 6269 1186 6335 1189
rect 24025 1186 24091 1189
rect 6269 1184 24091 1186
rect 6269 1128 6274 1184
rect 6330 1128 24030 1184
rect 24086 1128 24091 1184
rect 6269 1126 24091 1128
rect 6269 1123 6335 1126
rect 24025 1123 24091 1126
rect 9121 1050 9187 1053
rect 25497 1050 25563 1053
rect 9121 1048 25563 1050
rect 9121 992 9126 1048
rect 9182 992 25502 1048
rect 25558 992 25563 1048
rect 9121 990 25563 992
rect 9121 987 9187 990
rect 25497 987 25563 990
rect 0 914 480 944
rect 1577 914 1643 917
rect 0 912 1643 914
rect 0 856 1582 912
rect 1638 856 1643 912
rect 0 854 1643 856
rect 0 824 480 854
rect 1577 851 1643 854
rect 3509 914 3575 917
rect 16113 914 16179 917
rect 3509 912 16179 914
rect 3509 856 3514 912
rect 3570 856 16118 912
rect 16174 856 16179 912
rect 3509 854 16179 856
rect 3509 851 3575 854
rect 16113 851 16179 854
rect 23473 914 23539 917
rect 27520 914 28000 944
rect 23473 912 28000 914
rect 23473 856 23478 912
rect 23534 856 28000 912
rect 23473 854 28000 856
rect 23473 851 23539 854
rect 27520 824 28000 854
rect 0 370 480 400
rect 4245 370 4311 373
rect 0 368 4311 370
rect 0 312 4250 368
rect 4306 312 4311 368
rect 0 310 4311 312
rect 0 280 480 310
rect 4245 307 4311 310
rect 7097 370 7163 373
rect 17585 370 17651 373
rect 7097 368 17651 370
rect 7097 312 7102 368
rect 7158 312 17590 368
rect 17646 312 17651 368
rect 7097 310 17651 312
rect 7097 307 7163 310
rect 17585 307 17651 310
rect 26233 370 26299 373
rect 27520 370 28000 400
rect 26233 368 28000 370
rect 26233 312 26238 368
rect 26294 312 28000 368
rect 26233 310 28000 312
rect 26233 307 26299 310
rect 27520 280 28000 310
rect 7557 234 7623 237
rect 19425 234 19491 237
rect 7557 232 19491 234
rect 7557 176 7562 232
rect 7618 176 19430 232
rect 19486 176 19491 232
rect 7557 174 19491 176
rect 7557 171 7623 174
rect 19425 171 19491 174
rect 8477 98 8543 101
rect 9305 98 9371 101
rect 21081 98 21147 101
rect 8477 96 21147 98
rect 8477 40 8482 96
rect 8538 40 9310 96
rect 9366 40 21086 96
rect 21142 40 21147 96
rect 8477 38 21147 40
rect 8477 35 8543 38
rect 9305 35 9371 38
rect 21081 35 21147 38
<< via3 >>
rect 20116 26012 20180 26076
rect 14596 25876 14660 25940
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 14044 25468 14108 25532
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 11284 25196 11348 25260
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 13676 24924 13740 24988
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 15516 24788 15580 24852
rect 23612 24788 23676 24852
rect 20668 24516 20732 24580
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 13492 24380 13556 24444
rect 15700 24380 15764 24444
rect 23980 24108 24044 24172
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 15332 23700 15396 23764
rect 15884 23760 15948 23764
rect 15884 23704 15934 23760
rect 15934 23704 15948 23760
rect 15884 23700 15948 23704
rect 21404 23700 21468 23764
rect 19012 23564 19076 23628
rect 23060 23564 23124 23628
rect 25268 23564 25332 23628
rect 12388 23488 12452 23492
rect 12388 23432 12402 23488
rect 12402 23432 12452 23488
rect 12388 23428 12452 23432
rect 14780 23428 14844 23492
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 10916 23020 10980 23084
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 12020 22612 12084 22676
rect 12756 22476 12820 22540
rect 3924 22340 3988 22404
rect 17540 22340 17604 22404
rect 19380 22400 19444 22404
rect 19380 22344 19430 22400
rect 19430 22344 19444 22400
rect 19380 22340 19444 22344
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 13492 22128 13556 22132
rect 13492 22072 13506 22128
rect 13506 22072 13556 22128
rect 13492 22068 13556 22072
rect 9076 21932 9140 21996
rect 11100 21932 11164 21996
rect 15884 21932 15948 21996
rect 19012 21932 19076 21996
rect 22324 21992 22388 21996
rect 22324 21936 22338 21992
rect 22338 21936 22388 21992
rect 22324 21932 22388 21936
rect 23060 21992 23124 21996
rect 23060 21936 23074 21992
rect 23074 21936 23124 21992
rect 23060 21932 23124 21936
rect 16436 21796 16500 21860
rect 20300 21796 20364 21860
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 25820 21720 25884 21724
rect 25820 21664 25870 21720
rect 25870 21664 25884 21720
rect 25820 21660 25884 21664
rect 13308 21524 13372 21588
rect 10916 21388 10980 21452
rect 21036 21388 21100 21452
rect 24716 21388 24780 21452
rect 24716 21252 24780 21316
rect 25084 21312 25148 21316
rect 25084 21256 25098 21312
rect 25098 21256 25148 21312
rect 25084 21252 25148 21256
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 15332 20980 15396 21044
rect 18460 21040 18524 21044
rect 18460 20984 18474 21040
rect 18474 20984 18524 21040
rect 18460 20980 18524 20984
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14412 20708 14476 20772
rect 22324 20768 22388 20772
rect 22324 20712 22338 20768
rect 22338 20712 22388 20768
rect 22324 20708 22388 20712
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 11836 20436 11900 20500
rect 13308 20300 13372 20364
rect 23796 20300 23860 20364
rect 9628 20224 9692 20228
rect 9628 20168 9642 20224
rect 9642 20168 9692 20224
rect 9628 20164 9692 20168
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 9996 20028 10060 20092
rect 11468 20028 11532 20092
rect 14412 20028 14476 20092
rect 17540 19892 17604 19956
rect 20668 20028 20732 20092
rect 21772 20028 21836 20092
rect 23428 20028 23492 20092
rect 20484 19952 20548 19956
rect 20484 19896 20498 19952
rect 20498 19896 20548 19952
rect 20484 19892 20548 19896
rect 20852 19952 20916 19956
rect 20852 19896 20866 19952
rect 20866 19896 20916 19952
rect 20852 19892 20916 19896
rect 23060 19892 23124 19956
rect 10916 19816 10980 19820
rect 10916 19760 10966 19816
rect 10966 19760 10980 19816
rect 10916 19756 10980 19760
rect 16068 19756 16132 19820
rect 17908 19620 17972 19684
rect 20668 19620 20732 19684
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 16620 19408 16684 19412
rect 16620 19352 16670 19408
rect 16670 19352 16684 19408
rect 10916 19212 10980 19276
rect 11652 19212 11716 19276
rect 16620 19348 16684 19352
rect 20668 19348 20732 19412
rect 21036 19348 21100 19412
rect 25084 19348 25148 19412
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 21956 19212 22020 19276
rect 22876 19076 22940 19140
rect 25268 19076 25332 19140
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 6316 18804 6380 18868
rect 9812 18668 9876 18732
rect 10916 18728 10980 18732
rect 10916 18672 10966 18728
rect 10966 18672 10980 18728
rect 10916 18668 10980 18672
rect 11652 18668 11716 18732
rect 15700 18804 15764 18868
rect 17172 18668 17236 18732
rect 23244 18592 23308 18596
rect 23244 18536 23294 18592
rect 23294 18536 23308 18592
rect 23244 18532 23308 18536
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 3004 18260 3068 18324
rect 10916 18396 10980 18460
rect 10732 18260 10796 18324
rect 12388 18396 12452 18460
rect 2084 18048 2148 18052
rect 2084 17992 2098 18048
rect 2098 17992 2148 18048
rect 2084 17988 2148 17992
rect 3556 17988 3620 18052
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 20852 17988 20916 18052
rect 21220 18048 21284 18052
rect 21220 17992 21234 18048
rect 21234 17992 21284 18048
rect 21220 17988 21284 17992
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 12756 17852 12820 17916
rect 20116 17852 20180 17916
rect 25636 17852 25700 17916
rect 14596 17580 14660 17644
rect 15700 17580 15764 17644
rect 13676 17444 13740 17508
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 5212 17368 5276 17372
rect 5212 17312 5226 17368
rect 5226 17312 5276 17368
rect 5212 17308 5276 17312
rect 25084 17716 25148 17780
rect 25268 17444 25332 17508
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 25452 17368 25516 17372
rect 25452 17312 25466 17368
rect 25466 17312 25516 17368
rect 25452 17308 25516 17312
rect 15884 17172 15948 17236
rect 17540 17232 17604 17236
rect 17540 17176 17590 17232
rect 17590 17176 17604 17232
rect 17540 17172 17604 17176
rect 11468 17036 11532 17100
rect 14596 16900 14660 16964
rect 22692 16960 22756 16964
rect 22692 16904 22742 16960
rect 22742 16904 22756 16960
rect 22692 16900 22756 16904
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 8156 16628 8220 16692
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 15332 16628 15396 16692
rect 23612 16764 23676 16828
rect 23796 16764 23860 16828
rect 22692 16628 22756 16692
rect 22508 16492 22572 16556
rect 23428 16492 23492 16556
rect 16436 16356 16500 16420
rect 21588 16356 21652 16420
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 12756 16220 12820 16284
rect 14044 16220 14108 16284
rect 16252 16220 16316 16284
rect 9812 16084 9876 16148
rect 12388 16084 12452 16148
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 11836 15676 11900 15740
rect 12204 15676 12268 15740
rect 20852 15948 20916 16012
rect 21956 15948 22020 16012
rect 22140 15948 22204 16012
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 21588 15540 21652 15604
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 9996 15132 10060 15196
rect 11652 15192 11716 15196
rect 11652 15136 11666 15192
rect 11666 15136 11716 15192
rect 11652 15132 11716 15136
rect 21588 15404 21652 15468
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 18460 15132 18524 15196
rect 9812 14996 9876 15060
rect 9996 14996 10060 15060
rect 13492 14996 13556 15060
rect 23060 14996 23124 15060
rect 24716 14996 24780 15060
rect 12388 14860 12452 14924
rect 20300 14860 20364 14924
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 7052 14648 7116 14652
rect 7052 14592 7066 14648
rect 7066 14592 7116 14648
rect 7052 14588 7116 14592
rect 19012 14588 19076 14652
rect 25820 14588 25884 14652
rect 9812 14180 9876 14244
rect 16252 14180 16316 14244
rect 24716 14180 24780 14244
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 6868 13908 6932 13972
rect 11652 13908 11716 13972
rect 12388 13832 12452 13836
rect 12388 13776 12402 13832
rect 12402 13776 12452 13832
rect 12388 13772 12452 13776
rect 13308 13772 13372 13836
rect 14412 13832 14476 13836
rect 16804 14044 16868 14108
rect 15332 13968 15396 13972
rect 15332 13912 15346 13968
rect 15346 13912 15396 13968
rect 15332 13908 15396 13912
rect 14412 13776 14462 13832
rect 14462 13776 14476 13832
rect 14412 13772 14476 13776
rect 22692 13636 22756 13700
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 13676 13500 13740 13564
rect 25084 13500 25148 13564
rect 2452 13092 2516 13156
rect 6316 13152 6380 13156
rect 6316 13096 6366 13152
rect 6366 13096 6380 13152
rect 6316 13092 6380 13096
rect 16252 13228 16316 13292
rect 17724 13228 17788 13292
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 3372 12956 3436 13020
rect 14596 13016 14660 13020
rect 14596 12960 14646 13016
rect 14646 12960 14660 13016
rect 14596 12956 14660 12960
rect 24900 12956 24964 13020
rect 4844 12548 4908 12612
rect 9996 12548 10060 12612
rect 22324 12820 22388 12884
rect 23244 12820 23308 12884
rect 24900 12880 24964 12884
rect 24900 12824 24914 12880
rect 24914 12824 24964 12880
rect 24900 12820 24964 12824
rect 22876 12744 22940 12748
rect 22876 12688 22890 12744
rect 22890 12688 22940 12744
rect 22876 12684 22940 12688
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 6868 12412 6932 12476
rect 9996 12412 10060 12476
rect 13308 12412 13372 12476
rect 14596 12412 14660 12476
rect 13860 12276 13924 12340
rect 16252 12276 16316 12340
rect 16804 12336 16868 12340
rect 16804 12280 16818 12336
rect 16818 12280 16868 12336
rect 16804 12276 16868 12280
rect 11836 12140 11900 12204
rect 22508 12548 22572 12612
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 23612 12472 23676 12476
rect 23612 12416 23662 12472
rect 23662 12416 23676 12472
rect 23612 12412 23676 12416
rect 25452 12412 25516 12476
rect 22876 12276 22940 12340
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 12572 11868 12636 11932
rect 13676 11868 13740 11932
rect 11836 11792 11900 11796
rect 11836 11736 11850 11792
rect 11850 11736 11900 11792
rect 11836 11732 11900 11736
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 21036 11868 21100 11932
rect 23060 11868 23124 11932
rect 20484 11732 20548 11796
rect 11284 11656 11348 11660
rect 11284 11600 11298 11656
rect 11298 11600 11348 11656
rect 11284 11596 11348 11600
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 7420 11384 7484 11388
rect 7420 11328 7434 11384
rect 7434 11328 7484 11384
rect 7420 11324 7484 11328
rect 9996 11188 10060 11252
rect 17724 11460 17788 11524
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 10916 11324 10980 11388
rect 21956 11324 22020 11388
rect 3372 11052 3436 11116
rect 15700 11112 15764 11116
rect 15700 11056 15750 11112
rect 15750 11056 15764 11112
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 4844 10780 4908 10844
rect 15700 11052 15764 11056
rect 19380 11052 19444 11116
rect 17172 10916 17236 10980
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 15516 10780 15580 10844
rect 25268 10644 25332 10708
rect 7972 10568 8036 10572
rect 7972 10512 7986 10568
rect 7986 10512 8036 10568
rect 7972 10508 8036 10512
rect 10732 10508 10796 10572
rect 10916 10508 10980 10572
rect 13308 10508 13372 10572
rect 24900 10508 24964 10572
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 12572 10236 12636 10300
rect 23428 10236 23492 10300
rect 25636 10236 25700 10300
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 12756 9556 12820 9620
rect 14228 9556 14292 9620
rect 20852 9556 20916 9620
rect 21772 9556 21836 9620
rect 12388 9284 12452 9348
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 23060 9148 23124 9212
rect 15884 9012 15948 9076
rect 23612 9012 23676 9076
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 10916 8604 10980 8668
rect 11100 8664 11164 8668
rect 11100 8608 11150 8664
rect 11150 8608 11164 8664
rect 11100 8604 11164 8608
rect 13860 8604 13924 8668
rect 14596 8468 14660 8532
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 25084 8664 25148 8668
rect 25084 8608 25134 8664
rect 25134 8608 25148 8664
rect 25084 8604 25148 8608
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 9260 8120 9324 8124
rect 9260 8064 9274 8120
rect 9274 8064 9324 8120
rect 9260 8060 9324 8064
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 4292 7788 4356 7852
rect 21404 8060 21468 8124
rect 17724 7652 17788 7716
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 16068 7576 16132 7580
rect 16068 7520 16082 7576
rect 16082 7520 16132 7576
rect 16068 7516 16132 7520
rect 21588 7516 21652 7580
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 11100 7108 11164 7172
rect 23428 7168 23492 7172
rect 23428 7112 23478 7168
rect 23478 7112 23492 7168
rect 23428 7108 23492 7112
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 17540 6972 17604 7036
rect 17908 6836 17972 6900
rect 23796 6836 23860 6900
rect 3556 6700 3620 6764
rect 10732 6700 10796 6764
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 12388 6428 12452 6492
rect 11652 6292 11716 6356
rect 14412 6428 14476 6492
rect 15332 6700 15396 6764
rect 23980 6760 24044 6764
rect 23980 6704 24030 6760
rect 24030 6704 24044 6760
rect 23980 6700 24044 6704
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 12020 6080 12084 6084
rect 12020 6024 12070 6080
rect 12070 6024 12084 6080
rect 12020 6020 12084 6024
rect 20668 6020 20732 6084
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 11100 5884 11164 5948
rect 14596 5884 14660 5948
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 23428 5204 23492 5268
rect 24716 5204 24780 5268
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 14780 4932 14844 4996
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 8708 4584 8772 4588
rect 8708 4528 8722 4584
rect 8722 4528 8772 4584
rect 8708 4524 8772 4528
rect 23428 4524 23492 4588
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 21220 4252 21284 4316
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 3924 3708 3988 3772
rect 11836 3708 11900 3772
rect 23060 3844 23124 3908
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 23980 3708 24044 3772
rect 9628 3572 9692 3636
rect 10732 3300 10796 3364
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 3924 3088 3988 3092
rect 3924 3032 3974 3088
rect 3974 3032 3988 3088
rect 3924 3028 3988 3032
rect 19380 3028 19444 3092
rect 20668 3028 20732 3092
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 12388 2620 12452 2684
rect 23612 2408 23676 2412
rect 23612 2352 23662 2408
rect 23662 2352 23676 2408
rect 23612 2348 23676 2352
rect 15332 2212 15396 2276
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 25084 1804 25148 1868
rect 17908 1668 17972 1732
rect 11652 1532 11716 1596
<< metal4 >>
rect 20115 26076 20181 26077
rect 20115 26012 20116 26076
rect 20180 26012 20181 26076
rect 20115 26011 20181 26012
rect 14595 25940 14661 25941
rect 14595 25876 14596 25940
rect 14660 25876 14661 25940
rect 14595 25875 14661 25876
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 3923 22404 3989 22405
rect 3923 22340 3924 22404
rect 3988 22340 3989 22404
rect 3923 22339 3989 22340
rect 3003 18324 3069 18325
rect 3003 18260 3004 18324
rect 3068 18260 3069 18324
rect 3003 18259 3069 18260
rect 2083 18052 2149 18053
rect 2083 17988 2084 18052
rect 2148 17988 2149 18052
rect 2083 17987 2149 17988
rect 2086 5898 2146 17987
rect 2451 13156 2517 13157
rect 2451 13092 2452 13156
rect 2516 13092 2517 13156
rect 2451 13091 2517 13092
rect 2454 12698 2514 13091
rect 3006 1818 3066 18259
rect 3371 13020 3437 13021
rect 3371 12956 3372 13020
rect 3436 12956 3437 13020
rect 3371 12955 3437 12956
rect 3374 12018 3434 12955
rect 3374 11117 3434 11782
rect 3371 11116 3437 11117
rect 3371 11052 3372 11116
rect 3436 11052 3437 11116
rect 3371 11051 3437 11052
rect 3555 6764 3621 6765
rect 3555 6700 3556 6764
rect 3620 6700 3621 6764
rect 3555 6699 3621 6700
rect 3558 6578 3618 6699
rect 3926 3773 3986 22339
rect 5610 21792 5931 22816
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 14043 25532 14109 25533
rect 14043 25468 14044 25532
rect 14108 25468 14109 25532
rect 14043 25467 14109 25468
rect 11283 25260 11349 25261
rect 11283 25196 11284 25260
rect 11348 25196 11349 25260
rect 11283 25195 11349 25196
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10915 23084 10981 23085
rect 10915 23020 10916 23084
rect 10980 23020 10981 23084
rect 10915 23019 10981 23020
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 9075 21932 9076 21982
rect 9140 21932 9141 21982
rect 9075 21931 9141 21932
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 10277 21248 10597 22272
rect 10918 21453 10978 23019
rect 11099 21996 11165 21997
rect 11099 21932 11100 21996
rect 11164 21932 11165 21996
rect 11099 21931 11165 21932
rect 10915 21452 10981 21453
rect 10915 21388 10916 21452
rect 10980 21388 10981 21452
rect 10915 21387 10981 21388
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 9627 20228 9693 20229
rect 9627 20164 9628 20228
rect 9692 20164 9693 20228
rect 9627 20163 9693 20164
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 6315 18868 6381 18869
rect 6315 18804 6316 18868
rect 6380 18804 6381 18868
rect 6315 18803 6381 18804
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 4846 12613 4906 13142
rect 5610 13088 5931 14112
rect 6318 14058 6378 18803
rect 8155 16692 8221 16693
rect 8155 16628 8156 16692
rect 8220 16628 8221 16692
rect 8155 16627 8221 16628
rect 6867 13972 6933 13973
rect 6867 13908 6868 13972
rect 6932 13908 6933 13972
rect 6867 13907 6933 13908
rect 6318 13157 6378 13822
rect 6315 13156 6381 13157
rect 6315 13092 6316 13156
rect 6380 13092 6381 13156
rect 6315 13091 6381 13092
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 4843 12612 4909 12613
rect 4843 12548 4844 12612
rect 4908 12548 4909 12612
rect 4843 12547 4909 12548
rect 5610 12000 5931 13024
rect 6870 12477 6930 13907
rect 6867 12476 6933 12477
rect 6867 12412 6868 12476
rect 6932 12412 6933 12476
rect 6867 12411 6933 12412
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 7422 11389 7482 16542
rect 8158 16098 8218 16627
rect 9630 13378 9690 20163
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 9995 20092 10061 20093
rect 9995 20028 9996 20092
rect 10060 20028 10061 20092
rect 9995 20027 10061 20028
rect 9998 19498 10058 20027
rect 9811 18732 9877 18733
rect 9811 18668 9812 18732
rect 9876 18668 9877 18732
rect 9811 18667 9877 18668
rect 9814 16149 9874 18667
rect 9811 16148 9877 16149
rect 9811 16084 9812 16148
rect 9876 16084 9877 16148
rect 9811 16083 9877 16084
rect 9998 15197 10058 19262
rect 10277 19072 10597 20096
rect 10918 19821 10978 21387
rect 10915 19820 10981 19821
rect 10915 19756 10916 19820
rect 10980 19756 10981 19820
rect 10915 19755 10981 19756
rect 10915 19276 10981 19277
rect 10915 19212 10916 19276
rect 10980 19212 10981 19276
rect 10915 19211 10981 19212
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10918 18733 10978 19211
rect 10915 18732 10981 18733
rect 10915 18668 10916 18732
rect 10980 18668 10981 18732
rect 10915 18667 10981 18668
rect 10915 18460 10981 18461
rect 10915 18396 10916 18460
rect 10980 18396 10981 18460
rect 10915 18395 10981 18396
rect 10731 18324 10797 18325
rect 10731 18260 10732 18324
rect 10796 18260 10797 18324
rect 10731 18259 10797 18260
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 9995 15196 10061 15197
rect 9995 15132 9996 15196
rect 10060 15132 10061 15196
rect 9995 15131 10061 15132
rect 9811 15060 9877 15061
rect 9811 14996 9812 15060
rect 9876 14996 9877 15060
rect 9811 14995 9877 14996
rect 9995 15060 10061 15061
rect 9995 14996 9996 15060
rect 10060 14996 10061 15060
rect 9995 14995 10061 14996
rect 9814 14245 9874 14995
rect 9811 14244 9877 14245
rect 9811 14180 9812 14244
rect 9876 14180 9877 14244
rect 9811 14179 9877 14180
rect 7419 11388 7485 11389
rect 7419 11324 7420 11388
rect 7484 11324 7485 11388
rect 7419 11323 7485 11324
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 4843 10844 4909 10845
rect 4843 10780 4844 10844
rect 4908 10780 4909 10844
rect 4843 10779 4909 10780
rect 4846 9978 4906 10779
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 9259 8124 9325 8125
rect 9259 8060 9260 8124
rect 9324 8060 9325 8124
rect 9259 8059 9325 8060
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 9262 7258 9322 8059
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 8710 4589 8770 4982
rect 8707 4588 8773 4589
rect 8707 4524 8708 4588
rect 8772 4524 8773 4588
rect 8707 4523 8773 4524
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 3923 3772 3989 3773
rect 3923 3708 3924 3772
rect 3988 3708 3989 3772
rect 3923 3707 3989 3708
rect 5610 3296 5931 4320
rect 9630 3637 9690 13142
rect 9998 12613 10058 14995
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 9995 12612 10061 12613
rect 9995 12548 9996 12612
rect 10060 12548 10061 12612
rect 9995 12547 10061 12548
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 9995 12476 10061 12477
rect 9995 12412 9996 12476
rect 10060 12412 10061 12476
rect 9995 12411 10061 12412
rect 9998 11253 10058 12411
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 9995 11252 10061 11253
rect 9995 11188 9996 11252
rect 10060 11188 10061 11252
rect 9995 11187 10061 11188
rect 10277 10368 10597 11392
rect 10734 10573 10794 18259
rect 10918 11389 10978 18395
rect 10915 11388 10981 11389
rect 10915 11324 10916 11388
rect 10980 11324 10981 11388
rect 10915 11323 10981 11324
rect 10731 10572 10797 10573
rect 10731 10508 10732 10572
rect 10796 10508 10797 10572
rect 10731 10507 10797 10508
rect 10915 10572 10981 10573
rect 10915 10508 10916 10572
rect 10980 10508 10981 10572
rect 10915 10507 10981 10508
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10918 8669 10978 10507
rect 11102 8669 11162 21931
rect 11286 11661 11346 25195
rect 13675 24988 13741 24989
rect 13675 24924 13676 24988
rect 13740 24924 13741 24988
rect 13675 24923 13741 24924
rect 13491 24444 13557 24445
rect 13491 24380 13492 24444
rect 13556 24380 13557 24444
rect 13491 24379 13557 24380
rect 12387 23492 12453 23493
rect 12387 23428 12388 23492
rect 12452 23428 12453 23492
rect 12387 23427 12453 23428
rect 12019 22676 12085 22677
rect 12019 22612 12020 22676
rect 12084 22612 12085 22676
rect 12019 22611 12085 22612
rect 11835 20500 11901 20501
rect 11835 20436 11836 20500
rect 11900 20436 11901 20500
rect 11835 20435 11901 20436
rect 11467 20092 11533 20093
rect 11467 20028 11468 20092
rect 11532 20028 11533 20092
rect 11467 20027 11533 20028
rect 11470 17101 11530 20027
rect 11651 19276 11717 19277
rect 11651 19212 11652 19276
rect 11716 19212 11717 19276
rect 11651 19211 11717 19212
rect 11654 18733 11714 19211
rect 11651 18732 11717 18733
rect 11651 18668 11652 18732
rect 11716 18668 11717 18732
rect 11651 18667 11717 18668
rect 11838 18138 11898 20435
rect 11467 17100 11533 17101
rect 11467 17036 11468 17100
rect 11532 17036 11533 17100
rect 11467 17035 11533 17036
rect 11838 15741 11898 17902
rect 11835 15740 11901 15741
rect 11835 15676 11836 15740
rect 11900 15676 11901 15740
rect 11835 15675 11901 15676
rect 11651 15132 11652 15182
rect 11716 15132 11717 15182
rect 11651 15131 11717 15132
rect 11283 11660 11349 11661
rect 11283 11596 11284 11660
rect 11348 11596 11349 11660
rect 11283 11595 11349 11596
rect 11654 11338 11714 13822
rect 11835 12204 11901 12205
rect 11835 12140 11836 12204
rect 11900 12140 11901 12204
rect 11835 12139 11901 12140
rect 11838 11797 11898 12139
rect 11835 11796 11901 11797
rect 11835 11732 11836 11796
rect 11900 11732 11901 11796
rect 11835 11731 11901 11732
rect 10915 8668 10981 8669
rect 10915 8604 10916 8668
rect 10980 8604 10981 8668
rect 10915 8603 10981 8604
rect 11099 8668 11165 8669
rect 11099 8604 11100 8668
rect 11164 8604 11165 8668
rect 11099 8603 11165 8604
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 12022 7850 12082 22611
rect 12390 18461 12450 23427
rect 12755 22540 12821 22541
rect 12755 22476 12756 22540
rect 12820 22476 12821 22540
rect 12755 22475 12821 22476
rect 12387 18460 12453 18461
rect 12387 18396 12388 18460
rect 12452 18396 12453 18460
rect 12387 18395 12453 18396
rect 12758 17917 12818 22475
rect 13494 22133 13554 24379
rect 13491 22132 13557 22133
rect 13491 22068 13492 22132
rect 13556 22068 13557 22132
rect 13491 22067 13557 22068
rect 13307 21588 13373 21589
rect 13307 21524 13308 21588
rect 13372 21524 13373 21588
rect 13678 21538 13738 24923
rect 13307 21523 13373 21524
rect 13310 20365 13370 21523
rect 13307 20364 13373 20365
rect 13307 20300 13308 20364
rect 13372 20300 13373 20364
rect 13307 20299 13373 20300
rect 12755 17916 12821 17917
rect 12755 17852 12756 17916
rect 12820 17852 12821 17916
rect 12755 17851 12821 17852
rect 12758 16778 12818 17851
rect 12755 16284 12821 16285
rect 12755 16220 12756 16284
rect 12820 16220 12821 16284
rect 12755 16219 12821 16220
rect 12387 16148 12453 16149
rect 12387 16084 12388 16148
rect 12452 16084 12453 16148
rect 12387 16083 12453 16084
rect 12203 15740 12269 15741
rect 12203 15676 12204 15740
rect 12268 15676 12269 15740
rect 12203 15675 12269 15676
rect 11838 7790 12082 7850
rect 11102 7173 11162 7702
rect 11099 7172 11165 7173
rect 11099 7108 11100 7172
rect 11164 7108 11165 7172
rect 11838 7170 11898 7790
rect 12206 7170 12266 15675
rect 12390 14925 12450 16083
rect 12387 14924 12453 14925
rect 12387 14860 12388 14924
rect 12452 14860 12453 14924
rect 12387 14859 12453 14860
rect 12390 13970 12450 14859
rect 12758 14738 12818 16219
rect 12390 13910 12634 13970
rect 12387 13836 12453 13837
rect 12387 13772 12388 13836
rect 12452 13772 12453 13836
rect 12387 13771 12453 13772
rect 12390 9349 12450 13771
rect 12574 11933 12634 13910
rect 12571 11932 12637 11933
rect 12571 11868 12572 11932
rect 12636 11868 12637 11932
rect 12571 11867 12637 11868
rect 12574 10301 12634 11867
rect 12571 10300 12637 10301
rect 12571 10236 12572 10300
rect 12636 10236 12637 10300
rect 12571 10235 12637 10236
rect 12758 9621 12818 14502
rect 13310 13837 13370 20299
rect 13678 17642 13738 21302
rect 13494 17582 13738 17642
rect 13494 15061 13554 17582
rect 13675 17508 13741 17509
rect 13675 17444 13676 17508
rect 13740 17444 13741 17508
rect 14046 17458 14106 25467
rect 14411 20772 14477 20773
rect 14411 20708 14412 20772
rect 14476 20708 14477 20772
rect 14411 20707 14477 20708
rect 14414 20093 14474 20707
rect 14411 20092 14477 20093
rect 14411 20028 14412 20092
rect 14476 20028 14477 20092
rect 14411 20027 14477 20028
rect 14598 17645 14658 25875
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 15515 24852 15581 24853
rect 15515 24788 15516 24852
rect 15580 24788 15581 24852
rect 15515 24787 15581 24788
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14779 23492 14845 23493
rect 14779 23428 14780 23492
rect 14844 23428 14845 23492
rect 14779 23427 14845 23428
rect 14595 17644 14661 17645
rect 14595 17580 14596 17644
rect 14660 17580 14661 17644
rect 14595 17579 14661 17580
rect 13675 17443 13741 17444
rect 13491 15060 13557 15061
rect 13491 14996 13492 15060
rect 13556 14996 13557 15060
rect 13491 14995 13557 14996
rect 13307 13836 13373 13837
rect 13307 13772 13308 13836
rect 13372 13772 13373 13836
rect 13307 13771 13373 13772
rect 13678 13565 13738 17443
rect 14046 16285 14106 17222
rect 14595 16964 14661 16965
rect 14595 16900 14596 16964
rect 14660 16900 14661 16964
rect 14595 16899 14661 16900
rect 14043 16284 14109 16285
rect 14043 16220 14044 16284
rect 14108 16220 14109 16284
rect 14043 16219 14109 16220
rect 13675 13564 13741 13565
rect 13675 13500 13676 13564
rect 13740 13500 13741 13564
rect 13675 13499 13741 13500
rect 13307 12476 13373 12477
rect 13307 12412 13308 12476
rect 13372 12412 13373 12476
rect 13307 12411 13373 12412
rect 13310 10573 13370 12411
rect 13862 12341 13922 12462
rect 13859 12340 13925 12341
rect 13859 12276 13860 12340
rect 13924 12276 13925 12340
rect 13859 12275 13925 12276
rect 13307 10572 13373 10573
rect 13307 10508 13308 10572
rect 13372 10508 13373 10572
rect 13307 10507 13373 10508
rect 12755 9620 12821 9621
rect 12755 9556 12756 9620
rect 12820 9556 12821 9620
rect 12755 9555 12821 9556
rect 12387 9348 12453 9349
rect 12387 9284 12388 9348
rect 12452 9284 12453 9348
rect 12387 9283 12453 9284
rect 13862 8669 13922 9742
rect 14230 9621 14290 15862
rect 14411 13836 14477 13837
rect 14411 13772 14412 13836
rect 14476 13772 14477 13836
rect 14411 13771 14477 13772
rect 14227 9620 14293 9621
rect 14227 9556 14228 9620
rect 14292 9556 14293 9620
rect 14227 9555 14293 9556
rect 13859 8668 13925 8669
rect 13859 8604 13860 8668
rect 13924 8604 13925 8668
rect 13859 8603 13925 8604
rect 11838 7110 11944 7170
rect 11099 7107 11165 7108
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10731 6764 10797 6765
rect 10731 6700 10732 6764
rect 10796 6700 10797 6764
rect 10731 6699 10797 6700
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 9627 3636 9693 3637
rect 9627 3572 9628 3636
rect 9692 3572 9693 3636
rect 9627 3571 9693 3572
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 2752 10597 3776
rect 10734 3365 10794 6699
rect 11651 6292 11652 6342
rect 11716 6292 11717 6342
rect 11651 6291 11717 6292
rect 11099 5948 11165 5949
rect 11099 5898 11100 5948
rect 11164 5898 11165 5948
rect 11884 5810 11944 7110
rect 12022 7110 12266 7170
rect 12022 6085 12082 7110
rect 14414 6493 14474 13771
rect 14598 13021 14658 16899
rect 14595 13020 14661 13021
rect 14595 12956 14596 13020
rect 14660 12956 14661 13020
rect 14595 12955 14661 12956
rect 14595 12476 14661 12477
rect 14595 12412 14596 12476
rect 14660 12412 14661 12476
rect 14595 12411 14661 12412
rect 14598 8533 14658 12411
rect 14595 8532 14661 8533
rect 14595 8468 14596 8532
rect 14660 8468 14661 8532
rect 14595 8467 14661 8468
rect 14411 6492 14477 6493
rect 14411 6428 14412 6492
rect 14476 6428 14477 6492
rect 14411 6427 14477 6428
rect 12019 6084 12085 6085
rect 12019 6020 12020 6084
rect 12084 6020 12085 6084
rect 12019 6019 12085 6020
rect 14595 5948 14661 5949
rect 14595 5884 14596 5948
rect 14660 5884 14661 5948
rect 14595 5883 14661 5884
rect 11838 5750 11944 5810
rect 11838 3773 11898 5750
rect 14598 3858 14658 5883
rect 14782 4997 14842 23427
rect 14944 22880 15264 23904
rect 15331 23764 15397 23765
rect 15331 23700 15332 23764
rect 15396 23700 15397 23764
rect 15331 23699 15397 23700
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 15334 21045 15394 23699
rect 15331 21044 15397 21045
rect 15331 20980 15332 21044
rect 15396 20980 15397 21044
rect 15331 20979 15397 20980
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 15331 16692 15397 16693
rect 15331 16628 15332 16692
rect 15396 16628 15397 16692
rect 15331 16627 15397 16628
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 15334 13973 15394 16627
rect 15331 13972 15397 13973
rect 15331 13908 15332 13972
rect 15396 13908 15397 13972
rect 15331 13907 15397 13908
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 15518 10845 15578 24787
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 15699 24444 15765 24445
rect 15699 24380 15700 24444
rect 15764 24380 15765 24444
rect 15699 24379 15765 24380
rect 15702 18869 15762 24379
rect 15883 23764 15949 23765
rect 15883 23700 15884 23764
rect 15948 23700 15949 23764
rect 15883 23699 15949 23700
rect 15886 21997 15946 23699
rect 19011 23628 19077 23629
rect 19011 23564 19012 23628
rect 19076 23564 19077 23628
rect 19011 23563 19077 23564
rect 17539 22404 17605 22405
rect 17539 22340 17540 22404
rect 17604 22340 17605 22404
rect 17539 22339 17605 22340
rect 15883 21996 15949 21997
rect 15883 21932 15884 21996
rect 15948 21932 15949 21996
rect 15883 21931 15949 21932
rect 16435 21860 16501 21861
rect 16435 21796 16436 21860
rect 16500 21796 16501 21860
rect 16435 21795 16501 21796
rect 16067 19820 16133 19821
rect 16067 19756 16068 19820
rect 16132 19756 16133 19820
rect 16067 19755 16133 19756
rect 15699 18868 15765 18869
rect 15699 18804 15700 18868
rect 15764 18804 15765 18868
rect 15699 18803 15765 18804
rect 15699 17644 15765 17645
rect 15699 17580 15700 17644
rect 15764 17580 15765 17644
rect 15699 17579 15765 17580
rect 15702 11117 15762 17579
rect 15883 17236 15949 17237
rect 15883 17172 15884 17236
rect 15948 17172 15949 17236
rect 15883 17171 15949 17172
rect 15699 11116 15765 11117
rect 15699 11052 15700 11116
rect 15764 11052 15765 11116
rect 15699 11051 15765 11052
rect 15515 10844 15581 10845
rect 15515 10780 15516 10844
rect 15580 10780 15581 10844
rect 15515 10779 15581 10780
rect 15518 10658 15578 10779
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 15886 9077 15946 17171
rect 15883 9076 15949 9077
rect 15883 9012 15884 9076
rect 15948 9012 15949 9076
rect 15883 9011 15949 9012
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 16070 7581 16130 19755
rect 16438 16421 16498 21795
rect 17542 20178 17602 22339
rect 19014 21997 19074 23563
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19379 22404 19445 22405
rect 19379 22340 19380 22404
rect 19444 22340 19445 22404
rect 19379 22339 19445 22340
rect 19011 21996 19077 21997
rect 19011 21932 19012 21996
rect 19076 21932 19077 21996
rect 19011 21931 19077 21932
rect 18459 21044 18525 21045
rect 18459 20980 18460 21044
rect 18524 20980 18525 21044
rect 18459 20979 18525 20980
rect 17539 19892 17540 19942
rect 17604 19892 17605 19942
rect 17539 19891 17605 19892
rect 17907 19684 17973 19685
rect 17907 19620 17908 19684
rect 17972 19620 17973 19684
rect 17907 19619 17973 19620
rect 17910 19498 17970 19619
rect 16619 19412 16685 19413
rect 16619 19348 16620 19412
rect 16684 19410 16685 19412
rect 16684 19350 16866 19410
rect 16684 19348 16685 19350
rect 16619 19347 16685 19348
rect 16435 16420 16501 16421
rect 16435 16356 16436 16420
rect 16500 16356 16501 16420
rect 16435 16355 16501 16356
rect 16251 16284 16317 16285
rect 16251 16220 16252 16284
rect 16316 16220 16317 16284
rect 16251 16219 16317 16220
rect 16254 14245 16314 16219
rect 16251 14244 16317 14245
rect 16251 14180 16252 14244
rect 16316 14180 16317 14244
rect 16251 14179 16317 14180
rect 16806 14109 16866 19350
rect 17171 18732 17237 18733
rect 17171 18668 17172 18732
rect 17236 18668 17237 18732
rect 17171 18667 17237 18668
rect 16803 14108 16869 14109
rect 16803 14044 16804 14108
rect 16868 14044 16869 14108
rect 16803 14043 16869 14044
rect 16251 13292 16317 13293
rect 16251 13228 16252 13292
rect 16316 13228 16317 13292
rect 16251 13227 16317 13228
rect 16254 12341 16314 13227
rect 16806 12341 16866 14043
rect 16251 12340 16317 12341
rect 16251 12276 16252 12340
rect 16316 12276 16317 12340
rect 16251 12275 16317 12276
rect 16803 12340 16869 12341
rect 16803 12276 16804 12340
rect 16868 12276 16869 12340
rect 16803 12275 16869 12276
rect 17174 10981 17234 18667
rect 17539 17236 17605 17237
rect 17539 17172 17540 17236
rect 17604 17172 17605 17236
rect 17539 17171 17605 17172
rect 17171 10980 17237 10981
rect 17171 10916 17172 10980
rect 17236 10916 17237 10980
rect 17171 10915 17237 10916
rect 16067 7580 16133 7581
rect 16067 7516 16068 7580
rect 16132 7516 16133 7580
rect 16067 7515 16133 7516
rect 17542 7037 17602 17171
rect 18462 15197 18522 20979
rect 18459 15196 18525 15197
rect 18459 15132 18460 15196
rect 18524 15132 18525 15196
rect 18459 15131 18525 15132
rect 19014 14653 19074 21931
rect 19011 14652 19077 14653
rect 19011 14588 19012 14652
rect 19076 14588 19077 14652
rect 19011 14587 19077 14588
rect 17723 13292 17789 13293
rect 17723 13228 17724 13292
rect 17788 13228 17789 13292
rect 17723 13227 17789 13228
rect 17726 11525 17786 13227
rect 17723 11524 17789 11525
rect 17723 11460 17724 11524
rect 17788 11460 17789 11524
rect 17723 11459 17789 11460
rect 17726 7717 17786 11459
rect 19382 11338 19442 22339
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 20118 17917 20178 26011
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 23611 24852 23677 24853
rect 23611 24788 23612 24852
rect 23676 24788 23677 24852
rect 23611 24787 23677 24788
rect 20667 24580 20733 24581
rect 20667 24516 20668 24580
rect 20732 24516 20733 24580
rect 20667 24515 20733 24516
rect 20670 22218 20730 24515
rect 21403 23764 21469 23765
rect 21403 23700 21404 23764
rect 21468 23700 21469 23764
rect 21403 23699 21469 23700
rect 20299 21860 20365 21861
rect 20299 21796 20300 21860
rect 20364 21796 20365 21860
rect 20299 21795 20365 21796
rect 20115 17916 20181 17917
rect 20115 17852 20116 17916
rect 20180 17852 20181 17916
rect 20115 17851 20181 17852
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 20302 14925 20362 21795
rect 20667 20092 20733 20093
rect 20667 20028 20668 20092
rect 20732 20028 20733 20092
rect 20667 20027 20733 20028
rect 20483 19956 20549 19957
rect 20483 19892 20484 19956
rect 20548 19892 20549 19956
rect 20483 19891 20549 19892
rect 20299 14924 20365 14925
rect 20299 14860 20300 14924
rect 20364 14860 20365 14924
rect 20486 14922 20546 19891
rect 20670 19685 20730 20027
rect 20851 19956 20917 19957
rect 20851 19892 20852 19956
rect 20916 19892 20917 19956
rect 20851 19891 20917 19892
rect 20667 19684 20733 19685
rect 20667 19620 20668 19684
rect 20732 19620 20733 19684
rect 20667 19619 20733 19620
rect 20667 19412 20733 19413
rect 20667 19348 20668 19412
rect 20732 19348 20733 19412
rect 20667 19347 20733 19348
rect 20486 14862 20592 14922
rect 20299 14859 20365 14860
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 20532 14650 20592 14862
rect 20266 14590 20592 14650
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 20486 11797 20546 14590
rect 20483 11796 20549 11797
rect 20483 11732 20484 11796
rect 20548 11732 20549 11796
rect 20483 11731 20549 11732
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19379 11052 19380 11102
rect 19444 11052 19445 11102
rect 19379 11051 19445 11052
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 17723 7716 17789 7717
rect 17723 7652 17724 7716
rect 17788 7652 17789 7716
rect 17723 7651 17789 7652
rect 17539 7036 17605 7037
rect 17539 6972 17540 7036
rect 17604 6972 17605 7036
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 17539 6971 17605 6972
rect 17910 6901 17970 7022
rect 17907 6900 17973 6901
rect 17907 6836 17908 6900
rect 17972 6836 17973 6900
rect 17907 6835 17973 6836
rect 15331 6764 15397 6765
rect 15331 6700 15332 6764
rect 15396 6700 15397 6764
rect 15331 6699 15397 6700
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14779 4996 14845 4997
rect 14779 4932 14780 4996
rect 14844 4932 14845 4996
rect 14779 4931 14845 4932
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 11835 3772 11901 3773
rect 11835 3708 11836 3772
rect 11900 3708 11901 3772
rect 11835 3707 11901 3708
rect 10731 3364 10797 3365
rect 10731 3300 10732 3364
rect 10796 3300 10797 3364
rect 10731 3299 10797 3300
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 11654 1597 11714 2942
rect 12387 2684 12453 2685
rect 12387 2620 12388 2684
rect 12452 2620 12453 2684
rect 12387 2619 12453 2620
rect 12390 2498 12450 2619
rect 14944 2208 15264 3232
rect 15334 2277 15394 6699
rect 19610 6016 19930 7040
rect 20670 6085 20730 19347
rect 20854 18053 20914 19891
rect 21035 19412 21101 19413
rect 21035 19348 21036 19412
rect 21100 19348 21101 19412
rect 21035 19347 21101 19348
rect 20851 18052 20917 18053
rect 20851 17988 20852 18052
rect 20916 17988 20917 18052
rect 20851 17987 20917 17988
rect 20851 16012 20917 16013
rect 20851 15948 20852 16012
rect 20916 15948 20917 16012
rect 20851 15947 20917 15948
rect 20854 9621 20914 15947
rect 21038 11933 21098 19347
rect 21219 18052 21285 18053
rect 21219 17988 21220 18052
rect 21284 17988 21285 18052
rect 21219 17987 21285 17988
rect 21035 11932 21101 11933
rect 21035 11868 21036 11932
rect 21100 11868 21101 11932
rect 21035 11867 21101 11868
rect 20851 9620 20917 9621
rect 20851 9556 20852 9620
rect 20916 9556 20917 9620
rect 20851 9555 20917 9556
rect 20667 6084 20733 6085
rect 20667 6020 20668 6084
rect 20732 6020 20733 6084
rect 20667 6019 20733 6020
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 20670 3093 20730 4982
rect 21222 4317 21282 17987
rect 21406 8125 21466 23699
rect 23059 23628 23125 23629
rect 23059 23564 23060 23628
rect 23124 23564 23125 23628
rect 23059 23563 23125 23564
rect 23062 21997 23122 23563
rect 22323 21996 22389 21997
rect 22323 21932 22324 21996
rect 22388 21932 22389 21996
rect 22323 21931 22389 21932
rect 23059 21996 23125 21997
rect 23059 21932 23060 21996
rect 23124 21932 23125 21996
rect 23059 21931 23125 21932
rect 22326 20773 22386 21931
rect 22323 20772 22389 20773
rect 22323 20708 22324 20772
rect 22388 20708 22389 20772
rect 22323 20707 22389 20708
rect 21771 20092 21837 20093
rect 21771 20028 21772 20092
rect 21836 20028 21837 20092
rect 21771 20027 21837 20028
rect 21587 16420 21653 16421
rect 21587 16356 21588 16420
rect 21652 16356 21653 16420
rect 21587 16355 21653 16356
rect 21590 15605 21650 16355
rect 21587 15604 21653 15605
rect 21587 15540 21588 15604
rect 21652 15540 21653 15604
rect 21587 15539 21653 15540
rect 21587 15468 21653 15469
rect 21587 15404 21588 15468
rect 21652 15404 21653 15468
rect 21587 15403 21653 15404
rect 21403 8124 21469 8125
rect 21403 8060 21404 8124
rect 21468 8060 21469 8124
rect 21403 8059 21469 8060
rect 21590 7581 21650 15403
rect 21774 9621 21834 20027
rect 21955 19276 22021 19277
rect 21955 19212 21956 19276
rect 22020 19212 22021 19276
rect 21955 19211 22021 19212
rect 21958 18050 22018 19211
rect 21958 17990 22202 18050
rect 22142 16013 22202 17990
rect 21955 16012 22021 16013
rect 21955 15948 21956 16012
rect 22020 15948 22021 16012
rect 21955 15947 22021 15948
rect 22139 16012 22205 16013
rect 22139 15948 22140 16012
rect 22204 15948 22205 16012
rect 22139 15947 22205 15948
rect 21958 11389 22018 15947
rect 22326 12885 22386 20707
rect 23427 20092 23493 20093
rect 23427 20028 23428 20092
rect 23492 20028 23493 20092
rect 23427 20027 23493 20028
rect 23059 19956 23125 19957
rect 22694 16965 22754 19942
rect 23059 19892 23060 19956
rect 23124 19892 23125 19956
rect 23059 19891 23125 19892
rect 22875 19140 22941 19141
rect 22875 19076 22876 19140
rect 22940 19076 22941 19140
rect 22875 19075 22941 19076
rect 22691 16964 22757 16965
rect 22691 16900 22692 16964
rect 22756 16900 22757 16964
rect 22691 16899 22757 16900
rect 22691 16692 22757 16693
rect 22691 16628 22692 16692
rect 22756 16628 22757 16692
rect 22691 16627 22757 16628
rect 22507 16556 22573 16557
rect 22507 16492 22508 16556
rect 22572 16492 22573 16556
rect 22507 16491 22573 16492
rect 22323 12884 22389 12885
rect 22323 12820 22324 12884
rect 22388 12820 22389 12884
rect 22323 12819 22389 12820
rect 22510 12613 22570 16491
rect 22694 13701 22754 16627
rect 22691 13700 22757 13701
rect 22691 13636 22692 13700
rect 22756 13636 22757 13700
rect 22691 13635 22757 13636
rect 22878 12882 22938 19075
rect 23062 15061 23122 19891
rect 23243 18596 23309 18597
rect 23243 18532 23244 18596
rect 23308 18532 23309 18596
rect 23243 18531 23309 18532
rect 23059 15060 23125 15061
rect 23059 14996 23060 15060
rect 23124 14996 23125 15060
rect 23059 14995 23125 14996
rect 23246 12885 23306 18531
rect 23430 16690 23490 20027
rect 23614 16829 23674 24787
rect 23979 24172 24045 24173
rect 23979 24108 23980 24172
rect 24044 24108 24045 24172
rect 23979 24107 24045 24108
rect 23795 20364 23861 20365
rect 23795 20300 23796 20364
rect 23860 20300 23861 20364
rect 23795 20299 23861 20300
rect 23798 16829 23858 20299
rect 23611 16828 23677 16829
rect 23611 16764 23612 16828
rect 23676 16764 23677 16828
rect 23611 16763 23677 16764
rect 23795 16828 23861 16829
rect 23795 16764 23796 16828
rect 23860 16764 23861 16828
rect 23795 16763 23861 16764
rect 23430 16630 23674 16690
rect 23427 16556 23493 16557
rect 23427 16492 23428 16556
rect 23492 16492 23493 16556
rect 23427 16491 23493 16492
rect 23243 12884 23309 12885
rect 22878 12822 23122 12882
rect 22875 12748 22941 12749
rect 22875 12684 22876 12748
rect 22940 12684 22941 12748
rect 22875 12683 22941 12684
rect 22507 12612 22573 12613
rect 22507 12548 22508 12612
rect 22572 12548 22573 12612
rect 22507 12547 22573 12548
rect 22878 12341 22938 12683
rect 22875 12340 22941 12341
rect 22875 12276 22876 12340
rect 22940 12276 22941 12340
rect 22875 12275 22941 12276
rect 23062 11933 23122 12822
rect 23243 12820 23244 12884
rect 23308 12820 23309 12884
rect 23243 12819 23309 12820
rect 23059 11932 23125 11933
rect 23059 11868 23060 11932
rect 23124 11868 23125 11932
rect 23059 11867 23125 11868
rect 21955 11388 22021 11389
rect 21955 11324 21956 11388
rect 22020 11324 22021 11388
rect 21955 11323 22021 11324
rect 23430 10301 23490 16491
rect 23614 12477 23674 16630
rect 23611 12476 23677 12477
rect 23611 12412 23612 12476
rect 23676 12412 23677 12476
rect 23611 12411 23677 12412
rect 23427 10300 23493 10301
rect 23427 10236 23428 10300
rect 23492 10236 23493 10300
rect 23427 10235 23493 10236
rect 21771 9620 21837 9621
rect 21771 9556 21772 9620
rect 21836 9556 21837 9620
rect 21771 9555 21837 9556
rect 23059 9212 23125 9213
rect 23059 9148 23060 9212
rect 23124 9148 23125 9212
rect 23059 9147 23125 9148
rect 21587 7580 21653 7581
rect 21587 7516 21588 7580
rect 21652 7516 21653 7580
rect 21587 7515 21653 7516
rect 21219 4316 21285 4317
rect 21219 4252 21220 4316
rect 21284 4252 21285 4316
rect 21219 4251 21285 4252
rect 23062 3909 23122 9147
rect 23611 9076 23677 9077
rect 23611 9012 23612 9076
rect 23676 9012 23677 9076
rect 23611 9011 23677 9012
rect 23614 8618 23674 9011
rect 23795 6900 23861 6901
rect 23795 6836 23796 6900
rect 23860 6836 23861 6900
rect 23795 6835 23861 6836
rect 23798 6578 23858 6835
rect 23982 6765 24042 24107
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 25267 23628 25333 23629
rect 25267 23564 25268 23628
rect 25332 23564 25333 23628
rect 25267 23563 25333 23564
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24715 21452 24781 21453
rect 24715 21388 24716 21452
rect 24780 21450 24781 21452
rect 24780 21390 24962 21450
rect 24780 21388 24781 21390
rect 24715 21387 24781 21388
rect 24715 21316 24781 21317
rect 24715 21252 24716 21316
rect 24780 21252 24781 21316
rect 24715 21251 24781 21252
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24718 15061 24778 21251
rect 24715 15060 24781 15061
rect 24715 14996 24716 15060
rect 24780 14996 24781 15060
rect 24715 14995 24781 14996
rect 24715 14244 24781 14245
rect 24715 14180 24716 14244
rect 24780 14180 24781 14244
rect 24715 14179 24781 14180
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 23979 6764 24045 6765
rect 23979 6700 23980 6764
rect 24044 6700 24045 6764
rect 23979 6699 24045 6700
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 23427 5268 23493 5269
rect 23427 5204 23428 5268
rect 23492 5204 23493 5268
rect 23427 5203 23493 5204
rect 23430 4589 23490 5203
rect 23427 4588 23493 4589
rect 23427 4524 23428 4588
rect 23492 4524 23493 4588
rect 23427 4523 23493 4524
rect 24277 4384 24597 5408
rect 24718 5269 24778 14179
rect 24902 13021 24962 21390
rect 25083 21316 25149 21317
rect 25083 21252 25084 21316
rect 25148 21252 25149 21316
rect 25083 21251 25149 21252
rect 25086 19413 25146 21251
rect 25083 19412 25149 19413
rect 25083 19348 25084 19412
rect 25148 19348 25149 19412
rect 25083 19347 25149 19348
rect 25270 19141 25330 23563
rect 25819 21724 25885 21725
rect 25819 21660 25820 21724
rect 25884 21660 25885 21724
rect 25819 21659 25885 21660
rect 25267 19140 25333 19141
rect 25267 19076 25268 19140
rect 25332 19076 25333 19140
rect 25267 19075 25333 19076
rect 25635 17916 25701 17917
rect 25635 17852 25636 17916
rect 25700 17852 25701 17916
rect 25635 17851 25701 17852
rect 25083 17780 25149 17781
rect 25083 17716 25084 17780
rect 25148 17716 25149 17780
rect 25083 17715 25149 17716
rect 25086 13565 25146 17715
rect 25267 17508 25333 17509
rect 25267 17444 25268 17508
rect 25332 17444 25333 17508
rect 25267 17443 25333 17444
rect 25083 13564 25149 13565
rect 25083 13500 25084 13564
rect 25148 13500 25149 13564
rect 25083 13499 25149 13500
rect 24899 13020 24965 13021
rect 24899 12956 24900 13020
rect 24964 12956 24965 13020
rect 24899 12955 24965 12956
rect 24899 12884 24965 12885
rect 24899 12820 24900 12884
rect 24964 12820 24965 12884
rect 24899 12819 24965 12820
rect 24902 10573 24962 12819
rect 25270 10709 25330 17443
rect 25451 17372 25517 17373
rect 25451 17308 25452 17372
rect 25516 17308 25517 17372
rect 25451 17307 25517 17308
rect 25454 12477 25514 17307
rect 25451 12476 25517 12477
rect 25451 12412 25452 12476
rect 25516 12412 25517 12476
rect 25451 12411 25517 12412
rect 25267 10708 25333 10709
rect 25267 10644 25268 10708
rect 25332 10644 25333 10708
rect 25267 10643 25333 10644
rect 24899 10572 24965 10573
rect 24899 10508 24900 10572
rect 24964 10508 24965 10572
rect 24899 10507 24965 10508
rect 25638 10301 25698 17851
rect 25822 14653 25882 21659
rect 25819 14652 25885 14653
rect 25819 14588 25820 14652
rect 25884 14588 25885 14652
rect 25819 14587 25885 14588
rect 25635 10300 25701 10301
rect 25635 10236 25636 10300
rect 25700 10236 25701 10300
rect 25635 10235 25701 10236
rect 25083 8668 25149 8669
rect 25083 8604 25084 8668
rect 25148 8604 25149 8668
rect 25083 8603 25149 8604
rect 24715 5268 24781 5269
rect 24715 5204 24716 5268
rect 24780 5204 24781 5268
rect 24715 5203 24781 5204
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 23059 3908 23125 3909
rect 23059 3844 23060 3908
rect 23124 3844 23125 3908
rect 23059 3843 23125 3844
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 20667 3092 20733 3093
rect 20667 3028 20668 3092
rect 20732 3028 20733 3092
rect 20667 3027 20733 3028
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 15331 2276 15397 2277
rect 15331 2212 15332 2276
rect 15396 2212 15397 2276
rect 15331 2211 15397 2212
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 2128 19930 2688
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
rect 25086 1869 25146 8603
rect 25083 1868 25149 1869
rect 25083 1804 25084 1868
rect 25148 1804 25149 1868
rect 25083 1803 25149 1804
rect 11651 1596 11717 1597
rect 11651 1532 11652 1596
rect 11716 1532 11717 1596
rect 11651 1531 11717 1532
<< via4 >>
rect 2366 12462 2602 12698
rect 1998 5662 2234 5898
rect 3470 18052 3706 18138
rect 3470 17988 3556 18052
rect 3556 17988 3620 18052
rect 3620 17988 3706 18052
rect 3470 17902 3706 17988
rect 3286 11782 3522 12018
rect 3470 6342 3706 6578
rect 8990 21996 9226 22218
rect 8990 21982 9076 21996
rect 9076 21982 9140 21996
rect 9140 21982 9226 21996
rect 5126 17372 5362 17458
rect 5126 17308 5212 17372
rect 5212 17308 5276 17372
rect 5276 17308 5362 17372
rect 5126 17222 5362 17308
rect 4758 13142 4994 13378
rect 7334 16542 7570 16778
rect 6966 14652 7202 14738
rect 6966 14588 7052 14652
rect 7052 14588 7116 14652
rect 7116 14588 7202 14652
rect 6966 14502 7202 14588
rect 6230 13822 6466 14058
rect 8070 15862 8306 16098
rect 9910 19262 10146 19498
rect 9542 13142 9778 13378
rect 4758 9742 4994 9978
rect 7886 10572 8122 10658
rect 7886 10508 7972 10572
rect 7972 10508 8036 10572
rect 8036 10508 8122 10572
rect 7886 10422 8122 10508
rect 4206 7852 4442 7938
rect 4206 7788 4292 7852
rect 4292 7788 4356 7852
rect 4356 7788 4442 7852
rect 4206 7702 4442 7788
rect 9174 7022 9410 7258
rect 8622 4982 8858 5218
rect 11704 17902 11940 18138
rect 11566 15196 11802 15418
rect 11566 15182 11652 15196
rect 11652 15182 11716 15196
rect 11716 15182 11802 15196
rect 11566 13972 11802 14058
rect 11566 13908 11652 13972
rect 11652 13908 11716 13972
rect 11716 13908 11802 13972
rect 11566 13822 11802 13908
rect 11566 11102 11802 11338
rect 11014 7702 11250 7938
rect 13590 21302 13826 21538
rect 12670 16542 12906 16778
rect 12670 14502 12906 14738
rect 13958 17222 14194 17458
rect 14142 15862 14378 16098
rect 13774 12462 14010 12698
rect 13590 11932 13826 12018
rect 13590 11868 13676 11932
rect 13676 11868 13740 11932
rect 13740 11868 13826 11932
rect 13590 11782 13826 11868
rect 13774 9742 14010 9978
rect 3838 3092 4074 3178
rect 3838 3028 3924 3092
rect 3924 3028 3988 3092
rect 3988 3028 4074 3092
rect 3838 2942 4074 3028
rect 11566 6356 11802 6578
rect 11566 6342 11652 6356
rect 11652 6342 11716 6356
rect 11716 6342 11802 6356
rect 11014 5884 11100 5898
rect 11100 5884 11164 5898
rect 11164 5884 11250 5898
rect 11014 5662 11250 5884
rect 12302 6492 12538 6578
rect 12302 6428 12388 6492
rect 12388 6428 12452 6492
rect 12452 6428 12538 6492
rect 12302 6342 12538 6428
rect 15430 10422 15666 10658
rect 17454 19956 17690 20178
rect 17454 19942 17540 19956
rect 17540 19942 17604 19956
rect 17604 19942 17690 19956
rect 17822 19262 18058 19498
rect 20582 21982 20818 22218
rect 20950 21452 21186 21538
rect 20950 21388 21036 21452
rect 21036 21388 21100 21452
rect 21100 21388 21186 21452
rect 20950 21302 21186 21388
rect 20030 14502 20266 14738
rect 19294 11116 19530 11338
rect 19294 11102 19380 11116
rect 19380 11102 19444 11116
rect 19444 11102 19530 11116
rect 17822 7022 18058 7258
rect 14510 3622 14746 3858
rect 11566 2942 11802 3178
rect 2918 1582 3154 1818
rect 12302 2262 12538 2498
rect 20582 4982 20818 5218
rect 19294 3092 19530 3178
rect 19294 3028 19380 3092
rect 19380 3028 19444 3092
rect 19444 3028 19530 3092
rect 19294 2942 19530 3028
rect 22606 19942 22842 20178
rect 23526 8382 23762 8618
rect 23342 7172 23578 7258
rect 23342 7108 23428 7172
rect 23428 7108 23492 7172
rect 23492 7108 23578 7172
rect 23342 7022 23578 7108
rect 23710 6342 23946 6578
rect 23894 3772 24130 3858
rect 23894 3708 23980 3772
rect 23980 3708 24044 3772
rect 24044 3708 24130 3772
rect 23894 3622 24130 3708
rect 23526 2412 23762 2498
rect 23526 2348 23612 2412
rect 23612 2348 23676 2412
rect 23676 2348 23762 2412
rect 23526 2262 23762 2348
rect 17822 1732 18058 1818
rect 17822 1668 17908 1732
rect 17908 1668 17972 1732
rect 17972 1668 18058 1732
rect 17822 1582 18058 1668
<< metal5 >>
rect 8948 22218 20860 22260
rect 8948 21982 8990 22218
rect 9226 21982 20582 22218
rect 20818 21982 20860 22218
rect 8948 21940 20860 21982
rect 13548 21538 21228 21580
rect 13548 21302 13590 21538
rect 13826 21302 20950 21538
rect 21186 21302 21228 21538
rect 13548 21260 21228 21302
rect 17412 20178 22884 20220
rect 17412 19942 17454 20178
rect 17690 19942 22606 20178
rect 22842 19942 22884 20178
rect 17412 19900 22884 19942
rect 9868 19498 18100 19540
rect 9868 19262 9910 19498
rect 10146 19262 17822 19498
rect 18058 19262 18100 19498
rect 9868 19220 18100 19262
rect 3428 18138 11982 18180
rect 3428 17902 3470 18138
rect 3706 17902 11704 18138
rect 11940 17902 11982 18138
rect 3428 17860 11982 17902
rect 5084 17458 14236 17500
rect 5084 17222 5126 17458
rect 5362 17222 13958 17458
rect 14194 17222 14236 17458
rect 5084 17180 14236 17222
rect 7292 16778 12948 16820
rect 7292 16542 7334 16778
rect 7570 16542 12670 16778
rect 12906 16542 12948 16778
rect 7292 16500 12948 16542
rect 8028 16098 14420 16140
rect 8028 15862 8070 16098
rect 8306 15862 14142 16098
rect 14378 15862 14420 16098
rect 8028 15820 14420 15862
rect 11524 15418 13638 15460
rect 11524 15182 11566 15418
rect 11802 15182 13638 15418
rect 11524 15140 13638 15182
rect 13318 14780 13638 15140
rect 6924 14738 12948 14780
rect 6924 14502 6966 14738
rect 7202 14502 12670 14738
rect 12906 14502 12948 14738
rect 6924 14460 12948 14502
rect 13318 14738 20308 14780
rect 13318 14502 20030 14738
rect 20266 14502 20308 14738
rect 13318 14460 20308 14502
rect 6188 14058 11844 14100
rect 6188 13822 6230 14058
rect 6466 13822 11566 14058
rect 11802 13822 11844 14058
rect 6188 13780 11844 13822
rect 4716 13378 9820 13420
rect 4716 13142 4758 13378
rect 4994 13142 9542 13378
rect 9778 13142 9820 13378
rect 4716 13100 9820 13142
rect 2324 12698 14052 12740
rect 2324 12462 2366 12698
rect 2602 12462 13774 12698
rect 14010 12462 14052 12698
rect 2324 12420 14052 12462
rect 3244 12018 13868 12060
rect 3244 11782 3286 12018
rect 3522 11782 13590 12018
rect 13826 11782 13868 12018
rect 3244 11740 13868 11782
rect 11524 11338 19572 11380
rect 11524 11102 11566 11338
rect 11802 11102 19294 11338
rect 19530 11102 19572 11338
rect 11524 11060 19572 11102
rect 7844 10658 15708 10700
rect 7844 10422 7886 10658
rect 8122 10422 15430 10658
rect 15666 10422 15708 10658
rect 7844 10380 15708 10422
rect 4716 9978 14052 10020
rect 4716 9742 4758 9978
rect 4994 9742 13774 9978
rect 14010 9742 14052 9978
rect 4716 9700 14052 9742
rect 17044 8618 23804 8660
rect 17044 8382 23526 8618
rect 23762 8382 23804 8618
rect 17044 8340 23804 8382
rect 4164 7938 11292 7980
rect 4164 7702 4206 7938
rect 4442 7702 11014 7938
rect 11250 7702 11292 7938
rect 4164 7660 11292 7702
rect 17044 7300 17364 8340
rect 9132 7258 17364 7300
rect 9132 7022 9174 7258
rect 9410 7022 17364 7258
rect 9132 6980 17364 7022
rect 17780 7258 23620 7300
rect 17780 7022 17822 7258
rect 18058 7022 23342 7258
rect 23578 7022 23620 7258
rect 17780 6980 23620 7022
rect 3428 6578 11844 6620
rect 3428 6342 3470 6578
rect 3706 6342 11566 6578
rect 11802 6342 11844 6578
rect 3428 6300 11844 6342
rect 12260 6578 23988 6620
rect 12260 6342 12302 6578
rect 12538 6342 23710 6578
rect 23946 6342 23988 6578
rect 12260 6300 23988 6342
rect 1956 5898 11292 5940
rect 1956 5662 1998 5898
rect 2234 5662 11014 5898
rect 11250 5662 11292 5898
rect 1956 5620 11292 5662
rect 8580 5218 20860 5260
rect 8580 4982 8622 5218
rect 8858 4982 20582 5218
rect 20818 4982 20860 5218
rect 8580 4940 20860 4982
rect 14468 3858 24172 3900
rect 14468 3622 14510 3858
rect 14746 3622 23894 3858
rect 24130 3622 24172 3858
rect 14468 3580 24172 3622
rect 3796 3178 11108 3220
rect 3796 2942 3838 3178
rect 4074 2942 11108 3178
rect 3796 2900 11108 2942
rect 11524 3178 19572 3220
rect 11524 2942 11566 3178
rect 11802 2942 19294 3178
rect 19530 2942 19572 3178
rect 11524 2900 19572 2942
rect 10788 2540 11108 2900
rect 10788 2498 23804 2540
rect 10788 2262 12302 2498
rect 12538 2262 23526 2498
rect 23762 2262 23804 2498
rect 10788 2220 23804 2262
rect 2876 1818 18100 1860
rect 2876 1582 2918 1818
rect 3154 1582 17822 1818
rect 18058 1582 18100 1818
rect 2876 1540 18100 1582
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_6_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_5_
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_16 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2576 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_12
timestamp 1604681595
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16
timestamp 1604681595
transform 1 0 2576 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12
timestamp 1604681595
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_6__A0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_6__A1
timestamp 1604681595
transform 1 0 2392 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_5__A0
timestamp 1604681595
transform 1 0 2760 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_5__A1
timestamp 1604681595
transform 1 0 2392 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_20 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2944 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _054_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2944 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3496 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3312 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 3496 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23
timestamp 1604681595
transform 1 0 3220 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28
timestamp 1604681595
transform 1 0 3680 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_46
timestamp 1604681595
transform 1 0 5336 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_42
timestamp 1604681595
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5152 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48
timestamp 1604681595
transform 1 0 5520 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 5704 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604681595
transform 1 0 5704 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1604681595
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52
timestamp 1604681595
transform 1 0 5888 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_4__S
timestamp 1604681595
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1604681595
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_4__A1
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_62 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_72
timestamp 1604681595
transform 1 0 7728 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67
timestamp 1604681595
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_4__A0
timestamp 1604681595
transform 1 0 7084 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_4_
timestamp 1604681595
transform 1 0 6900 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_76
timestamp 1604681595
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7452 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8464 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1604681595
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_100
timestamp 1604681595
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_96
timestamp 1604681595
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 10672 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10304 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1604681595
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_5__A1
timestamp 1604681595
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_5__A0
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_117
timestamp 1604681595
transform 1 0 11868 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14444 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1604681595
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1604681595
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_136
timestamp 1604681595
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_140
timestamp 1604681595
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_144
timestamp 1604681595
transform 1 0 14352 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1604681595
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1604681595
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1604681595
transform 1 0 14904 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_163
timestamp 1604681595
transform 1 0 16100 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_159
timestamp 1604681595
transform 1 0 15732 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1604681595
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1604681595
transform 1 0 16284 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_3_
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_173
timestamp 1604681595
transform 1 0 17020 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1604681595
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 16468 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _115_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 17020 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 17480 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 17572 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_177
timestamp 1604681595
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_181
timestamp 1604681595
transform 1 0 17756 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_177
timestamp 1604681595
transform 1 0 17388 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_180
timestamp 1604681595
transform 1 0 17664 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_197
timestamp 1604681595
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_193
timestamp 1604681595
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_196
timestamp 1604681595
transform 1 0 19136 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_203
timestamp 1604681595
transform 1 0 19780 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_200
timestamp 1604681595
transform 1 0 19504 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 19596 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604681595
transform 1 0 19964 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20608 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1604681595
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_213
timestamp 1604681595
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_210
timestamp 1604681595
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 20976 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_214
timestamp 1604681595
transform 1 0 20792 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 21160 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_227
timestamp 1604681595
transform 1 0 21988 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_227
timestamp 1604681595
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 22172 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_234
timestamp 1604681595
transform 1 0 22632 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_231
timestamp 1604681595
transform 1 0 22356 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_231
timestamp 1604681595
transform 1 0 22356 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 22448 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1604681595
transform 1 0 22632 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604681595
transform 1 0 22816 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_240
timestamp 1604681595
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_244
timestamp 1604681595
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_240
timestamp 1604681595
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_4_
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_254
timestamp 1604681595
transform 1 0 24472 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 24656 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_258
timestamp 1604681595
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_262
timestamp 1604681595
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_258
timestamp 1604681595
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 25024 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_268
timestamp 1604681595
transform 1 0 25760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_269
timestamp 1604681595
transform 1 0 25852 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 25392 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1604681595
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 26036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 26312 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_273
timestamp 1604681595
transform 1 0 26220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_272
timestamp 1604681595
transform 1 0 26128 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_276
timestamp 1604681595
transform 1 0 26496 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_7_
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 2852 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_7__A0
timestamp 1604681595
transform 1 0 2392 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_12
timestamp 1604681595
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_16
timestamp 1604681595
transform 1 0 2576 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_5__S
timestamp 1604681595
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_21
timestamp 1604681595
transform 1 0 3036 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_25
timestamp 1604681595
transform 1 0 3404 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_41
timestamp 1604681595
transform 1 0 4876 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5888 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5428 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_45
timestamp 1604681595
transform 1 0 5244 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_49
timestamp 1604681595
transform 1 0 5612 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8280 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 7544 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 8096 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_68
timestamp 1604681595
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_72
timestamp 1604681595
transform 1 0 7728 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1604681595
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1604681595
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_88
timestamp 1604681595
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_102
timestamp 1604681595
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_5_
timestamp 1604681595
transform 1 0 11224 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_5__S
timestamp 1604681595
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_106
timestamp 1604681595
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_119
timestamp 1604681595
transform 1 0 12052 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_125
timestamp 1604681595
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12788 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 13800 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14260 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_136
timestamp 1604681595
transform 1 0 13616 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_140
timestamp 1604681595
transform 1 0 13984 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_145
timestamp 1604681595
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp 1604681595
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1604681595
transform 1 0 17480 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 17296 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 16928 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_170
timestamp 1604681595
transform 1 0 16744 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_174
timestamp 1604681595
transform 1 0 17112 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_187
timestamp 1604681595
transform 1 0 18308 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19044 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18492 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18860 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_191
timestamp 1604681595
transform 1 0 18676 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_204
timestamp 1604681595
transform 1 0 19872 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 21896 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_210
timestamp 1604681595
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_224
timestamp 1604681595
transform 1 0 21712 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_228
timestamp 1604681595
transform 1 0 22080 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 22448 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 24012 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 23644 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 22264 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_241
timestamp 1604681595
transform 1 0 23276 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_247
timestamp 1604681595
transform 1 0 23828 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 25024 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25392 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 25760 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_258
timestamp 1604681595
transform 1 0 24840 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_262
timestamp 1604681595
transform 1 0 25208 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_266
timestamp 1604681595
transform 1 0 25576 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_270
timestamp 1604681595
transform 1 0 25944 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 26128 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_274
timestamp 1604681595
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_7
timestamp 1604681595
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 1932 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_7__A1
timestamp 1604681595
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_11
timestamp 1604681595
transform 1 0 2116 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 2300 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 2852 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_4_
timestamp 1604681595
transform 1 0 4416 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 3864 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_28
timestamp 1604681595
transform 1 0 3680 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_32
timestamp 1604681595
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 5428 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6256 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_45
timestamp 1604681595
transform 1 0 5244 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_49
timestamp 1604681595
transform 1 0 5612 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1604681595
transform 1 0 6072 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_58
timestamp 1604681595
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 7820 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 7268 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_65
timestamp 1604681595
transform 1 0 7084 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_69
timestamp 1604681595
transform 1 0 7452 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l5_in_0_
timestamp 1604681595
transform 1 0 10028 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l5_in_0__S
timestamp 1604681595
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_2__S
timestamp 1604681595
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_89
timestamp 1604681595
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_93
timestamp 1604681595
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1604681595
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_106
timestamp 1604681595
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l5_in_0__A1
timestamp 1604681595
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604681595
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l5_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 14168 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_132
timestamp 1604681595
transform 1 0 13248 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_138
timestamp 1604681595
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_158
timestamp 1604681595
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_162
timestamp 1604681595
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 18308 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_175
timestamp 1604681595
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_179
timestamp 1604681595
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 19872 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 19688 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 19320 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_196
timestamp 1604681595
transform 1 0 19136 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_200
timestamp 1604681595
transform 1 0 19504 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1604681595
transform 1 0 21436 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_213
timestamp 1604681595
transform 1 0 20700 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_217
timestamp 1604681595
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 22448 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_230
timestamp 1604681595
transform 1 0 22264 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_234
timestamp 1604681595
transform 1 0 22632 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_238
timestamp 1604681595
transform 1 0 23000 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_254
timestamp 1604681595
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_258
timestamp 1604681595
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_268
timestamp 1604681595
transform 1 0 25760 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 26312 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_272
timestamp 1604681595
transform 1 0 26128 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_276
timestamp 1604681595
transform 1 0 26496 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_7__S
timestamp 1604681595
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_6__S
timestamp 1604681595
transform 1 0 1932 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_7
timestamp 1604681595
transform 1 0 1748 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_11
timestamp 1604681595
transform 1 0 2116 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_23
timestamp 1604681595
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_41
timestamp 1604681595
transform 1 0 4876 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5888 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 5428 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_45
timestamp 1604681595
transform 1 0 5244 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_49
timestamp 1604681595
transform 1 0 5612 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604681595
transform 1 0 8464 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 8004 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_68
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_73
timestamp 1604681595
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_77
timestamp 1604681595
transform 1 0 8188 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_2_
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_1__A0
timestamp 1604681595
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_2__A1
timestamp 1604681595
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_2__A0
timestamp 1604681595
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_84
timestamp 1604681595
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_88
timestamp 1604681595
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_102
timestamp 1604681595
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11408 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_106
timestamp 1604681595
transform 1 0 10856 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_128
timestamp 1604681595
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_132
timestamp 1604681595
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_145
timestamp 1604681595
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_149
timestamp 1604681595
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_163
timestamp 1604681595
transform 1 0 16100 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_4_
timestamp 1604681595
transform 1 0 17480 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 17296 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 16928 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_169
timestamp 1604681595
transform 1 0 16652 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_174
timestamp 1604681595
transform 1 0 17112 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_187
timestamp 1604681595
transform 1 0 18308 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 19044 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 18492 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 18860 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_191
timestamp 1604681595
transform 1 0 18676 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_204
timestamp 1604681595
transform 1 0 19872 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_210
timestamp 1604681595
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_224
timestamp 1604681595
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_228
timestamp 1604681595
transform 1 0 22080 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1604681595
transform 1 0 22448 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24012 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 23644 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 22264 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_241
timestamp 1604681595
transform 1 0 23276 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_247
timestamp 1604681595
transform 1 0 23828 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 25024 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 25392 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25760 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_258
timestamp 1604681595
transform 1 0 24840 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_262
timestamp 1604681595
transform 1 0 25208 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_266
timestamp 1604681595
transform 1 0 25576 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_270
timestamp 1604681595
transform 1 0 25944 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 26128 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_274
timestamp 1604681595
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604681595
transform 1 0 1840 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2852 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 2300 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 1656 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_11
timestamp 1604681595
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 4508 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_35
timestamp 1604681595
transform 1 0 4324 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_39
timestamp 1604681595
transform 1 0 4692 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5060 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6072 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_52
timestamp 1604681595
transform 1 0 5888 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_56
timestamp 1604681595
transform 1 0 6256 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 7728 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 7544 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_68
timestamp 1604681595
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_1_
timestamp 1604681595
transform 1 0 9936 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_1__S
timestamp 1604681595
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_4__D
timestamp 1604681595
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_88
timestamp 1604681595
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_92
timestamp 1604681595
transform 1 0 9568 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_109
timestamp 1604681595
transform 1 0 11132 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_105
timestamp 1604681595
transform 1 0 10764 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_1__A1
timestamp 1604681595
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1604681595
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_3_
timestamp 1604681595
transform 1 0 13524 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_127
timestamp 1604681595
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_131
timestamp 1604681595
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_144
timestamp 1604681595
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15088 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 14536 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_148
timestamp 1604681595
transform 1 0 14720 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_176
timestamp 1604681595
transform 1 0 17296 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_172
timestamp 1604681595
transform 1 0 16928 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_168
timestamp 1604681595
transform 1 0 16560 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_179
timestamp 1604681595
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 18216 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 19872 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_202
timestamp 1604681595
transform 1 0 19688 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_206
timestamp 1604681595
transform 1 0 20056 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 20792 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_210
timestamp 1604681595
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 22448 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_230
timestamp 1604681595
transform 1 0 22264 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_234
timestamp 1604681595
transform 1 0 22632 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_240
timestamp 1604681595
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604681595
transform 1 0 25208 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1604681595
transform 1 0 25760 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_254
timestamp 1604681595
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_258
timestamp 1604681595
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_266
timestamp 1604681595
transform 1 0 25576 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_270
timestamp 1604681595
transform 1 0 25944 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1604681595
transform 1 0 26128 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_274
timestamp 1604681595
transform 1 0 26312 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_10
timestamp 1604681595
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1604681595
transform 1 0 1748 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 1840 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_14
timestamp 1604681595
transform 1 0 2392 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 2576 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 2760 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 1748 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_23
timestamp 1604681595
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_38
timestamp 1604681595
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_34
timestamp 1604681595
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4416 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4600 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_51
timestamp 1604681595
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4968 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_55
timestamp 1604681595
transform 1 0 6164 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_58
timestamp 1604681595
transform 1 0 6440 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_54
timestamp 1604681595
transform 1 0 6072 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_3__A1
timestamp 1604681595
transform 1 0 6716 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_72
timestamp 1604681595
transform 1 0 7728 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_68
timestamp 1604681595
transform 1 0 7360 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_71
timestamp 1604681595
transform 1 0 7636 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_67
timestamp 1604681595
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1604681595
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7544 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1604681595
transform 1 0 6992 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604681595
transform 1 0 6900 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_3__S
timestamp 1604681595
transform 1 0 7912 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8096 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_91
timestamp 1604681595
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_85
timestamp 1604681595
transform 1 0 8924 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_88
timestamp 1604681595
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_84
timestamp 1604681595
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9844 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_111
timestamp 1604681595
transform 1 0 11316 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_113
timestamp 1604681595
transform 1 0 11500 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_109
timestamp 1604681595
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 11500 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_119
timestamp 1604681595
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_115
timestamp 1604681595
transform 1 0 11684 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_117
timestamp 1604681595
transform 1 0 11868 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11684 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12144 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 11868 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12604 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12328 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 13892 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 13340 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 13708 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 13984 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1604681595
transform 1 0 13800 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_142
timestamp 1604681595
transform 1 0 14168 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_131
timestamp 1604681595
transform 1 0 13156 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_135
timestamp 1604681595
transform 1 0 13524 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_155
timestamp 1604681595
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_149
timestamp 1604681595
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_146
timestamp 1604681595
transform 1 0 14536 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_159
timestamp 1604681595
transform 1 0 15732 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 15916 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_4_
timestamp 1604681595
transform 1 0 16100 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_7_176
timestamp 1604681595
transform 1 0 17296 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_172
timestamp 1604681595
transform 1 0 16928 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_175
timestamp 1604681595
transform 1 0 17204 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_170
timestamp 1604681595
transform 1 0 16744 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 17020 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17388 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_179
timestamp 1604681595
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_179
timestamp 1604681595
transform 1 0 17572 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 17756 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_197
timestamp 1604681595
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1604681595
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1604681595
transform 1 0 19228 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_206
timestamp 1604681595
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_201
timestamp 1604681595
transform 1 0 19596 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 19872 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19412 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 19596 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_217
timestamp 1604681595
transform 1 0 21068 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_218
timestamp 1604681595
transform 1 0 21160 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_210
timestamp 1604681595
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1604681595
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_222
timestamp 1604681595
transform 1 0 21528 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 21712 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21344 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 21252 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 21620 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21804 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 21896 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_7_238
timestamp 1604681595
transform 1 0 23000 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_234
timestamp 1604681595
transform 1 0 22632 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_247
timestamp 1604681595
transform 1 0 23828 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_242
timestamp 1604681595
transform 1 0 23368 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23644 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 24012 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_258
timestamp 1604681595
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_254
timestamp 1604681595
transform 1 0 24472 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_251
timestamp 1604681595
transform 1 0 24196 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 24656 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 24380 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_266
timestamp 1604681595
transform 1 0 25576 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_266
timestamp 1604681595
transform 1 0 25576 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_262
timestamp 1604681595
transform 1 0 25208 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 25760 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 25392 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 25024 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1604681595
transform 1 0 25760 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604681595
transform 1 0 25208 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_270
timestamp 1604681595
transform 1 0 25944 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_270
timestamp 1604681595
transform 1 0 25944 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 26128 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 26128 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_274
timestamp 1604681595
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_274
timestamp 1604681595
transform 1 0 26312 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2208 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_8
timestamp 1604681595
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_25
timestamp 1604681595
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_21
timestamp 1604681595
transform 1 0 3036 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1604681595
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_39
timestamp 1604681595
transform 1 0 4692 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_36
timestamp 1604681595
transform 1 0 4416 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4508 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5244 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_3__A0
timestamp 1604681595
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 6348 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_43
timestamp 1604681595
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_54
timestamp 1604681595
transform 1 0 6072 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_59
timestamp 1604681595
transform 1 0 6532 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1604681595
transform 1 0 6900 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_3_
timestamp 1604681595
transform 1 0 8004 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__S
timestamp 1604681595
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_67
timestamp 1604681595
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_71
timestamp 1604681595
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_7__A0
timestamp 1604681595
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1604681595
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_88
timestamp 1604681595
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_102
timestamp 1604681595
transform 1 0 10488 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1604681595
transform 1 0 11316 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12328 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 11132 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_107
timestamp 1604681595
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_120
timestamp 1604681595
transform 1 0 12144 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_124
timestamp 1604681595
transform 1 0 12512 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12880 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 13892 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 12696 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14260 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_137
timestamp 1604681595
transform 1 0 13708 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1604681595
transform 1 0 14076 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_145
timestamp 1604681595
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 16284 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_149
timestamp 1604681595
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1604681595
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 17388 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17204 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_167
timestamp 1604681595
transform 1 0 16468 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_172
timestamp 1604681595
transform 1 0 16928 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_186
timestamp 1604681595
transform 1 0 18216 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19044 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 18400 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 18768 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_190
timestamp 1604681595
transform 1 0 18584 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_194
timestamp 1604681595
transform 1 0 18952 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_204
timestamp 1604681595
transform 1 0 19872 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_208
timestamp 1604681595
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 21896 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1604681595
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_224
timestamp 1604681595
transform 1 0 21712 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_228
timestamp 1604681595
transform 1 0 22080 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1604681595
transform 1 0 22448 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 24012 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 23644 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 22264 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_241
timestamp 1604681595
transform 1 0 23276 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_247
timestamp 1604681595
transform 1 0 23828 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 25024 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 25392 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25760 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_258
timestamp 1604681595
transform 1 0 24840 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_262
timestamp 1604681595
transform 1 0 25208 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_266
timestamp 1604681595
transform 1 0 25576 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_270
timestamp 1604681595
transform 1 0 25944 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 26128 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_274
timestamp 1604681595
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_4_
timestamp 1604681595
transform 1 0 2024 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1604681595
transform 1 0 1748 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_19
timestamp 1604681595
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_23
timestamp 1604681595
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_36
timestamp 1604681595
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_40
timestamp 1604681595
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_53
timestamp 1604681595
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1604681595
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_7_
timestamp 1604681595
transform 1 0 8464 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_7__A1
timestamp 1604681595
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__A1
timestamp 1604681595
transform 1 0 7912 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_71
timestamp 1604681595
transform 1 0 7636 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_76
timestamp 1604681595
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__A0
timestamp 1604681595
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1604681595
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_89
timestamp 1604681595
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_93
timestamp 1604681595
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_97
timestamp 1604681595
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_101
timestamp 1604681595
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1604681595
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1604681595
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 14260 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 14076 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1604681595
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_136
timestamp 1604681595
transform 1 0 13616 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_140
timestamp 1604681595
transform 1 0 13984 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16284 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15916 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_159
timestamp 1604681595
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_163
timestamp 1604681595
transform 1 0 16100 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16468 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_173
timestamp 1604681595
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_177
timestamp 1604681595
transform 1 0 17388 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18584 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 20240 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_206
timestamp 1604681595
transform 1 0 20056 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1604681595
transform 1 0 20792 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 22172 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_210
timestamp 1604681595
transform 1 0 20424 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_223
timestamp 1604681595
transform 1 0 21620 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_227
timestamp 1604681595
transform 1 0 21988 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604681595
transform 1 0 22448 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1604681595
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_231
timestamp 1604681595
transform 1 0 22356 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_236
timestamp 1604681595
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_240
timestamp 1604681595
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604681595
transform 1 0 25208 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1604681595
transform 1 0 25760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_254
timestamp 1604681595
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_258
timestamp 1604681595
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_266
timestamp 1604681595
transform 1 0 25576 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_270
timestamp 1604681595
transform 1 0 25944 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 26128 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_274
timestamp 1604681595
transform 1 0 26312 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_8
timestamp 1604681595
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_12
timestamp 1604681595
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4876 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4692 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4324 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1604681595
transform 1 0 3220 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1604681595
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_37
timestamp 1604681595
transform 1 0 4508 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_57
timestamp 1604681595
transform 1 0 6348 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_61
timestamp 1604681595
transform 1 0 6716 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_6_
timestamp 1604681595
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7084 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7544 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_64
timestamp 1604681595
transform 1 0 6992 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_68
timestamp 1604681595
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_72
timestamp 1604681595
transform 1 0 7728 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_88
timestamp 1604681595
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_84
timestamp 1604681595
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_7__S
timestamp 1604681595
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604681595
transform 1 0 9844 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_99
timestamp 1604681595
transform 1 0 10212 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 10396 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_103
timestamp 1604681595
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10948 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_123
timestamp 1604681595
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13156 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14168 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_127
timestamp 1604681595
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_140
timestamp 1604681595
transform 1 0 13984 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_144
timestamp 1604681595
transform 1 0 14352 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 14536 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 16008 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_148
timestamp 1604681595
transform 1 0 14720 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_160
timestamp 1604681595
transform 1 0 15824 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_164
timestamp 1604681595
transform 1 0 16192 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 18308 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1604681595
transform 1 0 16744 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 16560 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_179
timestamp 1604681595
transform 1 0 17572 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_183
timestamp 1604681595
transform 1 0 17940 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_186
timestamp 1604681595
transform 1 0 18216 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19964 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_203
timestamp 1604681595
transform 1 0 19780 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_207
timestamp 1604681595
transform 1 0 20148 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 21804 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 21068 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 20516 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 21436 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1604681595
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_219
timestamp 1604681595
transform 1 0 21252 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_223
timestamp 1604681595
transform 1 0 21620 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24012 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_241
timestamp 1604681595
transform 1 0 23276 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_247
timestamp 1604681595
transform 1 0 23828 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25024 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 25392 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 25760 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_258
timestamp 1604681595
transform 1 0 24840 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_262
timestamp 1604681595
transform 1 0 25208 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_266
timestamp 1604681595
transform 1 0 25576 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_270
timestamp 1604681595
transform 1 0 25944 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 26128 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_274
timestamp 1604681595
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604681595
transform 1 0 1840 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2852 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 1656 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_11
timestamp 1604681595
transform 1 0 2116 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_16
timestamp 1604681595
transform 1 0 2576 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4508 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_35
timestamp 1604681595
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_39
timestamp 1604681595
transform 1 0 4692 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5060 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_52
timestamp 1604681595
transform 1 0 5888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1604681595
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8372 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_71
timestamp 1604681595
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_75
timestamp 1604681595
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 9936 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 9752 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_88
timestamp 1604681595
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_92
timestamp 1604681595
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_99
timestamp 1604681595
transform 1 0 10212 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_114
timestamp 1604681595
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_118
timestamp 1604681595
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_132
timestamp 1604681595
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_136
timestamp 1604681595
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_140
timestamp 1604681595
transform 1 0 13984 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 14904 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 14720 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_146
timestamp 1604681595
transform 1 0 14536 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_166
timestamp 1604681595
transform 1 0 16376 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 17204 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17664 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16652 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_171
timestamp 1604681595
transform 1 0 16836 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_178
timestamp 1604681595
transform 1 0 17480 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1604681595
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 19688 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_200
timestamp 1604681595
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_204
timestamp 1604681595
transform 1 0 19872 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_208
timestamp 1604681595
transform 1 0 20240 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 20516 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 20332 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 22172 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_227
timestamp 1604681595
transform 1 0 21988 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_231
timestamp 1604681595
transform 1 0 22356 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_236
timestamp 1604681595
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_240
timestamp 1604681595
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604681595
transform 1 0 25208 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1604681595
transform 1 0 24932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1604681595
transform 1 0 25760 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_254
timestamp 1604681595
transform 1 0 24472 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_258
timestamp 1604681595
transform 1 0 24840 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_261
timestamp 1604681595
transform 1 0 25116 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_266
timestamp 1604681595
transform 1 0 25576 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_270
timestamp 1604681595
transform 1 0 25944 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 26128 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_274
timestamp 1604681595
transform 1 0 26312 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1604681595
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_6
timestamp 1604681595
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_10
timestamp 1604681595
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_23
timestamp 1604681595
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_40
timestamp 1604681595
transform 1 0 4784 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_36
timestamp 1604681595
transform 1 0 4416 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 4600 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5428 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6440 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_46
timestamp 1604681595
transform 1 0 5336 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_56
timestamp 1604681595
transform 1 0 6256 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_60
timestamp 1604681595
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604681595
transform 1 0 8556 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1604681595
transform 1 0 6992 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 8004 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_73
timestamp 1604681595
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_77
timestamp 1604681595
transform 1 0 8188 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_84
timestamp 1604681595
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_88
timestamp 1604681595
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604681595
transform 1 0 9752 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_97
timestamp 1604681595
transform 1 0 10028 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_101
timestamp 1604681595
transform 1 0 10396 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 10212 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 10580 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10764 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_121
timestamp 1604681595
transform 1 0 12236 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_125
timestamp 1604681595
transform 1 0 12604 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1604681595
transform 1 0 12972 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1604681595
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_142
timestamp 1604681595
transform 1 0 14168 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_146
timestamp 1604681595
transform 1 0 14536 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_149
timestamp 1604681595
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_163
timestamp 1604681595
transform 1 0 16100 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 17112 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 16744 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 18124 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_168
timestamp 1604681595
transform 1 0 16560 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_172
timestamp 1604681595
transform 1 0 16928 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_183
timestamp 1604681595
transform 1 0 17940 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_187
timestamp 1604681595
transform 1 0 18308 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18676 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 20240 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 18492 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 19688 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_200
timestamp 1604681595
transform 1 0 19504 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_204
timestamp 1604681595
transform 1 0 19872 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_3_
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_211
timestamp 1604681595
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_224
timestamp 1604681595
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_228
timestamp 1604681595
transform 1 0 22080 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 22724 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 22264 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_232
timestamp 1604681595
transform 1 0 22448 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604681595
transform 1 0 24932 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 24380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 24748 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25484 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 25852 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_251
timestamp 1604681595
transform 1 0 24196 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_255
timestamp 1604681595
transform 1 0 24564 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_263
timestamp 1604681595
transform 1 0 25300 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_267
timestamp 1604681595
transform 1 0 25668 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_271
timestamp 1604681595
transform 1 0 26036 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_7
timestamp 1604681595
transform 1 0 1748 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_7
timestamp 1604681595
transform 1 0 1748 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 2024 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_11
timestamp 1604681595
transform 1 0 2116 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_16
timestamp 1604681595
transform 1 0 2576 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_12
timestamp 1604681595
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 2668 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1604681595
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_40
timestamp 1604681595
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_37
timestamp 1604681595
transform 1 0 4508 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_33
timestamp 1604681595
transform 1 0 4140 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4600 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_51
timestamp 1604681595
transform 1 0 5796 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_47
timestamp 1604681595
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 5612 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1604681595
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_53
timestamp 1604681595
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 5980 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 6164 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604681595
transform 1 0 8372 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 7452 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 7268 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_66
timestamp 1604681595
transform 1 0 7176 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_71
timestamp 1604681595
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_75
timestamp 1604681595
transform 1 0 8004 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_82
timestamp 1604681595
transform 1 0 8648 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_87
timestamp 1604681595
transform 1 0 9108 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_90
timestamp 1604681595
transform 1 0 9384 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_85
timestamp 1604681595
transform 1 0 8924 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9200 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 8924 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_102
timestamp 1604681595
transform 1 0 10488 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_101
timestamp 1604681595
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_97
timestamp 1604681595
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604681595
transform 1 0 9752 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_113
timestamp 1604681595
transform 1 0 11500 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_107
timestamp 1604681595
transform 1 0 10948 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_114
timestamp 1604681595
transform 1 0 11592 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 11316 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_13_119
timestamp 1604681595
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11868 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 11684 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11868 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_133
timestamp 1604681595
transform 1 0 13340 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_137
timestamp 1604681595
transform 1 0 13708 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_139
timestamp 1604681595
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 13892 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 13524 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_143
timestamp 1604681595
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1604681595
transform 1 0 14076 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604681595
transform 1 0 14076 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_145
timestamp 1604681595
transform 1 0 14444 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14444 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1604681595
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 14628 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_158
timestamp 1604681595
transform 1 0 15640 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_162
timestamp 1604681595
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_156
timestamp 1604681595
transform 1 0 15456 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 16008 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 15456 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 16192 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_4_
timestamp 1604681595
transform 1 0 16376 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_173
timestamp 1604681595
transform 1 0 17020 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_175
timestamp 1604681595
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17204 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_177
timestamp 1604681595
transform 1 0 17388 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_179
timestamp 1604681595
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 17572 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 18216 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 17756 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1604681595
transform 1 0 18952 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_190
timestamp 1604681595
transform 1 0 18584 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_188
timestamp 1604681595
transform 1 0 18400 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 19136 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 18768 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 18492 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_206
timestamp 1604681595
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_201
timestamp 1604681595
transform 1 0 19596 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_202
timestamp 1604681595
transform 1 0 19688 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_198
timestamp 1604681595
transform 1 0 19320 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1604681595
transform 1 0 19504 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 19320 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_3_
timestamp 1604681595
transform 1 0 20056 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604681595
transform 1 0 19688 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 20240 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_210
timestamp 1604681595
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_215
timestamp 1604681595
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21068 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_228
timestamp 1604681595
transform 1 0 22080 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_224
timestamp 1604681595
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_219
timestamp 1604681595
transform 1 0 21252 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21620 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_239
timestamp 1604681595
transform 1 0 23092 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_235
timestamp 1604681595
transform 1 0 22724 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_236
timestamp 1604681595
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_232
timestamp 1604681595
transform 1 0 22448 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 22908 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 22264 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_4__D
timestamp 1604681595
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 22632 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604681595
transform 1 0 22448 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_240
timestamp 1604681595
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23276 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 23460 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_259
timestamp 1604681595
transform 1 0 24932 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_261
timestamp 1604681595
transform 1 0 25116 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 25116 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_263
timestamp 1604681595
transform 1 0 25300 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25300 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_267
timestamp 1604681595
transform 1 0 25668 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_265
timestamp 1604681595
transform 1 0 25484 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 25668 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 25484 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_269
timestamp 1604681595
transform 1 0 25852 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1604681595
transform 1 0 26036 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_273
timestamp 1604681595
transform 1 0 26220 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_271
timestamp 1604681595
transform 1 0 26036 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_3_
timestamp 1604681595
transform 1 0 2208 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 2024 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 1656 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_8
timestamp 1604681595
transform 1 0 1840 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 3772 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 3588 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_21
timestamp 1604681595
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_25
timestamp 1604681595
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_49
timestamp 1604681595
transform 1 0 5612 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_45
timestamp 1604681595
transform 1 0 5244 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 5428 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1604681595
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_53
timestamp 1604681595
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 8372 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_71
timestamp 1604681595
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_75
timestamp 1604681595
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_82
timestamp 1604681595
transform 1 0 8648 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8924 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_101
timestamp 1604681595
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1604681595
transform 1 0 11316 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_105
timestamp 1604681595
transform 1 0 10764 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_114
timestamp 1604681595
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_118
timestamp 1604681595
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_132
timestamp 1604681595
transform 1 0 13248 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_138
timestamp 1604681595
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_142
timestamp 1604681595
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 14812 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_146
timestamp 1604681595
transform 1 0 14536 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_158
timestamp 1604681595
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_162
timestamp 1604681595
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 18216 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1604681595
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 1604681595
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604681595
transform 1 0 18400 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 19504 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1604681595
transform 1 0 18952 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 19320 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_192
timestamp 1604681595
transform 1 0 18768 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_196
timestamp 1604681595
transform 1 0 19136 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1604681595
transform 1 0 21712 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 21528 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_216
timestamp 1604681595
transform 1 0 20976 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_220
timestamp 1604681595
transform 1 0 21344 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1604681595
transform 1 0 22724 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_233
timestamp 1604681595
transform 1 0 22540 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_237
timestamp 1604681595
transform 1 0 22908 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_241
timestamp 1604681595
transform 1 0 23276 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 24656 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 25024 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_254
timestamp 1604681595
transform 1 0 24472 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_258
timestamp 1604681595
transform 1 0 24840 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_268
timestamp 1604681595
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 26312 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_272
timestamp 1604681595
transform 1 0 26128 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_276
timestamp 1604681595
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 1564 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1604681595
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_25
timestamp 1604681595
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_21
timestamp 1604681595
transform 1 0 3036 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l5_in_0__A1
timestamp 1604681595
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_36
timestamp 1604681595
transform 1 0 4416 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 4508 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4692 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 6716 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6348 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_55
timestamp 1604681595
transform 1 0 6164 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_59
timestamp 1604681595
transform 1 0 6532 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604681595
transform 1 0 8556 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6900 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 8004 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_72
timestamp 1604681595
transform 1 0 7728 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_77
timestamp 1604681595
transform 1 0 8188 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_3_
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_84
timestamp 1604681595
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_88
timestamp 1604681595
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_102
timestamp 1604681595
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1604681595
transform 1 0 11684 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 11500 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_106
timestamp 1604681595
transform 1 0 10856 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_111
timestamp 1604681595
transform 1 0 11316 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_124
timestamp 1604681595
transform 1 0 12512 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12788 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13616 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_145
timestamp 1604681595
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_149
timestamp 1604681595
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 17940 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16928 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 17296 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1604681595
transform 1 0 16744 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_174
timestamp 1604681595
transform 1 0 17112 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_178
timestamp 1604681595
transform 1 0 17480 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 19872 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_199
timestamp 1604681595
transform 1 0 19412 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_203
timestamp 1604681595
transform 1 0 19780 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_206
timestamp 1604681595
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_210
timestamp 1604681595
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_224
timestamp 1604681595
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_228
timestamp 1604681595
transform 1 0 22080 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1604681595
transform 1 0 22448 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 23552 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 22264 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 23000 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_236
timestamp 1604681595
transform 1 0 22816 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_240
timestamp 1604681595
transform 1 0 23184 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 25208 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 25576 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 25944 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_260
timestamp 1604681595
transform 1 0 25024 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_264
timestamp 1604681595
transform 1 0 25392 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_268
timestamp 1604681595
transform 1 0 25760 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_272
timestamp 1604681595
transform 1 0 26128 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2116 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_4__D
timestamp 1604681595
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l5_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_27
timestamp 1604681595
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_31
timestamp 1604681595
transform 1 0 3956 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_36
timestamp 1604681595
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_40
timestamp 1604681595
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_53
timestamp 1604681595
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1604681595
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8004 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_65
timestamp 1604681595
transform 1 0 7084 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_71
timestamp 1604681595
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_2_
timestamp 1604681595
transform 1 0 10212 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_91
timestamp 1604681595
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_95
timestamp 1604681595
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_108
timestamp 1604681595
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_112
timestamp 1604681595
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_116
timestamp 1604681595
transform 1 0 11776 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 14076 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_139
timestamp 1604681595
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_143
timestamp 1604681595
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_2_
timestamp 1604681595
transform 1 0 14628 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_156
timestamp 1604681595
transform 1 0 15456 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_162
timestamp 1604681595
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1604681595
transform 1 0 17480 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_175
timestamp 1604681595
transform 1 0 17204 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_180
timestamp 1604681595
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 20240 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 20056 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 19688 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_200
timestamp 1604681595
transform 1 0 19504 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_204
timestamp 1604681595
transform 1 0 19872 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1604681595
transform 1 0 21804 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 21620 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_217
timestamp 1604681595
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1604681595
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_234
timestamp 1604681595
transform 1 0 22632 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_238
timestamp 1604681595
transform 1 0 23000 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604681595
transform 1 0 25208 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 24656 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 25760 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_254
timestamp 1604681595
transform 1 0 24472 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_258
timestamp 1604681595
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_266
timestamp 1604681595
transform 1 0 25576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_270
timestamp 1604681595
transform 1 0 25944 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 26128 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_274
timestamp 1604681595
transform 1 0 26312 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 1748 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l5_in_0__S
timestamp 1604681595
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1604681595
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_36
timestamp 1604681595
transform 1 0 4416 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4232 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4692 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_41
timestamp 1604681595
transform 1 0 4876 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 6532 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4968 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5980 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 6348 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_51
timestamp 1604681595
transform 1 0 5796 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_55
timestamp 1604681595
transform 1 0 6164 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_75
timestamp 1604681595
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_79
timestamp 1604681595
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_83
timestamp 1604681595
transform 1 0 8740 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_88
timestamp 1604681595
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1604681595
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11132 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_106
timestamp 1604681595
transform 1 0 10856 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_118
timestamp 1604681595
transform 1 0 11960 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_122
timestamp 1604681595
transform 1 0 12328 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_125
timestamp 1604681595
transform 1 0 12604 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12696 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_146
timestamp 1604681595
transform 1 0 14536 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1604681595
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604681595
transform 1 0 17480 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 18032 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16928 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17296 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_170
timestamp 1604681595
transform 1 0 16744 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_174
timestamp 1604681595
transform 1 0 17112 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_182
timestamp 1604681595
transform 1 0 17848 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_186
timestamp 1604681595
transform 1 0 18216 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18584 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 19596 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_199
timestamp 1604681595
transform 1 0 19412 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_203
timestamp 1604681595
transform 1 0 19780 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_207
timestamp 1604681595
transform 1 0 20148 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 21988 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 21620 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1604681595
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_210
timestamp 1604681595
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_219
timestamp 1604681595
transform 1 0 21252 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_225
timestamp 1604681595
transform 1 0 21804 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 23644 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 24012 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_243
timestamp 1604681595
transform 1 0 23460 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_247
timestamp 1604681595
transform 1 0 23828 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l4_in_0_
timestamp 1604681595
transform 1 0 24196 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1604681595
transform 1 0 25208 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 25576 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 25944 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_260
timestamp 1604681595
transform 1 0 25024 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_264
timestamp 1604681595
transform 1 0 25392 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_268
timestamp 1604681595
transform 1 0 25760 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_272
timestamp 1604681595
transform 1 0 26128 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_7
timestamp 1604681595
transform 1 0 1748 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l5_in_0_
timestamp 1604681595
transform 1 0 1564 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_11
timestamp 1604681595
transform 1 0 2116 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_18
timestamp 1604681595
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_14
timestamp 1604681595
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 2944 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_1_
timestamp 1604681595
transform 1 0 3128 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_35
timestamp 1604681595
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_31
timestamp 1604681595
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4140 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4692 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_41
timestamp 1604681595
transform 1 0 4876 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_49
timestamp 1604681595
transform 1 0 5612 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_45
timestamp 1604681595
transform 1 0 5244 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_52
timestamp 1604681595
transform 1 0 5888 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_48
timestamp 1604681595
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 5428 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 5060 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 5704 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_53
timestamp 1604681595
transform 1 0 5980 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_60
timestamp 1604681595
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_56
timestamp 1604681595
transform 1 0 6256 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6256 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 6072 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 6440 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_2_
timestamp 1604681595
transform 1 0 6440 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8464 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_78
timestamp 1604681595
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_82
timestamp 1604681595
transform 1 0 8648 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_67
timestamp 1604681595
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_71
timestamp 1604681595
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_88
timestamp 1604681595
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1604681595
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8832 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9016 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_102
timestamp 1604681595
transform 1 0 10488 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_99
timestamp 1604681595
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_95
timestamp 1604681595
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10580 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_111
timestamp 1604681595
transform 1 0 11316 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_107
timestamp 1604681595
transform 1 0 10948 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_112
timestamp 1604681595
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11132 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_116
timestamp 1604681595
transform 1 0 11776 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 11408 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_132
timestamp 1604681595
transform 1 0 13248 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_128
timestamp 1604681595
transform 1 0 12880 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 13064 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_143
timestamp 1604681595
transform 1 0 14260 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_139
timestamp 1604681595
transform 1 0 13892 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14076 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_145
timestamp 1604681595
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 14444 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 14628 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 16284 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_163
timestamp 1604681595
transform 1 0 16100 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_149
timestamp 1604681595
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_170
timestamp 1604681595
transform 1 0 16744 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_171
timestamp 1604681595
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_167
timestamp 1604681595
transform 1 0 16468 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_174
timestamp 1604681595
transform 1 0 17112 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_175
timestamp 1604681595
transform 1 0 17204 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 17296 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 16928 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1604681595
transform 1 0 16928 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_180
timestamp 1604681595
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1604681595
transform 1 0 17480 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604681595
transform 1 0 17480 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_186
timestamp 1604681595
transform 1 0 18216 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_182
timestamp 1604681595
transform 1 0 17848 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 18216 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_197
timestamp 1604681595
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 18400 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18400 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_206
timestamp 1604681595
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_201
timestamp 1604681595
transform 1 0 19596 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1604681595
transform 1 0 19872 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604681595
transform 1 0 20056 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18584 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 20608 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_210
timestamp 1604681595
transform 1 0 20424 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_210
timestamp 1604681595
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 20976 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 21160 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_214
timestamp 1604681595
transform 1 0 20792 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1604681595
transform 1 0 21160 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_220
timestamp 1604681595
transform 1 0 21344 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_227
timestamp 1604681595
transform 1 0 21988 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21620 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 22172 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_236
timestamp 1604681595
transform 1 0 22816 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_232
timestamp 1604681595
transform 1 0 22448 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_239
timestamp 1604681595
transform 1 0 23092 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_235
timestamp 1604681595
transform 1 0 22724 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_231
timestamp 1604681595
transform 1 0 22356 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 22632 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 23000 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 22540 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_242
timestamp 1604681595
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 23184 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_256
timestamp 1604681595
transform 1 0 24656 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_260
timestamp 1604681595
transform 1 0 25024 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_261
timestamp 1604681595
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 24840 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_265
timestamp 1604681595
transform 1 0 25484 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25208 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604681595
transform 1 0 25392 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_267
timestamp 1604681595
transform 1 0 25668 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_269
timestamp 1604681595
transform 1 0 25852 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 25852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 25668 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 26220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 26036 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 26404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_273
timestamp 1604681595
transform 1 0 26220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_271
timestamp 1604681595
transform 1 0 26036 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 2760 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_1__S
timestamp 1604681595
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_10
timestamp 1604681595
transform 1 0 2024 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_14
timestamp 1604681595
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_34
timestamp 1604681595
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_38
timestamp 1604681595
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4968 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1604681595
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8556 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1604681595
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_75
timestamp 1604681595
transform 1 0 8004 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_97
timestamp 1604681595
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_101
timestamp 1604681595
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1604681595
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_2_
timestamp 1604681595
transform 1 0 13984 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1604681595
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_136
timestamp 1604681595
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_1_
timestamp 1604681595
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_149
timestamp 1604681595
transform 1 0 14812 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_153
timestamp 1604681595
transform 1 0 15180 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_156
timestamp 1604681595
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_160
timestamp 1604681595
transform 1 0 15824 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_175
timestamp 1604681595
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_179
timestamp 1604681595
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1604681595
transform 1 0 19688 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_200
timestamp 1604681595
transform 1 0 19504 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_204
timestamp 1604681595
transform 1 0 19872 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_208
timestamp 1604681595
transform 1 0 20240 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20700 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20332 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 21896 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_211
timestamp 1604681595
transform 1 0 20516 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_224
timestamp 1604681595
transform 1 0 21712 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_228
timestamp 1604681595
transform 1 0 22080 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604681595
transform 1 0 22448 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1604681595
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 22264 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_236
timestamp 1604681595
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_240
timestamp 1604681595
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 24656 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 25024 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_254
timestamp 1604681595
transform 1 0 24472 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_258
timestamp 1604681595
transform 1 0 24840 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_268
timestamp 1604681595
transform 1 0 25760 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 26312 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_272
timestamp 1604681595
transform 1 0 26128 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_276
timestamp 1604681595
transform 1 0 26496 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1604681595
transform 1 0 2944 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_1_
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2392 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 2760 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_12
timestamp 1604681595
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_16
timestamp 1604681595
transform 1 0 2576 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_1__A1
timestamp 1604681595
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_1__A0
timestamp 1604681595
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6716 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_3__A1
timestamp 1604681595
transform 1 0 5704 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_3__A0
timestamp 1604681595
transform 1 0 6072 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_48
timestamp 1604681595
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_52
timestamp 1604681595
transform 1 0 5888 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_56
timestamp 1604681595
transform 1 0 6256 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_77
timestamp 1604681595
transform 1 0 8188 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_81
timestamp 1604681595
transform 1 0 8556 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 8924 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_88
timestamp 1604681595
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_102
timestamp 1604681595
transform 1 0 10488 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1604681595
transform 1 0 11224 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10764 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_107
timestamp 1604681595
transform 1 0 10948 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_119
timestamp 1604681595
transform 1 0 12052 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_125
timestamp 1604681595
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_3_
timestamp 1604681595
transform 1 0 12788 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 13984 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 14352 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1604681595
transform 1 0 13616 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_142
timestamp 1604681595
transform 1 0 14168 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_3_
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 16376 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_146
timestamp 1604681595
transform 1 0 14536 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_150
timestamp 1604681595
transform 1 0 14904 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_163
timestamp 1604681595
transform 1 0 16100 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 17112 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 16836 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_168
timestamp 1604681595
transform 1 0 16560 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604681595
transform 1 0 19688 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 19412 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 18768 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 19228 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_190
timestamp 1604681595
transform 1 0 18584 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_194
timestamp 1604681595
transform 1 0 18952 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_206
timestamp 1604681595
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 21620 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21068 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21436 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_210
timestamp 1604681595
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_219
timestamp 1604681595
transform 1 0 21252 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23828 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 23644 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 23276 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_239
timestamp 1604681595
transform 1 0 23092 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_243
timestamp 1604681595
transform 1 0 23460 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1604681595
transform 1 0 25392 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25208 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 24840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 25852 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_256
timestamp 1604681595
transform 1 0 24656 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_260
timestamp 1604681595
transform 1 0 25024 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_267
timestamp 1604681595
transform 1 0 25668 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 26220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_271
timestamp 1604681595
transform 1 0 26036 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2392 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_4__S
timestamp 1604681595
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_3__S
timestamp 1604681595
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_7
timestamp 1604681595
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_11
timestamp 1604681595
transform 1 0 2116 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 4508 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 4324 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_23
timestamp 1604681595
transform 1 0 3220 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_29
timestamp 1604681595
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_33
timestamp 1604681595
transform 1 0 4140 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8372 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_71
timestamp 1604681595
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_75
timestamp 1604681595
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9936 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9752 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_88
timestamp 1604681595
transform 1 0 9200 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_92
timestamp 1604681595
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_105
timestamp 1604681595
transform 1 0 10764 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 10948 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_109
timestamp 1604681595
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 11500 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_116
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1604681595
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604681595
transform 1 0 12880 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13892 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 13708 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 12696 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_131
timestamp 1604681595
transform 1 0 13156 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_135
timestamp 1604681595
transform 1 0 13524 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_148
timestamp 1604681595
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_152
timestamp 1604681595
transform 1 0 15088 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_156
timestamp 1604681595
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_160
timestamp 1604681595
transform 1 0 15824 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_2_
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_175
timestamp 1604681595
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1604681595
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l4_in_0_
timestamp 1604681595
transform 1 0 19596 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_193
timestamp 1604681595
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_197
timestamp 1604681595
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21160 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 22172 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20976 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_210
timestamp 1604681595
transform 1 0 20424 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_214
timestamp 1604681595
transform 1 0 20792 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_227
timestamp 1604681595
transform 1 0 21988 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_2_
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 22632 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_231
timestamp 1604681595
transform 1 0 22356 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_236
timestamp 1604681595
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_240
timestamp 1604681595
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1604681595
transform 1 0 25944 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_254
timestamp 1604681595
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_258
timestamp 1604681595
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_268
timestamp 1604681595
transform 1 0 25760 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 26312 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_272
timestamp 1604681595
transform 1 0 26128 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_276
timestamp 1604681595
transform 1 0 26496 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_3_
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_2__S
timestamp 1604681595
transform 1 0 2392 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2944 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_12
timestamp 1604681595
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_16
timestamp 1604681595
transform 1 0 2576 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4324 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3312 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3680 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_22
timestamp 1604681595
transform 1 0 3128 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1604681595
transform 1 0 3496 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_30
timestamp 1604681595
transform 1 0 3864 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6532 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 5980 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_2__A1
timestamp 1604681595
transform 1 0 6348 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_51
timestamp 1604681595
transform 1 0 5796 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_55
timestamp 1604681595
transform 1 0 6164 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8096 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7912 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_68
timestamp 1604681595
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_72
timestamp 1604681595
transform 1 0 7728 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1604681595
transform 1 0 8648 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10212 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10580 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1604681595
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_86
timestamp 1604681595
transform 1 0 9016 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_97
timestamp 1604681595
transform 1 0 10028 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_101
timestamp 1604681595
transform 1 0 10396 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10856 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11868 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_105
timestamp 1604681595
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_115
timestamp 1604681595
transform 1 0 11684 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_119
timestamp 1604681595
transform 1 0 12052 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_125
timestamp 1604681595
transform 1 0 12604 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12880 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_144
timestamp 1604681595
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 16284 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14536 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_148
timestamp 1604681595
transform 1 0 14720 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_163
timestamp 1604681595
transform 1 0 16100 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_3_
timestamp 1604681595
transform 1 0 17020 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 16836 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_167
timestamp 1604681595
transform 1 0 16468 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_182
timestamp 1604681595
transform 1 0 17848 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_186
timestamp 1604681595
transform 1 0 18216 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18584 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18400 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1604681595
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 21344 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 21160 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_210
timestamp 1604681595
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23552 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 23368 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 23000 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_236
timestamp 1604681595
transform 1 0 22816 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_240
timestamp 1604681595
transform 1 0 23184 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604681595
transform 1 0 25116 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 24564 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 24932 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 25668 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1604681595
transform 1 0 24380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_257
timestamp 1604681595
transform 1 0 24748 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_265
timestamp 1604681595
transform 1 0 25484 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_269
timestamp 1604681595
transform 1 0 25852 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 26036 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_273
timestamp 1604681595
transform 1 0 26220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_2_
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2944 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_4__A1
timestamp 1604681595
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_4__A0
timestamp 1604681595
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_12
timestamp 1604681595
transform 1 0 2208 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_16
timestamp 1604681595
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4416 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_26
timestamp 1604681595
transform 1 0 3496 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_32
timestamp 1604681595
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 5612 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_45
timestamp 1604681595
transform 1 0 5244 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_51
timestamp 1604681595
transform 1 0 5796 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_55
timestamp 1604681595
transform 1 0 6164 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8280 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7544 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7912 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_68
timestamp 1604681595
transform 1 0 7360 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_72
timestamp 1604681595
transform 1 0 7728 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_76
timestamp 1604681595
transform 1 0 8096 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 10488 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_94
timestamp 1604681595
transform 1 0 9752 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_98
timestamp 1604681595
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12052 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_111
timestamp 1604681595
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_115
timestamp 1604681595
transform 1 0 11684 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1604681595
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 13708 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_126
timestamp 1604681595
transform 1 0 12696 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_130
timestamp 1604681595
transform 1 0 13064 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_134
timestamp 1604681595
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 15916 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 15732 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 15364 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_153
timestamp 1604681595
transform 1 0 15180 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_157
timestamp 1604681595
transform 1 0 15548 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 17480 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17296 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_170
timestamp 1604681595
transform 1 0 16744 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_174
timestamp 1604681595
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_181
timestamp 1604681595
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19596 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_193
timestamp 1604681595
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_197
timestamp 1604681595
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l4_in_0_
timestamp 1604681595
transform 1 0 21804 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 21620 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 21252 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_217
timestamp 1604681595
transform 1 0 21068 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1604681595
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_3_
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_234
timestamp 1604681595
transform 1 0 22632 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_240
timestamp 1604681595
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604681595
transform 1 0 25208 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1604681595
transform 1 0 25760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 24656 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 25024 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_254
timestamp 1604681595
transform 1 0 24472 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_258
timestamp 1604681595
transform 1 0 24840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_266
timestamp 1604681595
transform 1 0 25576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_270
timestamp 1604681595
transform 1 0 25944 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 26128 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_274
timestamp 1604681595
transform 1 0 26312 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_5_
timestamp 1604681595
transform 1 0 1564 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_4_
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_18
timestamp 1604681595
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_14
timestamp 1604681595
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_16
timestamp 1604681595
transform 1 0 2576 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_12
timestamp 1604681595
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__S
timestamp 1604681595
transform 1 0 2760 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A1
timestamp 1604681595
transform 1 0 2392 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A0
timestamp 1604681595
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A1
timestamp 1604681595
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604681595
transform 1 0 2944 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_23
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__S
timestamp 1604681595
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 3128 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_35
timestamp 1604681595
transform 1 0 4324 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_31
timestamp 1604681595
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4140 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4508 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4692 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_41
timestamp 1604681595
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_48
timestamp 1604681595
transform 1 0 5520 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_45
timestamp 1604681595
transform 1 0 5244 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5428 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_3__S
timestamp 1604681595
transform 1 0 5704 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5612 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_27_56
timestamp 1604681595
transform 1 0 6256 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_52
timestamp 1604681595
transform 1 0 5888 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_58
timestamp 1604681595
transform 1 0 6440 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_2__A0
timestamp 1604681595
transform 1 0 6624 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 6072 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_62
timestamp 1604681595
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_70
timestamp 1604681595
transform 1 0 7544 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_66
timestamp 1604681595
transform 1 0 7176 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1604681595
transform 1 0 7360 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7176 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_80
timestamp 1604681595
transform 1 0 8464 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_75
timestamp 1604681595
transform 1 0 8004 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7912 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 8280 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8096 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_89
timestamp 1604681595
transform 1 0 9292 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_85
timestamp 1604681595
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_88
timestamp 1604681595
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_84
timestamp 1604681595
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_3__A0
timestamp 1604681595
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_3__A1
timestamp 1604681595
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1604681595
transform 1 0 9108 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 9660 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1604681595
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_109
timestamp 1604681595
transform 1 0 11132 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_113
timestamp 1604681595
transform 1 0 11500 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_109
timestamp 1604681595
transform 1 0 11132 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11316 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11316 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_117
timestamp 1604681595
transform 1 0 11868 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_117
timestamp 1604681595
transform 1 0 11868 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 11684 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12052 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12696 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12880 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_141
timestamp 1604681595
transform 1 0 14076 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_137
timestamp 1604681595
transform 1 0 13708 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_139
timestamp 1604681595
transform 1 0 13892 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_135
timestamp 1604681595
transform 1 0 13524 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14260 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13708 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_145
timestamp 1604681595
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 14444 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_156
timestamp 1604681595
transform 1 0 15456 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_151
timestamp 1604681595
transform 1 0 14996 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_149
timestamp 1604681595
transform 1 0 14812 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1604681595
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1604681595
transform 1 0 14628 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15732 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1604681595
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_176
timestamp 1604681595
transform 1 0 17296 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_170
timestamp 1604681595
transform 1 0 16744 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 17112 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_179
timestamp 1604681595
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_186
timestamp 1604681595
transform 1 0 18216 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_181
timestamp 1604681595
transform 1 0 17756 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604681595
transform 1 0 17480 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18492 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_1_
timestamp 1604681595
transform 1 0 19596 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 19412 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_205
timestamp 1604681595
transform 1 0 19964 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_193
timestamp 1604681595
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_197
timestamp 1604681595
transform 1 0 19228 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_217
timestamp 1604681595
transform 1 0 21068 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_214
timestamp 1604681595
transform 1 0 20792 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_210
timestamp 1604681595
transform 1 0 20424 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_210
timestamp 1604681595
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21160 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1604681595
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 21620 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21252 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_1_
timestamp 1604681595
transform 1 0 21804 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 21344 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_27_234
timestamp 1604681595
transform 1 0 22632 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_236
timestamp 1604681595
transform 1 0 22816 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23000 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_240
timestamp 1604681595
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_240
timestamp 1604681595
transform 1 0 23184 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 23368 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23552 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_254
timestamp 1604681595
transform 1 0 24472 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1604681595
transform 1 0 24380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 24564 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 24656 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_258
timestamp 1604681595
transform 1 0 24840 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_257
timestamp 1604681595
transform 1 0 24748 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 24932 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 25024 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25116 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_268
timestamp 1604681595
transform 1 0 25760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_267
timestamp 1604681595
transform 1 0 25668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 26312 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 26220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_271
timestamp 1604681595
transform 1 0 26036 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_272
timestamp 1604681595
transform 1 0 26128 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_276
timestamp 1604681595
transform 1 0 26496 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_4_
timestamp 1604681595
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A0
timestamp 1604681595
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_7
timestamp 1604681595
transform 1 0 1748 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_12
timestamp 1604681595
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_3_
timestamp 1604681595
transform 1 0 4508 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A1
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__S
timestamp 1604681595
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_23
timestamp 1604681595
transform 1 0 3220 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1604681595
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_36
timestamp 1604681595
transform 1 0 4416 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6072 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 5520 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 5888 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_46
timestamp 1604681595
transform 1 0 5336 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_50
timestamp 1604681595
transform 1 0 5704 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604681595
transform 1 0 8280 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_4__D
timestamp 1604681595
transform 1 0 7728 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8096 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_70
timestamp 1604681595
transform 1 0 7544 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_74
timestamp 1604681595
transform 1 0 7912 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1604681595
transform 1 0 8648 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1604681595
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_86
timestamp 1604681595
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_2__A1
timestamp 1604681595
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_1__A1
timestamp 1604681595
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_100
timestamp 1604681595
transform 1 0 10304 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_96
timestamp 1604681595
transform 1 0 9936 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 10120 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10672 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12604 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 11684 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12052 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_113
timestamp 1604681595
transform 1 0 11500 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_117
timestamp 1604681595
transform 1 0 11868 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_121
timestamp 1604681595
transform 1 0 12236 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604681595
transform 1 0 14168 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 13984 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 13616 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_134
timestamp 1604681595
transform 1 0 13432 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1604681595
transform 1 0 13800 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_145
timestamp 1604681595
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 16284 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14628 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_149
timestamp 1604681595
transform 1 0 14812 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_163
timestamp 1604681595
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 17112 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 16744 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_167
timestamp 1604681595
transform 1 0 16468 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_172
timestamp 1604681595
transform 1 0 16928 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19320 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 18952 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_190
timestamp 1604681595
transform 1 0 18584 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_196
timestamp 1604681595
transform 1 0 19136 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_204
timestamp 1604681595
transform 1 0 19872 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_208
timestamp 1604681595
transform 1 0 20240 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21252 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21068 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_228
timestamp 1604681595
transform 1 0 22080 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1604681595
transform 1 0 22816 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 23828 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 22448 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_234
timestamp 1604681595
transform 1 0 22632 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_245
timestamp 1604681595
transform 1 0 23644 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_249
timestamp 1604681595
transform 1 0 24012 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_3_
timestamp 1604681595
transform 1 0 24380 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 24196 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_2__A0
timestamp 1604681595
transform 1 0 25392 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 25760 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_262
timestamp 1604681595
transform 1 0 25208 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_266
timestamp 1604681595
transform 1 0 25576 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_270
timestamp 1604681595
transform 1 0 25944 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 26128 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_274
timestamp 1604681595
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 2024 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_7
timestamp 1604681595
transform 1 0 1748 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_19
timestamp 1604681595
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_6_
timestamp 1604681595
transform 1 0 3588 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A0
timestamp 1604681595
transform 1 0 3404 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1604681595
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3036 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_23
timestamp 1604681595
transform 1 0 3220 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_36
timestamp 1604681595
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_40
timestamp 1604681595
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_2_
timestamp 1604681595
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_2__S
timestamp 1604681595
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_1__S
timestamp 1604681595
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1604681595
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1604681595
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8556 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6992 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 8372 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_73
timestamp 1604681595
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_77
timestamp 1604681595
transform 1 0 8188 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10120 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9936 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9568 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_90
timestamp 1604681595
transform 1 0 9384 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_94
timestamp 1604681595
transform 1 0 9752 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1604681595
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604681595
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13984 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_132
timestamp 1604681595
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_136
timestamp 1604681595
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_2_
timestamp 1604681595
transform 1 0 16192 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1604681595
transform 1 0 15640 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 16008 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 14996 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_149
timestamp 1604681595
transform 1 0 14812 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_153
timestamp 1604681595
transform 1 0 15180 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_157
timestamp 1604681595
transform 1 0 15548 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_160
timestamp 1604681595
transform 1 0 15824 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_173
timestamp 1604681595
transform 1 0 17020 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_179
timestamp 1604681595
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19596 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_193
timestamp 1604681595
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_197
timestamp 1604681595
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_3_
timestamp 1604681595
transform 1 0 21160 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 20976 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 20608 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_210
timestamp 1604681595
transform 1 0 20424 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_214
timestamp 1604681595
transform 1 0 20792 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_227
timestamp 1604681595
transform 1 0 21988 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 22448 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_231
timestamp 1604681595
transform 1 0 22356 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_234
timestamp 1604681595
transform 1 0 22632 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_238
timestamp 1604681595
transform 1 0 23000 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_2__S
timestamp 1604681595
transform 1 0 24656 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 25024 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_254
timestamp 1604681595
transform 1 0 24472 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_258
timestamp 1604681595
transform 1 0 24840 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_268
timestamp 1604681595
transform 1 0 25760 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 26312 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_272
timestamp 1604681595
transform 1 0 26128 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_276
timestamp 1604681595
transform 1 0 26496 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2208 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 1840 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_7
timestamp 1604681595
transform 1 0 1748 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_10
timestamp 1604681595
transform 1 0 2024 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4600 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_23
timestamp 1604681595
transform 1 0 3220 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1604681595
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_36
timestamp 1604681595
transform 1 0 4416 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_40
timestamp 1604681595
transform 1 0 4784 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_1_
timestamp 1604681595
transform 1 0 5336 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 5152 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 6348 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6716 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_55
timestamp 1604681595
transform 1 0 6164 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_59
timestamp 1604681595
transform 1 0 6532 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 6900 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 8556 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_79
timestamp 1604681595
transform 1 0 8372 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_83
timestamp 1604681595
transform 1 0 8740 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_87
timestamp 1604681595
transform 1 0 9108 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 8924 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 1604681595
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_2__A0
timestamp 1604681595
transform 1 0 9292 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_97
timestamp 1604681595
transform 1 0 10028 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9844 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_101
timestamp 1604681595
transform 1 0 10396 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 10212 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1604681595
transform 1 0 11132 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 10764 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_107
timestamp 1604681595
transform 1 0 10948 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_118
timestamp 1604681595
transform 1 0 11960 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_122
timestamp 1604681595
transform 1 0 12328 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_125
timestamp 1604681595
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12788 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_143
timestamp 1604681595
transform 1 0 14260 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_147
timestamp 1604681595
transform 1 0 14628 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 14812 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_151
timestamp 1604681595
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 15456 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604681595
transform 1 0 15640 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_162
timestamp 1604681595
transform 1 0 16008 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 16192 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_166
timestamp 1604681595
transform 1 0 16376 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16744 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 16560 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_186
timestamp 1604681595
transform 1 0 18216 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l4_in_0_
timestamp 1604681595
transform 1 0 18952 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 19964 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 18492 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_191
timestamp 1604681595
transform 1 0 18676 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_203
timestamp 1604681595
transform 1 0 19780 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_207
timestamp 1604681595
transform 1 0 20148 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21896 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_211
timestamp 1604681595
transform 1 0 20516 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_224
timestamp 1604681595
transform 1 0 21712 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_228
timestamp 1604681595
transform 1 0 22080 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_1_
timestamp 1604681595
transform 1 0 22448 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_2_
timestamp 1604681595
transform 1 0 24012 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 22264 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 23644 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_241
timestamp 1604681595
transform 1 0 23276 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_247
timestamp 1604681595
transform 1 0 23828 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_2__A1
timestamp 1604681595
transform 1 0 25024 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_3__A1
timestamp 1604681595
transform 1 0 25392 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 25760 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_258
timestamp 1604681595
transform 1 0 24840 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_262
timestamp 1604681595
transform 1 0 25208 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_266
timestamp 1604681595
transform 1 0 25576 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_270
timestamp 1604681595
transform 1 0 25944 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_274
timestamp 1604681595
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2024 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 1840 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_7
timestamp 1604681595
transform 1 0 1748 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_19
timestamp 1604681595
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3036 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_23
timestamp 1604681595
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_36
timestamp 1604681595
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_40
timestamp 1604681595
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_7_
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_7__A1
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_7__A0
timestamp 1604681595
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_53
timestamp 1604681595
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1604681595
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8556 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_71
timestamp 1604681595
transform 1 0 7636 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_77
timestamp 1604681595
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_97
timestamp 1604681595
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_101
timestamp 1604681595
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_4_
timestamp 1604681595
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_114
timestamp 1604681595
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1604681595
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13984 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_132
timestamp 1604681595
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_136
timestamp 1604681595
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 15732 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 15548 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15180 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_149
timestamp 1604681595
transform 1 0 14812 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_155
timestamp 1604681595
transform 1 0 15364 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_3_
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_175
timestamp 1604681595
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_179
timestamp 1604681595
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1604681595
transform 1 0 19596 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_193
timestamp 1604681595
transform 1 0 18860 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_197
timestamp 1604681595
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21160 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20976 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_210
timestamp 1604681595
transform 1 0 20424 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_214
timestamp 1604681595
transform 1 0 20792 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_227
timestamp 1604681595
transform 1 0 21988 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_3_
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 22448 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 22816 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_3__S
timestamp 1604681595
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_231
timestamp 1604681595
transform 1 0 22356 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_234
timestamp 1604681595
transform 1 0 22632 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_238
timestamp 1604681595
transform 1 0 23000 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604681595
transform 1 0 25208 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 24656 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1604681595
transform 1 0 25760 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 25024 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_254
timestamp 1604681595
transform 1 0 24472 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_258
timestamp 1604681595
transform 1 0 24840 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_266
timestamp 1604681595
transform 1 0 25576 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_270
timestamp 1604681595
transform 1 0 25944 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 26128 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_274
timestamp 1604681595
transform 1 0 26312 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1656 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 2392 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 2760 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_12
timestamp 1604681595
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_16
timestamp 1604681595
transform 1 0 2576 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_20
timestamp 1604681595
transform 1 0 2944 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4232 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3128 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_24
timestamp 1604681595
transform 1 0 3312 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1604681595
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 5796 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l5_in_0__S
timestamp 1604681595
transform 1 0 5244 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5612 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_43
timestamp 1604681595
transform 1 0 5060 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_47
timestamp 1604681595
transform 1 0 5428 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 8004 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 7820 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_7__S
timestamp 1604681595
transform 1 0 7452 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_67
timestamp 1604681595
transform 1 0 7268 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_71
timestamp 1604681595
transform 1 0 7636 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_88
timestamp 1604681595
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_84
timestamp 1604681595
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A
timestamp 1604681595
transform 1 0 9844 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604681595
transform 1 0 10028 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_100
timestamp 1604681595
transform 1 0 10304 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_104
timestamp 1604681595
transform 1 0 10672 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 11040 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 10764 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 12052 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_107
timestamp 1604681595
transform 1 0 10948 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_117
timestamp 1604681595
transform 1 0 11868 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_121
timestamp 1604681595
transform 1 0 12236 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_125
timestamp 1604681595
transform 1 0 12604 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12972 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 12788 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_145
timestamp 1604681595
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_149
timestamp 1604681595
transform 1 0 14812 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_161
timestamp 1604681595
transform 1 0 15916 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_157
timestamp 1604681595
transform 1 0 15548 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 16100 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 15732 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 16284 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 18124 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_181
timestamp 1604681595
transform 1 0 17756 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_187
timestamp 1604681595
transform 1 0 18308 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1604681595
transform 1 0 18492 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 19596 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19964 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_198
timestamp 1604681595
transform 1 0 19320 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_203
timestamp 1604681595
transform 1 0 19780 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_207
timestamp 1604681595
transform 1 0 20148 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l4_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 20332 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 21896 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_211
timestamp 1604681595
transform 1 0 20516 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_224
timestamp 1604681595
transform 1 0 21712 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_228
timestamp 1604681595
transform 1 0 22080 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 24012 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 22448 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_1__S
timestamp 1604681595
transform 1 0 23644 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 22264 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_241
timestamp 1604681595
transform 1 0 23276 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_247
timestamp 1604681595
transform 1 0 23828 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l5_in_0__A0
timestamp 1604681595
transform 1 0 25024 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_3__A0
timestamp 1604681595
transform 1 0 25392 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 25760 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_258
timestamp 1604681595
transform 1 0 24840 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_262
timestamp 1604681595
transform 1 0 25208 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_266
timestamp 1604681595
transform 1 0 25576 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_270
timestamp 1604681595
transform 1 0 25944 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_274
timestamp 1604681595
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_7
timestamp 1604681595
transform 1 0 1748 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_7
timestamp 1604681595
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A
timestamp 1604681595
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_13
timestamp 1604681595
transform 1 0 2300 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_11
timestamp 1604681595
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 2116 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1604681595
transform 1 0 2300 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_19
timestamp 1604681595
transform 1 0 2852 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_19
timestamp 1604681595
transform 1 0 2852 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_23
timestamp 1604681595
transform 1 0 3220 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_23
timestamp 1604681595
transform 1 0 3220 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1604681595
transform 1 0 3036 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1604681595
transform 1 0 3404 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1604681595
transform 1 0 3036 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1604681595
transform 1 0 4140 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_31
timestamp 1604681595
transform 1 0 3956 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4508 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l5_in_0__A0
timestamp 1604681595
transform 1 0 4324 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_35
timestamp 1604681595
transform 1 0 4324 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_37
timestamp 1604681595
transform 1 0 4508 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l5_in_0__A1
timestamp 1604681595
transform 1 0 4692 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_39
timestamp 1604681595
transform 1 0 4692 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4876 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4876 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_50
timestamp 1604681595
transform 1 0 5704 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_43
timestamp 1604681595
transform 1 0 5060 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l5_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_54
timestamp 1604681595
transform 1 0 6072 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1604681595
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_53
timestamp 1604681595
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_1__A0
timestamp 1604681595
transform 1 0 5888 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 6440 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_71
timestamp 1604681595
transform 1 0 7636 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_67
timestamp 1604681595
transform 1 0 7268 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_71
timestamp 1604681595
transform 1 0 7636 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 7452 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_77
timestamp 1604681595
transform 1 0 8188 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 7820 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 8004 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8372 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8556 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_88
timestamp 1604681595
transform 1 0 9200 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_84
timestamp 1604681595
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_90
timestamp 1604681595
transform 1 0 9384 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9016 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 9568 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _127_
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_101
timestamp 1604681595
transform 1 0 10396 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_97
timestamp 1604681595
transform 1 0 10028 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_94
timestamp 1604681595
transform 1 0 9752 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1604681595
transform 1 0 10580 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 10212 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 9936 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 10120 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_33_111
timestamp 1604681595
transform 1 0 11316 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_107
timestamp 1604681595
transform 1 0 10948 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11500 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11132 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_125
timestamp 1604681595
transform 1 0 12604 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_121
timestamp 1604681595
transform 1 0 12236 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_119
timestamp 1604681595
transform 1 0 12052 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_115
timestamp 1604681595
transform 1 0 11684 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10764 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_34_131
timestamp 1604681595
transform 1 0 13156 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_132
timestamp 1604681595
transform 1 0 13248 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12972 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 13340 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_135
timestamp 1604681595
transform 1 0 13524 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_138
timestamp 1604681595
transform 1 0 13800 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14168 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13616 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14352 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_145
timestamp 1604681595
transform 1 0 14444 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_149
timestamp 1604681595
transform 1 0 14812 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_153
timestamp 1604681595
transform 1 0 15180 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 15364 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14628 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_164
timestamp 1604681595
transform 1 0 16192 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_160
timestamp 1604681595
transform 1 0 15824 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_162
timestamp 1604681595
transform 1 0 16008 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_157
timestamp 1604681595
transform 1 0 15548 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 15824 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 16192 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 16008 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 16376 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_1_
timestamp 1604681595
transform 1 0 16376 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_33_175
timestamp 1604681595
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l4_in_0_
timestamp 1604681595
transform 1 0 16560 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17572 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_179
timestamp 1604681595
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_177
timestamp 1604681595
transform 1 0 17388 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_181
timestamp 1604681595
transform 1 0 17756 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 17940 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18124 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1604681595
transform 1 0 18952 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_197
timestamp 1604681595
transform 1 0 19228 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_193
timestamp 1604681595
transform 1 0 18860 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 19136 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_206
timestamp 1604681595
transform 1 0 20056 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_198
timestamp 1604681595
transform 1 0 19320 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19504 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1604681595
transform 1 0 19412 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19596 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604681595
transform 1 0 19688 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 20424 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_210
timestamp 1604681595
transform 1 0 20424 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_212
timestamp 1604681595
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20976 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_214
timestamp 1604681595
transform 1 0 20792 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21160 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20976 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_225
timestamp 1604681595
transform 1 0 21804 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_227
timestamp 1604681595
transform 1 0 21988 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 21988 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_229
timestamp 1604681595
transform 1 0 22172 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 22172 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_238
timestamp 1604681595
transform 1 0 23000 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_233
timestamp 1604681595
transform 1 0 22540 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_239
timestamp 1604681595
transform 1 0 23092 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_235
timestamp 1604681595
transform 1 0 22724 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_231
timestamp 1604681595
transform 1 0 22356 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_1__A0
timestamp 1604681595
transform 1 0 22816 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 22908 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 22356 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22540 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_1__A1
timestamp 1604681595
transform 1 0 23184 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l5_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l5_in_0_
timestamp 1604681595
transform 1 0 23368 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_255
timestamp 1604681595
transform 1 0 24564 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_251
timestamp 1604681595
transform 1 0 24196 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_258
timestamp 1604681595
transform 1 0 24840 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_254
timestamp 1604681595
transform 1 0 24472 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l5_in_0__A1
timestamp 1604681595
transform 1 0 24748 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 24380 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1604681595
transform 1 0 24932 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604681595
transform 1 0 24932 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_270 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 25944 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_266
timestamp 1604681595
transform 1 0 25576 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_261
timestamp 1604681595
transform 1 0 25116 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1604681595
transform 1 0 25760 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604681595
transform 1 0 25208 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_276
timestamp 1604681595
transform 1 0 26496 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A
timestamp 1604681595
transform 1 0 1932 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1604681595
transform 1 0 2300 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_7
timestamp 1604681595
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_11
timestamp 1604681595
transform 1 0 2116 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_19
timestamp 1604681595
transform 1 0 2852 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1604681595
transform 1 0 3036 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4600 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 4232 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 3864 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_23
timestamp 1604681595
transform 1 0 3220 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_29
timestamp 1604681595
transform 1 0 3772 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_32
timestamp 1604681595
transform 1 0 4048 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_36
timestamp 1604681595
transform 1 0 4416 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_40
timestamp 1604681595
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5152 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 4968 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_53
timestamp 1604681595
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1604681595
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7176 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6992 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_82
timestamp 1604681595
transform 1 0 8648 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 9384 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 9200 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 8832 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_86
timestamp 1604681595
transform 1 0 9016 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_106
timestamp 1604681595
transform 1 0 10856 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11040 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_110
timestamp 1604681595
transform 1 0 11224 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_115
timestamp 1604681595
transform 1 0 11684 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11500 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_119
timestamp 1604681595
transform 1 0 12052 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11868 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_123
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12604 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 13340 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13156 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_127
timestamp 1604681595
transform 1 0 12788 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15548 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 15364 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_149
timestamp 1604681595
transform 1 0 14812 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_153
timestamp 1604681595
transform 1 0 15180 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_173
timestamp 1604681595
transform 1 0 17020 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_179
timestamp 1604681595
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 19044 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 20240 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 19412 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 19780 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_193
timestamp 1604681595
transform 1 0 18860 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_197
timestamp 1604681595
transform 1 0 19228 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_201
timestamp 1604681595
transform 1 0 19596 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_205
timestamp 1604681595
transform 1 0 19964 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21988 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 20424 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 21804 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 21436 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_219
timestamp 1604681595
transform 1 0 21252 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_223
timestamp 1604681595
transform 1 0 21620 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 23828 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 23000 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_236
timestamp 1604681595
transform 1 0 22816 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_240
timestamp 1604681595
transform 1 0 23184 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_245
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604681595
transform 1 0 25392 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1604681595
transform 1 0 25944 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 24840 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 25208 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_256
timestamp 1604681595
transform 1 0 24656 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_260
timestamp 1604681595
transform 1 0 25024 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_268
timestamp 1604681595
transform 1 0 25760 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_272
timestamp 1604681595
transform 1 0 26128 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_276
timestamp 1604681595
transform 1 0 26496 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_7
timestamp 1604681595
transform 1 0 1748 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_19
timestamp 1604681595
transform 1 0 2852 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 4324 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 4692 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_32
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_37
timestamp 1604681595
transform 1 0 4508 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_41
timestamp 1604681595
transform 1 0 4876 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5060 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6808 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 5796 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 6440 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_49
timestamp 1604681595
transform 1 0 5612 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_53
timestamp 1604681595
transform 1 0 5980 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_57
timestamp 1604681595
transform 1 0 6348 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_60
timestamp 1604681595
transform 1 0 6624 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7084 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_36_64
timestamp 1604681595
transform 1 0 6992 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_81
timestamp 1604681595
transform 1 0 8556 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_85
timestamp 1604681595
transform 1 0 8924 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_88
timestamp 1604681595
transform 1 0 9200 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11868 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 11592 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_109
timestamp 1604681595
transform 1 0 11132 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_113
timestamp 1604681595
transform 1 0 11500 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_116
timestamp 1604681595
transform 1 0 11776 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13432 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 13248 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12880 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 14444 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_126
timestamp 1604681595
transform 1 0 12696 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_130
timestamp 1604681595
transform 1 0 13064 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_143
timestamp 1604681595
transform 1 0 14260 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16008 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 15456 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15824 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_147
timestamp 1604681595
transform 1 0 14628 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_154
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_158
timestamp 1604681595
transform 1 0 15640 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18216 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 18032 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 17664 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_178
timestamp 1604681595
transform 1 0 17480 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_182
timestamp 1604681595
transform 1 0 17848 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 19228 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 19596 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 20240 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_195
timestamp 1604681595
transform 1 0 19044 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_199
timestamp 1604681595
transform 1 0 19412 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_203
timestamp 1604681595
transform 1 0 19780 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_207
timestamp 1604681595
transform 1 0 20148 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21620 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 21436 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 21068 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_210
timestamp 1604681595
transform 1 0 20424 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_215
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_219
timestamp 1604681595
transform 1 0 21252 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1604681595
transform 1 0 23828 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_4__S
timestamp 1604681595
transform 1 0 22632 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 23644 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 23276 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_232
timestamp 1604681595
transform 1 0 22448 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_236
timestamp 1604681595
transform 1 0 22816 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_240
timestamp 1604681595
transform 1 0 23184 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_243
timestamp 1604681595
transform 1 0 23460 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 24840 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 25208 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 25576 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_256
timestamp 1604681595
transform 1 0 24656 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_260
timestamp 1604681595
transform 1 0 25024 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1604681595
transform 1 0 25392 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_268
timestamp 1604681595
transform 1 0 25760 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_274
timestamp 1604681595
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A
timestamp 1604681595
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2300 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_7
timestamp 1604681595
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_11
timestamp 1604681595
transform 1 0 2116 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1604681595
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1604681595
transform 1 0 4416 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_35
timestamp 1604681595
transform 1 0 4324 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_40
timestamp 1604681595
transform 1 0 4784 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_44
timestamp 1604681595
transform 1 0 5152 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1604681595
transform 1 0 4968 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_49
timestamp 1604681595
transform 1 0 5612 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 5428 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_53
timestamp 1604681595
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 5796 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1604681595
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7176 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6992 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_75
timestamp 1604681595
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_79
timestamp 1604681595
transform 1 0 8372 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_83
timestamp 1604681595
transform 1 0 8740 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10580 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 9016 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 8832 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10396 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10028 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_95
timestamp 1604681595
transform 1 0 9844 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_99
timestamp 1604681595
transform 1 0 10212 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_112
timestamp 1604681595
transform 1 0 11408 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_116
timestamp 1604681595
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_120
timestamp 1604681595
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_123
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13248 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 13064 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12696 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14352 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_128
timestamp 1604681595
transform 1 0 12880 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_141
timestamp 1604681595
transform 1 0 14076 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1604681595
transform 1 0 14904 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16008 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 15456 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1604681595
transform 1 0 14720 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 15824 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_146
timestamp 1604681595
transform 1 0 14536 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_154
timestamp 1604681595
transform 1 0 15272 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_158
timestamp 1604681595
transform 1 0 15640 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17020 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_171
timestamp 1604681595
transform 1 0 16836 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_175
timestamp 1604681595
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_179
timestamp 1604681595
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19596 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 19044 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 19412 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_193
timestamp 1604681595
transform 1 0 18860 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_197
timestamp 1604681595
transform 1 0 19228 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 21804 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_4__A1
timestamp 1604681595
transform 1 0 21620 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_4__A0
timestamp 1604681595
transform 1 0 21252 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 20608 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_210
timestamp 1604681595
transform 1 0 20424 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_214
timestamp 1604681595
transform 1 0 20792 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_218
timestamp 1604681595
transform 1 0 21160 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_221
timestamp 1604681595
transform 1 0 21436 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1604681595
transform 1 0 23828 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_234
timestamp 1604681595
transform 1 0 22632 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_240
timestamp 1604681595
transform 1 0 23184 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_245
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604681595
transform 1 0 25392 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1604681595
transform 1 0 25024 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1604681595
transform 1 0 25944 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_256
timestamp 1604681595
transform 1 0 24656 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_262
timestamp 1604681595
transform 1 0 25208 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_268
timestamp 1604681595
transform 1 0 25760 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_272
timestamp 1604681595
transform 1 0 26128 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_276
timestamp 1604681595
transform 1 0 26496 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2116 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__057__A
timestamp 1604681595
transform 1 0 1564 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_7
timestamp 1604681595
transform 1 0 1748 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_17
timestamp 1604681595
transform 1 0 2668 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1604681595
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6808 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1604681595
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_56
timestamp 1604681595
transform 1 0 6256 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 7544 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7176 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 8556 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_64
timestamp 1604681595
transform 1 0 6992 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_68
timestamp 1604681595
transform 1 0 7360 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_76
timestamp 1604681595
transform 1 0 8096 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_80
timestamp 1604681595
transform 1 0 8464 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_83
timestamp 1604681595
transform 1 0 8740 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10028 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9844 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 9016 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_88
timestamp 1604681595
transform 1 0 9200 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_3_
timestamp 1604681595
transform 1 0 11592 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 11316 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12604 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_106
timestamp 1604681595
transform 1 0 10856 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_110
timestamp 1604681595
transform 1 0 11224 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_113
timestamp 1604681595
transform 1 0 11500 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_123
timestamp 1604681595
transform 1 0 12420 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13156 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12972 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14168 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_127
timestamp 1604681595
transform 1 0 12788 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_140
timestamp 1604681595
transform 1 0 13984 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_144
timestamp 1604681595
transform 1 0 14352 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 14628 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16284 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_149
timestamp 1604681595
transform 1 0 14812 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_163
timestamp 1604681595
transform 1 0 16100 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16836 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18032 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 16652 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_167
timestamp 1604681595
transform 1 0 16468 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_180
timestamp 1604681595
transform 1 0 17664 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_186
timestamp 1604681595
transform 1 0 18216 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18400 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19596 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 20240 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_197
timestamp 1604681595
transform 1 0 19228 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_203
timestamp 1604681595
transform 1 0 19780 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_207
timestamp 1604681595
transform 1 0 20148 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_4_
timestamp 1604681595
transform 1 0 21896 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21068 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21436 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_210
timestamp 1604681595
transform 1 0 20424 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_215
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_219
timestamp 1604681595
transform 1 0 21252 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_223
timestamp 1604681595
transform 1 0 21620 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1604681595
transform 1 0 23460 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23092 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_235
timestamp 1604681595
transform 1 0 22724 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_241
timestamp 1604681595
transform 1 0 23276 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604681595
transform 1 0 25024 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 24656 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 25576 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_252
timestamp 1604681595
transform 1 0 24288 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_258
timestamp 1604681595
transform 1 0 24840 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1604681595
transform 1 0 25392 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_268
timestamp 1604681595
transform 1 0 25760 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_274
timestamp 1604681595
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_7
timestamp 1604681595
transform 1 0 1748 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__058__A
timestamp 1604681595
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_19
timestamp 1604681595
transform 1 0 2852 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_11
timestamp 1604681595
transform 1 0 2116 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_19
timestamp 1604681595
transform 1 0 2852 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_7
timestamp 1604681595
transform 1 0 1748 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__A
timestamp 1604681595
transform 1 0 3036 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_23
timestamp 1604681595
transform 1 0 3220 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_35
timestamp 1604681595
transform 1 0 4324 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_47
timestamp 1604681595
transform 1 0 5428 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1604681595
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_62
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1604681595
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1604681595
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1604681595
transform 1 0 7360 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1604681595
transform 1 0 7360 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_72
timestamp 1604681595
transform 1 0 7728 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_39_70
timestamp 1604681595
transform 1 0 7544 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _134_
timestamp 1604681595
transform 1 0 7820 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_81
timestamp 1604681595
transform 1 0 8556 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_77
timestamp 1604681595
transform 1 0 8188 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 8280 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A
timestamp 1604681595
transform 1 0 8740 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1604681595
transform 1 0 8372 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _133_
timestamp 1604681595
transform 1 0 8464 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_88
timestamp 1604681595
transform 1 0 9200 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_84
timestamp 1604681595
transform 1 0 8832 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1604681595
transform 1 0 8924 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_93
timestamp 1604681595
transform 1 0 9660 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_89
timestamp 1604681595
transform 1 0 9292 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__056__A
timestamp 1604681595
transform 1 0 9476 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_97
timestamp 1604681595
transform 1 0 10028 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_97
timestamp 1604681595
transform 1 0 10028 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 9844 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 9844 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_101
timestamp 1604681595
transform 1 0 10396 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1604681595
transform 1 0 10212 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _129_
timestamp 1604681595
transform 1 0 10212 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_103
timestamp 1604681595
transform 1 0 10580 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 10580 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_107
timestamp 1604681595
transform 1 0 10948 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_114
timestamp 1604681595
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 11132 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 10764 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1604681595
transform 1 0 10764 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_2_
timestamp 1604681595
transform 1 0 11316 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_40_120
timestamp 1604681595
transform 1 0 12144 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_123
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 1604681595
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_124
timestamp 1604681595
transform 1 0 12512 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 12604 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_131
timestamp 1604681595
transform 1 0 13156 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_127
timestamp 1604681595
transform 1 0 12788 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_128
timestamp 1604681595
transform 1 0 12880 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 12696 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 13064 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 12972 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1604681595
transform 1 0 13432 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1604681595
transform 1 0 13248 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_40_143
timestamp 1604681595
transform 1 0 14260 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_141
timestamp 1604681595
transform 1 0 14076 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 14260 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_145
timestamp 1604681595
transform 1 0 14444 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_150
timestamp 1604681595
transform 1 0 14904 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_147
timestamp 1604681595
transform 1 0 14628 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_149
timestamp 1604681595
transform 1 0 14812 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14720 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 14628 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 14996 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_2_
timestamp 1604681595
transform 1 0 15180 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_163
timestamp 1604681595
transform 1 0 16100 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_162
timestamp 1604681595
transform 1 0 16008 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16284 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 16192 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_166
timestamp 1604681595
transform 1 0 16376 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_167
timestamp 1604681595
transform 1 0 16468 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_175
timestamp 1604681595
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16652 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 16652 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1604681595
transform 1 0 16836 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1604681595
transform 1 0 16836 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_186
timestamp 1604681595
transform 1 0 18216 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_180
timestamp 1604681595
transform 1 0 17664 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_179
timestamp 1604681595
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18032 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1604681595
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_40_190
timestamp 1604681595
transform 1 0 18584 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_193
timestamp 1604681595
transform 1 0 18860 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 19044 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18400 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18860 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_203
timestamp 1604681595
transform 1 0 19780 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_199
timestamp 1604681595
transform 1 0 19412 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_197
timestamp 1604681595
transform 1 0 19228 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19596 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19412 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19596 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_207
timestamp 1604681595
transform 1 0 20148 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_215
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_211
timestamp 1604681595
transform 1 0 20516 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_211
timestamp 1604681595
transform 1 0 20516 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__A0
timestamp 1604681595
transform 1 0 20332 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__A1
timestamp 1604681595
transform 1 0 20700 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_5_
timestamp 1604681595
transform 1 0 20884 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20976 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_40_225
timestamp 1604681595
transform 1 0 21804 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_228
timestamp 1604681595
transform 1 0 22080 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_224
timestamp 1604681595
transform 1 0 21712 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 22080 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21896 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604681595
transform 1 0 22448 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__S
timestamp 1604681595
transform 1 0 22264 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 22448 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_230
timestamp 1604681595
transform 1 0 22264 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_234
timestamp 1604681595
transform 1 0 22632 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1604681595
transform 1 0 23000 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1604681595
transform 1 0 22816 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_236
timestamp 1604681595
transform 1 0 22816 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_238
timestamp 1604681595
transform 1 0 23000 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23092 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_248
timestamp 1604681595
transform 1 0 23920 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_240
timestamp 1604681595
transform 1 0 23184 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A1
timestamp 1604681595
transform 1 0 24104 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_252
timestamp 1604681595
transform 1 0 24288 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_258
timestamp 1604681595
transform 1 0 24840 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_254
timestamp 1604681595
transform 1 0 24472 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_7__A0
timestamp 1604681595
transform 1 0 24472 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 24656 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 24656 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_40_265
timestamp 1604681595
transform 1 0 25484 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_266
timestamp 1604681595
transform 1 0 25576 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 25024 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1604681595
transform 1 0 25760 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604681595
transform 1 0 25208 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_270
timestamp 1604681595
transform 1 0 25944 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 26128 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_274
timestamp 1604681595
transform 1 0 26312 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_273
timestamp 1604681595
transform 1 0 26220 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A
timestamp 1604681595
transform 1 0 1932 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_7
timestamp 1604681595
transform 1 0 1748 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_11
timestamp 1604681595
transform 1 0 2116 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_23
timestamp 1604681595
transform 1 0 3220 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_35
timestamp 1604681595
transform 1 0 4324 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_47
timestamp 1604681595
transform 1 0 5428 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_59
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 8556 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_74
timestamp 1604681595
transform 1 0 7912 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_80
timestamp 1604681595
transform 1 0 8464 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_83
timestamp 1604681595
transform 1 0 8740 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _131_
timestamp 1604681595
transform 1 0 10120 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _135_
timestamp 1604681595
transform 1 0 9016 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__A
timestamp 1604681595
transform 1 0 10672 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1604681595
transform 1 0 9568 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__A
timestamp 1604681595
transform 1 0 9936 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_90
timestamp 1604681595
transform 1 0 9384 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_94
timestamp 1604681595
transform 1 0 9752 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_102
timestamp 1604681595
transform 1 0 10488 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _128_
timestamp 1604681595
transform 1 0 11224 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__A
timestamp 1604681595
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__128__A
timestamp 1604681595
transform 1 0 11040 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_106
timestamp 1604681595
transform 1 0 10856 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_114
timestamp 1604681595
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_118
timestamp 1604681595
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_123
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12972 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 12788 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14168 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_138
timestamp 1604681595
transform 1 0 13800 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_144
timestamp 1604681595
transform 1 0 14352 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16284 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 14720 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 15732 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 16100 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 14536 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_157
timestamp 1604681595
transform 1 0 15548 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_161
timestamp 1604681595
transform 1 0 15916 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18308 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1604681595
transform 1 0 17296 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_174
timestamp 1604681595
transform 1 0 17112 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_178
timestamp 1604681595
transform 1 0 17480 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_184
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604681595
transform 1 0 20148 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1604681595
transform 1 0 19044 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1604681595
transform 1 0 19964 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_193
timestamp 1604681595
transform 1 0 18860 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_197
timestamp 1604681595
transform 1 0 19228 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _126_
timestamp 1604681595
transform 1 0 21252 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1604681595
transform 1 0 21804 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A
timestamp 1604681595
transform 1 0 21068 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1604681595
transform 1 0 20700 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_211
timestamp 1604681595
transform 1 0 20516 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_215
timestamp 1604681595
transform 1 0 20884 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_223
timestamp 1604681595
transform 1 0 21620 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_227
timestamp 1604681595
transform 1 0 21988 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604681595
transform 1 0 22448 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_6_
timestamp 1604681595
transform 1 0 23828 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1604681595
transform 1 0 23000 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A0
timestamp 1604681595
transform 1 0 23368 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_231
timestamp 1604681595
transform 1 0 22356 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_236
timestamp 1604681595
transform 1 0 22816 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_240
timestamp 1604681595
transform 1 0 23184 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604681595
transform 1 0 25392 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_7__A1
timestamp 1604681595
transform 1 0 24840 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1604681595
transform 1 0 25944 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_7__S
timestamp 1604681595
transform 1 0 25208 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_256
timestamp 1604681595
transform 1 0 24656 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_260
timestamp 1604681595
transform 1 0 25024 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_268
timestamp 1604681595
transform 1 0 25760 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_272
timestamp 1604681595
transform 1 0 26128 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_276
timestamp 1604681595
transform 1 0 26496 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1604681595
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604681595
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1604681595
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_56
timestamp 1604681595
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_63
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1604681595
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _132_
timestamp 1604681595
transform 1 0 10304 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 10120 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_87
timestamp 1604681595
transform 1 0 9108 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_92
timestamp 1604681595
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_94
timestamp 1604681595
transform 1 0 9752 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_104
timestamp 1604681595
transform 1 0 10672 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_108
timestamp 1604681595
transform 1 0 11040 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 10856 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 11224 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _130_
timestamp 1604681595
transform 1 0 11408 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_116
timestamp 1604681595
transform 1 0 11776 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11960 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_120
timestamp 1604681595
transform 1 0 12144 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 12328 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_125
timestamp 1604681595
transform 1 0 12604 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12788 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14076 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13524 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13892 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_133
timestamp 1604681595
transform 1 0 13340 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_137
timestamp 1604681595
transform 1 0 13708 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_4_
timestamp 1604681595
transform 1 0 15456 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14812 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 15180 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_147
timestamp 1604681595
transform 1 0 14628 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_151
timestamp 1604681595
transform 1 0 14996 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_165
timestamp 1604681595
transform 1 0 16284 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_173
timestamp 1604681595
transform 1 0 17020 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_169
timestamp 1604681595
transform 1 0 16652 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 16836 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16468 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_178
timestamp 1604681595
transform 1 0 17480 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 17664 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1604681595
transform 1 0 17112 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_187
timestamp 1604681595
transform 1 0 18308 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_182
timestamp 1604681595
transform 1 0 17848 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1604681595
transform 1 0 19964 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1604681595
transform 1 0 18860 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_197
timestamp 1604681595
transform 1 0 19228 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1604681595
transform 1 0 21712 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_209
timestamp 1604681595
transform 1 0 20332 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_218
timestamp 1604681595
transform 1 0 21160 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_228
timestamp 1604681595
transform 1 0 22080 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1604681595
transform 1 0 22816 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_7_
timestamp 1604681595
transform 1 0 24104 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__S
timestamp 1604681595
transform 1 0 23736 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_240
timestamp 1604681595
transform 1 0 23184 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_249
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_259
timestamp 1604681595
transform 1 0 24932 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_271
timestamp 1604681595
transform 1 0 26036 0 -1 25568
box -38 -48 590 592
<< labels >>
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_42_
port 0 nsew default input
rlabel metal2 s 662 0 718 480 6 bottom_left_grid_pin_43_
port 1 nsew default input
rlabel metal2 s 1214 0 1270 480 6 bottom_left_grid_pin_44_
port 2 nsew default input
rlabel metal2 s 1766 0 1822 480 6 bottom_left_grid_pin_45_
port 3 nsew default input
rlabel metal2 s 2318 0 2374 480 6 bottom_left_grid_pin_46_
port 4 nsew default input
rlabel metal2 s 2870 0 2926 480 6 bottom_left_grid_pin_47_
port 5 nsew default input
rlabel metal2 s 3422 0 3478 480 6 bottom_left_grid_pin_48_
port 6 nsew default input
rlabel metal2 s 3974 0 4030 480 6 bottom_left_grid_pin_49_
port 7 nsew default input
rlabel metal2 s 5078 0 5134 480 6 ccff_head
port 8 nsew default input
rlabel metal2 s 5630 0 5686 480 6 ccff_tail
port 9 nsew default tristate
rlabel metal3 s 0 4904 480 5024 6 chanx_left_in[0]
port 10 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[10]
port 11 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[11]
port 12 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_in[12]
port 13 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[13]
port 14 nsew default input
rlabel metal3 s 0 13064 480 13184 6 chanx_left_in[14]
port 15 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chanx_left_in[15]
port 16 nsew default input
rlabel metal3 s 0 14288 480 14408 6 chanx_left_in[16]
port 17 nsew default input
rlabel metal3 s 0 14832 480 14952 6 chanx_left_in[17]
port 18 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chanx_left_in[18]
port 19 nsew default input
rlabel metal3 s 0 15920 480 16040 6 chanx_left_in[19]
port 20 nsew default input
rlabel metal3 s 0 5448 480 5568 6 chanx_left_in[1]
port 21 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[2]
port 22 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[3]
port 23 nsew default input
rlabel metal3 s 0 7216 480 7336 6 chanx_left_in[4]
port 24 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[5]
port 25 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[6]
port 26 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[7]
port 27 nsew default input
rlabel metal3 s 0 9528 480 9648 6 chanx_left_in[8]
port 28 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[9]
port 29 nsew default input
rlabel metal3 s 0 16600 480 16720 6 chanx_left_out[0]
port 30 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[10]
port 31 nsew default tristate
rlabel metal3 s 0 22992 480 23112 6 chanx_left_out[11]
port 32 nsew default tristate
rlabel metal3 s 0 23536 480 23656 6 chanx_left_out[12]
port 33 nsew default tristate
rlabel metal3 s 0 24080 480 24200 6 chanx_left_out[13]
port 34 nsew default tristate
rlabel metal3 s 0 24760 480 24880 6 chanx_left_out[14]
port 35 nsew default tristate
rlabel metal3 s 0 25304 480 25424 6 chanx_left_out[15]
port 36 nsew default tristate
rlabel metal3 s 0 25848 480 25968 6 chanx_left_out[16]
port 37 nsew default tristate
rlabel metal3 s 0 26528 480 26648 6 chanx_left_out[17]
port 38 nsew default tristate
rlabel metal3 s 0 27072 480 27192 6 chanx_left_out[18]
port 39 nsew default tristate
rlabel metal3 s 0 27616 480 27736 6 chanx_left_out[19]
port 40 nsew default tristate
rlabel metal3 s 0 17144 480 17264 6 chanx_left_out[1]
port 41 nsew default tristate
rlabel metal3 s 0 17688 480 17808 6 chanx_left_out[2]
port 42 nsew default tristate
rlabel metal3 s 0 18368 480 18488 6 chanx_left_out[3]
port 43 nsew default tristate
rlabel metal3 s 0 18912 480 19032 6 chanx_left_out[4]
port 44 nsew default tristate
rlabel metal3 s 0 19456 480 19576 6 chanx_left_out[5]
port 45 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 chanx_left_out[6]
port 46 nsew default tristate
rlabel metal3 s 0 20680 480 20800 6 chanx_left_out[7]
port 47 nsew default tristate
rlabel metal3 s 0 21224 480 21344 6 chanx_left_out[8]
port 48 nsew default tristate
rlabel metal3 s 0 21768 480 21888 6 chanx_left_out[9]
port 49 nsew default tristate
rlabel metal3 s 27520 4904 28000 5024 6 chanx_right_in[0]
port 50 nsew default input
rlabel metal3 s 27520 10752 28000 10872 6 chanx_right_in[10]
port 51 nsew default input
rlabel metal3 s 27520 11296 28000 11416 6 chanx_right_in[11]
port 52 nsew default input
rlabel metal3 s 27520 11840 28000 11960 6 chanx_right_in[12]
port 53 nsew default input
rlabel metal3 s 27520 12520 28000 12640 6 chanx_right_in[13]
port 54 nsew default input
rlabel metal3 s 27520 13064 28000 13184 6 chanx_right_in[14]
port 55 nsew default input
rlabel metal3 s 27520 13608 28000 13728 6 chanx_right_in[15]
port 56 nsew default input
rlabel metal3 s 27520 14288 28000 14408 6 chanx_right_in[16]
port 57 nsew default input
rlabel metal3 s 27520 14832 28000 14952 6 chanx_right_in[17]
port 58 nsew default input
rlabel metal3 s 27520 15376 28000 15496 6 chanx_right_in[18]
port 59 nsew default input
rlabel metal3 s 27520 15920 28000 16040 6 chanx_right_in[19]
port 60 nsew default input
rlabel metal3 s 27520 5448 28000 5568 6 chanx_right_in[1]
port 61 nsew default input
rlabel metal3 s 27520 5992 28000 6112 6 chanx_right_in[2]
port 62 nsew default input
rlabel metal3 s 27520 6672 28000 6792 6 chanx_right_in[3]
port 63 nsew default input
rlabel metal3 s 27520 7216 28000 7336 6 chanx_right_in[4]
port 64 nsew default input
rlabel metal3 s 27520 7760 28000 7880 6 chanx_right_in[5]
port 65 nsew default input
rlabel metal3 s 27520 8440 28000 8560 6 chanx_right_in[6]
port 66 nsew default input
rlabel metal3 s 27520 8984 28000 9104 6 chanx_right_in[7]
port 67 nsew default input
rlabel metal3 s 27520 9528 28000 9648 6 chanx_right_in[8]
port 68 nsew default input
rlabel metal3 s 27520 10072 28000 10192 6 chanx_right_in[9]
port 69 nsew default input
rlabel metal3 s 27520 16600 28000 16720 6 chanx_right_out[0]
port 70 nsew default tristate
rlabel metal3 s 27520 22448 28000 22568 6 chanx_right_out[10]
port 71 nsew default tristate
rlabel metal3 s 27520 22992 28000 23112 6 chanx_right_out[11]
port 72 nsew default tristate
rlabel metal3 s 27520 23536 28000 23656 6 chanx_right_out[12]
port 73 nsew default tristate
rlabel metal3 s 27520 24080 28000 24200 6 chanx_right_out[13]
port 74 nsew default tristate
rlabel metal3 s 27520 24760 28000 24880 6 chanx_right_out[14]
port 75 nsew default tristate
rlabel metal3 s 27520 25304 28000 25424 6 chanx_right_out[15]
port 76 nsew default tristate
rlabel metal3 s 27520 25848 28000 25968 6 chanx_right_out[16]
port 77 nsew default tristate
rlabel metal3 s 27520 26528 28000 26648 6 chanx_right_out[17]
port 78 nsew default tristate
rlabel metal3 s 27520 27072 28000 27192 6 chanx_right_out[18]
port 79 nsew default tristate
rlabel metal3 s 27520 27616 28000 27736 6 chanx_right_out[19]
port 80 nsew default tristate
rlabel metal3 s 27520 17144 28000 17264 6 chanx_right_out[1]
port 81 nsew default tristate
rlabel metal3 s 27520 17688 28000 17808 6 chanx_right_out[2]
port 82 nsew default tristate
rlabel metal3 s 27520 18368 28000 18488 6 chanx_right_out[3]
port 83 nsew default tristate
rlabel metal3 s 27520 18912 28000 19032 6 chanx_right_out[4]
port 84 nsew default tristate
rlabel metal3 s 27520 19456 28000 19576 6 chanx_right_out[5]
port 85 nsew default tristate
rlabel metal3 s 27520 20000 28000 20120 6 chanx_right_out[6]
port 86 nsew default tristate
rlabel metal3 s 27520 20680 28000 20800 6 chanx_right_out[7]
port 87 nsew default tristate
rlabel metal3 s 27520 21224 28000 21344 6 chanx_right_out[8]
port 88 nsew default tristate
rlabel metal3 s 27520 21768 28000 21888 6 chanx_right_out[9]
port 89 nsew default tristate
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_in[0]
port 90 nsew default input
rlabel metal2 s 11702 0 11758 480 6 chany_bottom_in[10]
port 91 nsew default input
rlabel metal2 s 12254 0 12310 480 6 chany_bottom_in[11]
port 92 nsew default input
rlabel metal2 s 12806 0 12862 480 6 chany_bottom_in[12]
port 93 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[13]
port 94 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_in[14]
port 95 nsew default input
rlabel metal2 s 14370 0 14426 480 6 chany_bottom_in[15]
port 96 nsew default input
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_in[16]
port 97 nsew default input
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_in[17]
port 98 nsew default input
rlabel metal2 s 16026 0 16082 480 6 chany_bottom_in[18]
port 99 nsew default input
rlabel metal2 s 16578 0 16634 480 6 chany_bottom_in[19]
port 100 nsew default input
rlabel metal2 s 6734 0 6790 480 6 chany_bottom_in[1]
port 101 nsew default input
rlabel metal2 s 7286 0 7342 480 6 chany_bottom_in[2]
port 102 nsew default input
rlabel metal2 s 7838 0 7894 480 6 chany_bottom_in[3]
port 103 nsew default input
rlabel metal2 s 8390 0 8446 480 6 chany_bottom_in[4]
port 104 nsew default input
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_in[5]
port 105 nsew default input
rlabel metal2 s 9494 0 9550 480 6 chany_bottom_in[6]
port 106 nsew default input
rlabel metal2 s 10046 0 10102 480 6 chany_bottom_in[7]
port 107 nsew default input
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_in[8]
port 108 nsew default input
rlabel metal2 s 11150 0 11206 480 6 chany_bottom_in[9]
port 109 nsew default input
rlabel metal2 s 17130 0 17186 480 6 chany_bottom_out[0]
port 110 nsew default tristate
rlabel metal2 s 22650 0 22706 480 6 chany_bottom_out[10]
port 111 nsew default tristate
rlabel metal2 s 23202 0 23258 480 6 chany_bottom_out[11]
port 112 nsew default tristate
rlabel metal2 s 23754 0 23810 480 6 chany_bottom_out[12]
port 113 nsew default tristate
rlabel metal2 s 24306 0 24362 480 6 chany_bottom_out[13]
port 114 nsew default tristate
rlabel metal2 s 24858 0 24914 480 6 chany_bottom_out[14]
port 115 nsew default tristate
rlabel metal2 s 25410 0 25466 480 6 chany_bottom_out[15]
port 116 nsew default tristate
rlabel metal2 s 25962 0 26018 480 6 chany_bottom_out[16]
port 117 nsew default tristate
rlabel metal2 s 26514 0 26570 480 6 chany_bottom_out[17]
port 118 nsew default tristate
rlabel metal2 s 27066 0 27122 480 6 chany_bottom_out[18]
port 119 nsew default tristate
rlabel metal2 s 27618 0 27674 480 6 chany_bottom_out[19]
port 120 nsew default tristate
rlabel metal2 s 17682 0 17738 480 6 chany_bottom_out[1]
port 121 nsew default tristate
rlabel metal2 s 18234 0 18290 480 6 chany_bottom_out[2]
port 122 nsew default tristate
rlabel metal2 s 18786 0 18842 480 6 chany_bottom_out[3]
port 123 nsew default tristate
rlabel metal2 s 19338 0 19394 480 6 chany_bottom_out[4]
port 124 nsew default tristate
rlabel metal2 s 19890 0 19946 480 6 chany_bottom_out[5]
port 125 nsew default tristate
rlabel metal2 s 20442 0 20498 480 6 chany_bottom_out[6]
port 126 nsew default tristate
rlabel metal2 s 20994 0 21050 480 6 chany_bottom_out[7]
port 127 nsew default tristate
rlabel metal2 s 21546 0 21602 480 6 chany_bottom_out[8]
port 128 nsew default tristate
rlabel metal2 s 22098 0 22154 480 6 chany_bottom_out[9]
port 129 nsew default tristate
rlabel metal2 s 4894 27520 4950 28000 6 chany_top_in[0]
port 130 nsew default input
rlabel metal2 s 10782 27520 10838 28000 6 chany_top_in[10]
port 131 nsew default input
rlabel metal2 s 11334 27520 11390 28000 6 chany_top_in[11]
port 132 nsew default input
rlabel metal2 s 11886 27520 11942 28000 6 chany_top_in[12]
port 133 nsew default input
rlabel metal2 s 12530 27520 12586 28000 6 chany_top_in[13]
port 134 nsew default input
rlabel metal2 s 13082 27520 13138 28000 6 chany_top_in[14]
port 135 nsew default input
rlabel metal2 s 13634 27520 13690 28000 6 chany_top_in[15]
port 136 nsew default input
rlabel metal2 s 14278 27520 14334 28000 6 chany_top_in[16]
port 137 nsew default input
rlabel metal2 s 14830 27520 14886 28000 6 chany_top_in[17]
port 138 nsew default input
rlabel metal2 s 15382 27520 15438 28000 6 chany_top_in[18]
port 139 nsew default input
rlabel metal2 s 16026 27520 16082 28000 6 chany_top_in[19]
port 140 nsew default input
rlabel metal2 s 5538 27520 5594 28000 6 chany_top_in[1]
port 141 nsew default input
rlabel metal2 s 6090 27520 6146 28000 6 chany_top_in[2]
port 142 nsew default input
rlabel metal2 s 6642 27520 6698 28000 6 chany_top_in[3]
port 143 nsew default input
rlabel metal2 s 7286 27520 7342 28000 6 chany_top_in[4]
port 144 nsew default input
rlabel metal2 s 7838 27520 7894 28000 6 chany_top_in[5]
port 145 nsew default input
rlabel metal2 s 8390 27520 8446 28000 6 chany_top_in[6]
port 146 nsew default input
rlabel metal2 s 9034 27520 9090 28000 6 chany_top_in[7]
port 147 nsew default input
rlabel metal2 s 9586 27520 9642 28000 6 chany_top_in[8]
port 148 nsew default input
rlabel metal2 s 10138 27520 10194 28000 6 chany_top_in[9]
port 149 nsew default input
rlabel metal2 s 16578 27520 16634 28000 6 chany_top_out[0]
port 150 nsew default tristate
rlabel metal2 s 22374 27520 22430 28000 6 chany_top_out[10]
port 151 nsew default tristate
rlabel metal2 s 23018 27520 23074 28000 6 chany_top_out[11]
port 152 nsew default tristate
rlabel metal2 s 23570 27520 23626 28000 6 chany_top_out[12]
port 153 nsew default tristate
rlabel metal2 s 24122 27520 24178 28000 6 chany_top_out[13]
port 154 nsew default tristate
rlabel metal2 s 24766 27520 24822 28000 6 chany_top_out[14]
port 155 nsew default tristate
rlabel metal2 s 25318 27520 25374 28000 6 chany_top_out[15]
port 156 nsew default tristate
rlabel metal2 s 25870 27520 25926 28000 6 chany_top_out[16]
port 157 nsew default tristate
rlabel metal2 s 26514 27520 26570 28000 6 chany_top_out[17]
port 158 nsew default tristate
rlabel metal2 s 27066 27520 27122 28000 6 chany_top_out[18]
port 159 nsew default tristate
rlabel metal2 s 27618 27520 27674 28000 6 chany_top_out[19]
port 160 nsew default tristate
rlabel metal2 s 17130 27520 17186 28000 6 chany_top_out[1]
port 161 nsew default tristate
rlabel metal2 s 17774 27520 17830 28000 6 chany_top_out[2]
port 162 nsew default tristate
rlabel metal2 s 18326 27520 18382 28000 6 chany_top_out[3]
port 163 nsew default tristate
rlabel metal2 s 18878 27520 18934 28000 6 chany_top_out[4]
port 164 nsew default tristate
rlabel metal2 s 19522 27520 19578 28000 6 chany_top_out[5]
port 165 nsew default tristate
rlabel metal2 s 20074 27520 20130 28000 6 chany_top_out[6]
port 166 nsew default tristate
rlabel metal2 s 20626 27520 20682 28000 6 chany_top_out[7]
port 167 nsew default tristate
rlabel metal2 s 21270 27520 21326 28000 6 chany_top_out[8]
port 168 nsew default tristate
rlabel metal2 s 21822 27520 21878 28000 6 chany_top_out[9]
port 169 nsew default tristate
rlabel metal3 s 0 280 480 400 6 left_bottom_grid_pin_34_
port 170 nsew default input
rlabel metal3 s 0 824 480 944 6 left_bottom_grid_pin_35_
port 171 nsew default input
rlabel metal3 s 0 1368 480 1488 6 left_bottom_grid_pin_36_
port 172 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_37_
port 173 nsew default input
rlabel metal3 s 0 2592 480 2712 6 left_bottom_grid_pin_38_
port 174 nsew default input
rlabel metal3 s 0 3136 480 3256 6 left_bottom_grid_pin_39_
port 175 nsew default input
rlabel metal3 s 0 3680 480 3800 6 left_bottom_grid_pin_40_
port 176 nsew default input
rlabel metal3 s 0 4360 480 4480 6 left_bottom_grid_pin_41_
port 177 nsew default input
rlabel metal2 s 4526 0 4582 480 6 prog_clk
port 178 nsew default input
rlabel metal3 s 27520 280 28000 400 6 right_bottom_grid_pin_34_
port 179 nsew default input
rlabel metal3 s 27520 824 28000 944 6 right_bottom_grid_pin_35_
port 180 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 right_bottom_grid_pin_36_
port 181 nsew default input
rlabel metal3 s 27520 1912 28000 2032 6 right_bottom_grid_pin_37_
port 182 nsew default input
rlabel metal3 s 27520 2592 28000 2712 6 right_bottom_grid_pin_38_
port 183 nsew default input
rlabel metal3 s 27520 3136 28000 3256 6 right_bottom_grid_pin_39_
port 184 nsew default input
rlabel metal3 s 27520 3680 28000 3800 6 right_bottom_grid_pin_40_
port 185 nsew default input
rlabel metal3 s 27520 4360 28000 4480 6 right_bottom_grid_pin_41_
port 186 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_42_
port 187 nsew default input
rlabel metal2 s 846 27520 902 28000 6 top_left_grid_pin_43_
port 188 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 top_left_grid_pin_44_
port 189 nsew default input
rlabel metal2 s 2042 27520 2098 28000 6 top_left_grid_pin_45_
port 190 nsew default input
rlabel metal2 s 2594 27520 2650 28000 6 top_left_grid_pin_46_
port 191 nsew default input
rlabel metal2 s 3146 27520 3202 28000 6 top_left_grid_pin_47_
port 192 nsew default input
rlabel metal2 s 3790 27520 3846 28000 6 top_left_grid_pin_48_
port 193 nsew default input
rlabel metal2 s 4342 27520 4398 28000 6 top_left_grid_pin_49_
port 194 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 195 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 196 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
