VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__0_
  CLASS BLOCK ;
  FOREIGN sb_0__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 115.000 BY 114.280 ;
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.880 4.000 28.480 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.000 4.000 85.600 ;
    END
  END ccff_tail
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 20.400 115.000 21.000 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 43.520 115.000 44.120 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 45.560 115.000 46.160 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 47.600 115.000 48.200 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 50.320 115.000 50.920 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 52.360 115.000 52.960 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 55.080 115.000 55.680 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 57.120 115.000 57.720 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 59.160 115.000 59.760 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 61.880 115.000 62.480 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 63.920 115.000 64.520 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 22.440 115.000 23.040 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 25.160 115.000 25.760 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 27.200 115.000 27.800 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 29.240 115.000 29.840 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 31.960 115.000 32.560 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 34.000 115.000 34.600 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 36.720 115.000 37.320 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 38.760 115.000 39.360 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 40.800 115.000 41.400 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 66.640 115.000 67.240 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 89.080 115.000 89.680 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 91.800 115.000 92.400 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 93.840 115.000 94.440 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 95.880 115.000 96.480 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 98.600 115.000 99.200 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 100.640 115.000 101.240 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 103.360 115.000 103.960 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 105.400 115.000 106.000 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 107.440 115.000 108.040 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 110.160 115.000 110.760 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 68.680 115.000 69.280 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 70.720 115.000 71.320 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 73.440 115.000 74.040 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 75.480 115.000 76.080 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 77.520 115.000 78.120 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 80.240 115.000 80.840 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 82.280 115.000 82.880 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 85.000 115.000 85.600 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 87.040 115.000 87.640 ;
    END
  END chanx_right_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 110.280 4.510 114.280 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 110.280 32.570 114.280 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 110.280 35.330 114.280 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 110.280 38.090 114.280 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 110.280 40.850 114.280 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 110.280 43.610 114.280 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 110.280 46.370 114.280 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 110.280 49.130 114.280 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 110.280 51.890 114.280 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 110.280 54.650 114.280 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 110.280 57.410 114.280 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 110.280 7.270 114.280 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 110.280 10.030 114.280 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 110.280 12.790 114.280 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 110.280 15.550 114.280 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 110.280 18.310 114.280 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 110.280 21.070 114.280 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 110.280 23.830 114.280 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 110.280 26.590 114.280 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 110.280 29.350 114.280 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 110.280 60.630 114.280 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 110.280 88.690 114.280 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 110.280 91.450 114.280 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 110.280 94.210 114.280 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 110.280 96.970 114.280 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 110.280 99.730 114.280 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 110.280 102.490 114.280 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 110.280 105.250 114.280 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 110.280 108.010 114.280 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 110.280 110.770 114.280 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 110.280 113.530 114.280 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 110.280 63.390 114.280 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 110.280 66.150 114.280 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 110.280 68.910 114.280 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 110.280 71.670 114.280 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 110.280 74.430 114.280 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 110.280 77.190 114.280 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 110.280 79.950 114.280 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 110.280 82.710 114.280 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 110.280 85.470 114.280 ;
    END
  END chany_top_out[9]
  PIN prog_clk_0_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 112.200 115.000 112.800 ;
    END
  END prog_clk_0_E_in
  PIN right_bottom_grid_pin_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 10.880 115.000 11.480 ;
    END
  END right_bottom_grid_pin_11_
  PIN right_bottom_grid_pin_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 13.600 115.000 14.200 ;
    END
  END right_bottom_grid_pin_13_
  PIN right_bottom_grid_pin_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 15.640 115.000 16.240 ;
    END
  END right_bottom_grid_pin_15_
  PIN right_bottom_grid_pin_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 18.360 115.000 18.960 ;
    END
  END right_bottom_grid_pin_17_
  PIN right_bottom_grid_pin_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 0.000 115.000 0.600 ;
    END
  END right_bottom_grid_pin_1_
  PIN right_bottom_grid_pin_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 2.040 115.000 2.640 ;
    END
  END right_bottom_grid_pin_3_
  PIN right_bottom_grid_pin_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 4.080 115.000 4.680 ;
    END
  END right_bottom_grid_pin_5_
  PIN right_bottom_grid_pin_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 6.800 115.000 7.400 ;
    END
  END right_bottom_grid_pin_7_
  PIN right_bottom_grid_pin_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 8.840 115.000 9.440 ;
    END
  END right_bottom_grid_pin_9_
  PIN top_left_grid_pin_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 110.280 1.750 114.280 ;
    END
  END top_left_grid_pin_1_
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 91.355 9.920 92.955 102.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 56.700 9.920 58.300 102.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.045 9.920 23.645 102.880 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 74.025 9.920 75.625 102.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.375 9.920 40.975 102.880 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.075 110.255 102.725 ;
      LAYER met1 ;
        RECT 1.450 5.780 113.550 102.880 ;
      LAYER met2 ;
        RECT 2.030 110.000 3.950 112.685 ;
        RECT 4.790 110.000 6.710 112.685 ;
        RECT 7.550 110.000 9.470 112.685 ;
        RECT 10.310 110.000 12.230 112.685 ;
        RECT 13.070 110.000 14.990 112.685 ;
        RECT 15.830 110.000 17.750 112.685 ;
        RECT 18.590 110.000 20.510 112.685 ;
        RECT 21.350 110.000 23.270 112.685 ;
        RECT 24.110 110.000 26.030 112.685 ;
        RECT 26.870 110.000 28.790 112.685 ;
        RECT 29.630 110.000 32.010 112.685 ;
        RECT 32.850 110.000 34.770 112.685 ;
        RECT 35.610 110.000 37.530 112.685 ;
        RECT 38.370 110.000 40.290 112.685 ;
        RECT 41.130 110.000 43.050 112.685 ;
        RECT 43.890 110.000 45.810 112.685 ;
        RECT 46.650 110.000 48.570 112.685 ;
        RECT 49.410 110.000 51.330 112.685 ;
        RECT 52.170 110.000 54.090 112.685 ;
        RECT 54.930 110.000 56.850 112.685 ;
        RECT 57.690 110.000 60.070 112.685 ;
        RECT 60.910 110.000 62.830 112.685 ;
        RECT 63.670 110.000 65.590 112.685 ;
        RECT 66.430 110.000 68.350 112.685 ;
        RECT 69.190 110.000 71.110 112.685 ;
        RECT 71.950 110.000 73.870 112.685 ;
        RECT 74.710 110.000 76.630 112.685 ;
        RECT 77.470 110.000 79.390 112.685 ;
        RECT 80.230 110.000 82.150 112.685 ;
        RECT 82.990 110.000 84.910 112.685 ;
        RECT 85.750 110.000 88.130 112.685 ;
        RECT 88.970 110.000 90.890 112.685 ;
        RECT 91.730 110.000 93.650 112.685 ;
        RECT 94.490 110.000 96.410 112.685 ;
        RECT 97.250 110.000 99.170 112.685 ;
        RECT 100.010 110.000 101.930 112.685 ;
        RECT 102.770 110.000 104.690 112.685 ;
        RECT 105.530 110.000 107.450 112.685 ;
        RECT 108.290 110.000 110.210 112.685 ;
        RECT 111.050 110.000 112.970 112.685 ;
        RECT 1.480 0.115 113.520 110.000 ;
      LAYER met3 ;
        RECT 4.000 111.800 110.600 112.665 ;
        RECT 4.000 111.160 111.000 111.800 ;
        RECT 4.000 109.760 110.600 111.160 ;
        RECT 4.000 108.440 111.000 109.760 ;
        RECT 4.000 107.040 110.600 108.440 ;
        RECT 4.000 106.400 111.000 107.040 ;
        RECT 4.000 105.000 110.600 106.400 ;
        RECT 4.000 104.360 111.000 105.000 ;
        RECT 4.000 102.960 110.600 104.360 ;
        RECT 4.000 101.640 111.000 102.960 ;
        RECT 4.000 100.240 110.600 101.640 ;
        RECT 4.000 99.600 111.000 100.240 ;
        RECT 4.000 98.200 110.600 99.600 ;
        RECT 4.000 96.880 111.000 98.200 ;
        RECT 4.000 95.480 110.600 96.880 ;
        RECT 4.000 94.840 111.000 95.480 ;
        RECT 4.000 93.440 110.600 94.840 ;
        RECT 4.000 92.800 111.000 93.440 ;
        RECT 4.000 91.400 110.600 92.800 ;
        RECT 4.000 90.080 111.000 91.400 ;
        RECT 4.000 88.680 110.600 90.080 ;
        RECT 4.000 88.040 111.000 88.680 ;
        RECT 4.000 86.640 110.600 88.040 ;
        RECT 4.000 86.000 111.000 86.640 ;
        RECT 4.400 84.600 110.600 86.000 ;
        RECT 4.000 83.280 111.000 84.600 ;
        RECT 4.000 81.880 110.600 83.280 ;
        RECT 4.000 81.240 111.000 81.880 ;
        RECT 4.000 79.840 110.600 81.240 ;
        RECT 4.000 78.520 111.000 79.840 ;
        RECT 4.000 77.120 110.600 78.520 ;
        RECT 4.000 76.480 111.000 77.120 ;
        RECT 4.000 75.080 110.600 76.480 ;
        RECT 4.000 74.440 111.000 75.080 ;
        RECT 4.000 73.040 110.600 74.440 ;
        RECT 4.000 71.720 111.000 73.040 ;
        RECT 4.000 70.320 110.600 71.720 ;
        RECT 4.000 69.680 111.000 70.320 ;
        RECT 4.000 68.280 110.600 69.680 ;
        RECT 4.000 67.640 111.000 68.280 ;
        RECT 4.000 66.240 110.600 67.640 ;
        RECT 4.000 64.920 111.000 66.240 ;
        RECT 4.000 63.520 110.600 64.920 ;
        RECT 4.000 62.880 111.000 63.520 ;
        RECT 4.000 61.480 110.600 62.880 ;
        RECT 4.000 60.160 111.000 61.480 ;
        RECT 4.000 58.760 110.600 60.160 ;
        RECT 4.000 58.120 111.000 58.760 ;
        RECT 4.000 56.720 110.600 58.120 ;
        RECT 4.000 56.080 111.000 56.720 ;
        RECT 4.000 54.680 110.600 56.080 ;
        RECT 4.000 53.360 111.000 54.680 ;
        RECT 4.000 51.960 110.600 53.360 ;
        RECT 4.000 51.320 111.000 51.960 ;
        RECT 4.000 49.920 110.600 51.320 ;
        RECT 4.000 48.600 111.000 49.920 ;
        RECT 4.000 47.200 110.600 48.600 ;
        RECT 4.000 46.560 111.000 47.200 ;
        RECT 4.000 45.160 110.600 46.560 ;
        RECT 4.000 44.520 111.000 45.160 ;
        RECT 4.000 43.120 110.600 44.520 ;
        RECT 4.000 41.800 111.000 43.120 ;
        RECT 4.000 40.400 110.600 41.800 ;
        RECT 4.000 39.760 111.000 40.400 ;
        RECT 4.000 38.360 110.600 39.760 ;
        RECT 4.000 37.720 111.000 38.360 ;
        RECT 4.000 36.320 110.600 37.720 ;
        RECT 4.000 35.000 111.000 36.320 ;
        RECT 4.000 33.600 110.600 35.000 ;
        RECT 4.000 32.960 111.000 33.600 ;
        RECT 4.000 31.560 110.600 32.960 ;
        RECT 4.000 30.240 111.000 31.560 ;
        RECT 4.000 28.880 110.600 30.240 ;
        RECT 4.400 28.840 110.600 28.880 ;
        RECT 4.400 28.200 111.000 28.840 ;
        RECT 4.400 27.480 110.600 28.200 ;
        RECT 4.000 26.800 110.600 27.480 ;
        RECT 4.000 26.160 111.000 26.800 ;
        RECT 4.000 24.760 110.600 26.160 ;
        RECT 4.000 23.440 111.000 24.760 ;
        RECT 4.000 22.040 110.600 23.440 ;
        RECT 4.000 21.400 111.000 22.040 ;
        RECT 4.000 20.000 110.600 21.400 ;
        RECT 4.000 19.360 111.000 20.000 ;
        RECT 4.000 17.960 110.600 19.360 ;
        RECT 4.000 16.640 111.000 17.960 ;
        RECT 4.000 15.240 110.600 16.640 ;
        RECT 4.000 14.600 111.000 15.240 ;
        RECT 4.000 13.200 110.600 14.600 ;
        RECT 4.000 11.880 111.000 13.200 ;
        RECT 4.000 10.480 110.600 11.880 ;
        RECT 4.000 9.840 111.000 10.480 ;
        RECT 4.000 8.440 110.600 9.840 ;
        RECT 4.000 7.800 111.000 8.440 ;
        RECT 4.000 6.400 110.600 7.800 ;
        RECT 4.000 5.080 111.000 6.400 ;
        RECT 4.000 3.680 110.600 5.080 ;
        RECT 4.000 3.040 111.000 3.680 ;
        RECT 4.000 1.640 110.600 3.040 ;
        RECT 4.000 1.000 111.000 1.640 ;
        RECT 4.000 0.135 110.600 1.000 ;
      LAYER met4 ;
        RECT 41.375 9.920 56.300 102.880 ;
        RECT 58.700 9.920 73.625 102.880 ;
        RECT 76.025 9.920 90.955 102.880 ;
  END
END sb_0__0_
END LIBRARY

